magic
tech sky130A
magscale 1 2
timestamp 1682506875
<< viali >>
rect 18981 54281 19015 54315
rect 24501 54281 24535 54315
rect 18153 54213 18187 54247
rect 2237 54145 2271 54179
rect 4169 54145 4203 54179
rect 6745 54145 6779 54179
rect 13737 54145 13771 54179
rect 14105 54145 14139 54179
rect 15117 54145 15151 54179
rect 15393 54145 15427 54179
rect 17049 54145 17083 54179
rect 17325 54145 17359 54179
rect 17877 54145 17911 54179
rect 19717 54145 19751 54179
rect 23305 54145 23339 54179
rect 23765 54145 23799 54179
rect 24777 54145 24811 54179
rect 25053 54145 25087 54179
rect 2513 54077 2547 54111
rect 4445 54077 4479 54111
rect 7113 54077 7147 54111
rect 19441 54077 19475 54111
rect 23949 54009 23983 54043
rect 13553 53941 13587 53975
rect 14933 53941 14967 53975
rect 16865 53941 16899 53975
rect 17693 53941 17727 53975
rect 23121 53941 23155 53975
rect 25237 53941 25271 53975
rect 23489 53737 23523 53771
rect 2053 53601 2087 53635
rect 5733 53601 5767 53635
rect 1777 53533 1811 53567
rect 5457 53533 5491 53567
rect 23857 53533 23891 53567
rect 24409 53533 24443 53567
rect 24685 53533 24719 53567
rect 25053 53533 25087 53567
rect 23949 53397 23983 53431
rect 25237 53397 25271 53431
rect 4997 53193 5031 53227
rect 6561 53193 6595 53227
rect 5181 53057 5215 53091
rect 6745 53057 6779 53091
rect 24777 53057 24811 53091
rect 25053 53057 25087 53091
rect 25237 52853 25271 52887
rect 7665 52649 7699 52683
rect 7849 52445 7883 52479
rect 24593 52445 24627 52479
rect 25329 52445 25363 52479
rect 24961 52377 24995 52411
rect 8861 52105 8895 52139
rect 8769 51969 8803 52003
rect 25513 51765 25547 51799
rect 7665 51561 7699 51595
rect 8033 51561 8067 51595
rect 8493 51561 8527 51595
rect 7573 51357 7607 51391
rect 24961 51357 24995 51391
rect 25053 51221 25087 51255
rect 24593 50881 24627 50915
rect 24961 50881 24995 50915
rect 25053 50677 25087 50711
rect 25513 50133 25547 50167
rect 24501 49793 24535 49827
rect 24777 49725 24811 49759
rect 8401 49385 8435 49419
rect 9413 49385 9447 49419
rect 9781 49385 9815 49419
rect 10149 49317 10183 49351
rect 6653 49249 6687 49283
rect 9321 49181 9355 49215
rect 6929 49113 6963 49147
rect 8953 49113 8987 49147
rect 24777 49113 24811 49147
rect 25145 49113 25179 49147
rect 8769 49045 8803 49079
rect 25237 49045 25271 49079
rect 7941 48773 7975 48807
rect 10276 48705 10310 48739
rect 7757 48637 7791 48671
rect 8401 48637 8435 48671
rect 10379 48501 10413 48535
rect 25421 48501 25455 48535
rect 9781 48229 9815 48263
rect 9137 48093 9171 48127
rect 11564 48093 11598 48127
rect 25145 48093 25179 48127
rect 11667 47957 11701 47991
rect 25237 47957 25271 47991
rect 8861 47685 8895 47719
rect 12817 47685 12851 47719
rect 12633 47617 12667 47651
rect 24869 47617 24903 47651
rect 25329 47617 25363 47651
rect 8677 47549 8711 47583
rect 9321 47549 9355 47583
rect 14473 47549 14507 47583
rect 25145 47413 25179 47447
rect 10609 47209 10643 47243
rect 11161 47209 11195 47243
rect 10793 47141 10827 47175
rect 14289 47073 14323 47107
rect 10333 47005 10367 47039
rect 12576 47005 12610 47039
rect 13404 47005 13438 47039
rect 13507 47005 13541 47039
rect 12679 46937 12713 46971
rect 14473 46937 14507 46971
rect 16129 46937 16163 46971
rect 25421 46869 25455 46903
rect 10609 46665 10643 46699
rect 14657 46597 14691 46631
rect 25329 46529 25363 46563
rect 8861 46461 8895 46495
rect 9137 46461 9171 46495
rect 14473 46461 14507 46495
rect 16313 46461 16347 46495
rect 11069 46393 11103 46427
rect 10977 46325 11011 46359
rect 25145 46325 25179 46359
rect 25145 46053 25179 46087
rect 10609 45985 10643 46019
rect 12081 45985 12115 46019
rect 15853 45985 15887 46019
rect 10425 45917 10459 45951
rect 15669 45917 15703 45951
rect 24869 45917 24903 45951
rect 25329 45917 25363 45951
rect 17509 45849 17543 45883
rect 9505 45509 9539 45543
rect 9321 45373 9355 45407
rect 10885 45373 10919 45407
rect 25421 45237 25455 45271
rect 10609 45033 10643 45067
rect 11345 45033 11379 45067
rect 11529 45033 11563 45067
rect 20729 44897 20763 44931
rect 22477 44897 22511 44931
rect 9965 44829 9999 44863
rect 11069 44829 11103 44863
rect 11897 44829 11931 44863
rect 20453 44829 20487 44863
rect 25329 44829 25363 44863
rect 22201 44693 22235 44727
rect 25145 44693 25179 44727
rect 24777 44353 24811 44387
rect 25145 44353 25179 44387
rect 25329 44217 25363 44251
rect 25513 43605 25547 43639
rect 11161 43401 11195 43435
rect 25145 43333 25179 43367
rect 11713 43265 11747 43299
rect 9413 43197 9447 43231
rect 9689 43197 9723 43231
rect 25329 43129 25363 43163
rect 11621 43061 11655 43095
rect 24777 42585 24811 42619
rect 25145 42585 25179 42619
rect 25329 42585 25363 42619
rect 25421 41973 25455 42007
rect 25145 41565 25179 41599
rect 25329 41497 25363 41531
rect 24869 41089 24903 41123
rect 25329 41089 25363 41123
rect 25145 40885 25179 40919
rect 25421 40341 25455 40375
rect 12357 40137 12391 40171
rect 25145 40137 25179 40171
rect 11713 40001 11747 40035
rect 25329 40001 25363 40035
rect 9137 39593 9171 39627
rect 9321 39389 9355 39423
rect 24869 39389 24903 39423
rect 25329 39389 25363 39423
rect 25145 39253 25179 39287
rect 25421 38709 25455 38743
rect 17693 38301 17727 38335
rect 25329 38301 25363 38335
rect 18337 38165 18371 38199
rect 25145 38165 25179 38199
rect 24777 37825 24811 37859
rect 25145 37825 25179 37859
rect 25329 37689 25363 37723
rect 24869 37213 24903 37247
rect 25329 37213 25363 37247
rect 25145 37077 25179 37111
rect 11161 36873 11195 36907
rect 11713 36873 11747 36907
rect 24777 36737 24811 36771
rect 25145 36737 25179 36771
rect 9413 36669 9447 36703
rect 9689 36669 9723 36703
rect 25329 36601 25363 36635
rect 11621 36533 11655 36567
rect 9137 36329 9171 36363
rect 9321 36125 9355 36159
rect 25329 36125 25363 36159
rect 24869 35989 24903 36023
rect 25145 35989 25179 36023
rect 20361 35785 20395 35819
rect 21097 35785 21131 35819
rect 21189 35785 21223 35819
rect 22477 35785 22511 35819
rect 25145 35785 25179 35819
rect 22385 35649 22419 35683
rect 25329 35649 25363 35683
rect 21281 35581 21315 35615
rect 22569 35581 22603 35615
rect 20729 35513 20763 35547
rect 22017 35445 22051 35479
rect 24869 35445 24903 35479
rect 22385 35241 22419 35275
rect 24869 35241 24903 35275
rect 21373 35173 21407 35207
rect 21833 35173 21867 35207
rect 25145 35173 25179 35207
rect 23305 35105 23339 35139
rect 19625 35037 19659 35071
rect 23121 35037 23155 35071
rect 23213 35037 23247 35071
rect 25329 35037 25363 35071
rect 24501 34969 24535 35003
rect 20269 34901 20303 34935
rect 22753 34901 22787 34935
rect 24593 34901 24627 34935
rect 24501 34697 24535 34731
rect 15853 34629 15887 34663
rect 15117 34561 15151 34595
rect 19441 34561 19475 34595
rect 20821 34561 20855 34595
rect 22017 34561 22051 34595
rect 23121 34561 23155 34595
rect 24685 34561 24719 34595
rect 25329 34561 25363 34595
rect 16405 34493 16439 34527
rect 20085 34493 20119 34527
rect 21465 34493 21499 34527
rect 22661 34493 22695 34527
rect 24225 34493 24259 34527
rect 23765 34357 23799 34391
rect 25145 34357 25179 34391
rect 21189 34153 21223 34187
rect 23397 34153 23431 34187
rect 21649 34017 21683 34051
rect 18061 33949 18095 33983
rect 19441 33949 19475 33983
rect 24593 33949 24627 33983
rect 17233 33881 17267 33915
rect 19717 33881 19751 33915
rect 21925 33881 21959 33915
rect 25237 33881 25271 33915
rect 16865 33813 16899 33847
rect 23673 33813 23707 33847
rect 23857 33813 23891 33847
rect 24133 33813 24167 33847
rect 10057 33609 10091 33643
rect 21189 33609 21223 33643
rect 21465 33609 21499 33643
rect 24593 33609 24627 33643
rect 24685 33609 24719 33643
rect 25329 33541 25363 33575
rect 9413 33473 9447 33507
rect 19441 33473 19475 33507
rect 22017 33473 22051 33507
rect 19717 33405 19751 33439
rect 22293 33405 22327 33439
rect 24777 33405 24811 33439
rect 23765 33269 23799 33303
rect 24225 33269 24259 33303
rect 9137 33065 9171 33099
rect 21465 33065 21499 33099
rect 24041 33065 24075 33099
rect 19717 32929 19751 32963
rect 22293 32929 22327 32963
rect 25053 32929 25087 32963
rect 25145 32929 25179 32963
rect 9321 32861 9355 32895
rect 18153 32861 18187 32895
rect 19441 32861 19475 32895
rect 22569 32793 22603 32827
rect 24961 32793 24995 32827
rect 18797 32725 18831 32759
rect 21189 32725 21223 32759
rect 24593 32725 24627 32759
rect 8953 32521 8987 32555
rect 16037 32521 16071 32555
rect 16957 32521 16991 32555
rect 17141 32521 17175 32555
rect 15945 32453 15979 32487
rect 17693 32453 17727 32487
rect 20821 32453 20855 32487
rect 22845 32453 22879 32487
rect 9137 32385 9171 32419
rect 17417 32385 17451 32419
rect 19809 32385 19843 32419
rect 20085 32385 20119 32419
rect 21557 32385 21591 32419
rect 22109 32385 22143 32419
rect 23489 32385 23523 32419
rect 16221 32317 16255 32351
rect 16773 32317 16807 32351
rect 19533 32317 19567 32351
rect 23765 32317 23799 32351
rect 15577 32181 15611 32215
rect 19165 32181 19199 32215
rect 25237 32181 25271 32215
rect 18613 31977 18647 32011
rect 25237 31977 25271 32011
rect 15669 31909 15703 31943
rect 16129 31841 16163 31875
rect 16313 31841 16347 31875
rect 16865 31841 16899 31875
rect 19441 31841 19475 31875
rect 19717 31841 19751 31875
rect 22109 31841 22143 31875
rect 22201 31841 22235 31875
rect 15025 31773 15059 31807
rect 22845 31773 22879 31807
rect 23489 31773 23523 31807
rect 24593 31773 24627 31807
rect 14289 31705 14323 31739
rect 17141 31705 17175 31739
rect 18981 31705 19015 31739
rect 16037 31637 16071 31671
rect 21189 31637 21223 31671
rect 21649 31637 21683 31671
rect 22017 31637 22051 31671
rect 24133 31637 24167 31671
rect 17693 31433 17727 31467
rect 20637 31433 20671 31467
rect 21557 31433 21591 31467
rect 25329 31433 25363 31467
rect 21373 31365 21407 31399
rect 13277 31297 13311 31331
rect 17049 31297 17083 31331
rect 19073 31297 19107 31331
rect 20545 31297 20579 31331
rect 24685 31297 24719 31331
rect 13553 31229 13587 31263
rect 20729 31229 20763 31263
rect 22477 31229 22511 31263
rect 22753 31229 22787 31263
rect 20177 31161 20211 31195
rect 15025 31093 15059 31127
rect 15485 31093 15519 31127
rect 15669 31093 15703 31127
rect 16773 31093 16807 31127
rect 19717 31093 19751 31127
rect 24225 31093 24259 31127
rect 18613 30889 18647 30923
rect 18889 30889 18923 30923
rect 20361 30889 20395 30923
rect 23581 30889 23615 30923
rect 16865 30753 16899 30787
rect 20729 30753 20763 30787
rect 21005 30753 21039 30787
rect 14197 30685 14231 30719
rect 19441 30685 19475 30719
rect 22937 30685 22971 30719
rect 24593 30685 24627 30719
rect 14473 30617 14507 30651
rect 15209 30617 15243 30651
rect 17141 30617 17175 30651
rect 20085 30617 20119 30651
rect 25237 30617 25271 30651
rect 15761 30549 15795 30583
rect 22477 30549 22511 30583
rect 23949 30549 23983 30583
rect 24225 30549 24259 30583
rect 20361 30277 20395 30311
rect 22477 30277 22511 30311
rect 23581 30277 23615 30311
rect 25329 30277 25363 30311
rect 10057 30209 10091 30243
rect 14473 30209 14507 30243
rect 15945 30209 15979 30243
rect 17325 30209 17359 30243
rect 19257 30209 19291 30243
rect 20269 30209 20303 30243
rect 21281 30209 21315 30243
rect 22385 30209 22419 30243
rect 10149 30141 10183 30175
rect 10241 30141 10275 30175
rect 12265 30141 12299 30175
rect 12541 30141 12575 30175
rect 15117 30141 15151 30175
rect 16037 30141 16071 30175
rect 16129 30141 16163 30175
rect 20453 30141 20487 30175
rect 22661 30141 22695 30175
rect 23305 30141 23339 30175
rect 25053 30141 25087 30175
rect 9689 30073 9723 30107
rect 16865 30073 16899 30107
rect 14013 30005 14047 30039
rect 15577 30005 15611 30039
rect 16773 30005 16807 30039
rect 17969 30005 18003 30039
rect 19901 30005 19935 30039
rect 22017 30005 22051 30039
rect 11253 29801 11287 29835
rect 13277 29801 13311 29835
rect 19441 29801 19475 29835
rect 11529 29665 11563 29699
rect 14289 29665 14323 29699
rect 17141 29665 17175 29699
rect 17417 29665 17451 29699
rect 19901 29665 19935 29699
rect 19993 29665 20027 29699
rect 21097 29665 21131 29699
rect 21189 29665 21223 29699
rect 22109 29665 22143 29699
rect 24869 29665 24903 29699
rect 9137 29597 9171 29631
rect 22293 29597 22327 29631
rect 22753 29597 22787 29631
rect 24041 29597 24075 29631
rect 25329 29597 25363 29631
rect 9413 29529 9447 29563
rect 11805 29529 11839 29563
rect 14565 29529 14599 29563
rect 16405 29529 16439 29563
rect 21005 29529 21039 29563
rect 24501 29529 24535 29563
rect 10885 29461 10919 29495
rect 13553 29461 13587 29495
rect 16037 29461 16071 29495
rect 16589 29461 16623 29495
rect 18889 29461 18923 29495
rect 19809 29461 19843 29495
rect 20637 29461 20671 29495
rect 22569 29461 22603 29495
rect 23213 29461 23247 29495
rect 23857 29461 23891 29495
rect 24593 29461 24627 29495
rect 25145 29461 25179 29495
rect 13369 29257 13403 29291
rect 13461 29257 13495 29291
rect 14565 29257 14599 29291
rect 14657 29257 14691 29291
rect 15393 29257 15427 29291
rect 15853 29257 15887 29291
rect 16865 29257 16899 29291
rect 17969 29257 18003 29291
rect 18705 29257 18739 29291
rect 18889 29257 18923 29291
rect 19257 29257 19291 29291
rect 23121 29257 23155 29291
rect 23581 29257 23615 29291
rect 24869 29257 24903 29291
rect 20453 29189 20487 29223
rect 21557 29189 21591 29223
rect 23489 29189 23523 29223
rect 10517 29121 10551 29155
rect 11529 29121 11563 29155
rect 11897 29121 11931 29155
rect 15761 29121 15795 29155
rect 16405 29121 16439 29155
rect 17233 29121 17267 29155
rect 18061 29121 18095 29155
rect 22017 29121 22051 29155
rect 25329 29121 25363 29155
rect 13553 29053 13587 29087
rect 14749 29053 14783 29087
rect 15945 29053 15979 29087
rect 17325 29053 17359 29087
rect 17509 29053 17543 29087
rect 19901 29053 19935 29087
rect 23673 29053 23707 29087
rect 24317 29053 24351 29087
rect 11161 28985 11195 29019
rect 13001 28985 13035 29019
rect 14197 28985 14231 29019
rect 22661 28985 22695 29019
rect 25145 28985 25179 29019
rect 12541 28917 12575 28951
rect 11253 28713 11287 28747
rect 13921 28713 13955 28747
rect 18889 28713 18923 28747
rect 14197 28645 14231 28679
rect 24593 28645 24627 28679
rect 9505 28577 9539 28611
rect 11713 28577 11747 28611
rect 11989 28577 12023 28611
rect 15301 28577 15335 28611
rect 16497 28577 16531 28611
rect 17141 28577 17175 28611
rect 19993 28577 20027 28611
rect 20913 28577 20947 28611
rect 25053 28577 25087 28611
rect 25237 28577 25271 28611
rect 15117 28509 15151 28543
rect 19809 28509 19843 28543
rect 20637 28509 20671 28543
rect 9781 28441 9815 28475
rect 17417 28441 17451 28475
rect 22845 28441 22879 28475
rect 23581 28441 23615 28475
rect 24961 28441 24995 28475
rect 13461 28373 13495 28407
rect 14749 28373 14783 28407
rect 15209 28373 15243 28407
rect 15945 28373 15979 28407
rect 16313 28373 16347 28407
rect 16405 28373 16439 28407
rect 19441 28373 19475 28407
rect 19901 28373 19935 28407
rect 22385 28373 22419 28407
rect 24133 28373 24167 28407
rect 11161 28169 11195 28203
rect 12357 28169 12391 28203
rect 12725 28169 12759 28203
rect 13645 28169 13679 28203
rect 15025 28169 15059 28203
rect 19901 28169 19935 28203
rect 24685 28169 24719 28203
rect 25329 28169 25363 28203
rect 13553 28101 13587 28135
rect 18521 28101 18555 28135
rect 10517 28033 10551 28067
rect 11713 28033 11747 28067
rect 14381 28033 14415 28067
rect 15485 28033 15519 28067
rect 17233 28033 17267 28067
rect 17325 28033 17359 28067
rect 18429 28033 18463 28067
rect 19257 28033 19291 28067
rect 20545 28033 20579 28067
rect 24593 28033 24627 28067
rect 13737 27965 13771 27999
rect 17509 27965 17543 27999
rect 18613 27965 18647 27999
rect 21281 27965 21315 27999
rect 22017 27965 22051 27999
rect 22293 27965 22327 27999
rect 24777 27965 24811 27999
rect 16865 27897 16899 27931
rect 20177 27897 20211 27931
rect 24225 27897 24259 27931
rect 13185 27829 13219 27863
rect 16129 27829 16163 27863
rect 16405 27829 16439 27863
rect 18061 27829 18095 27863
rect 23765 27829 23799 27863
rect 25421 27829 25455 27863
rect 14657 27625 14691 27659
rect 20164 27625 20198 27659
rect 11989 27557 12023 27591
rect 25237 27557 25271 27591
rect 10517 27489 10551 27523
rect 13093 27489 13127 27523
rect 16037 27489 16071 27523
rect 18061 27489 18095 27523
rect 19349 27489 19383 27523
rect 22661 27489 22695 27523
rect 23949 27489 23983 27523
rect 10241 27421 10275 27455
rect 12449 27421 12483 27455
rect 15853 27421 15887 27455
rect 18889 27421 18923 27455
rect 19901 27421 19935 27455
rect 22477 27421 22511 27455
rect 23673 27421 23707 27455
rect 23765 27421 23799 27455
rect 24593 27421 24627 27455
rect 15945 27353 15979 27387
rect 16865 27353 16899 27387
rect 17233 27353 17267 27387
rect 22569 27353 22603 27387
rect 15485 27285 15519 27319
rect 16497 27285 16531 27319
rect 17049 27285 17083 27319
rect 17325 27285 17359 27319
rect 17509 27285 17543 27319
rect 17693 27285 17727 27319
rect 18705 27285 18739 27319
rect 21649 27285 21683 27319
rect 22109 27285 22143 27319
rect 23305 27285 23339 27319
rect 11529 27081 11563 27115
rect 12081 27081 12115 27115
rect 14473 27081 14507 27115
rect 21189 27081 21223 27115
rect 25237 27081 25271 27115
rect 25513 27081 25547 27115
rect 15485 27013 15519 27047
rect 9413 26945 9447 26979
rect 15393 26945 15427 26979
rect 16037 26945 16071 26979
rect 20453 26945 20487 26979
rect 21097 26945 21131 26979
rect 22017 26945 22051 26979
rect 9689 26877 9723 26911
rect 12725 26877 12759 26911
rect 13001 26877 13035 26911
rect 15577 26877 15611 26911
rect 17969 26877 18003 26911
rect 18245 26877 18279 26911
rect 21281 26877 21315 26911
rect 23213 26877 23247 26911
rect 23489 26877 23523 26911
rect 19717 26809 19751 26843
rect 19993 26809 20027 26843
rect 11161 26741 11195 26775
rect 15025 26741 15059 26775
rect 16221 26741 16255 26775
rect 20729 26741 20763 26775
rect 22661 26741 22695 26775
rect 24961 26741 24995 26775
rect 10885 26537 10919 26571
rect 15669 26537 15703 26571
rect 19704 26537 19738 26571
rect 11805 26469 11839 26503
rect 13001 26469 13035 26503
rect 24593 26469 24627 26503
rect 9137 26401 9171 26435
rect 9413 26401 9447 26435
rect 12357 26401 12391 26435
rect 13553 26401 13587 26435
rect 14197 26401 14231 26435
rect 15025 26401 15059 26435
rect 16129 26401 16163 26435
rect 16221 26401 16255 26435
rect 16681 26401 16715 26435
rect 18521 26401 18555 26435
rect 19441 26401 19475 26435
rect 21189 26401 21223 26435
rect 23213 26401 23247 26435
rect 25053 26401 25087 26435
rect 25145 26401 25179 26435
rect 11253 26333 11287 26367
rect 12265 26333 12299 26367
rect 16957 26333 16991 26367
rect 18245 26333 18279 26367
rect 23121 26333 23155 26367
rect 12173 26265 12207 26299
rect 13369 26265 13403 26299
rect 13461 26265 13495 26299
rect 14841 26265 14875 26299
rect 14933 26265 14967 26299
rect 21925 26265 21959 26299
rect 22109 26265 22143 26299
rect 23857 26265 23891 26299
rect 14473 26197 14507 26231
rect 16037 26197 16071 26231
rect 17877 26197 17911 26231
rect 18337 26197 18371 26231
rect 21557 26197 21591 26231
rect 22661 26197 22695 26231
rect 23029 26197 23063 26231
rect 24961 26197 24995 26231
rect 15761 25993 15795 26027
rect 16221 25993 16255 26027
rect 18245 25993 18279 26027
rect 20177 25993 20211 26027
rect 22477 25993 22511 26027
rect 25329 25993 25363 26027
rect 21465 25925 21499 25959
rect 23857 25925 23891 25959
rect 10517 25857 10551 25891
rect 12357 25857 12391 25891
rect 14933 25857 14967 25891
rect 17141 25857 17175 25891
rect 17785 25857 17819 25891
rect 19533 25857 19567 25891
rect 20821 25857 20855 25891
rect 22385 25857 22419 25891
rect 23213 25857 23247 25891
rect 12633 25789 12667 25823
rect 15025 25789 15059 25823
rect 15117 25789 15151 25823
rect 18889 25789 18923 25823
rect 22569 25789 22603 25823
rect 23029 25789 23063 25823
rect 23581 25789 23615 25823
rect 14565 25721 14599 25755
rect 16957 25721 16991 25755
rect 11161 25653 11195 25687
rect 14105 25653 14139 25687
rect 16497 25653 16531 25687
rect 17601 25653 17635 25687
rect 20545 25653 20579 25687
rect 22017 25653 22051 25687
rect 10333 25449 10367 25483
rect 13737 25449 13771 25483
rect 25237 25449 25271 25483
rect 11529 25381 11563 25415
rect 10885 25313 10919 25347
rect 12081 25313 12115 25347
rect 14841 25313 14875 25347
rect 18889 25313 18923 25347
rect 10701 25245 10735 25279
rect 13093 25245 13127 25279
rect 17325 25245 17359 25279
rect 18061 25245 18095 25279
rect 19717 25245 19751 25279
rect 20913 25245 20947 25279
rect 21557 25245 21591 25279
rect 22661 25245 22695 25279
rect 24593 25245 24627 25279
rect 11989 25177 12023 25211
rect 14657 25177 14691 25211
rect 15669 25177 15703 25211
rect 18705 25177 18739 25211
rect 23857 25177 23891 25211
rect 10793 25109 10827 25143
rect 11897 25109 11931 25143
rect 14289 25109 14323 25143
rect 14749 25109 14783 25143
rect 15393 25109 15427 25143
rect 17877 25109 17911 25143
rect 19349 25109 19383 25143
rect 20361 25109 20395 25143
rect 21005 25109 21039 25143
rect 22201 25109 22235 25143
rect 14289 24905 14323 24939
rect 15945 24905 15979 24939
rect 18429 24905 18463 24939
rect 19257 24905 19291 24939
rect 25329 24905 25363 24939
rect 8401 24837 8435 24871
rect 11989 24837 12023 24871
rect 17233 24837 17267 24871
rect 19993 24837 20027 24871
rect 22477 24837 22511 24871
rect 11253 24769 11287 24803
rect 14381 24769 14415 24803
rect 15301 24769 15335 24803
rect 22569 24769 22603 24803
rect 8493 24701 8527 24735
rect 8585 24701 8619 24735
rect 9229 24701 9263 24735
rect 9505 24701 9539 24735
rect 11713 24701 11747 24735
rect 14473 24701 14507 24735
rect 16037 24701 16071 24735
rect 16129 24701 16163 24735
rect 17325 24701 17359 24735
rect 17417 24701 17451 24735
rect 18521 24701 18555 24735
rect 18613 24701 18647 24735
rect 19717 24701 19751 24735
rect 21465 24701 21499 24735
rect 22753 24701 22787 24735
rect 23581 24701 23615 24735
rect 23857 24701 23891 24735
rect 8033 24565 8067 24599
rect 10977 24565 11011 24599
rect 13461 24565 13495 24599
rect 13921 24565 13955 24599
rect 15577 24565 15611 24599
rect 16865 24565 16899 24599
rect 18061 24565 18095 24599
rect 19073 24565 19107 24599
rect 22109 24565 22143 24599
rect 23213 24565 23247 24599
rect 8585 24361 8619 24395
rect 12357 24361 12391 24395
rect 13737 24361 13771 24395
rect 16405 24361 16439 24395
rect 16865 24361 16899 24395
rect 21189 24361 21223 24395
rect 21465 24361 21499 24395
rect 16129 24293 16163 24327
rect 23949 24293 23983 24327
rect 6837 24225 6871 24259
rect 10885 24225 10919 24259
rect 18613 24225 18647 24259
rect 18797 24225 18831 24259
rect 21925 24225 21959 24259
rect 9505 24157 9539 24191
rect 10609 24157 10643 24191
rect 12817 24157 12851 24191
rect 16313 24157 16347 24191
rect 17049 24157 17083 24191
rect 17693 24157 17727 24191
rect 18521 24157 18555 24191
rect 19441 24157 19475 24191
rect 24593 24157 24627 24191
rect 7113 24089 7147 24123
rect 8953 24089 8987 24123
rect 13461 24089 13495 24123
rect 19717 24089 19751 24123
rect 22201 24089 22235 24123
rect 9229 24021 9263 24055
rect 10149 24021 10183 24055
rect 17509 24021 17543 24055
rect 18153 24021 18187 24055
rect 23673 24021 23707 24055
rect 24133 24021 24167 24055
rect 25237 24021 25271 24055
rect 12541 23817 12575 23851
rect 13461 23817 13495 23851
rect 13921 23817 13955 23851
rect 15117 23817 15151 23851
rect 16405 23817 16439 23851
rect 18889 23817 18923 23851
rect 22661 23817 22695 23851
rect 8861 23749 8895 23783
rect 20913 23749 20947 23783
rect 23489 23749 23523 23783
rect 8585 23681 8619 23715
rect 13829 23681 13863 23715
rect 15025 23681 15059 23715
rect 15853 23681 15887 23715
rect 17233 23681 17267 23715
rect 18245 23681 18279 23715
rect 19625 23681 19659 23715
rect 19717 23681 19751 23715
rect 20821 23681 20855 23715
rect 22017 23681 22051 23715
rect 10333 23613 10367 23647
rect 14013 23613 14047 23647
rect 15209 23613 15243 23647
rect 17325 23613 17359 23647
rect 17417 23613 17451 23647
rect 18705 23613 18739 23647
rect 19901 23613 19935 23647
rect 21005 23613 21039 23647
rect 23213 23613 23247 23647
rect 24961 23613 24995 23647
rect 18521 23545 18555 23579
rect 10609 23477 10643 23511
rect 14657 23477 14691 23511
rect 16865 23477 16899 23511
rect 18061 23477 18095 23511
rect 19257 23477 19291 23511
rect 20453 23477 20487 23511
rect 21557 23477 21591 23511
rect 25237 23477 25271 23511
rect 25421 23477 25455 23511
rect 11253 23273 11287 23307
rect 14197 23273 14231 23307
rect 18981 23273 19015 23307
rect 14381 23205 14415 23239
rect 17877 23205 17911 23239
rect 20821 23205 20855 23239
rect 13553 23137 13587 23171
rect 15301 23137 15335 23171
rect 18337 23137 18371 23171
rect 18429 23137 18463 23171
rect 20085 23137 20119 23171
rect 23765 23137 23799 23171
rect 25053 23137 25087 23171
rect 25237 23137 25271 23171
rect 9505 23069 9539 23103
rect 10609 23069 10643 23103
rect 13461 23069 13495 23103
rect 19901 23069 19935 23103
rect 21005 23069 21039 23103
rect 21557 23069 21591 23103
rect 22845 23069 22879 23103
rect 24961 23069 24995 23103
rect 13369 23001 13403 23035
rect 18245 23001 18279 23035
rect 10149 22933 10183 22967
rect 13001 22933 13035 22967
rect 19533 22933 19567 22967
rect 19993 22933 20027 22967
rect 22201 22933 22235 22967
rect 24593 22933 24627 22967
rect 10241 22729 10275 22763
rect 11805 22729 11839 22763
rect 18705 22729 18739 22763
rect 21097 22729 21131 22763
rect 8493 22661 8527 22695
rect 15761 22661 15795 22695
rect 18429 22661 18463 22695
rect 21189 22661 21223 22695
rect 23305 22661 23339 22695
rect 8217 22593 8251 22627
rect 12173 22593 12207 22627
rect 17049 22593 17083 22627
rect 19993 22593 20027 22627
rect 22109 22593 22143 22627
rect 23949 22593 23983 22627
rect 12265 22525 12299 22559
rect 12357 22525 12391 22559
rect 13461 22525 13495 22559
rect 13737 22525 13771 22559
rect 15945 22525 15979 22559
rect 18613 22525 18647 22559
rect 19349 22525 19383 22559
rect 21281 22525 21315 22559
rect 24777 22525 24811 22559
rect 16865 22457 16899 22491
rect 9965 22389 9999 22423
rect 12817 22389 12851 22423
rect 15209 22389 15243 22423
rect 18245 22389 18279 22423
rect 18981 22389 19015 22423
rect 20729 22389 20763 22423
rect 7100 22185 7134 22219
rect 23305 22185 23339 22219
rect 23857 22185 23891 22219
rect 18429 22117 18463 22151
rect 6837 22049 6871 22083
rect 8953 22049 8987 22083
rect 10701 22049 10735 22083
rect 11897 22049 11931 22083
rect 13001 22049 13035 22083
rect 13185 22049 13219 22083
rect 15393 22049 15427 22083
rect 15485 22049 15519 22083
rect 16129 22049 16163 22083
rect 16405 22049 16439 22083
rect 20177 22049 20211 22083
rect 20361 22049 20395 22083
rect 20913 22049 20947 22083
rect 21557 22049 21591 22083
rect 25053 22049 25087 22083
rect 25237 22049 25271 22083
rect 11713 21981 11747 22015
rect 11805 21981 11839 22015
rect 18705 21981 18739 22015
rect 24041 21981 24075 22015
rect 10517 21913 10551 21947
rect 12909 21913 12943 21947
rect 21833 21913 21867 21947
rect 24961 21913 24995 21947
rect 8585 21845 8619 21879
rect 9505 21845 9539 21879
rect 10149 21845 10183 21879
rect 10609 21845 10643 21879
rect 11345 21845 11379 21879
rect 12541 21845 12575 21879
rect 14933 21845 14967 21879
rect 15301 21845 15335 21879
rect 17877 21845 17911 21879
rect 18245 21845 18279 21879
rect 19349 21845 19383 21879
rect 19717 21845 19751 21879
rect 20085 21845 20119 21879
rect 24593 21845 24627 21879
rect 10333 21641 10367 21675
rect 10701 21641 10735 21675
rect 15669 21641 15703 21675
rect 19257 21641 19291 21675
rect 22477 21641 22511 21675
rect 25053 21641 25087 21675
rect 9873 21573 9907 21607
rect 19349 21573 19383 21607
rect 11713 21505 11747 21539
rect 15025 21505 15059 21539
rect 16865 21505 16899 21539
rect 18429 21505 18463 21539
rect 20269 21505 20303 21539
rect 22385 21505 22419 21539
rect 23305 21505 23339 21539
rect 7573 21437 7607 21471
rect 7849 21437 7883 21471
rect 9597 21437 9631 21471
rect 10793 21437 10827 21471
rect 10885 21437 10919 21471
rect 12817 21437 12851 21471
rect 13093 21437 13127 21471
rect 14565 21437 14599 21471
rect 19533 21437 19567 21471
rect 21281 21437 21315 21471
rect 22661 21437 22695 21471
rect 23581 21437 23615 21471
rect 17877 21369 17911 21403
rect 12357 21301 12391 21335
rect 17509 21301 17543 21335
rect 18245 21301 18279 21335
rect 18889 21301 18923 21335
rect 22017 21301 22051 21335
rect 25329 21301 25363 21335
rect 8585 21097 8619 21131
rect 9689 21097 9723 21131
rect 16957 21097 16991 21131
rect 17647 21097 17681 21131
rect 21649 21097 21683 21131
rect 22017 21097 22051 21131
rect 10241 20961 10275 20995
rect 11161 20961 11195 20995
rect 13369 20961 13403 20995
rect 15485 20961 15519 20995
rect 17417 20961 17451 20995
rect 19993 20961 20027 20995
rect 21281 20961 21315 20995
rect 23857 20961 23891 20995
rect 25053 20961 25087 20995
rect 25145 20961 25179 20995
rect 7941 20893 7975 20927
rect 10057 20893 10091 20927
rect 15209 20893 15243 20927
rect 18889 20893 18923 20927
rect 19809 20893 19843 20927
rect 21005 20893 21039 20927
rect 22201 20893 22235 20927
rect 22661 20893 22695 20927
rect 11437 20825 11471 20859
rect 13829 20825 13863 20859
rect 14657 20825 14691 20859
rect 14841 20825 14875 20859
rect 9413 20757 9447 20791
rect 10149 20757 10183 20791
rect 12909 20757 12943 20791
rect 18705 20757 18739 20791
rect 19441 20757 19475 20791
rect 19901 20757 19935 20791
rect 20637 20757 20671 20791
rect 21097 20757 21131 20791
rect 24593 20757 24627 20791
rect 24961 20757 24995 20791
rect 8033 20553 8067 20587
rect 12357 20553 12391 20587
rect 15025 20553 15059 20587
rect 15485 20553 15519 20587
rect 19809 20553 19843 20587
rect 23121 20553 23155 20587
rect 25329 20553 25363 20587
rect 8493 20485 8527 20519
rect 13093 20485 13127 20519
rect 22017 20485 22051 20519
rect 6745 20417 6779 20451
rect 8401 20417 8435 20451
rect 11713 20417 11747 20451
rect 15393 20417 15427 20451
rect 19257 20417 19291 20451
rect 20085 20417 20119 20451
rect 21833 20417 21867 20451
rect 22477 20417 22511 20451
rect 8585 20349 8619 20383
rect 12817 20349 12851 20383
rect 14565 20349 14599 20383
rect 15577 20349 15611 20383
rect 16865 20349 16899 20383
rect 17141 20349 17175 20383
rect 21281 20349 21315 20383
rect 23581 20349 23615 20383
rect 23857 20349 23891 20383
rect 7389 20213 7423 20247
rect 18613 20213 18647 20247
rect 19073 20213 19107 20247
rect 19625 20213 19659 20247
rect 8493 20009 8527 20043
rect 11161 20009 11195 20043
rect 11897 20009 11931 20043
rect 18705 20009 18739 20043
rect 24225 20009 24259 20043
rect 25237 20009 25271 20043
rect 17509 19941 17543 19975
rect 6377 19873 6411 19907
rect 10885 19873 10919 19907
rect 12449 19873 12483 19907
rect 16037 19873 16071 19907
rect 17969 19873 18003 19907
rect 18061 19873 18095 19907
rect 19901 19873 19935 19907
rect 9137 19805 9171 19839
rect 12357 19805 12391 19839
rect 14289 19805 14323 19839
rect 16865 19805 16899 19839
rect 18889 19805 18923 19839
rect 22109 19805 22143 19839
rect 24593 19805 24627 19839
rect 6653 19737 6687 19771
rect 9413 19737 9447 19771
rect 12265 19737 12299 19771
rect 14565 19737 14599 19771
rect 20177 19737 20211 19771
rect 22385 19737 22419 19771
rect 8125 19669 8159 19703
rect 16313 19669 16347 19703
rect 16681 19669 16715 19703
rect 17877 19669 17911 19703
rect 19441 19669 19475 19703
rect 19625 19669 19659 19703
rect 21649 19669 21683 19703
rect 23857 19669 23891 19703
rect 9229 19465 9263 19499
rect 9505 19465 9539 19499
rect 10149 19465 10183 19499
rect 10609 19465 10643 19499
rect 14105 19465 14139 19499
rect 15669 19465 15703 19499
rect 16865 19465 16899 19499
rect 17325 19465 17359 19499
rect 18797 19465 18831 19499
rect 20085 19465 20119 19499
rect 20453 19465 20487 19499
rect 20545 19465 20579 19499
rect 22201 19465 22235 19499
rect 22661 19465 22695 19499
rect 7481 19329 7515 19363
rect 9873 19329 9907 19363
rect 10517 19329 10551 19363
rect 12357 19329 12391 19363
rect 14565 19329 14599 19363
rect 15209 19329 15243 19363
rect 15853 19329 15887 19363
rect 17233 19329 17267 19363
rect 18153 19329 18187 19363
rect 19441 19329 19475 19363
rect 21465 19329 21499 19363
rect 22569 19329 22603 19363
rect 7757 19261 7791 19295
rect 10701 19261 10735 19295
rect 11161 19261 11195 19295
rect 12633 19261 12667 19295
rect 17417 19261 17451 19295
rect 20729 19261 20763 19295
rect 22753 19261 22787 19295
rect 23397 19261 23431 19295
rect 23673 19261 23707 19295
rect 11529 19193 11563 19227
rect 21833 19193 21867 19227
rect 25421 19193 25455 19227
rect 19257 19125 19291 19159
rect 19717 19125 19751 19159
rect 21281 19125 21315 19159
rect 25145 19125 25179 19159
rect 9781 18921 9815 18955
rect 25329 18921 25363 18955
rect 10977 18853 11011 18887
rect 14289 18853 14323 18887
rect 17969 18853 18003 18887
rect 21373 18853 21407 18887
rect 6837 18785 6871 18819
rect 7113 18785 7147 18819
rect 10333 18785 10367 18819
rect 11529 18785 11563 18819
rect 14841 18785 14875 18819
rect 17233 18785 17267 18819
rect 17417 18785 17451 18819
rect 18521 18785 18555 18819
rect 21833 18785 21867 18819
rect 23489 18785 23523 18819
rect 16221 18717 16255 18751
rect 18429 18717 18463 18751
rect 19441 18717 19475 18751
rect 20729 18717 20763 18751
rect 22661 18717 22695 18751
rect 24685 18717 24719 18751
rect 10149 18649 10183 18683
rect 10241 18649 10275 18683
rect 11437 18649 11471 18683
rect 12173 18649 12207 18683
rect 12909 18649 12943 18683
rect 14749 18649 14783 18683
rect 8585 18581 8619 18615
rect 9137 18581 9171 18615
rect 11345 18581 11379 18615
rect 13461 18581 13495 18615
rect 13645 18581 13679 18615
rect 13921 18581 13955 18615
rect 14657 18581 14691 18615
rect 16037 18581 16071 18615
rect 16773 18581 16807 18615
rect 17141 18581 17175 18615
rect 18337 18581 18371 18615
rect 18981 18581 19015 18615
rect 20085 18581 20119 18615
rect 20453 18581 20487 18615
rect 22293 18581 22327 18615
rect 7941 18377 7975 18411
rect 11713 18377 11747 18411
rect 13185 18377 13219 18411
rect 13645 18377 13679 18411
rect 15025 18377 15059 18411
rect 22661 18377 22695 18411
rect 9413 18309 9447 18343
rect 11161 18309 11195 18343
rect 17141 18309 17175 18343
rect 18889 18309 18923 18343
rect 21281 18309 21315 18343
rect 23581 18309 23615 18343
rect 8309 18241 8343 18275
rect 13553 18241 13587 18275
rect 14381 18241 14415 18275
rect 15485 18241 15519 18275
rect 16865 18241 16899 18275
rect 19625 18241 19659 18275
rect 20269 18241 20303 18275
rect 22017 18241 22051 18275
rect 8401 18173 8435 18207
rect 8493 18173 8527 18207
rect 9137 18173 9171 18207
rect 13737 18173 13771 18207
rect 15761 18173 15795 18207
rect 23305 18173 23339 18207
rect 25329 18173 25363 18207
rect 12817 18105 12851 18139
rect 20729 18105 20763 18139
rect 22937 18105 22971 18139
rect 18613 18037 18647 18071
rect 19073 18037 19107 18071
rect 19441 18037 19475 18071
rect 20085 18037 20119 18071
rect 20913 18037 20947 18071
rect 21373 18037 21407 18071
rect 8769 17833 8803 17867
rect 9045 17833 9079 17867
rect 11805 17833 11839 17867
rect 21189 17833 21223 17867
rect 21649 17833 21683 17867
rect 7665 17765 7699 17799
rect 11621 17765 11655 17799
rect 13921 17765 13955 17799
rect 17969 17765 18003 17799
rect 8309 17697 8343 17731
rect 10977 17697 11011 17731
rect 14381 17697 14415 17731
rect 18429 17697 18463 17731
rect 18613 17697 18647 17731
rect 18981 17697 19015 17731
rect 23857 17697 23891 17731
rect 25053 17697 25087 17731
rect 25145 17697 25179 17731
rect 10241 17629 10275 17663
rect 12817 17629 12851 17663
rect 16865 17629 16899 17663
rect 19441 17629 19475 17663
rect 22017 17629 22051 17663
rect 22661 17629 22695 17663
rect 8125 17561 8159 17595
rect 17325 17561 17359 17595
rect 19717 17561 19751 17595
rect 7297 17493 7331 17527
rect 8033 17493 8067 17527
rect 11529 17493 11563 17527
rect 13461 17493 13495 17527
rect 15025 17493 15059 17527
rect 15669 17493 15703 17527
rect 16681 17493 16715 17527
rect 18337 17493 18371 17527
rect 22109 17493 22143 17527
rect 24593 17493 24627 17527
rect 24961 17493 24995 17527
rect 8033 17289 8067 17323
rect 9505 17289 9539 17323
rect 10333 17289 10367 17323
rect 11713 17289 11747 17323
rect 12909 17289 12943 17323
rect 13277 17289 13311 17323
rect 21097 17289 21131 17323
rect 21189 17289 21223 17323
rect 10793 17221 10827 17255
rect 17049 17221 17083 17255
rect 17325 17221 17359 17255
rect 19901 17221 19935 17255
rect 23305 17221 23339 17255
rect 6929 17153 6963 17187
rect 10701 17153 10735 17187
rect 12081 17153 12115 17187
rect 14473 17153 14507 17187
rect 18061 17153 18095 17187
rect 18705 17153 18739 17187
rect 20361 17153 20395 17187
rect 22201 17153 22235 17187
rect 23949 17153 23983 17187
rect 9597 17085 9631 17119
rect 9689 17085 9723 17119
rect 10885 17085 10919 17119
rect 12173 17085 12207 17119
rect 12265 17085 12299 17119
rect 13369 17085 13403 17119
rect 13553 17085 13587 17119
rect 14749 17085 14783 17119
rect 21281 17085 21315 17119
rect 24777 17085 24811 17119
rect 13921 17017 13955 17051
rect 16221 17017 16255 17051
rect 19349 17017 19383 17051
rect 7573 16949 7607 16983
rect 8861 16949 8895 16983
rect 9137 16949 9171 16983
rect 16681 16949 16715 16983
rect 19993 16949 20027 16983
rect 20729 16949 20763 16983
rect 7665 16745 7699 16779
rect 8033 16745 8067 16779
rect 11437 16745 11471 16779
rect 17049 16745 17083 16779
rect 18981 16745 19015 16779
rect 13001 16677 13035 16711
rect 14289 16677 14323 16711
rect 18153 16677 18187 16711
rect 5917 16609 5951 16643
rect 10701 16609 10735 16643
rect 10885 16609 10919 16643
rect 12357 16609 12391 16643
rect 13461 16609 13495 16643
rect 13553 16609 13587 16643
rect 14105 16609 14139 16643
rect 15025 16609 15059 16643
rect 15761 16609 15795 16643
rect 15945 16609 15979 16643
rect 15669 16541 15703 16575
rect 17785 16541 17819 16575
rect 18613 16541 18647 16575
rect 19441 16541 19475 16575
rect 20821 16541 20855 16575
rect 21925 16541 21959 16575
rect 22753 16541 22787 16575
rect 24593 16541 24627 16575
rect 25237 16541 25271 16575
rect 6193 16473 6227 16507
rect 9965 16473 9999 16507
rect 12173 16473 12207 16507
rect 16957 16473 16991 16507
rect 20177 16473 20211 16507
rect 23857 16473 23891 16507
rect 10241 16405 10275 16439
rect 10609 16405 10643 16439
rect 11805 16405 11839 16439
rect 12265 16405 12299 16439
rect 13369 16405 13403 16439
rect 15301 16405 15335 16439
rect 17601 16405 17635 16439
rect 18429 16405 18463 16439
rect 21465 16405 21499 16439
rect 14105 16201 14139 16235
rect 16313 16201 16347 16235
rect 19257 16201 19291 16235
rect 25145 16201 25179 16235
rect 7849 16133 7883 16167
rect 9873 16133 9907 16167
rect 16865 16133 16899 16167
rect 17233 16133 17267 16167
rect 17969 16133 18003 16167
rect 19993 16133 20027 16167
rect 25421 16133 25455 16167
rect 7573 16065 7607 16099
rect 11713 16065 11747 16099
rect 14473 16065 14507 16099
rect 15669 16065 15703 16099
rect 18613 16065 18647 16099
rect 24501 16065 24535 16099
rect 9597 15997 9631 16031
rect 11989 15997 12023 16031
rect 14565 15997 14599 16031
rect 14657 15997 14691 16031
rect 19717 15997 19751 16031
rect 22017 15997 22051 16031
rect 13737 15929 13771 15963
rect 21465 15929 21499 15963
rect 24133 15929 24167 15963
rect 13461 15861 13495 15895
rect 17325 15861 17359 15895
rect 22274 15861 22308 15895
rect 23765 15861 23799 15895
rect 8125 15657 8159 15691
rect 8493 15657 8527 15691
rect 13001 15657 13035 15691
rect 17969 15657 18003 15691
rect 9597 15589 9631 15623
rect 6653 15521 6687 15555
rect 11989 15521 12023 15555
rect 12357 15521 12391 15555
rect 13553 15521 13587 15555
rect 15301 15521 15335 15555
rect 16221 15521 16255 15555
rect 19441 15521 19475 15555
rect 22293 15521 22327 15555
rect 22569 15521 22603 15555
rect 25237 15521 25271 15555
rect 6377 15453 6411 15487
rect 9965 15453 9999 15487
rect 18705 15453 18739 15487
rect 21833 15453 21867 15487
rect 24593 15453 24627 15487
rect 10241 15385 10275 15419
rect 13461 15385 13495 15419
rect 14841 15385 14875 15419
rect 16497 15385 16531 15419
rect 19717 15385 19751 15419
rect 12725 15317 12759 15351
rect 13369 15317 13403 15351
rect 14289 15317 14323 15351
rect 15853 15317 15887 15351
rect 18521 15317 18555 15351
rect 21189 15317 21223 15351
rect 21649 15317 21683 15351
rect 24041 15317 24075 15351
rect 7297 15113 7331 15147
rect 10609 15113 10643 15147
rect 11345 15113 11379 15147
rect 13645 15113 13679 15147
rect 14013 15113 14047 15147
rect 19533 15113 19567 15147
rect 19993 15113 20027 15147
rect 21189 15113 21223 15147
rect 21925 15113 21959 15147
rect 22109 15113 22143 15147
rect 9781 15045 9815 15079
rect 12633 15045 12667 15079
rect 18061 15045 18095 15079
rect 18613 15045 18647 15079
rect 6653 14977 6687 15011
rect 11713 14977 11747 15011
rect 14105 14977 14139 15011
rect 14933 14977 14967 15011
rect 15945 14977 15979 15011
rect 19901 14977 19935 15011
rect 21097 14977 21131 15011
rect 22477 14977 22511 15011
rect 23949 14977 23983 15011
rect 7757 14909 7791 14943
rect 8033 14909 8067 14943
rect 10701 14909 10735 14943
rect 10793 14909 10827 14943
rect 13369 14909 13403 14943
rect 14289 14909 14323 14943
rect 16037 14909 16071 14943
rect 16221 14909 16255 14943
rect 16865 14909 16899 14943
rect 17141 14909 17175 14943
rect 20177 14909 20211 14943
rect 21373 14909 21407 14943
rect 24777 14909 24811 14943
rect 10241 14841 10275 14875
rect 12909 14841 12943 14875
rect 15577 14841 15611 14875
rect 12357 14773 12391 14807
rect 13185 14773 13219 14807
rect 18705 14773 18739 14807
rect 20729 14773 20763 14807
rect 23121 14773 23155 14807
rect 23489 14773 23523 14807
rect 23673 14773 23707 14807
rect 8585 14569 8619 14603
rect 9137 14569 9171 14603
rect 11713 14569 11747 14603
rect 14381 14569 14415 14603
rect 18337 14569 18371 14603
rect 19533 14569 19567 14603
rect 20913 14569 20947 14603
rect 15025 14501 15059 14535
rect 21833 14501 21867 14535
rect 9689 14433 9723 14467
rect 11069 14433 11103 14467
rect 12265 14433 12299 14467
rect 13461 14433 13495 14467
rect 13645 14433 13679 14467
rect 15577 14433 15611 14467
rect 17233 14433 17267 14467
rect 22569 14433 22603 14467
rect 7941 14365 7975 14399
rect 10333 14365 10367 14399
rect 14565 14365 14599 14399
rect 17509 14365 17543 14399
rect 18889 14365 18923 14399
rect 19717 14365 19751 14399
rect 20361 14365 20395 14399
rect 21097 14365 21131 14399
rect 22293 14365 22327 14399
rect 24777 14365 24811 14399
rect 12081 14297 12115 14331
rect 13369 14297 13403 14331
rect 21649 14297 21683 14331
rect 9505 14229 9539 14263
rect 9597 14229 9631 14263
rect 12173 14229 12207 14263
rect 13001 14229 13035 14263
rect 15393 14229 15427 14263
rect 15485 14229 15519 14263
rect 16037 14229 16071 14263
rect 16313 14229 16347 14263
rect 16589 14229 16623 14263
rect 18705 14229 18739 14263
rect 20177 14229 20211 14263
rect 24041 14229 24075 14263
rect 24593 14229 24627 14263
rect 25053 14229 25087 14263
rect 9137 14025 9171 14059
rect 10425 14025 10459 14059
rect 12357 14025 12391 14059
rect 12725 14025 12759 14059
rect 15853 14025 15887 14059
rect 18613 14025 18647 14059
rect 8677 13957 8711 13991
rect 10885 13957 10919 13991
rect 16129 13957 16163 13991
rect 19073 13957 19107 13991
rect 23305 13957 23339 13991
rect 25145 13957 25179 13991
rect 6561 13889 6595 13923
rect 9505 13889 9539 13923
rect 9597 13889 9631 13923
rect 10793 13889 10827 13923
rect 11713 13889 11747 13923
rect 12817 13889 12851 13923
rect 15577 13889 15611 13923
rect 20361 13889 20395 13923
rect 20821 13889 20855 13923
rect 21465 13889 21499 13923
rect 22109 13889 22143 13923
rect 23949 13889 23983 13923
rect 8309 13821 8343 13855
rect 9689 13821 9723 13855
rect 11069 13821 11103 13855
rect 12909 13821 12943 13855
rect 13553 13821 13587 13855
rect 15301 13821 15335 13855
rect 16865 13821 16899 13855
rect 19901 13821 19935 13855
rect 6824 13685 6858 13719
rect 13816 13685 13850 13719
rect 17128 13685 17162 13719
rect 20637 13685 20671 13719
rect 21281 13685 21315 13719
rect 7021 13481 7055 13515
rect 16405 13413 16439 13447
rect 7573 13345 7607 13379
rect 12817 13345 12851 13379
rect 14197 13345 14231 13379
rect 15761 13345 15795 13379
rect 16957 13345 16991 13379
rect 20729 13345 20763 13379
rect 22109 13345 22143 13379
rect 9781 13277 9815 13311
rect 11989 13277 12023 13311
rect 13185 13277 13219 13311
rect 13737 13277 13771 13311
rect 16773 13277 16807 13311
rect 17601 13277 17635 13311
rect 18889 13277 18923 13311
rect 22845 13277 22879 13311
rect 24593 13277 24627 13311
rect 7481 13209 7515 13243
rect 10057 13209 10091 13243
rect 14565 13209 14599 13243
rect 19533 13209 19567 13243
rect 21833 13209 21867 13243
rect 21925 13209 21959 13243
rect 23857 13209 23891 13243
rect 7389 13141 7423 13175
rect 9137 13141 9171 13175
rect 11529 13141 11563 13175
rect 13553 13141 13587 13175
rect 15209 13141 15243 13175
rect 15577 13141 15611 13175
rect 15669 13141 15703 13175
rect 16865 13141 16899 13175
rect 18245 13141 18279 13175
rect 18705 13141 18739 13175
rect 19625 13141 19659 13175
rect 20177 13141 20211 13175
rect 20545 13141 20579 13175
rect 20637 13141 20671 13175
rect 21465 13141 21499 13175
rect 25237 13141 25271 13175
rect 6561 12937 6595 12971
rect 10333 12937 10367 12971
rect 14105 12937 14139 12971
rect 16129 12937 16163 12971
rect 20913 12937 20947 12971
rect 22477 12937 22511 12971
rect 24777 12937 24811 12971
rect 9229 12869 9263 12903
rect 10701 12869 10735 12903
rect 19993 12869 20027 12903
rect 20453 12869 20487 12903
rect 20637 12869 20671 12903
rect 21465 12869 21499 12903
rect 23305 12869 23339 12903
rect 7205 12801 7239 12835
rect 10793 12801 10827 12835
rect 12173 12801 12207 12835
rect 13001 12801 13035 12835
rect 13093 12801 13127 12835
rect 14473 12801 14507 12835
rect 14565 12801 14599 12835
rect 15669 12801 15703 12835
rect 16313 12801 16347 12835
rect 16773 12801 16807 12835
rect 17233 12801 17267 12835
rect 19073 12801 19107 12835
rect 21281 12801 21315 12835
rect 22201 12801 22235 12835
rect 23029 12801 23063 12835
rect 7481 12733 7515 12767
rect 10885 12733 10919 12767
rect 13185 12733 13219 12767
rect 14749 12733 14783 12767
rect 17969 12733 18003 12767
rect 19165 12733 19199 12767
rect 19257 12733 19291 12767
rect 8953 12665 8987 12699
rect 12633 12665 12667 12699
rect 15209 12665 15243 12699
rect 22017 12665 22051 12699
rect 11621 12597 11655 12631
rect 11989 12597 12023 12631
rect 13737 12597 13771 12631
rect 15485 12597 15519 12631
rect 16957 12597 16991 12631
rect 18705 12597 18739 12631
rect 20085 12597 20119 12631
rect 22661 12597 22695 12631
rect 25145 12597 25179 12631
rect 7849 12393 7883 12427
rect 9781 12393 9815 12427
rect 11437 12393 11471 12427
rect 12633 12393 12667 12427
rect 14381 12393 14415 12427
rect 17969 12393 18003 12427
rect 20085 12393 20119 12427
rect 16865 12325 16899 12359
rect 8493 12257 8527 12291
rect 10425 12257 10459 12291
rect 11897 12257 11931 12291
rect 12081 12257 12115 12291
rect 13185 12257 13219 12291
rect 14933 12257 14967 12291
rect 17509 12257 17543 12291
rect 20361 12257 20395 12291
rect 8217 12189 8251 12223
rect 10241 12189 10275 12223
rect 13093 12189 13127 12223
rect 14841 12189 14875 12223
rect 16405 12189 16439 12223
rect 17325 12189 17359 12223
rect 19533 12189 19567 12223
rect 22661 12189 22695 12223
rect 24685 12189 24719 12223
rect 9413 12121 9447 12155
rect 10149 12121 10183 12155
rect 11805 12121 11839 12155
rect 18613 12121 18647 12155
rect 19717 12121 19751 12155
rect 20637 12121 20671 12155
rect 23857 12121 23891 12155
rect 8309 12053 8343 12087
rect 8953 12053 8987 12087
rect 13001 12053 13035 12087
rect 13645 12053 13679 12087
rect 13921 12053 13955 12087
rect 14749 12053 14783 12087
rect 15577 12053 15611 12087
rect 16221 12053 16255 12087
rect 17233 12053 17267 12087
rect 18245 12053 18279 12087
rect 18705 12053 18739 12087
rect 22109 12053 22143 12087
rect 25329 12053 25363 12087
rect 8953 11849 8987 11883
rect 9413 11849 9447 11883
rect 10149 11849 10183 11883
rect 11989 11849 12023 11883
rect 13185 11849 13219 11883
rect 13645 11849 13679 11883
rect 14381 11849 14415 11883
rect 14749 11849 14783 11883
rect 16221 11849 16255 11883
rect 17325 11849 17359 11883
rect 18061 11849 18095 11883
rect 19257 11849 19291 11883
rect 19625 11849 19659 11883
rect 22661 11849 22695 11883
rect 13553 11781 13587 11815
rect 19993 11781 20027 11815
rect 20913 11781 20947 11815
rect 21649 11781 21683 11815
rect 23397 11781 23431 11815
rect 7849 11713 7883 11747
rect 9321 11713 9355 11747
rect 10517 11713 10551 11747
rect 12357 11713 12391 11747
rect 12449 11713 12483 11747
rect 14841 11713 14875 11747
rect 15577 11713 15611 11747
rect 17233 11713 17267 11747
rect 18429 11713 18463 11747
rect 20085 11713 20119 11747
rect 21373 11713 21407 11747
rect 22005 11713 22039 11747
rect 23121 11713 23155 11747
rect 9597 11645 9631 11679
rect 10609 11645 10643 11679
rect 10793 11645 10827 11679
rect 12541 11645 12575 11679
rect 13829 11645 13863 11679
rect 14933 11645 14967 11679
rect 17417 11645 17451 11679
rect 18521 11645 18555 11679
rect 18705 11645 18739 11679
rect 20269 11645 20303 11679
rect 8493 11577 8527 11611
rect 19073 11577 19107 11611
rect 11253 11509 11287 11543
rect 16865 11509 16899 11543
rect 21005 11509 21039 11543
rect 24869 11509 24903 11543
rect 25145 11509 25179 11543
rect 8585 11305 8619 11339
rect 12633 11305 12667 11339
rect 16405 11305 16439 11339
rect 17785 11305 17819 11339
rect 18797 11305 18831 11339
rect 19073 11305 19107 11339
rect 19625 11305 19659 11339
rect 21557 11305 21591 11339
rect 13645 11237 13679 11271
rect 13921 11237 13955 11271
rect 22753 11237 22787 11271
rect 9137 11169 9171 11203
rect 10333 11169 10367 11203
rect 11805 11169 11839 11203
rect 11897 11169 11931 11203
rect 13277 11169 13311 11203
rect 14657 11169 14691 11203
rect 18337 11169 18371 11203
rect 23213 11169 23247 11203
rect 23397 11169 23431 11203
rect 7941 11101 7975 11135
rect 9413 11101 9447 11135
rect 11713 11101 11747 11135
rect 14197 11101 14231 11135
rect 17049 11101 17083 11135
rect 17417 11101 17451 11135
rect 19533 11101 19567 11135
rect 20453 11101 20487 11135
rect 21097 11101 21131 11135
rect 21741 11101 21775 11135
rect 24593 11101 24627 11135
rect 13001 11033 13035 11067
rect 13093 11033 13127 11067
rect 14381 11033 14415 11067
rect 14933 11033 14967 11067
rect 18245 11033 18279 11067
rect 20269 11033 20303 11067
rect 22477 11033 22511 11067
rect 23121 11033 23155 11067
rect 10701 10965 10735 10999
rect 11345 10965 11379 10999
rect 16865 10965 16899 10999
rect 18153 10965 18187 10999
rect 20913 10965 20947 10999
rect 25237 10965 25271 10999
rect 10977 10761 11011 10795
rect 11713 10761 11747 10795
rect 12173 10761 12207 10795
rect 12541 10761 12575 10795
rect 13921 10761 13955 10795
rect 14381 10761 14415 10795
rect 15209 10761 15243 10795
rect 15945 10761 15979 10795
rect 21465 10761 21499 10795
rect 23305 10761 23339 10795
rect 9505 10693 9539 10727
rect 13001 10693 13035 10727
rect 18061 10693 18095 10727
rect 9229 10625 9263 10659
rect 12909 10625 12943 10659
rect 14289 10625 14323 10659
rect 15853 10625 15887 10659
rect 16865 10625 16899 10659
rect 19073 10625 19107 10659
rect 19717 10625 19751 10659
rect 23489 10625 23523 10659
rect 23949 10625 23983 10659
rect 13185 10557 13219 10591
rect 14473 10557 14507 10591
rect 14933 10557 14967 10591
rect 16129 10557 16163 10591
rect 19993 10557 20027 10591
rect 22017 10557 22051 10591
rect 22293 10557 22327 10591
rect 24777 10557 24811 10591
rect 15485 10489 15519 10523
rect 13553 10421 13587 10455
rect 17509 10421 17543 10455
rect 18153 10421 18187 10455
rect 18705 10421 18739 10455
rect 19165 10421 19199 10455
rect 12725 10217 12759 10251
rect 15669 10217 15703 10251
rect 16865 10217 16899 10251
rect 20085 10217 20119 10251
rect 25145 10217 25179 10251
rect 14473 10149 14507 10183
rect 20361 10149 20395 10183
rect 20821 10149 20855 10183
rect 21925 10149 21959 10183
rect 9137 10081 9171 10115
rect 9413 10081 9447 10115
rect 11161 10081 11195 10115
rect 11989 10081 12023 10115
rect 12081 10081 12115 10115
rect 13369 10081 13403 10115
rect 15117 10081 15151 10115
rect 16129 10081 16163 10115
rect 16221 10081 16255 10115
rect 17417 10081 17451 10115
rect 18613 10081 18647 10115
rect 18797 10081 18831 10115
rect 21281 10081 21315 10115
rect 21465 10081 21499 10115
rect 22293 10081 22327 10115
rect 22569 10081 22603 10115
rect 8585 10013 8619 10047
rect 13185 10013 13219 10047
rect 14105 10013 14139 10047
rect 14841 10013 14875 10047
rect 18521 10013 18555 10047
rect 19441 10013 19475 10047
rect 17233 9945 17267 9979
rect 8401 9877 8435 9911
rect 10885 9877 10919 9911
rect 11529 9877 11563 9911
rect 11897 9877 11931 9911
rect 13093 9877 13127 9911
rect 13921 9877 13955 9911
rect 14933 9877 14967 9911
rect 16037 9877 16071 9911
rect 17325 9877 17359 9911
rect 18153 9877 18187 9911
rect 21189 9877 21223 9911
rect 24041 9877 24075 9911
rect 24593 9877 24627 9911
rect 15117 9605 15151 9639
rect 16957 9605 16991 9639
rect 20269 9605 20303 9639
rect 21189 9605 21223 9639
rect 23305 9605 23339 9639
rect 11713 9537 11747 9571
rect 15025 9537 15059 9571
rect 16129 9537 16163 9571
rect 22109 9537 22143 9571
rect 23949 9537 23983 9571
rect 8217 9469 8251 9503
rect 8493 9469 8527 9503
rect 9965 9469 9999 9503
rect 10609 9469 10643 9503
rect 11989 9469 12023 9503
rect 13921 9469 13955 9503
rect 15301 9469 15335 9503
rect 17693 9469 17727 9503
rect 17969 9469 18003 9503
rect 20361 9469 20395 9503
rect 20545 9469 20579 9503
rect 24685 9469 24719 9503
rect 14657 9401 14691 9435
rect 15669 9401 15703 9435
rect 16313 9401 16347 9435
rect 7849 9333 7883 9367
rect 11069 9333 11103 9367
rect 11253 9333 11287 9367
rect 13461 9333 13495 9367
rect 17049 9333 17083 9367
rect 19441 9333 19475 9367
rect 19901 9333 19935 9367
rect 21281 9333 21315 9367
rect 12357 9129 12391 9163
rect 18889 9129 18923 9163
rect 13001 9061 13035 9095
rect 10333 8993 10367 9027
rect 13553 8993 13587 9027
rect 15301 8993 15335 9027
rect 16221 8993 16255 9027
rect 20085 8993 20119 9027
rect 20269 8993 20303 9027
rect 9137 8925 9171 8959
rect 10609 8925 10643 8959
rect 11713 8925 11747 8959
rect 12541 8925 12575 8959
rect 13369 8925 13403 8959
rect 16037 8925 16071 8959
rect 16681 8925 16715 8959
rect 17141 8925 17175 8959
rect 18245 8925 18279 8959
rect 21005 8925 21039 8959
rect 22661 8925 22695 8959
rect 24593 8925 24627 8959
rect 14381 8857 14415 8891
rect 14565 8857 14599 8891
rect 19993 8857 20027 8891
rect 21833 8857 21867 8891
rect 23857 8857 23891 8891
rect 9781 8789 9815 8823
rect 13461 8789 13495 8823
rect 14841 8789 14875 8823
rect 15577 8789 15611 8823
rect 15945 8789 15979 8823
rect 16865 8789 16899 8823
rect 17785 8789 17819 8823
rect 19349 8789 19383 8823
rect 19625 8789 19659 8823
rect 25237 8789 25271 8823
rect 12081 8585 12115 8619
rect 15577 8585 15611 8619
rect 15945 8585 15979 8619
rect 17877 8585 17911 8619
rect 21833 8585 21867 8619
rect 22109 8585 22143 8619
rect 8861 8517 8895 8551
rect 16037 8517 16071 8551
rect 18705 8517 18739 8551
rect 19441 8517 19475 8551
rect 22661 8517 22695 8551
rect 8125 8449 8159 8483
rect 12909 8449 12943 8483
rect 17233 8449 17267 8483
rect 17325 8449 17359 8483
rect 19717 8449 19751 8483
rect 24593 8449 24627 8483
rect 8585 8381 8619 8415
rect 10977 8381 11011 8415
rect 12173 8381 12207 8415
rect 12357 8381 12391 8415
rect 14289 8381 14323 8415
rect 14565 8381 14599 8415
rect 16221 8381 16255 8415
rect 17509 8381 17543 8415
rect 18797 8381 18831 8415
rect 18981 8381 19015 8415
rect 19993 8381 20027 8415
rect 22385 8381 22419 8415
rect 24133 8381 24167 8415
rect 7941 8313 7975 8347
rect 10701 8313 10735 8347
rect 11713 8313 11747 8347
rect 18337 8313 18371 8347
rect 10333 8245 10367 8279
rect 13553 8245 13587 8279
rect 13829 8245 13863 8279
rect 16865 8245 16899 8279
rect 21465 8245 21499 8279
rect 25237 8245 25271 8279
rect 11805 8041 11839 8075
rect 14552 8041 14586 8075
rect 18889 8041 18923 8075
rect 10425 7973 10459 8007
rect 10885 7905 10919 7939
rect 10977 7905 11011 7939
rect 11529 7905 11563 7939
rect 12357 7905 12391 7939
rect 13553 7905 13587 7939
rect 14289 7905 14323 7939
rect 17141 7905 17175 7939
rect 17417 7905 17451 7939
rect 19993 7905 20027 7939
rect 22661 7905 22695 7939
rect 9321 7837 9355 7871
rect 12173 7837 12207 7871
rect 13369 7837 13403 7871
rect 16681 7837 16715 7871
rect 19533 7837 19567 7871
rect 20545 7837 20579 7871
rect 22201 7837 22235 7871
rect 24593 7837 24627 7871
rect 12265 7769 12299 7803
rect 13461 7769 13495 7803
rect 19717 7769 19751 7803
rect 21557 7769 21591 7803
rect 25237 7769 25271 7803
rect 9965 7701 9999 7735
rect 10793 7701 10827 7735
rect 13001 7701 13035 7735
rect 16037 7701 16071 7735
rect 16497 7701 16531 7735
rect 24133 7701 24167 7735
rect 10793 7497 10827 7531
rect 11713 7497 11747 7531
rect 15393 7497 15427 7531
rect 15485 7497 15519 7531
rect 16313 7497 16347 7531
rect 17509 7497 17543 7531
rect 9321 7429 9355 7463
rect 25145 7429 25179 7463
rect 12081 7361 12115 7395
rect 13461 7361 13495 7395
rect 14289 7361 14323 7395
rect 17417 7361 17451 7395
rect 18245 7361 18279 7395
rect 20085 7361 20119 7395
rect 22109 7361 22143 7395
rect 23949 7361 23983 7395
rect 9045 7293 9079 7327
rect 12173 7293 12207 7327
rect 12265 7293 12299 7327
rect 13553 7293 13587 7327
rect 13645 7293 13679 7327
rect 15577 7293 15611 7327
rect 17693 7293 17727 7327
rect 19441 7293 19475 7327
rect 21281 7293 21315 7327
rect 23305 7293 23339 7327
rect 12817 7225 12851 7259
rect 11161 7157 11195 7191
rect 13093 7157 13127 7191
rect 15025 7157 15059 7191
rect 16129 7157 16163 7191
rect 17049 7157 17083 7191
rect 12357 6953 12391 6987
rect 15209 6953 15243 6987
rect 20072 6953 20106 6987
rect 22280 6953 22314 6987
rect 21557 6885 21591 6919
rect 10609 6817 10643 6851
rect 12633 6817 12667 6851
rect 13461 6817 13495 6851
rect 13645 6817 13679 6851
rect 16957 6817 16991 6851
rect 19809 6817 19843 6851
rect 22017 6817 22051 6851
rect 23765 6817 23799 6851
rect 25053 6817 25087 6851
rect 25145 6817 25179 6851
rect 14289 6749 14323 6783
rect 16681 6749 16715 6783
rect 17509 6749 17543 6783
rect 10885 6681 10919 6715
rect 15669 6681 15703 6715
rect 15853 6681 15887 6715
rect 18705 6681 18739 6715
rect 13001 6613 13035 6647
rect 13369 6613 13403 6647
rect 14933 6613 14967 6647
rect 16313 6613 16347 6647
rect 16773 6613 16807 6647
rect 24041 6613 24075 6647
rect 24593 6613 24627 6647
rect 24961 6613 24995 6647
rect 12357 6409 12391 6443
rect 15577 6409 15611 6443
rect 19073 6409 19107 6443
rect 13277 6341 13311 6375
rect 15669 6341 15703 6375
rect 10517 6273 10551 6307
rect 11713 6273 11747 6307
rect 16405 6273 16439 6307
rect 16865 6273 16899 6307
rect 20085 6273 20119 6307
rect 22201 6273 22235 6307
rect 23949 6273 23983 6307
rect 13001 6205 13035 6239
rect 15761 6205 15795 6239
rect 17141 6205 17175 6239
rect 18613 6205 18647 6239
rect 21281 6205 21315 6239
rect 22477 6205 22511 6239
rect 24685 6205 24719 6239
rect 14749 6137 14783 6171
rect 11161 6069 11195 6103
rect 12633 6069 12667 6103
rect 15209 6069 15243 6103
rect 19533 6069 19567 6103
rect 11713 5865 11747 5899
rect 13737 5865 13771 5899
rect 24225 5865 24259 5899
rect 10241 5729 10275 5763
rect 19993 5729 20027 5763
rect 20821 5729 20855 5763
rect 22661 5729 22695 5763
rect 9965 5661 9999 5695
rect 12541 5661 12575 5695
rect 13093 5661 13127 5695
rect 14381 5661 14415 5695
rect 15669 5661 15703 5695
rect 17693 5661 17727 5695
rect 20545 5661 20579 5695
rect 22293 5661 22327 5695
rect 24593 5661 24627 5695
rect 16865 5593 16899 5627
rect 18705 5593 18739 5627
rect 19533 5593 19567 5627
rect 19717 5593 19751 5627
rect 11989 5525 12023 5559
rect 12357 5525 12391 5559
rect 15025 5525 15059 5559
rect 15301 5525 15335 5559
rect 23949 5525 23983 5559
rect 25237 5525 25271 5559
rect 10333 5321 10367 5355
rect 19073 5321 19107 5355
rect 14013 5253 14047 5287
rect 16129 5253 16163 5287
rect 19993 5253 20027 5287
rect 10885 5185 10919 5219
rect 11161 5185 11195 5219
rect 13185 5185 13219 5219
rect 13737 5185 13771 5219
rect 16865 5185 16899 5219
rect 19257 5185 19291 5219
rect 19717 5185 19751 5219
rect 22017 5185 22051 5219
rect 23949 5185 23983 5219
rect 11713 5117 11747 5151
rect 11989 5117 12023 5151
rect 17141 5117 17175 5151
rect 22477 5117 22511 5151
rect 24777 5117 24811 5151
rect 10977 4981 11011 5015
rect 13001 4981 13035 5015
rect 15485 4981 15519 5015
rect 16221 4981 16255 5015
rect 18613 4981 18647 5015
rect 21465 4981 21499 5015
rect 9045 4777 9079 4811
rect 16865 4777 16899 4811
rect 23765 4777 23799 4811
rect 9689 4709 9723 4743
rect 10333 4709 10367 4743
rect 14197 4709 14231 4743
rect 24869 4709 24903 4743
rect 5089 4641 5123 4675
rect 11621 4641 11655 4675
rect 11897 4641 11931 4675
rect 12909 4641 12943 4675
rect 13185 4641 13219 4675
rect 15117 4641 15151 4675
rect 19901 4641 19935 4675
rect 21741 4641 21775 4675
rect 7113 4573 7147 4607
rect 9873 4573 9907 4607
rect 10241 4573 10275 4607
rect 10517 4573 10551 4607
rect 11161 4573 11195 4607
rect 14657 4573 14691 4607
rect 17601 4573 17635 4607
rect 19625 4573 19659 4607
rect 21373 4573 21407 4607
rect 23121 4573 23155 4607
rect 5365 4505 5399 4539
rect 7389 4505 7423 4539
rect 15393 4505 15427 4539
rect 18337 4505 18371 4539
rect 24685 4505 24719 4539
rect 25145 4505 25179 4539
rect 1501 4437 1535 4471
rect 10977 4437 11011 4471
rect 14473 4437 14507 4471
rect 7297 4165 7331 4199
rect 20913 4165 20947 4199
rect 22937 4165 22971 4199
rect 1777 4097 1811 4131
rect 2421 4097 2455 4131
rect 2697 4097 2731 4131
rect 4353 4097 4387 4131
rect 4629 4097 4663 4131
rect 6745 4097 6779 4131
rect 7113 4097 7147 4131
rect 8861 4097 8895 4131
rect 9505 4097 9539 4131
rect 9781 4097 9815 4131
rect 10609 4097 10643 4131
rect 11897 4097 11931 4131
rect 13001 4097 13035 4131
rect 15117 4097 15151 4131
rect 17049 4097 17083 4131
rect 18705 4097 18739 4131
rect 21557 4097 21591 4131
rect 22109 4097 22143 4131
rect 23857 4097 23891 4131
rect 10333 4029 10367 4063
rect 13461 4029 13495 4063
rect 16129 4029 16163 4063
rect 17325 4029 17359 4063
rect 19165 4029 19199 4063
rect 21005 4029 21039 4063
rect 21189 4029 21223 4063
rect 24317 4029 24351 4063
rect 1593 3961 1627 3995
rect 6561 3961 6595 3995
rect 12541 3961 12575 3995
rect 2237 3893 2271 3927
rect 2881 3893 2915 3927
rect 4169 3893 4203 3927
rect 6101 3893 6135 3927
rect 7481 3893 7515 3927
rect 8677 3893 8711 3927
rect 9321 3893 9355 3927
rect 9965 3893 9999 3927
rect 11621 3893 11655 3927
rect 20545 3893 20579 3927
rect 2881 3689 2915 3723
rect 4261 3689 4295 3723
rect 18613 3689 18647 3723
rect 23305 3689 23339 3723
rect 23673 3689 23707 3723
rect 6377 3621 6411 3655
rect 10425 3621 10459 3655
rect 24869 3621 24903 3655
rect 1869 3553 1903 3587
rect 5181 3553 5215 3587
rect 8125 3553 8159 3587
rect 9781 3553 9815 3587
rect 11345 3553 11379 3587
rect 14749 3553 14783 3587
rect 16589 3553 16623 3587
rect 19901 3553 19935 3587
rect 21741 3553 21775 3587
rect 1593 3485 1627 3519
rect 3065 3485 3099 3519
rect 3525 3485 3559 3519
rect 4445 3485 4479 3519
rect 4905 3485 4939 3519
rect 6101 3485 6135 3519
rect 6561 3485 6595 3519
rect 7297 3485 7331 3519
rect 7941 3485 7975 3519
rect 8585 3485 8619 3519
rect 9321 3485 9355 3519
rect 10333 3485 10367 3519
rect 10609 3485 10643 3519
rect 11069 3485 11103 3519
rect 12541 3485 12575 3519
rect 14473 3485 14507 3519
rect 16313 3485 16347 3519
rect 17969 3485 18003 3519
rect 19625 3485 19659 3519
rect 21281 3485 21315 3519
rect 23581 3485 23615 3519
rect 24685 3485 24719 3519
rect 25145 3485 25179 3519
rect 13553 3417 13587 3451
rect 3341 3349 3375 3383
rect 7113 3349 7147 3383
rect 7757 3349 7791 3383
rect 8401 3349 8435 3383
rect 9137 3349 9171 3383
rect 18889 3349 18923 3383
rect 4537 3145 4571 3179
rect 4813 3145 4847 3179
rect 6561 3145 6595 3179
rect 7205 3145 7239 3179
rect 9229 3145 9263 3179
rect 10977 3145 11011 3179
rect 21281 3145 21315 3179
rect 22201 3145 22235 3179
rect 22937 3145 22971 3179
rect 24869 3145 24903 3179
rect 9413 3077 9447 3111
rect 20637 3077 20671 3111
rect 22109 3077 22143 3111
rect 22845 3077 22879 3111
rect 2145 3009 2179 3043
rect 3433 3009 3467 3043
rect 3709 3009 3743 3043
rect 5457 3009 5491 3043
rect 6745 3009 6779 3043
rect 7389 3009 7423 3043
rect 7849 3009 7883 3043
rect 9045 3009 9079 3043
rect 9873 3009 9907 3043
rect 10517 3009 10551 3043
rect 11161 3013 11195 3047
rect 11713 3009 11747 3043
rect 11989 3009 12023 3043
rect 13185 3009 13219 3043
rect 14841 3009 14875 3043
rect 17049 3009 17083 3043
rect 18889 3009 18923 3043
rect 20821 3009 20855 3043
rect 23581 3009 23615 3043
rect 2421 2941 2455 2975
rect 5181 2941 5215 2975
rect 8125 2941 8159 2975
rect 13645 2941 13679 2975
rect 15301 2941 15335 2975
rect 17417 2941 17451 2975
rect 19165 2941 19199 2975
rect 9689 2873 9723 2907
rect 10333 2805 10367 2839
rect 6653 2601 6687 2635
rect 10563 2601 10597 2635
rect 14105 2601 14139 2635
rect 18705 2601 18739 2635
rect 21281 2601 21315 2635
rect 23857 2601 23891 2635
rect 25421 2601 25455 2635
rect 4537 2533 4571 2567
rect 7757 2533 7791 2567
rect 5457 2465 5491 2499
rect 9689 2465 9723 2499
rect 11713 2465 11747 2499
rect 17325 2465 17359 2499
rect 19901 2465 19935 2499
rect 22477 2465 22511 2499
rect 2605 2397 2639 2431
rect 2881 2397 2915 2431
rect 4721 2397 4755 2431
rect 5181 2397 5215 2431
rect 6837 2397 6871 2431
rect 7297 2397 7331 2431
rect 7941 2397 7975 2431
rect 8585 2397 8619 2431
rect 9413 2397 9447 2431
rect 10333 2397 10367 2431
rect 12541 2397 12575 2431
rect 14473 2397 14507 2431
rect 17049 2397 17083 2431
rect 18889 2397 18923 2431
rect 19625 2397 19659 2431
rect 21465 2397 21499 2431
rect 22017 2397 22051 2431
rect 24041 2397 24075 2431
rect 3985 2329 4019 2363
rect 4261 2329 4295 2363
rect 9045 2329 9079 2363
rect 13277 2329 13311 2363
rect 15393 2329 15427 2363
rect 24685 2329 24719 2363
rect 25145 2329 25179 2363
rect 3801 2261 3835 2295
rect 6377 2261 6411 2295
rect 7113 2261 7147 2295
rect 8401 2261 8435 2295
rect 9229 2261 9263 2295
rect 16129 2261 16163 2295
rect 24777 2261 24811 2295
<< metal1 >>
rect 1104 54426 25852 54448
rect 1104 54374 7950 54426
rect 8002 54374 8014 54426
rect 8066 54374 8078 54426
rect 8130 54374 8142 54426
rect 8194 54374 8206 54426
rect 8258 54374 17950 54426
rect 18002 54374 18014 54426
rect 18066 54374 18078 54426
rect 18130 54374 18142 54426
rect 18194 54374 18206 54426
rect 18258 54374 25852 54426
rect 1104 54352 25852 54374
rect 18966 54272 18972 54324
rect 19024 54272 19030 54324
rect 24486 54272 24492 54324
rect 24544 54272 24550 54324
rect 18141 54247 18199 54253
rect 18141 54244 18153 54247
rect 17880 54216 18153 54244
rect 2225 54179 2283 54185
rect 2225 54145 2237 54179
rect 2271 54176 2283 54179
rect 3878 54176 3884 54188
rect 2271 54148 3884 54176
rect 2271 54145 2283 54148
rect 2225 54139 2283 54145
rect 3878 54136 3884 54148
rect 3936 54136 3942 54188
rect 4157 54179 4215 54185
rect 4157 54145 4169 54179
rect 4203 54176 4215 54179
rect 6546 54176 6552 54188
rect 4203 54148 6552 54176
rect 4203 54145 4215 54148
rect 4157 54139 4215 54145
rect 6546 54136 6552 54148
rect 6604 54136 6610 54188
rect 6730 54136 6736 54188
rect 6788 54136 6794 54188
rect 13446 54136 13452 54188
rect 13504 54176 13510 54188
rect 13725 54179 13783 54185
rect 13725 54176 13737 54179
rect 13504 54148 13737 54176
rect 13504 54136 13510 54148
rect 13725 54145 13737 54148
rect 13771 54176 13783 54179
rect 14093 54179 14151 54185
rect 14093 54176 14105 54179
rect 13771 54148 14105 54176
rect 13771 54145 13783 54148
rect 13725 54139 13783 54145
rect 14093 54145 14105 54148
rect 14139 54145 14151 54179
rect 14093 54139 14151 54145
rect 14826 54136 14832 54188
rect 14884 54176 14890 54188
rect 15105 54179 15163 54185
rect 15105 54176 15117 54179
rect 14884 54148 15117 54176
rect 14884 54136 14890 54148
rect 15105 54145 15117 54148
rect 15151 54176 15163 54179
rect 15381 54179 15439 54185
rect 15381 54176 15393 54179
rect 15151 54148 15393 54176
rect 15151 54145 15163 54148
rect 15105 54139 15163 54145
rect 15381 54145 15393 54148
rect 15427 54145 15439 54179
rect 15381 54139 15439 54145
rect 16574 54136 16580 54188
rect 16632 54176 16638 54188
rect 17037 54179 17095 54185
rect 17037 54176 17049 54179
rect 16632 54148 17049 54176
rect 16632 54136 16638 54148
rect 17037 54145 17049 54148
rect 17083 54176 17095 54179
rect 17313 54179 17371 54185
rect 17313 54176 17325 54179
rect 17083 54148 17325 54176
rect 17083 54145 17095 54148
rect 17037 54139 17095 54145
rect 17313 54145 17325 54148
rect 17359 54145 17371 54179
rect 17313 54139 17371 54145
rect 17586 54136 17592 54188
rect 17644 54176 17650 54188
rect 17880 54185 17908 54216
rect 18141 54213 18153 54216
rect 18187 54213 18199 54247
rect 18141 54207 18199 54213
rect 17865 54179 17923 54185
rect 17865 54176 17877 54179
rect 17644 54148 17877 54176
rect 17644 54136 17650 54148
rect 17865 54145 17877 54148
rect 17911 54145 17923 54179
rect 19705 54179 19763 54185
rect 19705 54176 19717 54179
rect 17865 54139 17923 54145
rect 18156 54148 19717 54176
rect 2406 54068 2412 54120
rect 2464 54108 2470 54120
rect 2501 54111 2559 54117
rect 2501 54108 2513 54111
rect 2464 54080 2513 54108
rect 2464 54068 2470 54080
rect 2501 54077 2513 54080
rect 2547 54077 2559 54111
rect 2501 54071 2559 54077
rect 4062 54068 4068 54120
rect 4120 54108 4126 54120
rect 4433 54111 4491 54117
rect 4433 54108 4445 54111
rect 4120 54080 4445 54108
rect 4120 54068 4126 54080
rect 4433 54077 4445 54080
rect 4479 54077 4491 54111
rect 4433 54071 4491 54077
rect 6914 54068 6920 54120
rect 6972 54108 6978 54120
rect 7101 54111 7159 54117
rect 7101 54108 7113 54111
rect 6972 54080 7113 54108
rect 6972 54068 6978 54080
rect 7101 54077 7113 54080
rect 7147 54077 7159 54111
rect 7101 54071 7159 54077
rect 8478 54068 8484 54120
rect 8536 54108 8542 54120
rect 18156 54108 18184 54148
rect 19705 54145 19717 54148
rect 19751 54145 19763 54179
rect 19705 54139 19763 54145
rect 23293 54179 23351 54185
rect 23293 54145 23305 54179
rect 23339 54176 23351 54179
rect 23474 54176 23480 54188
rect 23339 54148 23480 54176
rect 23339 54145 23351 54148
rect 23293 54139 23351 54145
rect 23474 54136 23480 54148
rect 23532 54136 23538 54188
rect 23753 54179 23811 54185
rect 23753 54145 23765 54179
rect 23799 54176 23811 54179
rect 24504 54176 24532 54272
rect 23799 54148 24532 54176
rect 23799 54145 23811 54148
rect 23753 54139 23811 54145
rect 24762 54136 24768 54188
rect 24820 54176 24826 54188
rect 25041 54179 25099 54185
rect 25041 54176 25053 54179
rect 24820 54148 25053 54176
rect 24820 54136 24826 54148
rect 25041 54145 25053 54148
rect 25087 54145 25099 54179
rect 25041 54139 25099 54145
rect 8536 54080 18184 54108
rect 8536 54068 8542 54080
rect 18966 54068 18972 54120
rect 19024 54108 19030 54120
rect 19429 54111 19487 54117
rect 19429 54108 19441 54111
rect 19024 54080 19441 54108
rect 19024 54068 19030 54080
rect 19429 54077 19441 54080
rect 19475 54077 19487 54111
rect 19429 54071 19487 54077
rect 18782 54000 18788 54052
rect 18840 54040 18846 54052
rect 23937 54043 23995 54049
rect 23937 54040 23949 54043
rect 18840 54012 23949 54040
rect 18840 54000 18846 54012
rect 23937 54009 23949 54012
rect 23983 54009 23995 54043
rect 23937 54003 23995 54009
rect 12618 53932 12624 53984
rect 12676 53972 12682 53984
rect 13541 53975 13599 53981
rect 13541 53972 13553 53975
rect 12676 53944 13553 53972
rect 12676 53932 12682 53944
rect 13541 53941 13553 53944
rect 13587 53941 13599 53975
rect 13541 53935 13599 53941
rect 14918 53932 14924 53984
rect 14976 53932 14982 53984
rect 15470 53932 15476 53984
rect 15528 53972 15534 53984
rect 16853 53975 16911 53981
rect 16853 53972 16865 53975
rect 15528 53944 16865 53972
rect 15528 53932 15534 53944
rect 16853 53941 16865 53944
rect 16899 53941 16911 53975
rect 16853 53935 16911 53941
rect 17126 53932 17132 53984
rect 17184 53972 17190 53984
rect 17681 53975 17739 53981
rect 17681 53972 17693 53975
rect 17184 53944 17693 53972
rect 17184 53932 17190 53944
rect 17681 53941 17693 53944
rect 17727 53941 17739 53975
rect 17681 53935 17739 53941
rect 20714 53932 20720 53984
rect 20772 53972 20778 53984
rect 23109 53975 23167 53981
rect 23109 53972 23121 53975
rect 20772 53944 23121 53972
rect 20772 53932 20778 53944
rect 23109 53941 23121 53944
rect 23155 53941 23167 53975
rect 23109 53935 23167 53941
rect 25225 53975 25283 53981
rect 25225 53941 25237 53975
rect 25271 53972 25283 53975
rect 26786 53972 26792 53984
rect 25271 53944 26792 53972
rect 25271 53941 25283 53944
rect 25225 53935 25283 53941
rect 26786 53932 26792 53944
rect 26844 53932 26850 53984
rect 1104 53882 25852 53904
rect 1104 53830 2950 53882
rect 3002 53830 3014 53882
rect 3066 53830 3078 53882
rect 3130 53830 3142 53882
rect 3194 53830 3206 53882
rect 3258 53830 12950 53882
rect 13002 53830 13014 53882
rect 13066 53830 13078 53882
rect 13130 53830 13142 53882
rect 13194 53830 13206 53882
rect 13258 53830 22950 53882
rect 23002 53830 23014 53882
rect 23066 53830 23078 53882
rect 23130 53830 23142 53882
rect 23194 53830 23206 53882
rect 23258 53830 25852 53882
rect 1104 53808 25852 53830
rect 23474 53728 23480 53780
rect 23532 53768 23538 53780
rect 25866 53768 25872 53780
rect 23532 53740 25872 53768
rect 23532 53728 23538 53740
rect 25866 53728 25872 53740
rect 25924 53728 25930 53780
rect 1026 53592 1032 53644
rect 1084 53632 1090 53644
rect 2041 53635 2099 53641
rect 2041 53632 2053 53635
rect 1084 53604 2053 53632
rect 1084 53592 1090 53604
rect 2041 53601 2053 53604
rect 2087 53601 2099 53635
rect 2041 53595 2099 53601
rect 5166 53592 5172 53644
rect 5224 53632 5230 53644
rect 5721 53635 5779 53641
rect 5721 53632 5733 53635
rect 5224 53604 5733 53632
rect 5224 53592 5230 53604
rect 5721 53601 5733 53604
rect 5767 53601 5779 53635
rect 5721 53595 5779 53601
rect 1765 53567 1823 53573
rect 1765 53533 1777 53567
rect 1811 53533 1823 53567
rect 1765 53527 1823 53533
rect 5445 53567 5503 53573
rect 5445 53533 5457 53567
rect 5491 53564 5503 53567
rect 7650 53564 7656 53576
rect 5491 53536 7656 53564
rect 5491 53533 5503 53536
rect 5445 53527 5503 53533
rect 1780 53496 1808 53527
rect 7650 53524 7656 53536
rect 7708 53524 7714 53576
rect 23382 53524 23388 53576
rect 23440 53564 23446 53576
rect 23845 53567 23903 53573
rect 23845 53564 23857 53567
rect 23440 53536 23857 53564
rect 23440 53524 23446 53536
rect 23845 53533 23857 53536
rect 23891 53564 23903 53567
rect 24397 53567 24455 53573
rect 24397 53564 24409 53567
rect 23891 53536 24409 53564
rect 23891 53533 23903 53536
rect 23845 53527 23903 53533
rect 24397 53533 24409 53536
rect 24443 53533 24455 53567
rect 24397 53527 24455 53533
rect 24670 53524 24676 53576
rect 24728 53564 24734 53576
rect 25041 53567 25099 53573
rect 25041 53564 25053 53567
rect 24728 53536 25053 53564
rect 24728 53524 24734 53536
rect 25041 53533 25053 53536
rect 25087 53533 25099 53567
rect 25041 53527 25099 53533
rect 7558 53496 7564 53508
rect 1780 53468 7564 53496
rect 7558 53456 7564 53468
rect 7616 53456 7622 53508
rect 23934 53388 23940 53440
rect 23992 53388 23998 53440
rect 24854 53388 24860 53440
rect 24912 53428 24918 53440
rect 25225 53431 25283 53437
rect 25225 53428 25237 53431
rect 24912 53400 25237 53428
rect 24912 53388 24918 53400
rect 25225 53397 25237 53400
rect 25271 53397 25283 53431
rect 25225 53391 25283 53397
rect 1104 53338 25852 53360
rect 1104 53286 7950 53338
rect 8002 53286 8014 53338
rect 8066 53286 8078 53338
rect 8130 53286 8142 53338
rect 8194 53286 8206 53338
rect 8258 53286 17950 53338
rect 18002 53286 18014 53338
rect 18066 53286 18078 53338
rect 18130 53286 18142 53338
rect 18194 53286 18206 53338
rect 18258 53286 25852 53338
rect 1104 53264 25852 53286
rect 3878 53184 3884 53236
rect 3936 53224 3942 53236
rect 4985 53227 5043 53233
rect 4985 53224 4997 53227
rect 3936 53196 4997 53224
rect 3936 53184 3942 53196
rect 4985 53193 4997 53196
rect 5031 53193 5043 53227
rect 4985 53187 5043 53193
rect 6546 53184 6552 53236
rect 6604 53184 6610 53236
rect 5169 53091 5227 53097
rect 5169 53057 5181 53091
rect 5215 53057 5227 53091
rect 5169 53051 5227 53057
rect 6733 53091 6791 53097
rect 6733 53057 6745 53091
rect 6779 53088 6791 53091
rect 9582 53088 9588 53100
rect 6779 53060 9588 53088
rect 6779 53057 6791 53060
rect 6733 53051 6791 53057
rect 5184 53020 5212 53051
rect 9582 53048 9588 53060
rect 9640 53048 9646 53100
rect 24765 53091 24823 53097
rect 24765 53057 24777 53091
rect 24811 53088 24823 53091
rect 25038 53088 25044 53100
rect 24811 53060 25044 53088
rect 24811 53057 24823 53060
rect 24765 53051 24823 53057
rect 25038 53048 25044 53060
rect 25096 53048 25102 53100
rect 7742 53020 7748 53032
rect 5184 52992 7748 53020
rect 7742 52980 7748 52992
rect 7800 52980 7806 53032
rect 25225 52887 25283 52893
rect 25225 52853 25237 52887
rect 25271 52884 25283 52887
rect 26050 52884 26056 52896
rect 25271 52856 26056 52884
rect 25271 52853 25283 52856
rect 25225 52847 25283 52853
rect 26050 52844 26056 52856
rect 26108 52844 26114 52896
rect 1104 52794 25852 52816
rect 1104 52742 2950 52794
rect 3002 52742 3014 52794
rect 3066 52742 3078 52794
rect 3130 52742 3142 52794
rect 3194 52742 3206 52794
rect 3258 52742 12950 52794
rect 13002 52742 13014 52794
rect 13066 52742 13078 52794
rect 13130 52742 13142 52794
rect 13194 52742 13206 52794
rect 13258 52742 22950 52794
rect 23002 52742 23014 52794
rect 23066 52742 23078 52794
rect 23130 52742 23142 52794
rect 23194 52742 23206 52794
rect 23258 52742 25852 52794
rect 1104 52720 25852 52742
rect 7650 52640 7656 52692
rect 7708 52640 7714 52692
rect 7834 52572 7840 52624
rect 7892 52612 7898 52624
rect 8386 52612 8392 52624
rect 7892 52584 8392 52612
rect 7892 52572 7898 52584
rect 8386 52572 8392 52584
rect 8444 52572 8450 52624
rect 7837 52479 7895 52485
rect 7837 52445 7849 52479
rect 7883 52476 7895 52479
rect 9490 52476 9496 52488
rect 7883 52448 9496 52476
rect 7883 52445 7895 52448
rect 7837 52439 7895 52445
rect 9490 52436 9496 52448
rect 9548 52436 9554 52488
rect 16942 52436 16948 52488
rect 17000 52476 17006 52488
rect 20346 52476 20352 52488
rect 17000 52448 20352 52476
rect 17000 52436 17006 52448
rect 20346 52436 20352 52448
rect 20404 52436 20410 52488
rect 24581 52479 24639 52485
rect 24581 52445 24593 52479
rect 24627 52476 24639 52479
rect 25317 52479 25375 52485
rect 24627 52448 24992 52476
rect 24627 52445 24639 52448
rect 24581 52439 24639 52445
rect 24964 52420 24992 52448
rect 25317 52445 25329 52479
rect 25363 52476 25375 52479
rect 26510 52476 26516 52488
rect 25363 52448 26516 52476
rect 25363 52445 25375 52448
rect 25317 52439 25375 52445
rect 26510 52436 26516 52448
rect 26568 52436 26574 52488
rect 24946 52368 24952 52420
rect 25004 52368 25010 52420
rect 1104 52250 25852 52272
rect 1104 52198 7950 52250
rect 8002 52198 8014 52250
rect 8066 52198 8078 52250
rect 8130 52198 8142 52250
rect 8194 52198 8206 52250
rect 8258 52198 17950 52250
rect 18002 52198 18014 52250
rect 18066 52198 18078 52250
rect 18130 52198 18142 52250
rect 18194 52198 18206 52250
rect 18258 52198 25852 52250
rect 1104 52176 25852 52198
rect 6730 52096 6736 52148
rect 6788 52136 6794 52148
rect 8849 52139 8907 52145
rect 8849 52136 8861 52139
rect 6788 52108 8861 52136
rect 6788 52096 6794 52108
rect 8849 52105 8861 52108
rect 8895 52105 8907 52139
rect 8849 52099 8907 52105
rect 8757 52003 8815 52009
rect 8757 51969 8769 52003
rect 8803 52000 8815 52003
rect 10318 52000 10324 52012
rect 8803 51972 10324 52000
rect 8803 51969 8815 51972
rect 8757 51963 8815 51969
rect 10318 51960 10324 51972
rect 10376 51960 10382 52012
rect 25498 51756 25504 51808
rect 25556 51756 25562 51808
rect 1104 51706 25852 51728
rect 1104 51654 2950 51706
rect 3002 51654 3014 51706
rect 3066 51654 3078 51706
rect 3130 51654 3142 51706
rect 3194 51654 3206 51706
rect 3258 51654 12950 51706
rect 13002 51654 13014 51706
rect 13066 51654 13078 51706
rect 13130 51654 13142 51706
rect 13194 51654 13206 51706
rect 13258 51654 22950 51706
rect 23002 51654 23014 51706
rect 23066 51654 23078 51706
rect 23130 51654 23142 51706
rect 23194 51654 23206 51706
rect 23258 51654 25852 51706
rect 1104 51632 25852 51654
rect 7650 51552 7656 51604
rect 7708 51552 7714 51604
rect 7742 51552 7748 51604
rect 7800 51592 7806 51604
rect 8021 51595 8079 51601
rect 8021 51592 8033 51595
rect 7800 51564 8033 51592
rect 7800 51552 7806 51564
rect 8021 51561 8033 51564
rect 8067 51561 8079 51595
rect 8021 51555 8079 51561
rect 8478 51552 8484 51604
rect 8536 51552 8542 51604
rect 7561 51391 7619 51397
rect 7561 51357 7573 51391
rect 7607 51388 7619 51391
rect 8478 51388 8484 51400
rect 7607 51360 8484 51388
rect 7607 51357 7619 51360
rect 7561 51351 7619 51357
rect 8478 51348 8484 51360
rect 8536 51348 8542 51400
rect 24949 51391 25007 51397
rect 24949 51357 24961 51391
rect 24995 51388 25007 51391
rect 25498 51388 25504 51400
rect 24995 51360 25504 51388
rect 24995 51357 25007 51360
rect 24949 51351 25007 51357
rect 25498 51348 25504 51360
rect 25556 51348 25562 51400
rect 21358 51212 21364 51264
rect 21416 51252 21422 51264
rect 25041 51255 25099 51261
rect 25041 51252 25053 51255
rect 21416 51224 25053 51252
rect 21416 51212 21422 51224
rect 25041 51221 25053 51224
rect 25087 51221 25099 51255
rect 25041 51215 25099 51221
rect 1104 51162 25852 51184
rect 1104 51110 7950 51162
rect 8002 51110 8014 51162
rect 8066 51110 8078 51162
rect 8130 51110 8142 51162
rect 8194 51110 8206 51162
rect 8258 51110 17950 51162
rect 18002 51110 18014 51162
rect 18066 51110 18078 51162
rect 18130 51110 18142 51162
rect 18194 51110 18206 51162
rect 18258 51110 25852 51162
rect 1104 51088 25852 51110
rect 24581 50915 24639 50921
rect 24581 50881 24593 50915
rect 24627 50912 24639 50915
rect 24946 50912 24952 50924
rect 24627 50884 24952 50912
rect 24627 50881 24639 50884
rect 24581 50875 24639 50881
rect 24946 50872 24952 50884
rect 25004 50872 25010 50924
rect 25038 50668 25044 50720
rect 25096 50668 25102 50720
rect 1104 50618 25852 50640
rect 1104 50566 2950 50618
rect 3002 50566 3014 50618
rect 3066 50566 3078 50618
rect 3130 50566 3142 50618
rect 3194 50566 3206 50618
rect 3258 50566 12950 50618
rect 13002 50566 13014 50618
rect 13066 50566 13078 50618
rect 13130 50566 13142 50618
rect 13194 50566 13206 50618
rect 13258 50566 22950 50618
rect 23002 50566 23014 50618
rect 23066 50566 23078 50618
rect 23130 50566 23142 50618
rect 23194 50566 23206 50618
rect 23258 50566 25852 50618
rect 1104 50544 25852 50566
rect 16022 50464 16028 50516
rect 16080 50504 16086 50516
rect 25038 50504 25044 50516
rect 16080 50476 25044 50504
rect 16080 50464 16086 50476
rect 25038 50464 25044 50476
rect 25096 50464 25102 50516
rect 17218 50396 17224 50448
rect 17276 50436 17282 50448
rect 24394 50436 24400 50448
rect 17276 50408 24400 50436
rect 17276 50396 17282 50408
rect 24394 50396 24400 50408
rect 24452 50396 24458 50448
rect 25498 50124 25504 50176
rect 25556 50124 25562 50176
rect 1104 50074 25852 50096
rect 1104 50022 7950 50074
rect 8002 50022 8014 50074
rect 8066 50022 8078 50074
rect 8130 50022 8142 50074
rect 8194 50022 8206 50074
rect 8258 50022 17950 50074
rect 18002 50022 18014 50074
rect 18066 50022 18078 50074
rect 18130 50022 18142 50074
rect 18194 50022 18206 50074
rect 18258 50022 25852 50074
rect 1104 50000 25852 50022
rect 24489 49827 24547 49833
rect 24489 49793 24501 49827
rect 24535 49824 24547 49827
rect 25498 49824 25504 49836
rect 24535 49796 25504 49824
rect 24535 49793 24547 49796
rect 24489 49787 24547 49793
rect 25498 49784 25504 49796
rect 25556 49784 25562 49836
rect 20898 49716 20904 49768
rect 20956 49756 20962 49768
rect 24765 49759 24823 49765
rect 24765 49756 24777 49759
rect 20956 49728 24777 49756
rect 20956 49716 20962 49728
rect 24765 49725 24777 49728
rect 24811 49725 24823 49759
rect 24765 49719 24823 49725
rect 1104 49530 25852 49552
rect 1104 49478 2950 49530
rect 3002 49478 3014 49530
rect 3066 49478 3078 49530
rect 3130 49478 3142 49530
rect 3194 49478 3206 49530
rect 3258 49478 12950 49530
rect 13002 49478 13014 49530
rect 13066 49478 13078 49530
rect 13130 49478 13142 49530
rect 13194 49478 13206 49530
rect 13258 49478 22950 49530
rect 23002 49478 23014 49530
rect 23066 49478 23078 49530
rect 23130 49478 23142 49530
rect 23194 49478 23206 49530
rect 23258 49478 25852 49530
rect 1104 49456 25852 49478
rect 7650 49376 7656 49428
rect 7708 49416 7714 49428
rect 8389 49419 8447 49425
rect 8389 49416 8401 49419
rect 7708 49388 8401 49416
rect 7708 49376 7714 49388
rect 8389 49385 8401 49388
rect 8435 49385 8447 49419
rect 8389 49379 8447 49385
rect 9122 49376 9128 49428
rect 9180 49416 9186 49428
rect 9401 49419 9459 49425
rect 9401 49416 9413 49419
rect 9180 49388 9413 49416
rect 9180 49376 9186 49388
rect 9401 49385 9413 49388
rect 9447 49385 9459 49419
rect 9401 49379 9459 49385
rect 9582 49376 9588 49428
rect 9640 49416 9646 49428
rect 9769 49419 9827 49425
rect 9769 49416 9781 49419
rect 9640 49388 9781 49416
rect 9640 49376 9646 49388
rect 9769 49385 9781 49388
rect 9815 49385 9827 49419
rect 9769 49379 9827 49385
rect 8478 49308 8484 49360
rect 8536 49348 8542 49360
rect 10137 49351 10195 49357
rect 10137 49348 10149 49351
rect 8536 49320 10149 49348
rect 8536 49308 8542 49320
rect 6641 49283 6699 49289
rect 6641 49249 6653 49283
rect 6687 49280 6699 49283
rect 8754 49280 8760 49292
rect 6687 49252 8760 49280
rect 6687 49249 6699 49252
rect 6641 49243 6699 49249
rect 8754 49240 8760 49252
rect 8812 49240 8818 49292
rect 9324 49221 9352 49320
rect 10137 49317 10149 49320
rect 10183 49348 10195 49351
rect 10962 49348 10968 49360
rect 10183 49320 10968 49348
rect 10183 49317 10195 49320
rect 10137 49311 10195 49317
rect 10962 49308 10968 49320
rect 11020 49308 11026 49360
rect 9309 49215 9367 49221
rect 9309 49181 9321 49215
rect 9355 49181 9367 49215
rect 9309 49175 9367 49181
rect 6917 49147 6975 49153
rect 6917 49113 6929 49147
rect 6963 49113 6975 49147
rect 8941 49147 8999 49153
rect 8941 49144 8953 49147
rect 8142 49116 8953 49144
rect 6917 49107 6975 49113
rect 8941 49113 8953 49116
rect 8987 49144 8999 49147
rect 9674 49144 9680 49156
rect 8987 49116 9680 49144
rect 8987 49113 8999 49116
rect 8941 49107 8999 49113
rect 6932 49076 6960 49107
rect 9674 49104 9680 49116
rect 9732 49104 9738 49156
rect 24765 49147 24823 49153
rect 24765 49113 24777 49147
rect 24811 49144 24823 49147
rect 25130 49144 25136 49156
rect 24811 49116 25136 49144
rect 24811 49113 24823 49116
rect 24765 49107 24823 49113
rect 25130 49104 25136 49116
rect 25188 49104 25194 49156
rect 8294 49076 8300 49088
rect 6932 49048 8300 49076
rect 8294 49036 8300 49048
rect 8352 49036 8358 49088
rect 8754 49036 8760 49088
rect 8812 49036 8818 49088
rect 25222 49036 25228 49088
rect 25280 49036 25286 49088
rect 1104 48986 25852 49008
rect 1104 48934 7950 48986
rect 8002 48934 8014 48986
rect 8066 48934 8078 48986
rect 8130 48934 8142 48986
rect 8194 48934 8206 48986
rect 8258 48934 17950 48986
rect 18002 48934 18014 48986
rect 18066 48934 18078 48986
rect 18130 48934 18142 48986
rect 18194 48934 18206 48986
rect 18258 48934 25852 48986
rect 1104 48912 25852 48934
rect 7742 48764 7748 48816
rect 7800 48804 7806 48816
rect 7929 48807 7987 48813
rect 7929 48804 7941 48807
rect 7800 48776 7941 48804
rect 7800 48764 7806 48776
rect 7929 48773 7941 48776
rect 7975 48804 7987 48807
rect 7975 48776 9168 48804
rect 7975 48773 7987 48776
rect 7929 48767 7987 48773
rect 9140 48736 9168 48776
rect 10264 48739 10322 48745
rect 10264 48736 10276 48739
rect 9140 48708 10276 48736
rect 10264 48705 10276 48708
rect 10310 48705 10322 48739
rect 10264 48699 10322 48705
rect 7742 48628 7748 48680
rect 7800 48628 7806 48680
rect 8386 48628 8392 48680
rect 8444 48628 8450 48680
rect 10367 48535 10425 48541
rect 10367 48501 10379 48535
rect 10413 48532 10425 48535
rect 12342 48532 12348 48544
rect 10413 48504 12348 48532
rect 10413 48501 10425 48504
rect 10367 48495 10425 48501
rect 12342 48492 12348 48504
rect 12400 48492 12406 48544
rect 25130 48492 25136 48544
rect 25188 48532 25194 48544
rect 25409 48535 25467 48541
rect 25409 48532 25421 48535
rect 25188 48504 25421 48532
rect 25188 48492 25194 48504
rect 25409 48501 25421 48504
rect 25455 48501 25467 48535
rect 25409 48495 25467 48501
rect 1104 48442 25852 48464
rect 1104 48390 2950 48442
rect 3002 48390 3014 48442
rect 3066 48390 3078 48442
rect 3130 48390 3142 48442
rect 3194 48390 3206 48442
rect 3258 48390 12950 48442
rect 13002 48390 13014 48442
rect 13066 48390 13078 48442
rect 13130 48390 13142 48442
rect 13194 48390 13206 48442
rect 13258 48390 22950 48442
rect 23002 48390 23014 48442
rect 23066 48390 23078 48442
rect 23130 48390 23142 48442
rect 23194 48390 23206 48442
rect 23258 48390 25852 48442
rect 1104 48368 25852 48390
rect 9582 48288 9588 48340
rect 9640 48328 9646 48340
rect 9640 48300 11100 48328
rect 9640 48288 9646 48300
rect 8294 48220 8300 48272
rect 8352 48260 8358 48272
rect 9769 48263 9827 48269
rect 9769 48260 9781 48263
rect 8352 48232 9781 48260
rect 8352 48220 8358 48232
rect 9769 48229 9781 48232
rect 9815 48229 9827 48263
rect 9769 48223 9827 48229
rect 9122 48084 9128 48136
rect 9180 48084 9186 48136
rect 11072 48124 11100 48300
rect 11552 48127 11610 48133
rect 11552 48124 11564 48127
rect 11072 48096 11564 48124
rect 11552 48093 11564 48096
rect 11598 48093 11610 48127
rect 11552 48087 11610 48093
rect 25130 48084 25136 48136
rect 25188 48084 25194 48136
rect 11655 47991 11713 47997
rect 11655 47957 11667 47991
rect 11701 47988 11713 47991
rect 14458 47988 14464 48000
rect 11701 47960 14464 47988
rect 11701 47957 11713 47960
rect 11655 47951 11713 47957
rect 14458 47948 14464 47960
rect 14516 47948 14522 48000
rect 17586 47948 17592 48000
rect 17644 47988 17650 48000
rect 25225 47991 25283 47997
rect 25225 47988 25237 47991
rect 17644 47960 25237 47988
rect 17644 47948 17650 47960
rect 25225 47957 25237 47960
rect 25271 47957 25283 47991
rect 25225 47951 25283 47957
rect 1104 47898 25852 47920
rect 1104 47846 7950 47898
rect 8002 47846 8014 47898
rect 8066 47846 8078 47898
rect 8130 47846 8142 47898
rect 8194 47846 8206 47898
rect 8258 47846 17950 47898
rect 18002 47846 18014 47898
rect 18066 47846 18078 47898
rect 18130 47846 18142 47898
rect 18194 47846 18206 47898
rect 18258 47846 25852 47898
rect 1104 47824 25852 47846
rect 8849 47719 8907 47725
rect 8849 47685 8861 47719
rect 8895 47716 8907 47719
rect 9582 47716 9588 47728
rect 8895 47688 9588 47716
rect 8895 47685 8907 47688
rect 8849 47679 8907 47685
rect 9582 47676 9588 47688
rect 9640 47676 9646 47728
rect 12342 47676 12348 47728
rect 12400 47716 12406 47728
rect 12805 47719 12863 47725
rect 12805 47716 12817 47719
rect 12400 47688 12817 47716
rect 12400 47676 12406 47688
rect 12805 47685 12817 47688
rect 12851 47685 12863 47719
rect 12805 47679 12863 47685
rect 12618 47608 12624 47660
rect 12676 47608 12682 47660
rect 24857 47651 24915 47657
rect 24857 47617 24869 47651
rect 24903 47648 24915 47651
rect 25314 47648 25320 47660
rect 24903 47620 25320 47648
rect 24903 47617 24915 47620
rect 24857 47611 24915 47617
rect 25314 47608 25320 47620
rect 25372 47608 25378 47660
rect 8665 47583 8723 47589
rect 8665 47549 8677 47583
rect 8711 47549 8723 47583
rect 8665 47543 8723 47549
rect 8680 47512 8708 47543
rect 9306 47540 9312 47592
rect 9364 47540 9370 47592
rect 14461 47583 14519 47589
rect 14461 47549 14473 47583
rect 14507 47580 14519 47583
rect 14826 47580 14832 47592
rect 14507 47552 14832 47580
rect 14507 47549 14519 47552
rect 14461 47543 14519 47549
rect 14826 47540 14832 47552
rect 14884 47540 14890 47592
rect 9030 47512 9036 47524
rect 8680 47484 9036 47512
rect 9030 47472 9036 47484
rect 9088 47472 9094 47524
rect 25133 47447 25191 47453
rect 25133 47413 25145 47447
rect 25179 47444 25191 47447
rect 25958 47444 25964 47456
rect 25179 47416 25964 47444
rect 25179 47413 25191 47416
rect 25133 47407 25191 47413
rect 25958 47404 25964 47416
rect 26016 47404 26022 47456
rect 1104 47354 25852 47376
rect 1104 47302 2950 47354
rect 3002 47302 3014 47354
rect 3066 47302 3078 47354
rect 3130 47302 3142 47354
rect 3194 47302 3206 47354
rect 3258 47302 12950 47354
rect 13002 47302 13014 47354
rect 13066 47302 13078 47354
rect 13130 47302 13142 47354
rect 13194 47302 13206 47354
rect 13258 47302 22950 47354
rect 23002 47302 23014 47354
rect 23066 47302 23078 47354
rect 23130 47302 23142 47354
rect 23194 47302 23206 47354
rect 23258 47302 25852 47354
rect 1104 47280 25852 47302
rect 10597 47243 10655 47249
rect 10597 47209 10609 47243
rect 10643 47240 10655 47243
rect 10686 47240 10692 47252
rect 10643 47212 10692 47240
rect 10643 47209 10655 47212
rect 10597 47203 10655 47209
rect 10686 47200 10692 47212
rect 10744 47200 10750 47252
rect 10962 47200 10968 47252
rect 11020 47240 11026 47252
rect 11149 47243 11207 47249
rect 11149 47240 11161 47243
rect 11020 47212 11161 47240
rect 11020 47200 11026 47212
rect 11149 47209 11161 47212
rect 11195 47209 11207 47243
rect 11149 47203 11207 47209
rect 18966 47200 18972 47252
rect 19024 47240 19030 47252
rect 25222 47240 25228 47252
rect 19024 47212 25228 47240
rect 19024 47200 19030 47212
rect 25222 47200 25228 47212
rect 25280 47200 25286 47252
rect 9490 47132 9496 47184
rect 9548 47172 9554 47184
rect 10781 47175 10839 47181
rect 10781 47172 10793 47175
rect 9548 47144 10793 47172
rect 9548 47132 9554 47144
rect 10781 47141 10793 47144
rect 10827 47141 10839 47175
rect 10781 47135 10839 47141
rect 10321 47039 10379 47045
rect 10321 47005 10333 47039
rect 10367 47005 10379 47039
rect 10796 47036 10824 47135
rect 11514 47064 11520 47116
rect 11572 47104 11578 47116
rect 14277 47107 14335 47113
rect 11572 47076 12756 47104
rect 11572 47064 11578 47076
rect 12564 47039 12622 47045
rect 12564 47036 12576 47039
rect 10796 47008 12576 47036
rect 10321 46999 10379 47005
rect 12564 47005 12576 47008
rect 12610 47005 12622 47039
rect 12728 47036 12756 47076
rect 14277 47073 14289 47107
rect 14323 47104 14335 47107
rect 14918 47104 14924 47116
rect 14323 47076 14924 47104
rect 14323 47073 14335 47076
rect 14277 47067 14335 47073
rect 14918 47064 14924 47076
rect 14976 47064 14982 47116
rect 13392 47039 13450 47045
rect 13392 47036 13404 47039
rect 12728 47008 13404 47036
rect 12564 46999 12622 47005
rect 13392 47005 13404 47008
rect 13438 47005 13450 47039
rect 13392 46999 13450 47005
rect 13495 47039 13553 47045
rect 13495 47005 13507 47039
rect 13541 47036 13553 47039
rect 14182 47036 14188 47048
rect 13541 47008 14188 47036
rect 13541 47005 13553 47008
rect 13495 46999 13553 47005
rect 10336 46968 10364 46999
rect 14182 46996 14188 47008
rect 14240 46996 14246 47048
rect 10962 46968 10968 46980
rect 10336 46940 10968 46968
rect 10962 46928 10968 46940
rect 11020 46928 11026 46980
rect 12667 46971 12725 46977
rect 12667 46937 12679 46971
rect 12713 46968 12725 46971
rect 14274 46968 14280 46980
rect 12713 46940 14280 46968
rect 12713 46937 12725 46940
rect 12667 46931 12725 46937
rect 14274 46928 14280 46940
rect 14332 46928 14338 46980
rect 14458 46928 14464 46980
rect 14516 46928 14522 46980
rect 16114 46928 16120 46980
rect 16172 46928 16178 46980
rect 25314 46860 25320 46912
rect 25372 46900 25378 46912
rect 25409 46903 25467 46909
rect 25409 46900 25421 46903
rect 25372 46872 25421 46900
rect 25372 46860 25378 46872
rect 25409 46869 25421 46872
rect 25455 46869 25467 46903
rect 25409 46863 25467 46869
rect 1104 46810 25852 46832
rect 1104 46758 7950 46810
rect 8002 46758 8014 46810
rect 8066 46758 8078 46810
rect 8130 46758 8142 46810
rect 8194 46758 8206 46810
rect 8258 46758 17950 46810
rect 18002 46758 18014 46810
rect 18066 46758 18078 46810
rect 18130 46758 18142 46810
rect 18194 46758 18206 46810
rect 18258 46758 25852 46810
rect 1104 46736 25852 46758
rect 9122 46656 9128 46708
rect 9180 46696 9186 46708
rect 10597 46699 10655 46705
rect 10597 46696 10609 46699
rect 9180 46668 10609 46696
rect 9180 46656 9186 46668
rect 10597 46665 10609 46668
rect 10643 46665 10655 46699
rect 10597 46659 10655 46665
rect 9674 46588 9680 46640
rect 9732 46588 9738 46640
rect 14274 46588 14280 46640
rect 14332 46628 14338 46640
rect 14645 46631 14703 46637
rect 14645 46628 14657 46631
rect 14332 46600 14657 46628
rect 14332 46588 14338 46600
rect 14645 46597 14657 46600
rect 14691 46597 14703 46631
rect 14645 46591 14703 46597
rect 25314 46520 25320 46572
rect 25372 46520 25378 46572
rect 8754 46452 8760 46504
rect 8812 46492 8818 46504
rect 8849 46495 8907 46501
rect 8849 46492 8861 46495
rect 8812 46464 8861 46492
rect 8812 46452 8818 46464
rect 8849 46461 8861 46464
rect 8895 46461 8907 46495
rect 8849 46455 8907 46461
rect 9125 46495 9183 46501
rect 9125 46461 9137 46495
rect 9171 46492 9183 46495
rect 10594 46492 10600 46504
rect 9171 46464 10600 46492
rect 9171 46461 9183 46464
rect 9125 46455 9183 46461
rect 8864 46356 8892 46455
rect 10594 46452 10600 46464
rect 10652 46452 10658 46504
rect 14461 46495 14519 46501
rect 14461 46461 14473 46495
rect 14507 46492 14519 46495
rect 15470 46492 15476 46504
rect 14507 46464 15476 46492
rect 14507 46461 14519 46464
rect 14461 46455 14519 46461
rect 15470 46452 15476 46464
rect 15528 46452 15534 46504
rect 16298 46452 16304 46504
rect 16356 46452 16362 46504
rect 11057 46427 11115 46433
rect 11057 46424 11069 46427
rect 10336 46396 11069 46424
rect 9214 46356 9220 46368
rect 8864 46328 9220 46356
rect 9214 46316 9220 46328
rect 9272 46316 9278 46368
rect 9674 46316 9680 46368
rect 9732 46356 9738 46368
rect 10336 46356 10364 46396
rect 11057 46393 11069 46396
rect 11103 46424 11115 46427
rect 11146 46424 11152 46436
rect 11103 46396 11152 46424
rect 11103 46393 11115 46396
rect 11057 46387 11115 46393
rect 11146 46384 11152 46396
rect 11204 46384 11210 46436
rect 9732 46328 10364 46356
rect 9732 46316 9738 46328
rect 10962 46316 10968 46368
rect 11020 46316 11026 46368
rect 23290 46316 23296 46368
rect 23348 46356 23354 46368
rect 25133 46359 25191 46365
rect 25133 46356 25145 46359
rect 23348 46328 25145 46356
rect 23348 46316 23354 46328
rect 25133 46325 25145 46328
rect 25179 46325 25191 46359
rect 25133 46319 25191 46325
rect 1104 46266 25852 46288
rect 1104 46214 2950 46266
rect 3002 46214 3014 46266
rect 3066 46214 3078 46266
rect 3130 46214 3142 46266
rect 3194 46214 3206 46266
rect 3258 46214 12950 46266
rect 13002 46214 13014 46266
rect 13066 46214 13078 46266
rect 13130 46214 13142 46266
rect 13194 46214 13206 46266
rect 13258 46214 22950 46266
rect 23002 46214 23014 46266
rect 23066 46214 23078 46266
rect 23130 46214 23142 46266
rect 23194 46214 23206 46266
rect 23258 46214 25852 46266
rect 1104 46192 25852 46214
rect 24210 46044 24216 46096
rect 24268 46084 24274 46096
rect 25133 46087 25191 46093
rect 25133 46084 25145 46087
rect 24268 46056 25145 46084
rect 24268 46044 24274 46056
rect 25133 46053 25145 46056
rect 25179 46053 25191 46087
rect 25133 46047 25191 46053
rect 10318 45976 10324 46028
rect 10376 46016 10382 46028
rect 10597 46019 10655 46025
rect 10597 46016 10609 46019
rect 10376 45988 10609 46016
rect 10376 45976 10382 45988
rect 10597 45985 10609 45988
rect 10643 46016 10655 46019
rect 11514 46016 11520 46028
rect 10643 45988 11520 46016
rect 10643 45985 10655 45988
rect 10597 45979 10655 45985
rect 11514 45976 11520 45988
rect 11572 45976 11578 46028
rect 12066 45976 12072 46028
rect 12124 45976 12130 46028
rect 14182 45976 14188 46028
rect 14240 46016 14246 46028
rect 15841 46019 15899 46025
rect 15841 46016 15853 46019
rect 14240 45988 15853 46016
rect 14240 45976 14246 45988
rect 15841 45985 15853 45988
rect 15887 45985 15899 46019
rect 15841 45979 15899 45985
rect 10410 45908 10416 45960
rect 10468 45908 10474 45960
rect 15657 45951 15715 45957
rect 15657 45917 15669 45951
rect 15703 45917 15715 45951
rect 15657 45911 15715 45917
rect 24857 45951 24915 45957
rect 24857 45917 24869 45951
rect 24903 45948 24915 45951
rect 25314 45948 25320 45960
rect 24903 45920 25320 45948
rect 24903 45917 24915 45920
rect 24857 45911 24915 45917
rect 15672 45812 15700 45911
rect 25314 45908 25320 45920
rect 25372 45908 25378 45960
rect 17126 45880 17132 45892
rect 16546 45852 17132 45880
rect 16546 45812 16574 45852
rect 17126 45840 17132 45852
rect 17184 45840 17190 45892
rect 17494 45840 17500 45892
rect 17552 45840 17558 45892
rect 15672 45784 16574 45812
rect 1104 45722 25852 45744
rect 1104 45670 7950 45722
rect 8002 45670 8014 45722
rect 8066 45670 8078 45722
rect 8130 45670 8142 45722
rect 8194 45670 8206 45722
rect 8258 45670 17950 45722
rect 18002 45670 18014 45722
rect 18066 45670 18078 45722
rect 18130 45670 18142 45722
rect 18194 45670 18206 45722
rect 18258 45670 25852 45722
rect 1104 45648 25852 45670
rect 9490 45500 9496 45552
rect 9548 45500 9554 45552
rect 8938 45364 8944 45416
rect 8996 45404 9002 45416
rect 9309 45407 9367 45413
rect 9309 45404 9321 45407
rect 8996 45376 9321 45404
rect 8996 45364 9002 45376
rect 9309 45373 9321 45376
rect 9355 45373 9367 45407
rect 9309 45367 9367 45373
rect 10870 45364 10876 45416
rect 10928 45364 10934 45416
rect 25314 45228 25320 45280
rect 25372 45268 25378 45280
rect 25409 45271 25467 45277
rect 25409 45268 25421 45271
rect 25372 45240 25421 45268
rect 25372 45228 25378 45240
rect 25409 45237 25421 45240
rect 25455 45237 25467 45271
rect 25409 45231 25467 45237
rect 1104 45178 25852 45200
rect 1104 45126 2950 45178
rect 3002 45126 3014 45178
rect 3066 45126 3078 45178
rect 3130 45126 3142 45178
rect 3194 45126 3206 45178
rect 3258 45126 12950 45178
rect 13002 45126 13014 45178
rect 13066 45126 13078 45178
rect 13130 45126 13142 45178
rect 13194 45126 13206 45178
rect 13258 45126 22950 45178
rect 23002 45126 23014 45178
rect 23066 45126 23078 45178
rect 23130 45126 23142 45178
rect 23194 45126 23206 45178
rect 23258 45126 25852 45178
rect 1104 45104 25852 45126
rect 10594 45024 10600 45076
rect 10652 45024 10658 45076
rect 11330 45024 11336 45076
rect 11388 45024 11394 45076
rect 11514 45024 11520 45076
rect 11572 45024 11578 45076
rect 15746 45024 15752 45076
rect 15804 45064 15810 45076
rect 21358 45064 21364 45076
rect 15804 45036 21364 45064
rect 15804 45024 15810 45036
rect 21358 45024 21364 45036
rect 21416 45024 21422 45076
rect 20714 44888 20720 44940
rect 20772 44888 20778 44940
rect 21266 44888 21272 44940
rect 21324 44928 21330 44940
rect 22465 44931 22523 44937
rect 22465 44928 22477 44931
rect 21324 44900 22477 44928
rect 21324 44888 21330 44900
rect 22465 44897 22477 44900
rect 22511 44897 22523 44931
rect 22465 44891 22523 44897
rect 9950 44820 9956 44872
rect 10008 44860 10014 44872
rect 10686 44860 10692 44872
rect 10008 44832 10692 44860
rect 10008 44820 10014 44832
rect 10686 44820 10692 44832
rect 10744 44820 10750 44872
rect 11054 44820 11060 44872
rect 11112 44860 11118 44872
rect 11885 44863 11943 44869
rect 11885 44860 11897 44863
rect 11112 44832 11897 44860
rect 11112 44820 11118 44832
rect 11885 44829 11897 44832
rect 11931 44829 11943 44863
rect 11885 44823 11943 44829
rect 19426 44820 19432 44872
rect 19484 44860 19490 44872
rect 20441 44863 20499 44869
rect 20441 44860 20453 44863
rect 19484 44832 20453 44860
rect 19484 44820 19490 44832
rect 20441 44829 20453 44832
rect 20487 44829 20499 44863
rect 20441 44823 20499 44829
rect 25314 44820 25320 44872
rect 25372 44820 25378 44872
rect 21266 44752 21272 44804
rect 21324 44752 21330 44804
rect 22186 44684 22192 44736
rect 22244 44684 22250 44736
rect 23474 44684 23480 44736
rect 23532 44724 23538 44736
rect 25133 44727 25191 44733
rect 25133 44724 25145 44727
rect 23532 44696 25145 44724
rect 23532 44684 23538 44696
rect 25133 44693 25145 44696
rect 25179 44693 25191 44727
rect 25133 44687 25191 44693
rect 1104 44634 25852 44656
rect 1104 44582 7950 44634
rect 8002 44582 8014 44634
rect 8066 44582 8078 44634
rect 8130 44582 8142 44634
rect 8194 44582 8206 44634
rect 8258 44582 17950 44634
rect 18002 44582 18014 44634
rect 18066 44582 18078 44634
rect 18130 44582 18142 44634
rect 18194 44582 18206 44634
rect 18258 44582 25852 44634
rect 1104 44560 25852 44582
rect 24762 44344 24768 44396
rect 24820 44384 24826 44396
rect 25133 44387 25191 44393
rect 25133 44384 25145 44387
rect 24820 44356 25145 44384
rect 24820 44344 24826 44356
rect 25133 44353 25145 44356
rect 25179 44353 25191 44387
rect 25133 44347 25191 44353
rect 25317 44251 25375 44257
rect 25317 44217 25329 44251
rect 25363 44248 25375 44251
rect 25774 44248 25780 44260
rect 25363 44220 25780 44248
rect 25363 44217 25375 44220
rect 25317 44211 25375 44217
rect 25774 44208 25780 44220
rect 25832 44208 25838 44260
rect 1104 44090 25852 44112
rect 1104 44038 2950 44090
rect 3002 44038 3014 44090
rect 3066 44038 3078 44090
rect 3130 44038 3142 44090
rect 3194 44038 3206 44090
rect 3258 44038 12950 44090
rect 13002 44038 13014 44090
rect 13066 44038 13078 44090
rect 13130 44038 13142 44090
rect 13194 44038 13206 44090
rect 13258 44038 22950 44090
rect 23002 44038 23014 44090
rect 23066 44038 23078 44090
rect 23130 44038 23142 44090
rect 23194 44038 23206 44090
rect 23258 44038 25852 44090
rect 1104 44016 25852 44038
rect 25498 43596 25504 43648
rect 25556 43596 25562 43648
rect 1104 43546 25852 43568
rect 1104 43494 7950 43546
rect 8002 43494 8014 43546
rect 8066 43494 8078 43546
rect 8130 43494 8142 43546
rect 8194 43494 8206 43546
rect 8258 43494 17950 43546
rect 18002 43494 18014 43546
rect 18066 43494 18078 43546
rect 18130 43494 18142 43546
rect 18194 43494 18206 43546
rect 18258 43494 25852 43546
rect 1104 43472 25852 43494
rect 9950 43392 9956 43444
rect 10008 43432 10014 43444
rect 11149 43435 11207 43441
rect 11149 43432 11161 43435
rect 10008 43404 11161 43432
rect 10008 43392 10014 43404
rect 11149 43401 11161 43404
rect 11195 43401 11207 43435
rect 11149 43395 11207 43401
rect 25133 43367 25191 43373
rect 25133 43333 25145 43367
rect 25179 43364 25191 43367
rect 25498 43364 25504 43376
rect 25179 43336 25504 43364
rect 25179 43333 25191 43336
rect 25133 43327 25191 43333
rect 25498 43324 25504 43336
rect 25556 43324 25562 43376
rect 11146 43296 11152 43308
rect 10810 43268 11152 43296
rect 11146 43256 11152 43268
rect 11204 43296 11210 43308
rect 11698 43296 11704 43308
rect 11204 43268 11704 43296
rect 11204 43256 11210 43268
rect 11698 43256 11704 43268
rect 11756 43256 11762 43308
rect 9214 43188 9220 43240
rect 9272 43228 9278 43240
rect 9401 43231 9459 43237
rect 9401 43228 9413 43231
rect 9272 43200 9413 43228
rect 9272 43188 9278 43200
rect 9401 43197 9413 43200
rect 9447 43197 9459 43231
rect 9401 43191 9459 43197
rect 9677 43231 9735 43237
rect 9677 43197 9689 43231
rect 9723 43228 9735 43231
rect 12342 43228 12348 43240
rect 9723 43200 12348 43228
rect 9723 43197 9735 43200
rect 9677 43191 9735 43197
rect 9416 43092 9444 43191
rect 12342 43188 12348 43200
rect 12400 43188 12406 43240
rect 11054 43160 11060 43172
rect 10704 43132 11060 43160
rect 10704 43092 10732 43132
rect 11054 43120 11060 43132
rect 11112 43160 11118 43172
rect 25317 43163 25375 43169
rect 11112 43132 11652 43160
rect 11112 43120 11118 43132
rect 11624 43104 11652 43132
rect 25317 43129 25329 43163
rect 25363 43160 25375 43163
rect 25590 43160 25596 43172
rect 25363 43132 25596 43160
rect 25363 43129 25375 43132
rect 25317 43123 25375 43129
rect 25590 43120 25596 43132
rect 25648 43120 25654 43172
rect 9416 43064 10732 43092
rect 11606 43052 11612 43104
rect 11664 43052 11670 43104
rect 1104 43002 25852 43024
rect 1104 42950 2950 43002
rect 3002 42950 3014 43002
rect 3066 42950 3078 43002
rect 3130 42950 3142 43002
rect 3194 42950 3206 43002
rect 3258 42950 12950 43002
rect 13002 42950 13014 43002
rect 13066 42950 13078 43002
rect 13130 42950 13142 43002
rect 13194 42950 13206 43002
rect 13258 42950 22950 43002
rect 23002 42950 23014 43002
rect 23066 42950 23078 43002
rect 23130 42950 23142 43002
rect 23194 42950 23206 43002
rect 23258 42950 25852 43002
rect 1104 42928 25852 42950
rect 24765 42619 24823 42625
rect 24765 42585 24777 42619
rect 24811 42616 24823 42619
rect 25130 42616 25136 42628
rect 24811 42588 25136 42616
rect 24811 42585 24823 42588
rect 24765 42579 24823 42585
rect 25130 42576 25136 42588
rect 25188 42576 25194 42628
rect 25317 42619 25375 42625
rect 25317 42585 25329 42619
rect 25363 42616 25375 42619
rect 26142 42616 26148 42628
rect 25363 42588 26148 42616
rect 25363 42585 25375 42588
rect 25317 42579 25375 42585
rect 26142 42576 26148 42588
rect 26200 42576 26206 42628
rect 1104 42458 25852 42480
rect 1104 42406 7950 42458
rect 8002 42406 8014 42458
rect 8066 42406 8078 42458
rect 8130 42406 8142 42458
rect 8194 42406 8206 42458
rect 8258 42406 17950 42458
rect 18002 42406 18014 42458
rect 18066 42406 18078 42458
rect 18130 42406 18142 42458
rect 18194 42406 18206 42458
rect 18258 42406 25852 42458
rect 1104 42384 25852 42406
rect 25130 41964 25136 42016
rect 25188 42004 25194 42016
rect 25409 42007 25467 42013
rect 25409 42004 25421 42007
rect 25188 41976 25421 42004
rect 25188 41964 25194 41976
rect 25409 41973 25421 41976
rect 25455 41973 25467 42007
rect 25409 41967 25467 41973
rect 1104 41914 25852 41936
rect 1104 41862 2950 41914
rect 3002 41862 3014 41914
rect 3066 41862 3078 41914
rect 3130 41862 3142 41914
rect 3194 41862 3206 41914
rect 3258 41862 12950 41914
rect 13002 41862 13014 41914
rect 13066 41862 13078 41914
rect 13130 41862 13142 41914
rect 13194 41862 13206 41914
rect 13258 41862 22950 41914
rect 23002 41862 23014 41914
rect 23066 41862 23078 41914
rect 23130 41862 23142 41914
rect 23194 41862 23206 41914
rect 23258 41862 25852 41914
rect 1104 41840 25852 41862
rect 25130 41556 25136 41608
rect 25188 41556 25194 41608
rect 25317 41531 25375 41537
rect 25317 41497 25329 41531
rect 25363 41528 25375 41531
rect 25866 41528 25872 41540
rect 25363 41500 25872 41528
rect 25363 41497 25375 41500
rect 25317 41491 25375 41497
rect 25866 41488 25872 41500
rect 25924 41488 25930 41540
rect 16850 41420 16856 41472
rect 16908 41460 16914 41472
rect 23934 41460 23940 41472
rect 16908 41432 23940 41460
rect 16908 41420 16914 41432
rect 23934 41420 23940 41432
rect 23992 41420 23998 41472
rect 1104 41370 25852 41392
rect 1104 41318 7950 41370
rect 8002 41318 8014 41370
rect 8066 41318 8078 41370
rect 8130 41318 8142 41370
rect 8194 41318 8206 41370
rect 8258 41318 17950 41370
rect 18002 41318 18014 41370
rect 18066 41318 18078 41370
rect 18130 41318 18142 41370
rect 18194 41318 18206 41370
rect 18258 41318 25852 41370
rect 1104 41296 25852 41318
rect 24857 41123 24915 41129
rect 24857 41089 24869 41123
rect 24903 41120 24915 41123
rect 25314 41120 25320 41132
rect 24903 41092 25320 41120
rect 24903 41089 24915 41092
rect 24857 41083 24915 41089
rect 25314 41080 25320 41092
rect 25372 41080 25378 41132
rect 25133 40919 25191 40925
rect 25133 40885 25145 40919
rect 25179 40916 25191 40919
rect 25222 40916 25228 40928
rect 25179 40888 25228 40916
rect 25179 40885 25191 40888
rect 25133 40879 25191 40885
rect 25222 40876 25228 40888
rect 25280 40876 25286 40928
rect 1104 40826 25852 40848
rect 1104 40774 2950 40826
rect 3002 40774 3014 40826
rect 3066 40774 3078 40826
rect 3130 40774 3142 40826
rect 3194 40774 3206 40826
rect 3258 40774 12950 40826
rect 13002 40774 13014 40826
rect 13066 40774 13078 40826
rect 13130 40774 13142 40826
rect 13194 40774 13206 40826
rect 13258 40774 22950 40826
rect 23002 40774 23014 40826
rect 23066 40774 23078 40826
rect 23130 40774 23142 40826
rect 23194 40774 23206 40826
rect 23258 40774 25852 40826
rect 1104 40752 25852 40774
rect 25406 40332 25412 40384
rect 25464 40332 25470 40384
rect 1104 40282 25852 40304
rect 1104 40230 7950 40282
rect 8002 40230 8014 40282
rect 8066 40230 8078 40282
rect 8130 40230 8142 40282
rect 8194 40230 8206 40282
rect 8258 40230 17950 40282
rect 18002 40230 18014 40282
rect 18066 40230 18078 40282
rect 18130 40230 18142 40282
rect 18194 40230 18206 40282
rect 18258 40230 25852 40282
rect 1104 40208 25852 40230
rect 12342 40128 12348 40180
rect 12400 40128 12406 40180
rect 25038 40128 25044 40180
rect 25096 40168 25102 40180
rect 25133 40171 25191 40177
rect 25133 40168 25145 40171
rect 25096 40140 25145 40168
rect 25096 40128 25102 40140
rect 25133 40137 25145 40140
rect 25179 40137 25191 40171
rect 25133 40131 25191 40137
rect 25406 40100 25412 40112
rect 25332 40072 25412 40100
rect 11330 39992 11336 40044
rect 11388 40032 11394 40044
rect 11701 40035 11759 40041
rect 11701 40032 11713 40035
rect 11388 40004 11713 40032
rect 11388 39992 11394 40004
rect 11701 40001 11713 40004
rect 11747 40001 11759 40035
rect 11701 39995 11759 40001
rect 21174 39992 21180 40044
rect 21232 40032 21238 40044
rect 23290 40032 23296 40044
rect 21232 40004 23296 40032
rect 21232 39992 21238 40004
rect 23290 39992 23296 40004
rect 23348 39992 23354 40044
rect 25332 40041 25360 40072
rect 25406 40060 25412 40072
rect 25464 40060 25470 40112
rect 25317 40035 25375 40041
rect 25317 40001 25329 40035
rect 25363 40001 25375 40035
rect 25317 39995 25375 40001
rect 1104 39738 25852 39760
rect 1104 39686 2950 39738
rect 3002 39686 3014 39738
rect 3066 39686 3078 39738
rect 3130 39686 3142 39738
rect 3194 39686 3206 39738
rect 3258 39686 12950 39738
rect 13002 39686 13014 39738
rect 13066 39686 13078 39738
rect 13130 39686 13142 39738
rect 13194 39686 13206 39738
rect 13258 39686 22950 39738
rect 23002 39686 23014 39738
rect 23066 39686 23078 39738
rect 23130 39686 23142 39738
rect 23194 39686 23206 39738
rect 23258 39686 25852 39738
rect 1104 39664 25852 39686
rect 7742 39584 7748 39636
rect 7800 39624 7806 39636
rect 9125 39627 9183 39633
rect 9125 39624 9137 39627
rect 7800 39596 9137 39624
rect 7800 39584 7806 39596
rect 9125 39593 9137 39596
rect 9171 39593 9183 39627
rect 9125 39587 9183 39593
rect 9309 39423 9367 39429
rect 9309 39389 9321 39423
rect 9355 39420 9367 39423
rect 9766 39420 9772 39432
rect 9355 39392 9772 39420
rect 9355 39389 9367 39392
rect 9309 39383 9367 39389
rect 9766 39380 9772 39392
rect 9824 39380 9830 39432
rect 24857 39423 24915 39429
rect 24857 39389 24869 39423
rect 24903 39420 24915 39423
rect 25314 39420 25320 39432
rect 24903 39392 25320 39420
rect 24903 39389 24915 39392
rect 24857 39383 24915 39389
rect 25314 39380 25320 39392
rect 25372 39380 25378 39432
rect 22002 39244 22008 39296
rect 22060 39284 22066 39296
rect 25133 39287 25191 39293
rect 25133 39284 25145 39287
rect 22060 39256 25145 39284
rect 22060 39244 22066 39256
rect 25133 39253 25145 39256
rect 25179 39253 25191 39287
rect 25133 39247 25191 39253
rect 1104 39194 25852 39216
rect 1104 39142 7950 39194
rect 8002 39142 8014 39194
rect 8066 39142 8078 39194
rect 8130 39142 8142 39194
rect 8194 39142 8206 39194
rect 8258 39142 17950 39194
rect 18002 39142 18014 39194
rect 18066 39142 18078 39194
rect 18130 39142 18142 39194
rect 18194 39142 18206 39194
rect 18258 39142 25852 39194
rect 1104 39120 25852 39142
rect 25314 38700 25320 38752
rect 25372 38740 25378 38752
rect 25409 38743 25467 38749
rect 25409 38740 25421 38743
rect 25372 38712 25421 38740
rect 25372 38700 25378 38712
rect 25409 38709 25421 38712
rect 25455 38709 25467 38743
rect 25409 38703 25467 38709
rect 1104 38650 25852 38672
rect 1104 38598 2950 38650
rect 3002 38598 3014 38650
rect 3066 38598 3078 38650
rect 3130 38598 3142 38650
rect 3194 38598 3206 38650
rect 3258 38598 12950 38650
rect 13002 38598 13014 38650
rect 13066 38598 13078 38650
rect 13130 38598 13142 38650
rect 13194 38598 13206 38650
rect 13258 38598 22950 38650
rect 23002 38598 23014 38650
rect 23066 38598 23078 38650
rect 23130 38598 23142 38650
rect 23194 38598 23206 38650
rect 23258 38598 25852 38650
rect 1104 38576 25852 38598
rect 22462 38496 22468 38548
rect 22520 38536 22526 38548
rect 24210 38536 24216 38548
rect 22520 38508 24216 38536
rect 22520 38496 22526 38508
rect 24210 38496 24216 38508
rect 24268 38496 24274 38548
rect 16666 38292 16672 38344
rect 16724 38332 16730 38344
rect 17681 38335 17739 38341
rect 17681 38332 17693 38335
rect 16724 38304 17693 38332
rect 16724 38292 16730 38304
rect 17681 38301 17693 38304
rect 17727 38332 17739 38335
rect 22186 38332 22192 38344
rect 17727 38304 22192 38332
rect 17727 38301 17739 38304
rect 17681 38295 17739 38301
rect 22186 38292 22192 38304
rect 22244 38292 22250 38344
rect 25314 38292 25320 38344
rect 25372 38292 25378 38344
rect 16758 38156 16764 38208
rect 16816 38196 16822 38208
rect 18325 38199 18383 38205
rect 18325 38196 18337 38199
rect 16816 38168 18337 38196
rect 16816 38156 16822 38168
rect 18325 38165 18337 38168
rect 18371 38165 18383 38199
rect 18325 38159 18383 38165
rect 20530 38156 20536 38208
rect 20588 38196 20594 38208
rect 25133 38199 25191 38205
rect 25133 38196 25145 38199
rect 20588 38168 25145 38196
rect 20588 38156 20594 38168
rect 25133 38165 25145 38168
rect 25179 38165 25191 38199
rect 25133 38159 25191 38165
rect 1104 38106 25852 38128
rect 1104 38054 7950 38106
rect 8002 38054 8014 38106
rect 8066 38054 8078 38106
rect 8130 38054 8142 38106
rect 8194 38054 8206 38106
rect 8258 38054 17950 38106
rect 18002 38054 18014 38106
rect 18066 38054 18078 38106
rect 18130 38054 18142 38106
rect 18194 38054 18206 38106
rect 18258 38054 25852 38106
rect 1104 38032 25852 38054
rect 24765 37859 24823 37865
rect 24765 37825 24777 37859
rect 24811 37856 24823 37859
rect 25130 37856 25136 37868
rect 24811 37828 25136 37856
rect 24811 37825 24823 37828
rect 24765 37819 24823 37825
rect 25130 37816 25136 37828
rect 25188 37816 25194 37868
rect 25317 37723 25375 37729
rect 25317 37689 25329 37723
rect 25363 37720 25375 37723
rect 26602 37720 26608 37732
rect 25363 37692 26608 37720
rect 25363 37689 25375 37692
rect 25317 37683 25375 37689
rect 26602 37680 26608 37692
rect 26660 37680 26666 37732
rect 1104 37562 25852 37584
rect 1104 37510 2950 37562
rect 3002 37510 3014 37562
rect 3066 37510 3078 37562
rect 3130 37510 3142 37562
rect 3194 37510 3206 37562
rect 3258 37510 12950 37562
rect 13002 37510 13014 37562
rect 13066 37510 13078 37562
rect 13130 37510 13142 37562
rect 13194 37510 13206 37562
rect 13258 37510 22950 37562
rect 23002 37510 23014 37562
rect 23066 37510 23078 37562
rect 23130 37510 23142 37562
rect 23194 37510 23206 37562
rect 23258 37510 25852 37562
rect 1104 37488 25852 37510
rect 24857 37247 24915 37253
rect 24857 37213 24869 37247
rect 24903 37244 24915 37247
rect 25314 37244 25320 37256
rect 24903 37216 25320 37244
rect 24903 37213 24915 37216
rect 24857 37207 24915 37213
rect 25314 37204 25320 37216
rect 25372 37204 25378 37256
rect 25133 37111 25191 37117
rect 25133 37077 25145 37111
rect 25179 37108 25191 37111
rect 25682 37108 25688 37120
rect 25179 37080 25688 37108
rect 25179 37077 25191 37080
rect 25133 37071 25191 37077
rect 25682 37068 25688 37080
rect 25740 37068 25746 37120
rect 1104 37018 25852 37040
rect 1104 36966 7950 37018
rect 8002 36966 8014 37018
rect 8066 36966 8078 37018
rect 8130 36966 8142 37018
rect 8194 36966 8206 37018
rect 8258 36966 17950 37018
rect 18002 36966 18014 37018
rect 18066 36966 18078 37018
rect 18130 36966 18142 37018
rect 18194 36966 18206 37018
rect 18258 36966 25852 37018
rect 1104 36944 25852 36966
rect 11149 36907 11207 36913
rect 11149 36873 11161 36907
rect 11195 36904 11207 36907
rect 11330 36904 11336 36916
rect 11195 36876 11336 36904
rect 11195 36873 11207 36876
rect 11149 36867 11207 36873
rect 11330 36864 11336 36876
rect 11388 36864 11394 36916
rect 11698 36864 11704 36916
rect 11756 36864 11762 36916
rect 11238 36836 11244 36848
rect 10902 36808 11244 36836
rect 11238 36796 11244 36808
rect 11296 36836 11302 36848
rect 11716 36836 11744 36864
rect 11296 36808 11744 36836
rect 11296 36796 11302 36808
rect 24765 36771 24823 36777
rect 24765 36737 24777 36771
rect 24811 36768 24823 36771
rect 25130 36768 25136 36780
rect 24811 36740 25136 36768
rect 24811 36737 24823 36740
rect 24765 36731 24823 36737
rect 25130 36728 25136 36740
rect 25188 36728 25194 36780
rect 9401 36703 9459 36709
rect 9401 36669 9413 36703
rect 9447 36669 9459 36703
rect 9401 36663 9459 36669
rect 9416 36564 9444 36663
rect 9674 36660 9680 36712
rect 9732 36660 9738 36712
rect 25317 36635 25375 36641
rect 10704 36604 11652 36632
rect 10704 36564 10732 36604
rect 11624 36576 11652 36604
rect 25317 36601 25329 36635
rect 25363 36632 25375 36635
rect 26694 36632 26700 36644
rect 25363 36604 26700 36632
rect 25363 36601 25375 36604
rect 25317 36595 25375 36601
rect 26694 36592 26700 36604
rect 26752 36592 26758 36644
rect 9416 36536 10732 36564
rect 11606 36524 11612 36576
rect 11664 36524 11670 36576
rect 1104 36474 25852 36496
rect 1104 36422 2950 36474
rect 3002 36422 3014 36474
rect 3066 36422 3078 36474
rect 3130 36422 3142 36474
rect 3194 36422 3206 36474
rect 3258 36422 12950 36474
rect 13002 36422 13014 36474
rect 13066 36422 13078 36474
rect 13130 36422 13142 36474
rect 13194 36422 13206 36474
rect 13258 36422 22950 36474
rect 23002 36422 23014 36474
rect 23066 36422 23078 36474
rect 23130 36422 23142 36474
rect 23194 36422 23206 36474
rect 23258 36422 25852 36474
rect 1104 36400 25852 36422
rect 9030 36320 9036 36372
rect 9088 36360 9094 36372
rect 9125 36363 9183 36369
rect 9125 36360 9137 36363
rect 9088 36332 9137 36360
rect 9088 36320 9094 36332
rect 9125 36329 9137 36332
rect 9171 36329 9183 36363
rect 9125 36323 9183 36329
rect 9214 36116 9220 36168
rect 9272 36156 9278 36168
rect 9309 36159 9367 36165
rect 9309 36156 9321 36159
rect 9272 36128 9321 36156
rect 9272 36116 9278 36128
rect 9309 36125 9321 36128
rect 9355 36125 9367 36159
rect 25317 36159 25375 36165
rect 25317 36156 25329 36159
rect 9309 36119 9367 36125
rect 24872 36128 25329 36156
rect 24762 35980 24768 36032
rect 24820 36020 24826 36032
rect 24872 36029 24900 36128
rect 25317 36125 25329 36128
rect 25363 36125 25375 36159
rect 25317 36119 25375 36125
rect 24857 36023 24915 36029
rect 24857 36020 24869 36023
rect 24820 35992 24869 36020
rect 24820 35980 24826 35992
rect 24857 35989 24869 35992
rect 24903 35989 24915 36023
rect 24857 35983 24915 35989
rect 25133 36023 25191 36029
rect 25133 35989 25145 36023
rect 25179 36020 25191 36023
rect 25498 36020 25504 36032
rect 25179 35992 25504 36020
rect 25179 35989 25191 35992
rect 25133 35983 25191 35989
rect 25498 35980 25504 35992
rect 25556 35980 25562 36032
rect 1104 35930 25852 35952
rect 1104 35878 7950 35930
rect 8002 35878 8014 35930
rect 8066 35878 8078 35930
rect 8130 35878 8142 35930
rect 8194 35878 8206 35930
rect 8258 35878 17950 35930
rect 18002 35878 18014 35930
rect 18066 35878 18078 35930
rect 18130 35878 18142 35930
rect 18194 35878 18206 35930
rect 18258 35878 25852 35930
rect 1104 35856 25852 35878
rect 16114 35776 16120 35828
rect 16172 35816 16178 35828
rect 20349 35819 20407 35825
rect 20349 35816 20361 35819
rect 16172 35788 20361 35816
rect 16172 35776 16178 35788
rect 20349 35785 20361 35788
rect 20395 35816 20407 35819
rect 21085 35819 21143 35825
rect 21085 35816 21097 35819
rect 20395 35788 21097 35816
rect 20395 35785 20407 35788
rect 20349 35779 20407 35785
rect 21085 35785 21097 35788
rect 21131 35785 21143 35819
rect 21085 35779 21143 35785
rect 21100 35748 21128 35779
rect 21174 35776 21180 35828
rect 21232 35776 21238 35828
rect 22462 35776 22468 35828
rect 22520 35776 22526 35828
rect 22830 35776 22836 35828
rect 22888 35816 22894 35828
rect 25133 35819 25191 35825
rect 25133 35816 25145 35819
rect 22888 35788 25145 35816
rect 22888 35776 22894 35788
rect 25133 35785 25145 35788
rect 25179 35785 25191 35819
rect 25133 35779 25191 35785
rect 24946 35748 24952 35760
rect 21100 35720 24952 35748
rect 24946 35708 24952 35720
rect 25004 35708 25010 35760
rect 16298 35640 16304 35692
rect 16356 35680 16362 35692
rect 21818 35680 21824 35692
rect 16356 35652 21824 35680
rect 16356 35640 16362 35652
rect 21818 35640 21824 35652
rect 21876 35680 21882 35692
rect 22373 35683 22431 35689
rect 22373 35680 22385 35683
rect 21876 35652 22385 35680
rect 21876 35640 21882 35652
rect 22373 35649 22385 35652
rect 22419 35649 22431 35683
rect 25317 35683 25375 35689
rect 25317 35680 25329 35683
rect 22373 35643 22431 35649
rect 24872 35652 25329 35680
rect 21266 35572 21272 35624
rect 21324 35572 21330 35624
rect 22094 35572 22100 35624
rect 22152 35612 22158 35624
rect 22557 35615 22615 35621
rect 22557 35612 22569 35615
rect 22152 35584 22569 35612
rect 22152 35572 22158 35584
rect 22557 35581 22569 35584
rect 22603 35581 22615 35615
rect 22557 35575 22615 35581
rect 19886 35504 19892 35556
rect 19944 35544 19950 35556
rect 20717 35547 20775 35553
rect 20717 35544 20729 35547
rect 19944 35516 20729 35544
rect 19944 35504 19950 35516
rect 20717 35513 20729 35516
rect 20763 35513 20775 35547
rect 20717 35507 20775 35513
rect 20622 35436 20628 35488
rect 20680 35476 20686 35488
rect 22005 35479 22063 35485
rect 22005 35476 22017 35479
rect 20680 35448 22017 35476
rect 20680 35436 20686 35448
rect 22005 35445 22017 35448
rect 22051 35445 22063 35479
rect 22005 35439 22063 35445
rect 24762 35436 24768 35488
rect 24820 35476 24826 35488
rect 24872 35485 24900 35652
rect 25317 35649 25329 35652
rect 25363 35649 25375 35683
rect 25317 35643 25375 35649
rect 24857 35479 24915 35485
rect 24857 35476 24869 35479
rect 24820 35448 24869 35476
rect 24820 35436 24826 35448
rect 24857 35445 24869 35448
rect 24903 35445 24915 35479
rect 24857 35439 24915 35445
rect 1104 35386 25852 35408
rect 1104 35334 2950 35386
rect 3002 35334 3014 35386
rect 3066 35334 3078 35386
rect 3130 35334 3142 35386
rect 3194 35334 3206 35386
rect 3258 35334 12950 35386
rect 13002 35334 13014 35386
rect 13066 35334 13078 35386
rect 13130 35334 13142 35386
rect 13194 35334 13206 35386
rect 13258 35334 22950 35386
rect 23002 35334 23014 35386
rect 23066 35334 23078 35386
rect 23130 35334 23142 35386
rect 23194 35334 23206 35386
rect 23258 35334 25852 35386
rect 1104 35312 25852 35334
rect 17494 35232 17500 35284
rect 17552 35272 17558 35284
rect 22373 35275 22431 35281
rect 22373 35272 22385 35275
rect 17552 35244 22385 35272
rect 17552 35232 17558 35244
rect 22373 35241 22385 35244
rect 22419 35241 22431 35275
rect 22373 35235 22431 35241
rect 24857 35275 24915 35281
rect 24857 35241 24869 35275
rect 24903 35272 24915 35275
rect 24946 35272 24952 35284
rect 24903 35244 24952 35272
rect 24903 35241 24915 35244
rect 24857 35235 24915 35241
rect 21358 35164 21364 35216
rect 21416 35164 21422 35216
rect 21818 35164 21824 35216
rect 21876 35164 21882 35216
rect 19610 35028 19616 35080
rect 19668 35028 19674 35080
rect 22186 35028 22192 35080
rect 22244 35068 22250 35080
rect 22388 35068 22416 35235
rect 24946 35232 24952 35244
rect 25004 35272 25010 35284
rect 25314 35272 25320 35284
rect 25004 35244 25320 35272
rect 25004 35232 25010 35244
rect 25314 35232 25320 35244
rect 25372 35232 25378 35284
rect 24118 35164 24124 35216
rect 24176 35204 24182 35216
rect 25133 35207 25191 35213
rect 25133 35204 25145 35207
rect 24176 35176 25145 35204
rect 24176 35164 24182 35176
rect 25133 35173 25145 35176
rect 25179 35173 25191 35207
rect 25133 35167 25191 35173
rect 23290 35096 23296 35148
rect 23348 35096 23354 35148
rect 23109 35071 23167 35077
rect 23109 35068 23121 35071
rect 22244 35040 23121 35068
rect 22244 35028 22250 35040
rect 23109 35037 23121 35040
rect 23155 35037 23167 35071
rect 23109 35031 23167 35037
rect 23201 35071 23259 35077
rect 23201 35037 23213 35071
rect 23247 35068 23259 35071
rect 23382 35068 23388 35080
rect 23247 35040 23388 35068
rect 23247 35037 23259 35040
rect 23201 35031 23259 35037
rect 23382 35028 23388 35040
rect 23440 35028 23446 35080
rect 24578 35028 24584 35080
rect 24636 35068 24642 35080
rect 25317 35071 25375 35077
rect 25317 35068 25329 35071
rect 24636 35040 25329 35068
rect 24636 35028 24642 35040
rect 25317 35037 25329 35040
rect 25363 35037 25375 35071
rect 25317 35031 25375 35037
rect 24489 35003 24547 35009
rect 24489 34969 24501 35003
rect 24535 35000 24547 35003
rect 24670 35000 24676 35012
rect 24535 34972 24676 35000
rect 24535 34969 24547 34972
rect 24489 34963 24547 34969
rect 24670 34960 24676 34972
rect 24728 34960 24734 35012
rect 19702 34892 19708 34944
rect 19760 34932 19766 34944
rect 20257 34935 20315 34941
rect 20257 34932 20269 34935
rect 19760 34904 20269 34932
rect 19760 34892 19766 34904
rect 20257 34901 20269 34904
rect 20303 34901 20315 34935
rect 20257 34895 20315 34901
rect 22462 34892 22468 34944
rect 22520 34932 22526 34944
rect 22741 34935 22799 34941
rect 22741 34932 22753 34935
rect 22520 34904 22753 34932
rect 22520 34892 22526 34904
rect 22741 34901 22753 34904
rect 22787 34901 22799 34935
rect 22741 34895 22799 34901
rect 24578 34892 24584 34944
rect 24636 34892 24642 34944
rect 1104 34842 25852 34864
rect 1104 34790 7950 34842
rect 8002 34790 8014 34842
rect 8066 34790 8078 34842
rect 8130 34790 8142 34842
rect 8194 34790 8206 34842
rect 8258 34790 17950 34842
rect 18002 34790 18014 34842
rect 18066 34790 18078 34842
rect 18130 34790 18142 34842
rect 18194 34790 18206 34842
rect 18258 34790 25852 34842
rect 1104 34768 25852 34790
rect 23658 34688 23664 34740
rect 23716 34728 23722 34740
rect 24489 34731 24547 34737
rect 24489 34728 24501 34731
rect 23716 34700 24501 34728
rect 23716 34688 23722 34700
rect 24489 34697 24501 34700
rect 24535 34697 24547 34731
rect 24489 34691 24547 34697
rect 11606 34620 11612 34672
rect 11664 34660 11670 34672
rect 15841 34663 15899 34669
rect 15841 34660 15853 34663
rect 11664 34632 15853 34660
rect 11664 34620 11670 34632
rect 15841 34629 15853 34632
rect 15887 34629 15899 34663
rect 15841 34623 15899 34629
rect 15105 34595 15163 34601
rect 15105 34561 15117 34595
rect 15151 34561 15163 34595
rect 15105 34555 15163 34561
rect 15120 34524 15148 34555
rect 19334 34552 19340 34604
rect 19392 34592 19398 34604
rect 19429 34595 19487 34601
rect 19429 34592 19441 34595
rect 19392 34564 19441 34592
rect 19392 34552 19398 34564
rect 19429 34561 19441 34564
rect 19475 34561 19487 34595
rect 19429 34555 19487 34561
rect 20809 34595 20867 34601
rect 20809 34561 20821 34595
rect 20855 34592 20867 34595
rect 21266 34592 21272 34604
rect 20855 34564 21272 34592
rect 20855 34561 20867 34564
rect 20809 34555 20867 34561
rect 21266 34552 21272 34564
rect 21324 34552 21330 34604
rect 22005 34595 22063 34601
rect 22005 34561 22017 34595
rect 22051 34592 22063 34595
rect 22094 34592 22100 34604
rect 22051 34564 22100 34592
rect 22051 34561 22063 34564
rect 22005 34555 22063 34561
rect 22094 34552 22100 34564
rect 22152 34552 22158 34604
rect 23109 34595 23167 34601
rect 23109 34561 23121 34595
rect 23155 34592 23167 34595
rect 23290 34592 23296 34604
rect 23155 34564 23296 34592
rect 23155 34561 23167 34564
rect 23109 34555 23167 34561
rect 23290 34552 23296 34564
rect 23348 34552 23354 34604
rect 24670 34552 24676 34604
rect 24728 34552 24734 34604
rect 25317 34595 25375 34601
rect 25317 34561 25329 34595
rect 25363 34561 25375 34595
rect 25317 34555 25375 34561
rect 16393 34527 16451 34533
rect 16393 34524 16405 34527
rect 15120 34496 16405 34524
rect 16393 34493 16405 34496
rect 16439 34524 16451 34527
rect 16439 34496 16574 34524
rect 16439 34493 16451 34496
rect 16393 34487 16451 34493
rect 16546 34468 16574 34496
rect 20070 34484 20076 34536
rect 20128 34484 20134 34536
rect 20254 34484 20260 34536
rect 20312 34524 20318 34536
rect 21453 34527 21511 34533
rect 21453 34524 21465 34527
rect 20312 34496 21465 34524
rect 20312 34484 20318 34496
rect 21453 34493 21465 34496
rect 21499 34493 21511 34527
rect 21453 34487 21511 34493
rect 21542 34484 21548 34536
rect 21600 34524 21606 34536
rect 22649 34527 22707 34533
rect 22649 34524 22661 34527
rect 21600 34496 22661 34524
rect 21600 34484 21606 34496
rect 22649 34493 22661 34496
rect 22695 34493 22707 34527
rect 22649 34487 22707 34493
rect 24213 34527 24271 34533
rect 24213 34493 24225 34527
rect 24259 34524 24271 34527
rect 24486 34524 24492 34536
rect 24259 34496 24492 34524
rect 24259 34493 24271 34496
rect 24213 34487 24271 34493
rect 24486 34484 24492 34496
rect 24544 34524 24550 34536
rect 25332 34524 25360 34555
rect 24544 34496 25360 34524
rect 24544 34484 24550 34496
rect 16546 34428 16580 34468
rect 16574 34416 16580 34428
rect 16632 34416 16638 34468
rect 23750 34348 23756 34400
rect 23808 34348 23814 34400
rect 25130 34348 25136 34400
rect 25188 34348 25194 34400
rect 1104 34298 25852 34320
rect 1104 34246 2950 34298
rect 3002 34246 3014 34298
rect 3066 34246 3078 34298
rect 3130 34246 3142 34298
rect 3194 34246 3206 34298
rect 3258 34246 12950 34298
rect 13002 34246 13014 34298
rect 13066 34246 13078 34298
rect 13130 34246 13142 34298
rect 13194 34246 13206 34298
rect 13258 34246 22950 34298
rect 23002 34246 23014 34298
rect 23066 34246 23078 34298
rect 23130 34246 23142 34298
rect 23194 34246 23206 34298
rect 23258 34246 25852 34298
rect 1104 34224 25852 34246
rect 21177 34187 21235 34193
rect 21177 34153 21189 34187
rect 21223 34184 21235 34187
rect 21266 34184 21272 34196
rect 21223 34156 21272 34184
rect 21223 34153 21235 34156
rect 21177 34147 21235 34153
rect 21266 34144 21272 34156
rect 21324 34144 21330 34196
rect 22094 34144 22100 34196
rect 22152 34184 22158 34196
rect 23385 34187 23443 34193
rect 23385 34184 23397 34187
rect 22152 34156 23397 34184
rect 22152 34144 22158 34156
rect 23385 34153 23397 34156
rect 23431 34153 23443 34187
rect 23385 34147 23443 34153
rect 19426 34076 19432 34128
rect 19484 34076 19490 34128
rect 19444 34048 19472 34076
rect 21637 34051 21695 34057
rect 21637 34048 21649 34051
rect 19444 34020 21649 34048
rect 21637 34017 21649 34020
rect 21683 34048 21695 34051
rect 22278 34048 22284 34060
rect 21683 34020 22284 34048
rect 21683 34017 21695 34020
rect 21637 34011 21695 34017
rect 22278 34008 22284 34020
rect 22336 34008 22342 34060
rect 17402 33940 17408 33992
rect 17460 33980 17466 33992
rect 18049 33983 18107 33989
rect 18049 33980 18061 33983
rect 17460 33952 18061 33980
rect 17460 33940 17466 33952
rect 18049 33949 18061 33952
rect 18095 33980 18107 33983
rect 19429 33983 19487 33989
rect 19429 33980 19441 33983
rect 18095 33952 19441 33980
rect 18095 33949 18107 33952
rect 18049 33943 18107 33949
rect 19429 33949 19441 33952
rect 19475 33949 19487 33983
rect 19429 33943 19487 33949
rect 23474 33940 23480 33992
rect 23532 33980 23538 33992
rect 24581 33983 24639 33989
rect 24581 33980 24593 33983
rect 23532 33952 24593 33980
rect 23532 33940 23538 33952
rect 24581 33949 24593 33952
rect 24627 33949 24639 33983
rect 24581 33943 24639 33949
rect 17221 33915 17279 33921
rect 17221 33912 17233 33915
rect 16868 33884 17233 33912
rect 16574 33804 16580 33856
rect 16632 33844 16638 33856
rect 16868 33853 16896 33884
rect 17221 33881 17233 33884
rect 17267 33881 17279 33915
rect 17221 33875 17279 33881
rect 19702 33872 19708 33924
rect 19760 33872 19766 33924
rect 21358 33912 21364 33924
rect 20930 33884 21364 33912
rect 21358 33872 21364 33884
rect 21416 33872 21422 33924
rect 21913 33915 21971 33921
rect 21913 33881 21925 33915
rect 21959 33912 21971 33915
rect 21959 33884 22094 33912
rect 21959 33881 21971 33884
rect 21913 33875 21971 33881
rect 16853 33847 16911 33853
rect 16853 33844 16865 33847
rect 16632 33816 16865 33844
rect 16632 33804 16638 33816
rect 16853 33813 16865 33816
rect 16899 33813 16911 33847
rect 22066 33844 22094 33884
rect 22370 33872 22376 33924
rect 22428 33872 22434 33924
rect 25225 33915 25283 33921
rect 25225 33912 25237 33915
rect 23308 33884 25237 33912
rect 23308 33844 23336 33884
rect 25225 33881 25237 33884
rect 25271 33881 25283 33915
rect 25225 33875 25283 33881
rect 22066 33816 23336 33844
rect 16853 33807 16911 33813
rect 23566 33804 23572 33856
rect 23624 33844 23630 33856
rect 23661 33847 23719 33853
rect 23661 33844 23673 33847
rect 23624 33816 23673 33844
rect 23624 33804 23630 33816
rect 23661 33813 23673 33816
rect 23707 33844 23719 33847
rect 23845 33847 23903 33853
rect 23845 33844 23857 33847
rect 23707 33816 23857 33844
rect 23707 33813 23719 33816
rect 23661 33807 23719 33813
rect 23845 33813 23857 33816
rect 23891 33813 23903 33847
rect 23845 33807 23903 33813
rect 24121 33847 24179 33853
rect 24121 33813 24133 33847
rect 24167 33844 24179 33847
rect 24394 33844 24400 33856
rect 24167 33816 24400 33844
rect 24167 33813 24179 33816
rect 24121 33807 24179 33813
rect 24394 33804 24400 33816
rect 24452 33804 24458 33856
rect 1104 33754 25852 33776
rect 1104 33702 7950 33754
rect 8002 33702 8014 33754
rect 8066 33702 8078 33754
rect 8130 33702 8142 33754
rect 8194 33702 8206 33754
rect 8258 33702 17950 33754
rect 18002 33702 18014 33754
rect 18066 33702 18078 33754
rect 18130 33702 18142 33754
rect 18194 33702 18206 33754
rect 18258 33702 25852 33754
rect 1104 33680 25852 33702
rect 9674 33600 9680 33652
rect 9732 33640 9738 33652
rect 10045 33643 10103 33649
rect 10045 33640 10057 33643
rect 9732 33612 10057 33640
rect 9732 33600 9738 33612
rect 10045 33609 10057 33612
rect 10091 33609 10103 33643
rect 10045 33603 10103 33609
rect 19610 33600 19616 33652
rect 19668 33640 19674 33652
rect 20438 33640 20444 33652
rect 19668 33612 20444 33640
rect 19668 33600 19674 33612
rect 20438 33600 20444 33612
rect 20496 33640 20502 33652
rect 21177 33643 21235 33649
rect 21177 33640 21189 33643
rect 20496 33612 21189 33640
rect 20496 33600 20502 33612
rect 21177 33609 21189 33612
rect 21223 33609 21235 33643
rect 21177 33603 21235 33609
rect 21358 33600 21364 33652
rect 21416 33640 21422 33652
rect 21453 33643 21511 33649
rect 21453 33640 21465 33643
rect 21416 33612 21465 33640
rect 21416 33600 21422 33612
rect 21453 33609 21465 33612
rect 21499 33640 21511 33643
rect 22370 33640 22376 33652
rect 21499 33612 22376 33640
rect 21499 33609 21511 33612
rect 21453 33603 21511 33609
rect 22370 33600 22376 33612
rect 22428 33640 22434 33652
rect 23566 33640 23572 33652
rect 22428 33612 23572 33640
rect 22428 33600 22434 33612
rect 21376 33572 21404 33600
rect 22278 33572 22284 33584
rect 20930 33544 21404 33572
rect 22020 33544 22284 33572
rect 9401 33507 9459 33513
rect 9401 33473 9413 33507
rect 9447 33504 9459 33507
rect 10226 33504 10232 33516
rect 9447 33476 10232 33504
rect 9447 33473 9459 33476
rect 9401 33467 9459 33473
rect 10226 33464 10232 33476
rect 10284 33464 10290 33516
rect 19426 33464 19432 33516
rect 19484 33464 19490 33516
rect 22020 33513 22048 33544
rect 22278 33532 22284 33544
rect 22336 33532 22342 33584
rect 22664 33572 22692 33612
rect 23566 33600 23572 33612
rect 23624 33600 23630 33652
rect 24394 33600 24400 33652
rect 24452 33640 24458 33652
rect 24581 33643 24639 33649
rect 24581 33640 24593 33643
rect 24452 33612 24593 33640
rect 24452 33600 24458 33612
rect 24581 33609 24593 33612
rect 24627 33609 24639 33643
rect 24581 33603 24639 33609
rect 24673 33643 24731 33649
rect 24673 33609 24685 33643
rect 24719 33640 24731 33643
rect 25222 33640 25228 33652
rect 24719 33612 25228 33640
rect 24719 33609 24731 33612
rect 24673 33603 24731 33609
rect 25222 33600 25228 33612
rect 25280 33600 25286 33652
rect 23584 33572 23612 33600
rect 25317 33575 25375 33581
rect 25317 33572 25329 33575
rect 22664 33544 22770 33572
rect 23584 33544 25329 33572
rect 25317 33541 25329 33544
rect 25363 33541 25375 33575
rect 25317 33535 25375 33541
rect 22005 33507 22063 33513
rect 22005 33473 22017 33507
rect 22051 33473 22063 33507
rect 22005 33467 22063 33473
rect 19705 33439 19763 33445
rect 19705 33405 19717 33439
rect 19751 33436 19763 33439
rect 21542 33436 21548 33448
rect 19751 33408 21548 33436
rect 19751 33405 19763 33408
rect 19705 33399 19763 33405
rect 21542 33396 21548 33408
rect 21600 33396 21606 33448
rect 22281 33439 22339 33445
rect 22281 33405 22293 33439
rect 22327 33436 22339 33439
rect 23750 33436 23756 33448
rect 22327 33408 23756 33436
rect 22327 33405 22339 33408
rect 22281 33399 22339 33405
rect 23750 33396 23756 33408
rect 23808 33396 23814 33448
rect 24762 33396 24768 33448
rect 24820 33396 24826 33448
rect 23474 33260 23480 33312
rect 23532 33300 23538 33312
rect 23753 33303 23811 33309
rect 23753 33300 23765 33303
rect 23532 33272 23765 33300
rect 23532 33260 23538 33272
rect 23753 33269 23765 33272
rect 23799 33269 23811 33303
rect 23753 33263 23811 33269
rect 24213 33303 24271 33309
rect 24213 33269 24225 33303
rect 24259 33300 24271 33303
rect 24946 33300 24952 33312
rect 24259 33272 24952 33300
rect 24259 33269 24271 33272
rect 24213 33263 24271 33269
rect 24946 33260 24952 33272
rect 25004 33260 25010 33312
rect 1104 33210 25852 33232
rect 1104 33158 2950 33210
rect 3002 33158 3014 33210
rect 3066 33158 3078 33210
rect 3130 33158 3142 33210
rect 3194 33158 3206 33210
rect 3258 33158 12950 33210
rect 13002 33158 13014 33210
rect 13066 33158 13078 33210
rect 13130 33158 13142 33210
rect 13194 33158 13206 33210
rect 13258 33158 22950 33210
rect 23002 33158 23014 33210
rect 23066 33158 23078 33210
rect 23130 33158 23142 33210
rect 23194 33158 23206 33210
rect 23258 33158 25852 33210
rect 1104 33136 25852 33158
rect 9125 33099 9183 33105
rect 9125 33065 9137 33099
rect 9171 33096 9183 33099
rect 10410 33096 10416 33108
rect 9171 33068 10416 33096
rect 9171 33065 9183 33068
rect 9125 33059 9183 33065
rect 10410 33056 10416 33068
rect 10468 33056 10474 33108
rect 21358 33056 21364 33108
rect 21416 33096 21422 33108
rect 21453 33099 21511 33105
rect 21453 33096 21465 33099
rect 21416 33068 21465 33096
rect 21416 33056 21422 33068
rect 21453 33065 21465 33068
rect 21499 33065 21511 33099
rect 21453 33059 21511 33065
rect 23290 33056 23296 33108
rect 23348 33096 23354 33108
rect 24029 33099 24087 33105
rect 24029 33096 24041 33099
rect 23348 33068 24041 33096
rect 23348 33056 23354 33068
rect 24029 33065 24041 33068
rect 24075 33065 24087 33099
rect 24029 33059 24087 33065
rect 19705 32963 19763 32969
rect 19705 32929 19717 32963
rect 19751 32960 19763 32963
rect 20254 32960 20260 32972
rect 19751 32932 20260 32960
rect 19751 32929 19763 32932
rect 19705 32923 19763 32929
rect 20254 32920 20260 32932
rect 20312 32920 20318 32972
rect 22278 32920 22284 32972
rect 22336 32920 22342 32972
rect 25038 32920 25044 32972
rect 25096 32920 25102 32972
rect 25133 32963 25191 32969
rect 25133 32929 25145 32963
rect 25179 32929 25191 32963
rect 25133 32923 25191 32929
rect 9306 32852 9312 32904
rect 9364 32852 9370 32904
rect 18141 32895 18199 32901
rect 18141 32861 18153 32895
rect 18187 32892 18199 32895
rect 18598 32892 18604 32904
rect 18187 32864 18604 32892
rect 18187 32861 18199 32864
rect 18141 32855 18199 32861
rect 18598 32852 18604 32864
rect 18656 32852 18662 32904
rect 19426 32852 19432 32904
rect 19484 32852 19490 32904
rect 23934 32852 23940 32904
rect 23992 32892 23998 32904
rect 25148 32892 25176 32923
rect 26050 32920 26056 32972
rect 26108 32960 26114 32972
rect 26234 32960 26240 32972
rect 26108 32932 26240 32960
rect 26108 32920 26114 32932
rect 26234 32920 26240 32932
rect 26292 32920 26298 32972
rect 23992 32864 25176 32892
rect 23992 32852 23998 32864
rect 21358 32824 21364 32836
rect 20930 32796 21364 32824
rect 21358 32784 21364 32796
rect 21416 32784 21422 32836
rect 22554 32784 22560 32836
rect 22612 32784 22618 32836
rect 23566 32784 23572 32836
rect 23624 32784 23630 32836
rect 24949 32827 25007 32833
rect 24949 32793 24961 32827
rect 24995 32824 25007 32827
rect 25314 32824 25320 32836
rect 24995 32796 25320 32824
rect 24995 32793 25007 32796
rect 24949 32787 25007 32793
rect 25314 32784 25320 32796
rect 25372 32824 25378 32836
rect 26050 32824 26056 32836
rect 25372 32796 26056 32824
rect 25372 32784 25378 32796
rect 26050 32784 26056 32796
rect 26108 32784 26114 32836
rect 17678 32716 17684 32768
rect 17736 32756 17742 32768
rect 18785 32759 18843 32765
rect 18785 32756 18797 32759
rect 17736 32728 18797 32756
rect 17736 32716 17742 32728
rect 18785 32725 18797 32728
rect 18831 32725 18843 32759
rect 18785 32719 18843 32725
rect 19518 32716 19524 32768
rect 19576 32756 19582 32768
rect 21177 32759 21235 32765
rect 21177 32756 21189 32759
rect 19576 32728 21189 32756
rect 19576 32716 19582 32728
rect 21177 32725 21189 32728
rect 21223 32725 21235 32759
rect 21177 32719 21235 32725
rect 24026 32716 24032 32768
rect 24084 32756 24090 32768
rect 24581 32759 24639 32765
rect 24581 32756 24593 32759
rect 24084 32728 24593 32756
rect 24084 32716 24090 32728
rect 24581 32725 24593 32728
rect 24627 32725 24639 32759
rect 24581 32719 24639 32725
rect 1104 32666 25852 32688
rect 1104 32614 7950 32666
rect 8002 32614 8014 32666
rect 8066 32614 8078 32666
rect 8130 32614 8142 32666
rect 8194 32614 8206 32666
rect 8258 32614 17950 32666
rect 18002 32614 18014 32666
rect 18066 32614 18078 32666
rect 18130 32614 18142 32666
rect 18194 32614 18206 32666
rect 18258 32614 25852 32666
rect 1104 32592 25852 32614
rect 8938 32512 8944 32564
rect 8996 32512 9002 32564
rect 16025 32555 16083 32561
rect 16025 32521 16037 32555
rect 16071 32552 16083 32555
rect 16945 32555 17003 32561
rect 16945 32552 16957 32555
rect 16071 32524 16957 32552
rect 16071 32521 16083 32524
rect 16025 32515 16083 32521
rect 16945 32521 16957 32524
rect 16991 32552 17003 32555
rect 17034 32552 17040 32564
rect 16991 32524 17040 32552
rect 16991 32521 17003 32524
rect 16945 32515 17003 32521
rect 17034 32512 17040 32524
rect 17092 32512 17098 32564
rect 17126 32512 17132 32564
rect 17184 32512 17190 32564
rect 18414 32512 18420 32564
rect 18472 32552 18478 32564
rect 18472 32524 18828 32552
rect 18472 32512 18478 32524
rect 15933 32487 15991 32493
rect 15933 32453 15945 32487
rect 15979 32484 15991 32487
rect 17144 32484 17172 32512
rect 15979 32456 17172 32484
rect 15979 32453 15991 32456
rect 15933 32447 15991 32453
rect 17678 32444 17684 32496
rect 17736 32444 17742 32496
rect 8662 32376 8668 32428
rect 8720 32416 8726 32428
rect 9125 32419 9183 32425
rect 9125 32416 9137 32419
rect 8720 32388 9137 32416
rect 8720 32376 8726 32388
rect 9125 32385 9137 32388
rect 9171 32385 9183 32419
rect 9125 32379 9183 32385
rect 16850 32376 16856 32428
rect 16908 32416 16914 32428
rect 17402 32416 17408 32428
rect 16908 32388 17408 32416
rect 16908 32376 16914 32388
rect 17402 32376 17408 32388
rect 17460 32376 17466 32428
rect 18800 32416 18828 32524
rect 18966 32512 18972 32564
rect 19024 32552 19030 32564
rect 19024 32524 20944 32552
rect 19024 32512 19030 32524
rect 19426 32444 19432 32496
rect 19484 32484 19490 32496
rect 20809 32487 20867 32493
rect 20809 32484 20821 32487
rect 19484 32456 20821 32484
rect 19484 32444 19490 32456
rect 20809 32453 20821 32456
rect 20855 32453 20867 32487
rect 20916 32484 20944 32524
rect 21082 32512 21088 32564
rect 21140 32552 21146 32564
rect 26510 32552 26516 32564
rect 21140 32524 26516 32552
rect 21140 32512 21146 32524
rect 26510 32512 26516 32524
rect 26568 32512 26574 32564
rect 20916 32456 22232 32484
rect 20809 32447 20867 32453
rect 19797 32419 19855 32425
rect 18800 32402 19104 32416
rect 18814 32388 19104 32402
rect 16209 32351 16267 32357
rect 16209 32317 16221 32351
rect 16255 32348 16267 32351
rect 16666 32348 16672 32360
rect 16255 32320 16672 32348
rect 16255 32317 16267 32320
rect 16209 32311 16267 32317
rect 16666 32308 16672 32320
rect 16724 32308 16730 32360
rect 16761 32351 16819 32357
rect 16761 32317 16773 32351
rect 16807 32348 16819 32351
rect 17310 32348 17316 32360
rect 16807 32320 17316 32348
rect 16807 32317 16819 32320
rect 16761 32311 16819 32317
rect 17310 32308 17316 32320
rect 17368 32348 17374 32360
rect 18966 32348 18972 32360
rect 17368 32320 18972 32348
rect 17368 32308 17374 32320
rect 18966 32308 18972 32320
rect 19024 32308 19030 32360
rect 19076 32348 19104 32388
rect 19797 32385 19809 32419
rect 19843 32416 19855 32419
rect 20073 32419 20131 32425
rect 20073 32416 20085 32419
rect 19843 32388 20085 32416
rect 19843 32385 19855 32388
rect 19797 32379 19855 32385
rect 20073 32385 20085 32388
rect 20119 32416 20131 32419
rect 21545 32419 21603 32425
rect 21545 32416 21557 32419
rect 20119 32388 21557 32416
rect 20119 32385 20131 32388
rect 20073 32379 20131 32385
rect 21545 32385 21557 32388
rect 21591 32385 21603 32419
rect 21545 32379 21603 32385
rect 19521 32351 19579 32357
rect 19521 32348 19533 32351
rect 19076 32320 19533 32348
rect 19521 32317 19533 32320
rect 19567 32348 19579 32351
rect 21358 32348 21364 32360
rect 19567 32320 21364 32348
rect 19567 32317 19579 32320
rect 19521 32311 19579 32317
rect 21358 32308 21364 32320
rect 21416 32308 21422 32360
rect 21082 32280 21088 32292
rect 18708 32252 21088 32280
rect 13446 32172 13452 32224
rect 13504 32212 13510 32224
rect 15565 32215 15623 32221
rect 15565 32212 15577 32215
rect 13504 32184 15577 32212
rect 13504 32172 13510 32184
rect 15565 32181 15577 32184
rect 15611 32181 15623 32215
rect 15565 32175 15623 32181
rect 17862 32172 17868 32224
rect 17920 32212 17926 32224
rect 18708 32212 18736 32252
rect 21082 32240 21088 32252
rect 21140 32240 21146 32292
rect 17920 32184 18736 32212
rect 19153 32215 19211 32221
rect 17920 32172 17926 32184
rect 19153 32181 19165 32215
rect 19199 32212 19211 32215
rect 19334 32212 19340 32224
rect 19199 32184 19340 32212
rect 19199 32181 19211 32184
rect 19153 32175 19211 32181
rect 19334 32172 19340 32184
rect 19392 32172 19398 32224
rect 21560 32212 21588 32379
rect 22094 32376 22100 32428
rect 22152 32376 22158 32428
rect 22094 32212 22100 32224
rect 21560 32184 22100 32212
rect 22094 32172 22100 32184
rect 22152 32172 22158 32224
rect 22204 32212 22232 32456
rect 22278 32444 22284 32496
rect 22336 32484 22342 32496
rect 22833 32487 22891 32493
rect 22833 32484 22845 32487
rect 22336 32456 22845 32484
rect 22336 32444 22342 32456
rect 22833 32453 22845 32456
rect 22879 32484 22891 32487
rect 22879 32456 23520 32484
rect 22879 32453 22891 32456
rect 22833 32447 22891 32453
rect 23492 32425 23520 32456
rect 23750 32444 23756 32496
rect 23808 32484 23814 32496
rect 23808 32456 24242 32484
rect 23808 32444 23814 32456
rect 23477 32419 23535 32425
rect 23477 32385 23489 32419
rect 23523 32385 23535 32419
rect 23477 32379 23535 32385
rect 23753 32351 23811 32357
rect 23753 32317 23765 32351
rect 23799 32348 23811 32351
rect 25314 32348 25320 32360
rect 23799 32320 25320 32348
rect 23799 32317 23811 32320
rect 23753 32311 23811 32317
rect 25314 32308 25320 32320
rect 25372 32308 25378 32360
rect 24854 32212 24860 32224
rect 22204 32184 24860 32212
rect 24854 32172 24860 32184
rect 24912 32172 24918 32224
rect 25222 32172 25228 32224
rect 25280 32172 25286 32224
rect 1104 32122 25852 32144
rect 1104 32070 2950 32122
rect 3002 32070 3014 32122
rect 3066 32070 3078 32122
rect 3130 32070 3142 32122
rect 3194 32070 3206 32122
rect 3258 32070 12950 32122
rect 13002 32070 13014 32122
rect 13066 32070 13078 32122
rect 13130 32070 13142 32122
rect 13194 32070 13206 32122
rect 13258 32070 22950 32122
rect 23002 32070 23014 32122
rect 23066 32070 23078 32122
rect 23130 32070 23142 32122
rect 23194 32070 23206 32122
rect 23258 32070 25852 32122
rect 1104 32048 25852 32070
rect 17862 32008 17868 32020
rect 16132 31980 17868 32008
rect 13354 31900 13360 31952
rect 13412 31940 13418 31952
rect 15657 31943 15715 31949
rect 15657 31940 15669 31943
rect 13412 31912 15669 31940
rect 13412 31900 13418 31912
rect 15657 31909 15669 31912
rect 15703 31909 15715 31943
rect 15657 31903 15715 31909
rect 16132 31881 16160 31980
rect 17862 31968 17868 31980
rect 17920 31968 17926 32020
rect 18598 31968 18604 32020
rect 18656 31968 18662 32020
rect 19334 31968 19340 32020
rect 19392 32008 19398 32020
rect 19392 31980 22094 32008
rect 19392 31968 19398 31980
rect 21174 31900 21180 31952
rect 21232 31940 21238 31952
rect 22066 31940 22094 31980
rect 22554 31968 22560 32020
rect 22612 32008 22618 32020
rect 25225 32011 25283 32017
rect 25225 32008 25237 32011
rect 22612 31980 25237 32008
rect 22612 31968 22618 31980
rect 25225 31977 25237 31980
rect 25271 31977 25283 32011
rect 25225 31971 25283 31977
rect 21232 31912 21680 31940
rect 22066 31912 22232 31940
rect 21232 31900 21238 31912
rect 16117 31875 16175 31881
rect 16117 31841 16129 31875
rect 16163 31841 16175 31875
rect 16117 31835 16175 31841
rect 16301 31875 16359 31881
rect 16301 31841 16313 31875
rect 16347 31872 16359 31875
rect 16666 31872 16672 31884
rect 16347 31844 16672 31872
rect 16347 31841 16359 31844
rect 16301 31835 16359 31841
rect 16666 31832 16672 31844
rect 16724 31832 16730 31884
rect 16850 31832 16856 31884
rect 16908 31832 16914 31884
rect 19426 31832 19432 31884
rect 19484 31832 19490 31884
rect 19705 31875 19763 31881
rect 19705 31841 19717 31875
rect 19751 31872 19763 31875
rect 20070 31872 20076 31884
rect 19751 31844 20076 31872
rect 19751 31841 19763 31844
rect 19705 31835 19763 31841
rect 20070 31832 20076 31844
rect 20128 31832 20134 31884
rect 11514 31764 11520 31816
rect 11572 31804 11578 31816
rect 15013 31807 15071 31813
rect 15013 31804 15025 31807
rect 11572 31776 15025 31804
rect 11572 31764 11578 31776
rect 15013 31773 15025 31776
rect 15059 31773 15071 31807
rect 21652 31804 21680 31912
rect 22002 31832 22008 31884
rect 22060 31872 22066 31884
rect 22204 31881 22232 31912
rect 22097 31875 22155 31881
rect 22097 31872 22109 31875
rect 22060 31844 22109 31872
rect 22060 31832 22066 31844
rect 22097 31841 22109 31844
rect 22143 31841 22155 31875
rect 22097 31835 22155 31841
rect 22189 31875 22247 31881
rect 22189 31841 22201 31875
rect 22235 31841 22247 31875
rect 22189 31835 22247 31841
rect 22833 31807 22891 31813
rect 22833 31804 22845 31807
rect 21652 31776 22845 31804
rect 15013 31767 15071 31773
rect 22833 31773 22845 31776
rect 22879 31773 22891 31807
rect 22833 31767 22891 31773
rect 23290 31764 23296 31816
rect 23348 31804 23354 31816
rect 23477 31807 23535 31813
rect 23477 31804 23489 31807
rect 23348 31776 23489 31804
rect 23348 31764 23354 31776
rect 23477 31773 23489 31776
rect 23523 31773 23535 31807
rect 23477 31767 23535 31773
rect 24581 31807 24639 31813
rect 24581 31773 24593 31807
rect 24627 31804 24639 31807
rect 25222 31804 25228 31816
rect 24627 31776 25228 31804
rect 24627 31773 24639 31776
rect 24581 31767 24639 31773
rect 25222 31764 25228 31776
rect 25280 31764 25286 31816
rect 14274 31696 14280 31748
rect 14332 31696 14338 31748
rect 17126 31696 17132 31748
rect 17184 31696 17190 31748
rect 18414 31736 18420 31748
rect 18354 31708 18420 31736
rect 18414 31696 18420 31708
rect 18472 31736 18478 31748
rect 18874 31736 18880 31748
rect 18472 31708 18880 31736
rect 18472 31696 18478 31708
rect 18874 31696 18880 31708
rect 18932 31736 18938 31748
rect 18969 31739 19027 31745
rect 18969 31736 18981 31739
rect 18932 31708 18981 31736
rect 18932 31696 18938 31708
rect 18969 31705 18981 31708
rect 19015 31736 19027 31739
rect 19015 31708 20194 31736
rect 19015 31705 19027 31708
rect 18969 31699 19027 31705
rect 16025 31671 16083 31677
rect 16025 31637 16037 31671
rect 16071 31668 16083 31671
rect 16666 31668 16672 31680
rect 16071 31640 16672 31668
rect 16071 31637 16083 31640
rect 16025 31631 16083 31637
rect 16666 31628 16672 31640
rect 16724 31668 16730 31680
rect 17310 31668 17316 31680
rect 16724 31640 17316 31668
rect 16724 31628 16730 31640
rect 17310 31628 17316 31640
rect 17368 31628 17374 31680
rect 20070 31628 20076 31680
rect 20128 31668 20134 31680
rect 21174 31668 21180 31680
rect 20128 31640 21180 31668
rect 20128 31628 20134 31640
rect 21174 31628 21180 31640
rect 21232 31628 21238 31680
rect 21266 31628 21272 31680
rect 21324 31668 21330 31680
rect 21637 31671 21695 31677
rect 21637 31668 21649 31671
rect 21324 31640 21649 31668
rect 21324 31628 21330 31640
rect 21637 31637 21649 31640
rect 21683 31637 21695 31671
rect 21637 31631 21695 31637
rect 22002 31628 22008 31680
rect 22060 31628 22066 31680
rect 23842 31628 23848 31680
rect 23900 31668 23906 31680
rect 24121 31671 24179 31677
rect 24121 31668 24133 31671
rect 23900 31640 24133 31668
rect 23900 31628 23906 31640
rect 24121 31637 24133 31640
rect 24167 31637 24179 31671
rect 24121 31631 24179 31637
rect 1104 31578 25852 31600
rect 1104 31526 7950 31578
rect 8002 31526 8014 31578
rect 8066 31526 8078 31578
rect 8130 31526 8142 31578
rect 8194 31526 8206 31578
rect 8258 31526 17950 31578
rect 18002 31526 18014 31578
rect 18066 31526 18078 31578
rect 18130 31526 18142 31578
rect 18194 31526 18206 31578
rect 18258 31526 25852 31578
rect 1104 31504 25852 31526
rect 16850 31464 16856 31476
rect 13280 31436 16856 31464
rect 13280 31337 13308 31436
rect 16850 31424 16856 31436
rect 16908 31424 16914 31476
rect 17126 31424 17132 31476
rect 17184 31464 17190 31476
rect 17681 31467 17739 31473
rect 17681 31464 17693 31467
rect 17184 31436 17693 31464
rect 17184 31424 17190 31436
rect 17681 31433 17693 31436
rect 17727 31433 17739 31467
rect 17681 31427 17739 31433
rect 20530 31424 20536 31476
rect 20588 31464 20594 31476
rect 20625 31467 20683 31473
rect 20625 31464 20637 31467
rect 20588 31436 20637 31464
rect 20588 31424 20594 31436
rect 20625 31433 20637 31436
rect 20671 31433 20683 31467
rect 20625 31427 20683 31433
rect 21545 31467 21603 31473
rect 21545 31433 21557 31467
rect 21591 31464 21603 31467
rect 22002 31464 22008 31476
rect 21591 31436 22008 31464
rect 21591 31433 21603 31436
rect 21545 31427 21603 31433
rect 22002 31424 22008 31436
rect 22060 31464 22066 31476
rect 22278 31464 22284 31476
rect 22060 31436 22284 31464
rect 22060 31424 22066 31436
rect 22278 31424 22284 31436
rect 22336 31424 22342 31476
rect 23124 31436 23888 31464
rect 15470 31396 15476 31408
rect 14766 31368 15476 31396
rect 15470 31356 15476 31368
rect 15528 31356 15534 31408
rect 21358 31356 21364 31408
rect 21416 31396 21422 31408
rect 21726 31396 21732 31408
rect 21416 31368 21732 31396
rect 21416 31356 21422 31368
rect 21726 31356 21732 31368
rect 21784 31396 21790 31408
rect 23124 31396 23152 31436
rect 21784 31368 23152 31396
rect 21784 31356 21790 31368
rect 13265 31331 13323 31337
rect 13265 31297 13277 31331
rect 13311 31297 13323 31331
rect 13265 31291 13323 31297
rect 17037 31331 17095 31337
rect 17037 31297 17049 31331
rect 17083 31297 17095 31331
rect 17037 31291 17095 31297
rect 19061 31331 19119 31337
rect 19061 31297 19073 31331
rect 19107 31328 19119 31331
rect 19518 31328 19524 31340
rect 19107 31300 19524 31328
rect 19107 31297 19119 31300
rect 19061 31291 19119 31297
rect 13541 31263 13599 31269
rect 13541 31229 13553 31263
rect 13587 31260 13599 31263
rect 16758 31260 16764 31272
rect 13587 31232 16764 31260
rect 13587 31229 13599 31232
rect 13541 31223 13599 31229
rect 16758 31220 16764 31232
rect 16816 31220 16822 31272
rect 17052 31260 17080 31291
rect 19518 31288 19524 31300
rect 19576 31328 19582 31340
rect 19978 31328 19984 31340
rect 19576 31300 19984 31328
rect 19576 31288 19582 31300
rect 19978 31288 19984 31300
rect 20036 31288 20042 31340
rect 20346 31288 20352 31340
rect 20404 31328 20410 31340
rect 20533 31331 20591 31337
rect 20533 31328 20545 31331
rect 20404 31300 20545 31328
rect 20404 31288 20410 31300
rect 20533 31297 20545 31300
rect 20579 31328 20591 31331
rect 22186 31328 22192 31340
rect 20579 31300 22192 31328
rect 20579 31297 20591 31300
rect 20533 31291 20591 31297
rect 22186 31288 22192 31300
rect 22244 31328 22250 31340
rect 22370 31328 22376 31340
rect 22244 31300 22376 31328
rect 22244 31288 22250 31300
rect 22370 31288 22376 31300
rect 22428 31288 22434 31340
rect 23750 31288 23756 31340
rect 23808 31328 23814 31340
rect 23860 31328 23888 31436
rect 25314 31424 25320 31476
rect 25372 31424 25378 31476
rect 23808 31314 23888 31328
rect 24673 31331 24731 31337
rect 23808 31300 23874 31314
rect 23808 31288 23814 31300
rect 24673 31297 24685 31331
rect 24719 31328 24731 31331
rect 24762 31328 24768 31340
rect 24719 31300 24768 31328
rect 24719 31297 24731 31300
rect 24673 31291 24731 31297
rect 24762 31288 24768 31300
rect 24820 31288 24826 31340
rect 18690 31260 18696 31272
rect 17052 31232 18696 31260
rect 18690 31220 18696 31232
rect 18748 31260 18754 31272
rect 20717 31263 20775 31269
rect 20717 31260 20729 31263
rect 18748 31232 20729 31260
rect 18748 31220 18754 31232
rect 20717 31229 20729 31232
rect 20763 31229 20775 31263
rect 22465 31263 22523 31269
rect 22465 31260 22477 31263
rect 20717 31223 20775 31229
rect 22066 31232 22477 31260
rect 19426 31152 19432 31204
rect 19484 31192 19490 31204
rect 20165 31195 20223 31201
rect 20165 31192 20177 31195
rect 19484 31164 20177 31192
rect 19484 31152 19490 31164
rect 20165 31161 20177 31164
rect 20211 31161 20223 31195
rect 20165 31155 20223 31161
rect 20530 31152 20536 31204
rect 20588 31192 20594 31204
rect 22066 31192 22094 31232
rect 22465 31229 22477 31232
rect 22511 31229 22523 31263
rect 22465 31223 22523 31229
rect 22738 31220 22744 31272
rect 22796 31220 22802 31272
rect 20588 31164 22094 31192
rect 20588 31152 20594 31164
rect 13906 31084 13912 31136
rect 13964 31124 13970 31136
rect 15013 31127 15071 31133
rect 15013 31124 15025 31127
rect 13964 31096 15025 31124
rect 13964 31084 13970 31096
rect 15013 31093 15025 31096
rect 15059 31093 15071 31127
rect 15013 31087 15071 31093
rect 15470 31084 15476 31136
rect 15528 31084 15534 31136
rect 15657 31127 15715 31133
rect 15657 31093 15669 31127
rect 15703 31124 15715 31127
rect 16574 31124 16580 31136
rect 15703 31096 16580 31124
rect 15703 31093 15715 31096
rect 15657 31087 15715 31093
rect 16574 31084 16580 31096
rect 16632 31084 16638 31136
rect 16761 31127 16819 31133
rect 16761 31093 16773 31127
rect 16807 31124 16819 31127
rect 17678 31124 17684 31136
rect 16807 31096 17684 31124
rect 16807 31093 16819 31096
rect 16761 31087 16819 31093
rect 17678 31084 17684 31096
rect 17736 31084 17742 31136
rect 19705 31127 19763 31133
rect 19705 31093 19717 31127
rect 19751 31124 19763 31127
rect 20070 31124 20076 31136
rect 19751 31096 20076 31124
rect 19751 31093 19763 31096
rect 19705 31087 19763 31093
rect 20070 31084 20076 31096
rect 20128 31084 20134 31136
rect 23934 31084 23940 31136
rect 23992 31124 23998 31136
rect 24213 31127 24271 31133
rect 24213 31124 24225 31127
rect 23992 31096 24225 31124
rect 23992 31084 23998 31096
rect 24213 31093 24225 31096
rect 24259 31093 24271 31127
rect 24213 31087 24271 31093
rect 1104 31034 25852 31056
rect 1104 30982 2950 31034
rect 3002 30982 3014 31034
rect 3066 30982 3078 31034
rect 3130 30982 3142 31034
rect 3194 30982 3206 31034
rect 3258 30982 12950 31034
rect 13002 30982 13014 31034
rect 13066 30982 13078 31034
rect 13130 30982 13142 31034
rect 13194 30982 13206 31034
rect 13258 30982 22950 31034
rect 23002 30982 23014 31034
rect 23066 30982 23078 31034
rect 23130 30982 23142 31034
rect 23194 30982 23206 31034
rect 23258 30982 25852 31034
rect 1104 30960 25852 30982
rect 18601 30923 18659 30929
rect 18601 30889 18613 30923
rect 18647 30920 18659 30923
rect 18690 30920 18696 30932
rect 18647 30892 18696 30920
rect 18647 30889 18659 30892
rect 18601 30883 18659 30889
rect 18690 30880 18696 30892
rect 18748 30880 18754 30932
rect 18874 30880 18880 30932
rect 18932 30880 18938 30932
rect 20346 30880 20352 30932
rect 20404 30880 20410 30932
rect 22738 30880 22744 30932
rect 22796 30920 22802 30932
rect 23569 30923 23627 30929
rect 23569 30920 23581 30923
rect 22796 30892 23581 30920
rect 22796 30880 22802 30892
rect 23569 30889 23581 30892
rect 23615 30889 23627 30923
rect 23569 30883 23627 30889
rect 16853 30787 16911 30793
rect 16853 30753 16865 30787
rect 16899 30784 16911 30787
rect 19334 30784 19340 30796
rect 16899 30756 19340 30784
rect 16899 30753 16911 30756
rect 16853 30747 16911 30753
rect 19334 30744 19340 30756
rect 19392 30784 19398 30796
rect 20530 30784 20536 30796
rect 19392 30756 20536 30784
rect 19392 30744 19398 30756
rect 20530 30744 20536 30756
rect 20588 30784 20594 30796
rect 20717 30787 20775 30793
rect 20717 30784 20729 30787
rect 20588 30756 20729 30784
rect 20588 30744 20594 30756
rect 20717 30753 20729 30756
rect 20763 30753 20775 30787
rect 20717 30747 20775 30753
rect 20993 30787 21051 30793
rect 20993 30753 21005 30787
rect 21039 30784 21051 30787
rect 23290 30784 23296 30796
rect 21039 30756 23296 30784
rect 21039 30753 21051 30756
rect 20993 30747 21051 30753
rect 23290 30744 23296 30756
rect 23348 30744 23354 30796
rect 14185 30719 14243 30725
rect 14185 30685 14197 30719
rect 14231 30716 14243 30719
rect 15470 30716 15476 30728
rect 14231 30688 15476 30716
rect 14231 30685 14243 30688
rect 14185 30679 14243 30685
rect 15470 30676 15476 30688
rect 15528 30676 15534 30728
rect 18874 30676 18880 30728
rect 18932 30716 18938 30728
rect 19429 30719 19487 30725
rect 19429 30716 19441 30719
rect 18932 30688 19441 30716
rect 18932 30676 18938 30688
rect 19429 30685 19441 30688
rect 19475 30685 19487 30719
rect 19429 30679 19487 30685
rect 22925 30719 22983 30725
rect 22925 30685 22937 30719
rect 22971 30716 22983 30719
rect 23842 30716 23848 30728
rect 22971 30688 23848 30716
rect 22971 30685 22983 30688
rect 22925 30679 22983 30685
rect 14274 30608 14280 30660
rect 14332 30648 14338 30660
rect 14461 30651 14519 30657
rect 14461 30648 14473 30651
rect 14332 30620 14473 30648
rect 14332 30608 14338 30620
rect 14461 30617 14473 30620
rect 14507 30617 14519 30651
rect 14461 30611 14519 30617
rect 14476 30580 14504 30611
rect 15102 30608 15108 30660
rect 15160 30648 15166 30660
rect 15197 30651 15255 30657
rect 15197 30648 15209 30651
rect 15160 30620 15209 30648
rect 15160 30608 15166 30620
rect 15197 30617 15209 30620
rect 15243 30617 15255 30651
rect 15197 30611 15255 30617
rect 17129 30651 17187 30657
rect 17129 30617 17141 30651
rect 17175 30648 17187 30651
rect 18414 30648 18420 30660
rect 17175 30620 17540 30648
rect 18354 30620 18420 30648
rect 17175 30617 17187 30620
rect 17129 30611 17187 30617
rect 15749 30583 15807 30589
rect 15749 30580 15761 30583
rect 14476 30552 15761 30580
rect 15749 30549 15761 30552
rect 15795 30580 15807 30583
rect 16574 30580 16580 30592
rect 15795 30552 16580 30580
rect 15795 30549 15807 30552
rect 15749 30543 15807 30549
rect 16574 30540 16580 30552
rect 16632 30580 16638 30592
rect 17310 30580 17316 30592
rect 16632 30552 17316 30580
rect 16632 30540 16638 30552
rect 17310 30540 17316 30552
rect 17368 30540 17374 30592
rect 17512 30580 17540 30620
rect 18414 30608 18420 30620
rect 18472 30608 18478 30660
rect 20073 30651 20131 30657
rect 20073 30648 20085 30651
rect 18524 30620 20085 30648
rect 18524 30580 18552 30620
rect 20073 30617 20085 30620
rect 20119 30617 20131 30651
rect 20073 30611 20131 30617
rect 21726 30608 21732 30660
rect 21784 30608 21790 30660
rect 17512 30552 18552 30580
rect 22465 30583 22523 30589
rect 22465 30549 22477 30583
rect 22511 30580 22523 30583
rect 22940 30580 22968 30679
rect 23842 30676 23848 30688
rect 23900 30676 23906 30728
rect 23934 30676 23940 30728
rect 23992 30716 23998 30728
rect 24581 30719 24639 30725
rect 24581 30716 24593 30719
rect 23992 30688 24593 30716
rect 23992 30676 23998 30688
rect 24581 30685 24593 30688
rect 24627 30685 24639 30719
rect 24581 30679 24639 30685
rect 23566 30608 23572 30660
rect 23624 30648 23630 30660
rect 25225 30651 25283 30657
rect 25225 30648 25237 30651
rect 23624 30620 25237 30648
rect 23624 30608 23630 30620
rect 25225 30617 25237 30620
rect 25271 30617 25283 30651
rect 25225 30611 25283 30617
rect 22511 30552 22968 30580
rect 22511 30549 22523 30552
rect 22465 30543 22523 30549
rect 23750 30540 23756 30592
rect 23808 30580 23814 30592
rect 23937 30583 23995 30589
rect 23937 30580 23949 30583
rect 23808 30552 23949 30580
rect 23808 30540 23814 30552
rect 23937 30549 23949 30552
rect 23983 30580 23995 30583
rect 24213 30583 24271 30589
rect 24213 30580 24225 30583
rect 23983 30552 24225 30580
rect 23983 30549 23995 30552
rect 23937 30543 23995 30549
rect 24213 30549 24225 30552
rect 24259 30580 24271 30583
rect 24578 30580 24584 30592
rect 24259 30552 24584 30580
rect 24259 30549 24271 30552
rect 24213 30543 24271 30549
rect 24578 30540 24584 30552
rect 24636 30540 24642 30592
rect 1104 30490 25852 30512
rect 1104 30438 7950 30490
rect 8002 30438 8014 30490
rect 8066 30438 8078 30490
rect 8130 30438 8142 30490
rect 8194 30438 8206 30490
rect 8258 30438 17950 30490
rect 18002 30438 18014 30490
rect 18066 30438 18078 30490
rect 18130 30438 18142 30490
rect 18194 30438 18206 30490
rect 18258 30438 25852 30490
rect 1104 30416 25852 30438
rect 20254 30336 20260 30388
rect 20312 30376 20318 30388
rect 21266 30376 21272 30388
rect 20312 30348 21272 30376
rect 20312 30336 20318 30348
rect 21266 30336 21272 30348
rect 21324 30336 21330 30388
rect 22370 30336 22376 30388
rect 22428 30376 22434 30388
rect 24486 30376 24492 30388
rect 22428 30348 24492 30376
rect 22428 30336 22434 30348
rect 24486 30336 24492 30348
rect 24544 30336 24550 30388
rect 24578 30336 24584 30388
rect 24636 30376 24642 30388
rect 24636 30348 24900 30376
rect 24636 30336 24642 30348
rect 11238 30268 11244 30320
rect 11296 30308 11302 30320
rect 20349 30311 20407 30317
rect 11296 30280 13018 30308
rect 14476 30280 16160 30308
rect 11296 30268 11302 30280
rect 10045 30243 10103 30249
rect 10045 30209 10057 30243
rect 10091 30240 10103 30243
rect 10318 30240 10324 30252
rect 10091 30212 10324 30240
rect 10091 30209 10103 30212
rect 10045 30203 10103 30209
rect 10318 30200 10324 30212
rect 10376 30200 10382 30252
rect 14366 30200 14372 30252
rect 14424 30240 14430 30252
rect 14476 30249 14504 30280
rect 14461 30243 14519 30249
rect 14461 30240 14473 30243
rect 14424 30212 14473 30240
rect 14424 30200 14430 30212
rect 14461 30209 14473 30212
rect 14507 30209 14519 30243
rect 14461 30203 14519 30209
rect 15838 30200 15844 30252
rect 15896 30240 15902 30252
rect 15933 30243 15991 30249
rect 15933 30240 15945 30243
rect 15896 30212 15945 30240
rect 15896 30200 15902 30212
rect 15933 30209 15945 30212
rect 15979 30209 15991 30243
rect 15933 30203 15991 30209
rect 10137 30175 10195 30181
rect 10137 30172 10149 30175
rect 10060 30144 10149 30172
rect 10060 30116 10088 30144
rect 10137 30141 10149 30144
rect 10183 30141 10195 30175
rect 10137 30135 10195 30141
rect 10226 30132 10232 30184
rect 10284 30132 10290 30184
rect 12253 30175 12311 30181
rect 12253 30141 12265 30175
rect 12299 30141 12311 30175
rect 12253 30135 12311 30141
rect 12529 30175 12587 30181
rect 12529 30141 12541 30175
rect 12575 30172 12587 30175
rect 15105 30175 15163 30181
rect 15105 30172 15117 30175
rect 12575 30144 15117 30172
rect 12575 30141 12587 30144
rect 12529 30135 12587 30141
rect 15105 30141 15117 30144
rect 15151 30141 15163 30175
rect 15105 30135 15163 30141
rect 9677 30107 9735 30113
rect 9677 30073 9689 30107
rect 9723 30104 9735 30107
rect 9766 30104 9772 30116
rect 9723 30076 9772 30104
rect 9723 30073 9735 30076
rect 9677 30067 9735 30073
rect 9766 30064 9772 30076
rect 9824 30064 9830 30116
rect 10042 30064 10048 30116
rect 10100 30064 10106 30116
rect 12268 30036 12296 30135
rect 15948 30104 15976 30203
rect 16132 30184 16160 30280
rect 20349 30277 20361 30311
rect 20395 30308 20407 30311
rect 20622 30308 20628 30320
rect 20395 30280 20628 30308
rect 20395 30277 20407 30280
rect 20349 30271 20407 30277
rect 20622 30268 20628 30280
rect 20680 30268 20686 30320
rect 22462 30268 22468 30320
rect 22520 30268 22526 30320
rect 23474 30308 23480 30320
rect 23032 30280 23480 30308
rect 17313 30243 17371 30249
rect 17313 30209 17325 30243
rect 17359 30240 17371 30243
rect 18782 30240 18788 30252
rect 17359 30212 18788 30240
rect 17359 30209 17371 30212
rect 17313 30203 17371 30209
rect 18782 30200 18788 30212
rect 18840 30200 18846 30252
rect 19245 30243 19303 30249
rect 19245 30209 19257 30243
rect 19291 30240 19303 30243
rect 20257 30243 20315 30249
rect 20257 30240 20269 30243
rect 19291 30212 20269 30240
rect 19291 30209 19303 30212
rect 19245 30203 19303 30209
rect 20257 30209 20269 30212
rect 20303 30209 20315 30243
rect 20257 30203 20315 30209
rect 21269 30243 21327 30249
rect 21269 30209 21281 30243
rect 21315 30240 21327 30243
rect 22373 30243 22431 30249
rect 22373 30240 22385 30243
rect 21315 30212 22385 30240
rect 21315 30209 21327 30212
rect 21269 30203 21327 30209
rect 22373 30209 22385 30212
rect 22419 30209 22431 30243
rect 22373 30203 22431 30209
rect 16022 30132 16028 30184
rect 16080 30132 16086 30184
rect 16114 30132 16120 30184
rect 16172 30132 16178 30184
rect 20438 30132 20444 30184
rect 20496 30132 20502 30184
rect 22649 30175 22707 30181
rect 22649 30141 22661 30175
rect 22695 30172 22707 30175
rect 23032 30172 23060 30280
rect 23474 30268 23480 30280
rect 23532 30268 23538 30320
rect 23566 30268 23572 30320
rect 23624 30268 23630 30320
rect 24872 30308 24900 30348
rect 25317 30311 25375 30317
rect 25317 30308 25329 30311
rect 24794 30280 25329 30308
rect 25317 30277 25329 30280
rect 25363 30277 25375 30311
rect 25317 30271 25375 30277
rect 22695 30144 23060 30172
rect 22695 30141 22707 30144
rect 22649 30135 22707 30141
rect 23290 30132 23296 30184
rect 23348 30132 23354 30184
rect 24762 30132 24768 30184
rect 24820 30172 24826 30184
rect 25041 30175 25099 30181
rect 25041 30172 25053 30175
rect 24820 30144 25053 30172
rect 24820 30132 24826 30144
rect 25041 30141 25053 30144
rect 25087 30141 25099 30175
rect 25041 30135 25099 30141
rect 16853 30107 16911 30113
rect 16853 30104 16865 30107
rect 15948 30076 16865 30104
rect 16853 30073 16865 30076
rect 16899 30104 16911 30107
rect 16942 30104 16948 30116
rect 16899 30076 16948 30104
rect 16899 30073 16911 30076
rect 16853 30067 16911 30073
rect 16942 30064 16948 30076
rect 17000 30064 17006 30116
rect 17052 30076 23428 30104
rect 12526 30036 12532 30048
rect 12268 30008 12532 30036
rect 12526 29996 12532 30008
rect 12584 29996 12590 30048
rect 13722 29996 13728 30048
rect 13780 30036 13786 30048
rect 14001 30039 14059 30045
rect 14001 30036 14013 30039
rect 13780 30008 14013 30036
rect 13780 29996 13786 30008
rect 14001 30005 14013 30008
rect 14047 30005 14059 30039
rect 14001 29999 14059 30005
rect 14550 29996 14556 30048
rect 14608 30036 14614 30048
rect 15565 30039 15623 30045
rect 15565 30036 15577 30039
rect 14608 30008 15577 30036
rect 14608 29996 14614 30008
rect 15565 30005 15577 30008
rect 15611 30005 15623 30039
rect 15565 29999 15623 30005
rect 16022 29996 16028 30048
rect 16080 30036 16086 30048
rect 16206 30036 16212 30048
rect 16080 30008 16212 30036
rect 16080 29996 16086 30008
rect 16206 29996 16212 30008
rect 16264 30036 16270 30048
rect 16761 30039 16819 30045
rect 16761 30036 16773 30039
rect 16264 30008 16773 30036
rect 16264 29996 16270 30008
rect 16761 30005 16773 30008
rect 16807 30036 16819 30039
rect 17052 30036 17080 30076
rect 16807 30008 17080 30036
rect 16807 30005 16819 30008
rect 16761 29999 16819 30005
rect 17402 29996 17408 30048
rect 17460 30036 17466 30048
rect 17957 30039 18015 30045
rect 17957 30036 17969 30039
rect 17460 30008 17969 30036
rect 17460 29996 17466 30008
rect 17957 30005 17969 30008
rect 18003 30005 18015 30039
rect 17957 29999 18015 30005
rect 19610 29996 19616 30048
rect 19668 30036 19674 30048
rect 19889 30039 19947 30045
rect 19889 30036 19901 30039
rect 19668 30008 19901 30036
rect 19668 29996 19674 30008
rect 19889 30005 19901 30008
rect 19935 30005 19947 30039
rect 19889 29999 19947 30005
rect 21450 29996 21456 30048
rect 21508 30036 21514 30048
rect 22005 30039 22063 30045
rect 22005 30036 22017 30039
rect 21508 30008 22017 30036
rect 21508 29996 21514 30008
rect 22005 30005 22017 30008
rect 22051 30005 22063 30039
rect 23400 30036 23428 30076
rect 26786 30036 26792 30048
rect 23400 30008 26792 30036
rect 22005 29999 22063 30005
rect 26786 29996 26792 30008
rect 26844 29996 26850 30048
rect 1104 29946 25852 29968
rect 1104 29894 2950 29946
rect 3002 29894 3014 29946
rect 3066 29894 3078 29946
rect 3130 29894 3142 29946
rect 3194 29894 3206 29946
rect 3258 29894 12950 29946
rect 13002 29894 13014 29946
rect 13066 29894 13078 29946
rect 13130 29894 13142 29946
rect 13194 29894 13206 29946
rect 13258 29894 22950 29946
rect 23002 29894 23014 29946
rect 23066 29894 23078 29946
rect 23130 29894 23142 29946
rect 23194 29894 23206 29946
rect 23258 29894 25852 29946
rect 1104 29872 25852 29894
rect 11238 29792 11244 29844
rect 11296 29792 11302 29844
rect 13265 29835 13323 29841
rect 13265 29801 13277 29835
rect 13311 29832 13323 29835
rect 14366 29832 14372 29844
rect 13311 29804 14372 29832
rect 13311 29801 13323 29804
rect 13265 29795 13323 29801
rect 14366 29792 14372 29804
rect 14424 29792 14430 29844
rect 16298 29792 16304 29844
rect 16356 29832 16362 29844
rect 19429 29835 19487 29841
rect 19429 29832 19441 29835
rect 16356 29804 19441 29832
rect 16356 29792 16362 29804
rect 19429 29801 19441 29804
rect 19475 29801 19487 29835
rect 22646 29832 22652 29844
rect 19429 29795 19487 29801
rect 19536 29804 22652 29832
rect 11514 29656 11520 29708
rect 11572 29656 11578 29708
rect 12526 29656 12532 29708
rect 12584 29696 12590 29708
rect 14277 29699 14335 29705
rect 14277 29696 14289 29699
rect 12584 29668 14289 29696
rect 12584 29656 12590 29668
rect 14277 29665 14289 29668
rect 14323 29696 14335 29699
rect 15102 29696 15108 29708
rect 14323 29668 15108 29696
rect 14323 29665 14335 29668
rect 14277 29659 14335 29665
rect 15102 29656 15108 29668
rect 15160 29696 15166 29708
rect 17129 29699 17187 29705
rect 17129 29696 17141 29699
rect 15160 29668 17141 29696
rect 15160 29656 15166 29668
rect 17129 29665 17141 29668
rect 17175 29665 17187 29699
rect 17129 29659 17187 29665
rect 17402 29656 17408 29708
rect 17460 29656 17466 29708
rect 19536 29696 19564 29804
rect 22646 29792 22652 29804
rect 22704 29792 22710 29844
rect 22830 29764 22836 29776
rect 21100 29736 22836 29764
rect 18708 29668 19564 29696
rect 9122 29588 9128 29640
rect 9180 29588 9186 29640
rect 9401 29563 9459 29569
rect 9401 29529 9413 29563
rect 9447 29529 9459 29563
rect 11238 29560 11244 29572
rect 10626 29532 11244 29560
rect 9401 29523 9459 29529
rect 9416 29492 9444 29523
rect 11238 29520 11244 29532
rect 11296 29520 11302 29572
rect 11790 29520 11796 29572
rect 11848 29520 11854 29572
rect 14553 29563 14611 29569
rect 11900 29532 12282 29560
rect 9582 29492 9588 29504
rect 9416 29464 9588 29492
rect 9582 29452 9588 29464
rect 9640 29452 9646 29504
rect 10226 29452 10232 29504
rect 10284 29492 10290 29504
rect 10873 29495 10931 29501
rect 10873 29492 10885 29495
rect 10284 29464 10885 29492
rect 10284 29452 10290 29464
rect 10873 29461 10885 29464
rect 10919 29461 10931 29495
rect 11256 29492 11284 29520
rect 11900 29492 11928 29532
rect 11256 29464 11928 29492
rect 12176 29492 12204 29532
rect 14553 29529 14565 29563
rect 14599 29560 14611 29563
rect 14826 29560 14832 29572
rect 14599 29532 14832 29560
rect 14599 29529 14611 29532
rect 14553 29523 14611 29529
rect 14826 29520 14832 29532
rect 14884 29520 14890 29572
rect 16393 29563 16451 29569
rect 16393 29560 16405 29563
rect 15778 29532 16405 29560
rect 13538 29492 13544 29504
rect 12176 29464 13544 29492
rect 10873 29455 10931 29461
rect 13538 29452 13544 29464
rect 13596 29452 13602 29504
rect 15194 29452 15200 29504
rect 15252 29492 15258 29504
rect 15470 29492 15476 29504
rect 15252 29464 15476 29492
rect 15252 29452 15258 29464
rect 15470 29452 15476 29464
rect 15528 29492 15534 29504
rect 15856 29492 15884 29532
rect 16393 29529 16405 29532
rect 16439 29560 16451 29563
rect 16439 29532 17894 29560
rect 16439 29529 16451 29532
rect 16393 29523 16451 29529
rect 18414 29520 18420 29572
rect 18472 29520 18478 29572
rect 15528 29464 15884 29492
rect 15528 29452 15534 29464
rect 16022 29452 16028 29504
rect 16080 29452 16086 29504
rect 16574 29452 16580 29504
rect 16632 29492 16638 29504
rect 16850 29492 16856 29504
rect 16632 29464 16856 29492
rect 16632 29452 16638 29464
rect 16850 29452 16856 29464
rect 16908 29492 16914 29504
rect 18708 29492 18736 29668
rect 19886 29656 19892 29708
rect 19944 29656 19950 29708
rect 19978 29656 19984 29708
rect 20036 29656 20042 29708
rect 21100 29705 21128 29736
rect 22830 29724 22836 29736
rect 22888 29724 22894 29776
rect 21085 29699 21143 29705
rect 21085 29665 21097 29699
rect 21131 29665 21143 29699
rect 21085 29659 21143 29665
rect 21177 29699 21235 29705
rect 21177 29665 21189 29699
rect 21223 29665 21235 29699
rect 21177 29659 21235 29665
rect 18782 29588 18788 29640
rect 18840 29628 18846 29640
rect 21192 29628 21220 29659
rect 22094 29656 22100 29708
rect 22152 29656 22158 29708
rect 24857 29699 24915 29705
rect 24857 29665 24869 29699
rect 24903 29665 24915 29699
rect 24857 29659 24915 29665
rect 18840 29600 21220 29628
rect 22281 29631 22339 29637
rect 18840 29588 18846 29600
rect 22281 29597 22293 29631
rect 22327 29628 22339 29631
rect 22462 29628 22468 29640
rect 22327 29600 22468 29628
rect 22327 29597 22339 29600
rect 22281 29591 22339 29597
rect 22462 29588 22468 29600
rect 22520 29628 22526 29640
rect 22741 29631 22799 29637
rect 22741 29628 22753 29631
rect 22520 29600 22753 29628
rect 22520 29588 22526 29600
rect 22741 29597 22753 29600
rect 22787 29597 22799 29631
rect 22741 29591 22799 29597
rect 24029 29631 24087 29637
rect 24029 29597 24041 29631
rect 24075 29597 24087 29631
rect 24872 29628 24900 29659
rect 25314 29628 25320 29640
rect 24872 29600 25320 29628
rect 24029 29591 24087 29597
rect 20438 29520 20444 29572
rect 20496 29560 20502 29572
rect 20993 29563 21051 29569
rect 20993 29560 21005 29563
rect 20496 29532 21005 29560
rect 20496 29520 20502 29532
rect 20993 29529 21005 29532
rect 21039 29529 21051 29563
rect 24044 29560 24072 29591
rect 25314 29588 25320 29600
rect 25372 29588 25378 29640
rect 24489 29563 24547 29569
rect 24489 29560 24501 29563
rect 24044 29532 24501 29560
rect 20993 29523 21051 29529
rect 24489 29529 24501 29532
rect 24535 29560 24547 29563
rect 24854 29560 24860 29572
rect 24535 29532 24860 29560
rect 24535 29529 24547 29532
rect 24489 29523 24547 29529
rect 24854 29520 24860 29532
rect 24912 29520 24918 29572
rect 16908 29464 18736 29492
rect 16908 29452 16914 29464
rect 18874 29452 18880 29504
rect 18932 29452 18938 29504
rect 19794 29452 19800 29504
rect 19852 29452 19858 29504
rect 19978 29452 19984 29504
rect 20036 29492 20042 29504
rect 20625 29495 20683 29501
rect 20625 29492 20637 29495
rect 20036 29464 20637 29492
rect 20036 29452 20042 29464
rect 20625 29461 20637 29464
rect 20671 29461 20683 29495
rect 20625 29455 20683 29461
rect 22554 29452 22560 29504
rect 22612 29452 22618 29504
rect 23201 29495 23259 29501
rect 23201 29461 23213 29495
rect 23247 29492 23259 29495
rect 23658 29492 23664 29504
rect 23247 29464 23664 29492
rect 23247 29461 23259 29464
rect 23201 29455 23259 29461
rect 23658 29452 23664 29464
rect 23716 29452 23722 29504
rect 23750 29452 23756 29504
rect 23808 29492 23814 29504
rect 23845 29495 23903 29501
rect 23845 29492 23857 29495
rect 23808 29464 23857 29492
rect 23808 29452 23814 29464
rect 23845 29461 23857 29464
rect 23891 29461 23903 29495
rect 23845 29455 23903 29461
rect 24578 29452 24584 29504
rect 24636 29452 24642 29504
rect 25038 29452 25044 29504
rect 25096 29492 25102 29504
rect 25133 29495 25191 29501
rect 25133 29492 25145 29495
rect 25096 29464 25145 29492
rect 25096 29452 25102 29464
rect 25133 29461 25145 29464
rect 25179 29461 25191 29495
rect 25133 29455 25191 29461
rect 1104 29402 25852 29424
rect 1104 29350 7950 29402
rect 8002 29350 8014 29402
rect 8066 29350 8078 29402
rect 8130 29350 8142 29402
rect 8194 29350 8206 29402
rect 8258 29350 17950 29402
rect 18002 29350 18014 29402
rect 18066 29350 18078 29402
rect 18130 29350 18142 29402
rect 18194 29350 18206 29402
rect 18258 29350 25852 29402
rect 1104 29328 25852 29350
rect 13354 29248 13360 29300
rect 13412 29248 13418 29300
rect 13446 29248 13452 29300
rect 13504 29248 13510 29300
rect 14550 29248 14556 29300
rect 14608 29248 14614 29300
rect 14645 29291 14703 29297
rect 14645 29257 14657 29291
rect 14691 29288 14703 29291
rect 15381 29291 15439 29297
rect 15381 29288 15393 29291
rect 14691 29260 15393 29288
rect 14691 29257 14703 29260
rect 14645 29251 14703 29257
rect 15381 29257 15393 29260
rect 15427 29257 15439 29291
rect 15381 29251 15439 29257
rect 15841 29291 15899 29297
rect 15841 29257 15853 29291
rect 15887 29288 15899 29291
rect 16482 29288 16488 29300
rect 15887 29260 16488 29288
rect 15887 29257 15899 29260
rect 15841 29251 15899 29257
rect 16482 29248 16488 29260
rect 16540 29248 16546 29300
rect 16574 29248 16580 29300
rect 16632 29288 16638 29300
rect 16853 29291 16911 29297
rect 16853 29288 16865 29291
rect 16632 29260 16865 29288
rect 16632 29248 16638 29260
rect 16853 29257 16865 29260
rect 16899 29257 16911 29291
rect 16853 29251 16911 29257
rect 17034 29248 17040 29300
rect 17092 29288 17098 29300
rect 17957 29291 18015 29297
rect 17957 29288 17969 29291
rect 17092 29260 17969 29288
rect 17092 29248 17098 29260
rect 17957 29257 17969 29260
rect 18003 29257 18015 29291
rect 17957 29251 18015 29257
rect 18414 29248 18420 29300
rect 18472 29288 18478 29300
rect 18693 29291 18751 29297
rect 18693 29288 18705 29291
rect 18472 29260 18705 29288
rect 18472 29248 18478 29260
rect 18693 29257 18705 29260
rect 18739 29288 18751 29291
rect 18877 29291 18935 29297
rect 18877 29288 18889 29291
rect 18739 29260 18889 29288
rect 18739 29257 18751 29260
rect 18693 29251 18751 29257
rect 18877 29257 18889 29260
rect 18923 29257 18935 29291
rect 18877 29251 18935 29257
rect 19245 29291 19303 29297
rect 19245 29257 19257 29291
rect 19291 29288 19303 29291
rect 19794 29288 19800 29300
rect 19291 29260 19800 29288
rect 19291 29257 19303 29260
rect 19245 29251 19303 29257
rect 19794 29248 19800 29260
rect 19852 29248 19858 29300
rect 23106 29248 23112 29300
rect 23164 29248 23170 29300
rect 23569 29291 23627 29297
rect 23569 29257 23581 29291
rect 23615 29288 23627 29291
rect 24857 29291 24915 29297
rect 24857 29288 24869 29291
rect 23615 29260 24869 29288
rect 23615 29257 23627 29260
rect 23569 29251 23627 29257
rect 24857 29257 24869 29260
rect 24903 29288 24915 29291
rect 25958 29288 25964 29300
rect 24903 29260 25964 29288
rect 24903 29257 24915 29260
rect 24857 29251 24915 29257
rect 25958 29248 25964 29260
rect 26016 29248 26022 29300
rect 14918 29180 14924 29232
rect 14976 29220 14982 29232
rect 20438 29220 20444 29232
rect 14976 29192 20444 29220
rect 14976 29180 14982 29192
rect 20438 29180 20444 29192
rect 20496 29220 20502 29232
rect 21545 29223 21603 29229
rect 21545 29220 21557 29223
rect 20496 29192 21557 29220
rect 20496 29180 20502 29192
rect 21545 29189 21557 29192
rect 21591 29220 21603 29223
rect 23477 29223 23535 29229
rect 23477 29220 23489 29223
rect 21591 29192 23489 29220
rect 21591 29189 21603 29192
rect 21545 29183 21603 29189
rect 23477 29189 23489 29192
rect 23523 29220 23535 29223
rect 24394 29220 24400 29232
rect 23523 29192 24400 29220
rect 23523 29189 23535 29192
rect 23477 29183 23535 29189
rect 24394 29180 24400 29192
rect 24452 29180 24458 29232
rect 10505 29155 10563 29161
rect 10505 29121 10517 29155
rect 10551 29152 10563 29155
rect 10778 29152 10784 29164
rect 10551 29124 10784 29152
rect 10551 29121 10563 29124
rect 10505 29115 10563 29121
rect 10778 29112 10784 29124
rect 10836 29152 10842 29164
rect 11517 29155 11575 29161
rect 11517 29152 11529 29155
rect 10836 29124 11529 29152
rect 10836 29112 10842 29124
rect 11517 29121 11529 29124
rect 11563 29121 11575 29155
rect 11517 29115 11575 29121
rect 11885 29155 11943 29161
rect 11885 29121 11897 29155
rect 11931 29152 11943 29155
rect 12618 29152 12624 29164
rect 11931 29124 12624 29152
rect 11931 29121 11943 29124
rect 11885 29115 11943 29121
rect 11532 29084 11560 29115
rect 12618 29112 12624 29124
rect 12676 29152 12682 29164
rect 13722 29152 13728 29164
rect 12676 29124 13728 29152
rect 12676 29112 12682 29124
rect 13722 29112 13728 29124
rect 13780 29152 13786 29164
rect 13780 29124 14780 29152
rect 13780 29112 13786 29124
rect 13541 29087 13599 29093
rect 13541 29084 13553 29087
rect 11532 29056 13553 29084
rect 13541 29053 13553 29056
rect 13587 29084 13599 29087
rect 13906 29084 13912 29096
rect 13587 29056 13912 29084
rect 13587 29053 13599 29056
rect 13541 29047 13599 29053
rect 13906 29044 13912 29056
rect 13964 29044 13970 29096
rect 14752 29093 14780 29124
rect 15378 29112 15384 29164
rect 15436 29152 15442 29164
rect 15746 29152 15752 29164
rect 15436 29124 15752 29152
rect 15436 29112 15442 29124
rect 15746 29112 15752 29124
rect 15804 29152 15810 29164
rect 16393 29155 16451 29161
rect 16393 29152 16405 29155
rect 15804 29124 16405 29152
rect 15804 29112 15810 29124
rect 16393 29121 16405 29124
rect 16439 29121 16451 29155
rect 16393 29115 16451 29121
rect 17218 29112 17224 29164
rect 17276 29152 17282 29164
rect 18049 29155 18107 29161
rect 18049 29152 18061 29155
rect 17276 29124 18061 29152
rect 17276 29112 17282 29124
rect 18049 29121 18061 29124
rect 18095 29121 18107 29155
rect 18049 29115 18107 29121
rect 22005 29155 22063 29161
rect 22005 29121 22017 29155
rect 22051 29152 22063 29155
rect 22646 29152 22652 29164
rect 22051 29124 22652 29152
rect 22051 29121 22063 29124
rect 22005 29115 22063 29121
rect 22646 29112 22652 29124
rect 22704 29112 22710 29164
rect 25317 29155 25375 29161
rect 25317 29121 25329 29155
rect 25363 29152 25375 29155
rect 25406 29152 25412 29164
rect 25363 29124 25412 29152
rect 25363 29121 25375 29124
rect 25317 29115 25375 29121
rect 25406 29112 25412 29124
rect 25464 29112 25470 29164
rect 14737 29087 14795 29093
rect 14737 29053 14749 29087
rect 14783 29053 14795 29087
rect 14737 29047 14795 29053
rect 15933 29087 15991 29093
rect 15933 29053 15945 29087
rect 15979 29084 15991 29087
rect 16114 29084 16120 29096
rect 15979 29056 16120 29084
rect 15979 29053 15991 29056
rect 15933 29047 15991 29053
rect 16114 29044 16120 29056
rect 16172 29044 16178 29096
rect 17034 29044 17040 29096
rect 17092 29084 17098 29096
rect 17313 29087 17371 29093
rect 17313 29084 17325 29087
rect 17092 29056 17325 29084
rect 17092 29044 17098 29056
rect 17313 29053 17325 29056
rect 17359 29053 17371 29087
rect 17313 29047 17371 29053
rect 17402 29044 17408 29096
rect 17460 29084 17466 29096
rect 17497 29087 17555 29093
rect 17497 29084 17509 29087
rect 17460 29056 17509 29084
rect 17460 29044 17466 29056
rect 17497 29053 17509 29056
rect 17543 29053 17555 29087
rect 17497 29047 17555 29053
rect 19794 29044 19800 29096
rect 19852 29084 19858 29096
rect 19889 29087 19947 29093
rect 19889 29084 19901 29087
rect 19852 29056 19901 29084
rect 19852 29044 19858 29056
rect 19889 29053 19901 29056
rect 19935 29053 19947 29087
rect 23661 29087 23719 29093
rect 23661 29084 23673 29087
rect 19889 29047 19947 29053
rect 22756 29056 23673 29084
rect 9490 28976 9496 29028
rect 9548 29016 9554 29028
rect 11149 29019 11207 29025
rect 11149 29016 11161 29019
rect 9548 28988 11161 29016
rect 9548 28976 9554 28988
rect 11149 28985 11161 28988
rect 11195 28985 11207 29019
rect 11149 28979 11207 28985
rect 12158 28976 12164 29028
rect 12216 29016 12222 29028
rect 12989 29019 13047 29025
rect 12989 29016 13001 29019
rect 12216 28988 13001 29016
rect 12216 28976 12222 28988
rect 12989 28985 13001 28988
rect 13035 28985 13047 29019
rect 12989 28979 13047 28985
rect 13630 28976 13636 29028
rect 13688 29016 13694 29028
rect 14185 29019 14243 29025
rect 14185 29016 14197 29019
rect 13688 28988 14197 29016
rect 13688 28976 13694 28988
rect 14185 28985 14197 28988
rect 14231 28985 14243 29019
rect 14185 28979 14243 28985
rect 21174 28976 21180 29028
rect 21232 29016 21238 29028
rect 22649 29019 22707 29025
rect 22649 29016 22661 29019
rect 21232 28988 22661 29016
rect 21232 28976 21238 28988
rect 22649 28985 22661 28988
rect 22695 28985 22707 29019
rect 22649 28979 22707 28985
rect 12434 28908 12440 28960
rect 12492 28948 12498 28960
rect 12529 28951 12587 28957
rect 12529 28948 12541 28951
rect 12492 28920 12541 28948
rect 12492 28908 12498 28920
rect 12529 28917 12541 28920
rect 12575 28917 12587 28951
rect 12529 28911 12587 28917
rect 22554 28908 22560 28960
rect 22612 28948 22618 28960
rect 22756 28948 22784 29056
rect 23661 29053 23673 29056
rect 23707 29053 23719 29087
rect 23661 29047 23719 29053
rect 24305 29087 24363 29093
rect 24305 29053 24317 29087
rect 24351 29084 24363 29087
rect 24854 29084 24860 29096
rect 24351 29056 24860 29084
rect 24351 29053 24363 29056
rect 24305 29047 24363 29053
rect 24854 29044 24860 29056
rect 24912 29044 24918 29096
rect 25133 29019 25191 29025
rect 25133 28985 25145 29019
rect 25179 29016 25191 29019
rect 25314 29016 25320 29028
rect 25179 28988 25320 29016
rect 25179 28985 25191 28988
rect 25133 28979 25191 28985
rect 25314 28976 25320 28988
rect 25372 28976 25378 29028
rect 22612 28920 22784 28948
rect 22612 28908 22618 28920
rect 1104 28858 25852 28880
rect 1104 28806 2950 28858
rect 3002 28806 3014 28858
rect 3066 28806 3078 28858
rect 3130 28806 3142 28858
rect 3194 28806 3206 28858
rect 3258 28806 12950 28858
rect 13002 28806 13014 28858
rect 13066 28806 13078 28858
rect 13130 28806 13142 28858
rect 13194 28806 13206 28858
rect 13258 28806 22950 28858
rect 23002 28806 23014 28858
rect 23066 28806 23078 28858
rect 23130 28806 23142 28858
rect 23194 28806 23206 28858
rect 23258 28806 25852 28858
rect 1104 28784 25852 28806
rect 10226 28704 10232 28756
rect 10284 28744 10290 28756
rect 11241 28747 11299 28753
rect 11241 28744 11253 28747
rect 10284 28716 11253 28744
rect 10284 28704 10290 28716
rect 11241 28713 11253 28716
rect 11287 28713 11299 28747
rect 11241 28707 11299 28713
rect 13906 28704 13912 28756
rect 13964 28704 13970 28756
rect 18782 28704 18788 28756
rect 18840 28744 18846 28756
rect 18877 28747 18935 28753
rect 18877 28744 18889 28747
rect 18840 28716 18889 28744
rect 18840 28704 18846 28716
rect 18877 28713 18889 28716
rect 18923 28713 18935 28747
rect 18877 28707 18935 28713
rect 13538 28676 13544 28688
rect 13096 28648 13544 28676
rect 9122 28568 9128 28620
rect 9180 28608 9186 28620
rect 9398 28608 9404 28620
rect 9180 28580 9404 28608
rect 9180 28568 9186 28580
rect 9398 28568 9404 28580
rect 9456 28608 9462 28620
rect 9493 28611 9551 28617
rect 9493 28608 9505 28611
rect 9456 28580 9505 28608
rect 9456 28568 9462 28580
rect 9493 28577 9505 28580
rect 9539 28608 9551 28611
rect 11514 28608 11520 28620
rect 9539 28580 11520 28608
rect 9539 28577 9551 28580
rect 9493 28571 9551 28577
rect 11514 28568 11520 28580
rect 11572 28608 11578 28620
rect 11701 28611 11759 28617
rect 11701 28608 11713 28611
rect 11572 28580 11713 28608
rect 11572 28568 11578 28580
rect 11701 28577 11713 28580
rect 11747 28577 11759 28611
rect 11701 28571 11759 28577
rect 11977 28611 12035 28617
rect 11977 28577 11989 28611
rect 12023 28608 12035 28611
rect 12434 28608 12440 28620
rect 12023 28580 12440 28608
rect 12023 28577 12035 28580
rect 11977 28571 12035 28577
rect 12434 28568 12440 28580
rect 12492 28568 12498 28620
rect 13096 28552 13124 28648
rect 13538 28636 13544 28648
rect 13596 28676 13602 28688
rect 14185 28679 14243 28685
rect 14185 28676 14197 28679
rect 13596 28648 14197 28676
rect 13596 28636 13602 28648
rect 14185 28645 14197 28648
rect 14231 28676 14243 28679
rect 15102 28676 15108 28688
rect 14231 28648 15108 28676
rect 14231 28645 14243 28648
rect 14185 28639 14243 28645
rect 15102 28636 15108 28648
rect 15160 28636 15166 28688
rect 20162 28676 20168 28688
rect 19996 28648 20168 28676
rect 19996 28617 20024 28648
rect 20162 28636 20168 28648
rect 20220 28636 20226 28688
rect 22830 28636 22836 28688
rect 22888 28676 22894 28688
rect 24581 28679 24639 28685
rect 24581 28676 24593 28679
rect 22888 28648 24593 28676
rect 22888 28636 22894 28648
rect 24581 28645 24593 28648
rect 24627 28645 24639 28679
rect 24581 28639 24639 28645
rect 15289 28611 15347 28617
rect 15289 28608 15301 28611
rect 13372 28580 15301 28608
rect 13078 28500 13084 28552
rect 13136 28500 13142 28552
rect 9766 28432 9772 28484
rect 9824 28432 9830 28484
rect 10152 28444 10258 28472
rect 10152 28416 10180 28444
rect 10134 28364 10140 28416
rect 10192 28364 10198 28416
rect 11974 28364 11980 28416
rect 12032 28404 12038 28416
rect 13372 28404 13400 28580
rect 15289 28577 15301 28580
rect 15335 28608 15347 28611
rect 16485 28611 16543 28617
rect 16485 28608 16497 28611
rect 15335 28580 16497 28608
rect 15335 28577 15347 28580
rect 15289 28571 15347 28577
rect 16485 28577 16497 28580
rect 16531 28577 16543 28611
rect 16485 28571 16543 28577
rect 17129 28611 17187 28617
rect 17129 28577 17141 28611
rect 17175 28608 17187 28611
rect 19981 28611 20039 28617
rect 17175 28580 19932 28608
rect 17175 28577 17187 28580
rect 17129 28571 17187 28577
rect 19904 28552 19932 28580
rect 19981 28577 19993 28611
rect 20027 28577 20039 28611
rect 19981 28571 20039 28577
rect 20070 28568 20076 28620
rect 20128 28608 20134 28620
rect 20901 28611 20959 28617
rect 20901 28608 20913 28611
rect 20128 28580 20913 28608
rect 20128 28568 20134 28580
rect 20901 28577 20913 28580
rect 20947 28577 20959 28611
rect 20901 28571 20959 28577
rect 24946 28568 24952 28620
rect 25004 28608 25010 28620
rect 25041 28611 25099 28617
rect 25041 28608 25053 28611
rect 25004 28580 25053 28608
rect 25004 28568 25010 28580
rect 25041 28577 25053 28580
rect 25087 28577 25099 28611
rect 25041 28571 25099 28577
rect 25222 28568 25228 28620
rect 25280 28568 25286 28620
rect 15105 28543 15163 28549
rect 15105 28509 15117 28543
rect 15151 28540 15163 28543
rect 15930 28540 15936 28552
rect 15151 28512 15936 28540
rect 15151 28509 15163 28512
rect 15105 28503 15163 28509
rect 15930 28500 15936 28512
rect 15988 28540 15994 28552
rect 16390 28540 16396 28552
rect 15988 28512 16396 28540
rect 15988 28500 15994 28512
rect 16390 28500 16396 28512
rect 16448 28500 16454 28552
rect 19794 28500 19800 28552
rect 19852 28500 19858 28552
rect 19886 28500 19892 28552
rect 19944 28540 19950 28552
rect 20625 28543 20683 28549
rect 20625 28540 20637 28543
rect 19944 28512 20637 28540
rect 19944 28500 19950 28512
rect 20625 28509 20637 28512
rect 20671 28509 20683 28543
rect 22034 28512 24164 28540
rect 20625 28503 20683 28509
rect 17402 28432 17408 28484
rect 17460 28432 17466 28484
rect 18414 28432 18420 28484
rect 18472 28432 18478 28484
rect 22186 28432 22192 28484
rect 22244 28472 22250 28484
rect 22833 28475 22891 28481
rect 22833 28472 22845 28475
rect 22244 28444 22845 28472
rect 22244 28432 22250 28444
rect 22833 28441 22845 28444
rect 22879 28441 22891 28475
rect 22833 28435 22891 28441
rect 23290 28432 23296 28484
rect 23348 28472 23354 28484
rect 23569 28475 23627 28481
rect 23569 28472 23581 28475
rect 23348 28444 23581 28472
rect 23348 28432 23354 28444
rect 23569 28441 23581 28444
rect 23615 28441 23627 28475
rect 23569 28435 23627 28441
rect 12032 28376 13400 28404
rect 12032 28364 12038 28376
rect 13446 28364 13452 28416
rect 13504 28364 13510 28416
rect 14734 28364 14740 28416
rect 14792 28364 14798 28416
rect 15194 28364 15200 28416
rect 15252 28364 15258 28416
rect 15930 28364 15936 28416
rect 15988 28364 15994 28416
rect 16206 28364 16212 28416
rect 16264 28404 16270 28416
rect 16301 28407 16359 28413
rect 16301 28404 16313 28407
rect 16264 28376 16313 28404
rect 16264 28364 16270 28376
rect 16301 28373 16313 28376
rect 16347 28373 16359 28407
rect 16301 28367 16359 28373
rect 16393 28407 16451 28413
rect 16393 28373 16405 28407
rect 16439 28404 16451 28407
rect 16482 28404 16488 28416
rect 16439 28376 16488 28404
rect 16439 28373 16451 28376
rect 16393 28367 16451 28373
rect 16482 28364 16488 28376
rect 16540 28364 16546 28416
rect 19150 28364 19156 28416
rect 19208 28404 19214 28416
rect 19429 28407 19487 28413
rect 19429 28404 19441 28407
rect 19208 28376 19441 28404
rect 19208 28364 19214 28376
rect 19429 28373 19441 28376
rect 19475 28373 19487 28407
rect 19429 28367 19487 28373
rect 19889 28407 19947 28413
rect 19889 28373 19901 28407
rect 19935 28404 19947 28407
rect 20254 28404 20260 28416
rect 19935 28376 20260 28404
rect 19935 28373 19947 28376
rect 19889 28367 19947 28373
rect 20254 28364 20260 28376
rect 20312 28364 20318 28416
rect 22373 28407 22431 28413
rect 22373 28373 22385 28407
rect 22419 28404 22431 28407
rect 22554 28404 22560 28416
rect 22419 28376 22560 28404
rect 22419 28373 22431 28376
rect 22373 28367 22431 28373
rect 22554 28364 22560 28376
rect 22612 28364 22618 28416
rect 24136 28413 24164 28512
rect 24854 28432 24860 28484
rect 24912 28472 24918 28484
rect 24949 28475 25007 28481
rect 24949 28472 24961 28475
rect 24912 28444 24961 28472
rect 24912 28432 24918 28444
rect 24949 28441 24961 28444
rect 24995 28441 25007 28475
rect 24949 28435 25007 28441
rect 24121 28407 24179 28413
rect 24121 28373 24133 28407
rect 24167 28404 24179 28407
rect 24302 28404 24308 28416
rect 24167 28376 24308 28404
rect 24167 28373 24179 28376
rect 24121 28367 24179 28373
rect 24302 28364 24308 28376
rect 24360 28364 24366 28416
rect 1104 28314 25852 28336
rect 1104 28262 7950 28314
rect 8002 28262 8014 28314
rect 8066 28262 8078 28314
rect 8130 28262 8142 28314
rect 8194 28262 8206 28314
rect 8258 28262 17950 28314
rect 18002 28262 18014 28314
rect 18066 28262 18078 28314
rect 18130 28262 18142 28314
rect 18194 28262 18206 28314
rect 18258 28262 25852 28314
rect 1104 28240 25852 28262
rect 9766 28160 9772 28212
rect 9824 28200 9830 28212
rect 11149 28203 11207 28209
rect 11149 28200 11161 28203
rect 9824 28172 11161 28200
rect 9824 28160 9830 28172
rect 11149 28169 11161 28172
rect 11195 28169 11207 28203
rect 11149 28163 11207 28169
rect 11790 28160 11796 28212
rect 11848 28200 11854 28212
rect 12345 28203 12403 28209
rect 12345 28200 12357 28203
rect 11848 28172 12357 28200
rect 11848 28160 11854 28172
rect 12345 28169 12357 28172
rect 12391 28169 12403 28203
rect 12345 28163 12403 28169
rect 12710 28160 12716 28212
rect 12768 28200 12774 28212
rect 13078 28200 13084 28212
rect 12768 28172 13084 28200
rect 12768 28160 12774 28172
rect 13078 28160 13084 28172
rect 13136 28160 13142 28212
rect 13633 28203 13691 28209
rect 13633 28169 13645 28203
rect 13679 28200 13691 28203
rect 14734 28200 14740 28212
rect 13679 28172 14740 28200
rect 13679 28169 13691 28172
rect 13633 28163 13691 28169
rect 14734 28160 14740 28172
rect 14792 28160 14798 28212
rect 14826 28160 14832 28212
rect 14884 28200 14890 28212
rect 15013 28203 15071 28209
rect 15013 28200 15025 28203
rect 14884 28172 15025 28200
rect 14884 28160 14890 28172
rect 15013 28169 15025 28172
rect 15059 28169 15071 28203
rect 15013 28163 15071 28169
rect 17402 28160 17408 28212
rect 17460 28200 17466 28212
rect 19889 28203 19947 28209
rect 19889 28200 19901 28203
rect 17460 28172 19901 28200
rect 17460 28160 17466 28172
rect 19889 28169 19901 28172
rect 19935 28169 19947 28203
rect 19889 28163 19947 28169
rect 20162 28160 20168 28212
rect 20220 28200 20226 28212
rect 23198 28200 23204 28212
rect 20220 28172 23204 28200
rect 20220 28160 20226 28172
rect 23198 28160 23204 28172
rect 23256 28160 23262 28212
rect 24673 28203 24731 28209
rect 24673 28169 24685 28203
rect 24719 28200 24731 28203
rect 25130 28200 25136 28212
rect 24719 28172 25136 28200
rect 24719 28169 24731 28172
rect 24673 28163 24731 28169
rect 25130 28160 25136 28172
rect 25188 28160 25194 28212
rect 25317 28203 25375 28209
rect 25317 28169 25329 28203
rect 25363 28200 25375 28203
rect 25406 28200 25412 28212
rect 25363 28172 25412 28200
rect 25363 28169 25375 28172
rect 25317 28163 25375 28169
rect 25406 28160 25412 28172
rect 25464 28160 25470 28212
rect 11974 28132 11980 28144
rect 10520 28104 11980 28132
rect 10520 28073 10548 28104
rect 11974 28092 11980 28104
rect 12032 28092 12038 28144
rect 13541 28135 13599 28141
rect 13541 28101 13553 28135
rect 13587 28132 13599 28135
rect 15930 28132 15936 28144
rect 13587 28104 15936 28132
rect 13587 28101 13599 28104
rect 13541 28095 13599 28101
rect 15930 28092 15936 28104
rect 15988 28092 15994 28144
rect 18509 28135 18567 28141
rect 18509 28101 18521 28135
rect 18555 28132 18567 28135
rect 19426 28132 19432 28144
rect 18555 28104 19432 28132
rect 18555 28101 18567 28104
rect 18509 28095 18567 28101
rect 19426 28092 19432 28104
rect 19484 28092 19490 28144
rect 22186 28132 22192 28144
rect 20548 28104 22192 28132
rect 10505 28067 10563 28073
rect 10505 28033 10517 28067
rect 10551 28033 10563 28067
rect 10505 28027 10563 28033
rect 11146 28024 11152 28076
rect 11204 28064 11210 28076
rect 11701 28067 11759 28073
rect 11701 28064 11713 28067
rect 11204 28036 11713 28064
rect 11204 28024 11210 28036
rect 11701 28033 11713 28036
rect 11747 28033 11759 28067
rect 11701 28027 11759 28033
rect 13446 28024 13452 28076
rect 13504 28064 13510 28076
rect 14369 28067 14427 28073
rect 14369 28064 14381 28067
rect 13504 28036 14381 28064
rect 13504 28024 13510 28036
rect 14369 28033 14381 28036
rect 14415 28033 14427 28067
rect 14369 28027 14427 28033
rect 15473 28067 15531 28073
rect 15473 28033 15485 28067
rect 15519 28064 15531 28067
rect 16022 28064 16028 28076
rect 15519 28036 16028 28064
rect 15519 28033 15531 28036
rect 15473 28027 15531 28033
rect 16022 28024 16028 28036
rect 16080 28024 16086 28076
rect 16666 28024 16672 28076
rect 16724 28064 16730 28076
rect 17221 28067 17279 28073
rect 17221 28064 17233 28067
rect 16724 28036 17233 28064
rect 16724 28024 16730 28036
rect 17221 28033 17233 28036
rect 17267 28033 17279 28067
rect 17221 28027 17279 28033
rect 17313 28067 17371 28073
rect 17313 28033 17325 28067
rect 17359 28064 17371 28067
rect 17678 28064 17684 28076
rect 17359 28036 17684 28064
rect 17359 28033 17371 28036
rect 17313 28027 17371 28033
rect 13725 27999 13783 28005
rect 13725 27965 13737 27999
rect 13771 27965 13783 27999
rect 17236 27996 17264 28027
rect 17678 28024 17684 28036
rect 17736 28024 17742 28076
rect 18414 28024 18420 28076
rect 18472 28024 18478 28076
rect 19242 28024 19248 28076
rect 19300 28024 19306 28076
rect 20548 28073 20576 28104
rect 22186 28092 22192 28104
rect 22244 28092 22250 28144
rect 24302 28132 24308 28144
rect 23506 28104 24308 28132
rect 24302 28092 24308 28104
rect 24360 28092 24366 28144
rect 20533 28067 20591 28073
rect 20533 28064 20545 28067
rect 19812 28036 20545 28064
rect 17402 27996 17408 28008
rect 17236 27968 17408 27996
rect 13725 27959 13783 27965
rect 10226 27888 10232 27940
rect 10284 27928 10290 27940
rect 13740 27928 13768 27959
rect 17402 27956 17408 27968
rect 17460 27956 17466 28008
rect 17494 27956 17500 28008
rect 17552 27956 17558 28008
rect 18598 27956 18604 28008
rect 18656 27956 18662 28008
rect 10284 27900 13768 27928
rect 10284 27888 10290 27900
rect 14826 27888 14832 27940
rect 14884 27928 14890 27940
rect 16853 27931 16911 27937
rect 16853 27928 16865 27931
rect 14884 27900 16865 27928
rect 14884 27888 14890 27900
rect 16853 27897 16865 27900
rect 16899 27897 16911 27931
rect 19812 27928 19840 28036
rect 20533 28033 20545 28036
rect 20579 28033 20591 28067
rect 20533 28027 20591 28033
rect 24578 28024 24584 28076
rect 24636 28024 24642 28076
rect 19886 27956 19892 28008
rect 19944 27996 19950 28008
rect 21269 27999 21327 28005
rect 21269 27996 21281 27999
rect 19944 27968 21281 27996
rect 19944 27956 19950 27968
rect 21269 27965 21281 27968
rect 21315 27965 21327 27999
rect 21269 27959 21327 27965
rect 21910 27956 21916 28008
rect 21968 27956 21974 28008
rect 22005 27999 22063 28005
rect 22005 27965 22017 27999
rect 22051 27965 22063 27999
rect 22005 27959 22063 27965
rect 22281 27999 22339 28005
rect 22281 27965 22293 27999
rect 22327 27996 22339 27999
rect 22327 27968 24716 27996
rect 22327 27965 22339 27968
rect 22281 27959 22339 27965
rect 20165 27931 20223 27937
rect 20165 27928 20177 27931
rect 16853 27891 16911 27897
rect 17328 27900 20177 27928
rect 17328 27872 17356 27900
rect 20165 27897 20177 27900
rect 20211 27897 20223 27931
rect 21928 27928 21956 27956
rect 20165 27891 20223 27897
rect 20272 27900 21956 27928
rect 12802 27820 12808 27872
rect 12860 27860 12866 27872
rect 13173 27863 13231 27869
rect 13173 27860 13185 27863
rect 12860 27832 13185 27860
rect 12860 27820 12866 27832
rect 13173 27829 13185 27832
rect 13219 27829 13231 27863
rect 13173 27823 13231 27829
rect 13998 27820 14004 27872
rect 14056 27860 14062 27872
rect 16117 27863 16175 27869
rect 16117 27860 16129 27863
rect 14056 27832 16129 27860
rect 14056 27820 14062 27832
rect 16117 27829 16129 27832
rect 16163 27829 16175 27863
rect 16117 27823 16175 27829
rect 16390 27820 16396 27872
rect 16448 27820 16454 27872
rect 17310 27820 17316 27872
rect 17368 27820 17374 27872
rect 17954 27820 17960 27872
rect 18012 27860 18018 27872
rect 18049 27863 18107 27869
rect 18049 27860 18061 27863
rect 18012 27832 18061 27860
rect 18012 27820 18018 27832
rect 18049 27829 18061 27832
rect 18095 27829 18107 27863
rect 18049 27823 18107 27829
rect 19058 27820 19064 27872
rect 19116 27860 19122 27872
rect 20272 27860 20300 27900
rect 19116 27832 20300 27860
rect 19116 27820 19122 27832
rect 20438 27820 20444 27872
rect 20496 27860 20502 27872
rect 22020 27860 22048 27959
rect 23474 27888 23480 27940
rect 23532 27928 23538 27940
rect 24213 27931 24271 27937
rect 24213 27928 24225 27931
rect 23532 27900 24225 27928
rect 23532 27888 23538 27900
rect 24213 27897 24225 27900
rect 24259 27897 24271 27931
rect 24688 27928 24716 27968
rect 24762 27956 24768 28008
rect 24820 27956 24826 28008
rect 25222 27928 25228 27940
rect 24688 27900 25228 27928
rect 24213 27891 24271 27897
rect 25222 27888 25228 27900
rect 25280 27888 25286 27940
rect 23290 27860 23296 27872
rect 20496 27832 23296 27860
rect 20496 27820 20502 27832
rect 23290 27820 23296 27832
rect 23348 27820 23354 27872
rect 23382 27820 23388 27872
rect 23440 27860 23446 27872
rect 23753 27863 23811 27869
rect 23753 27860 23765 27863
rect 23440 27832 23765 27860
rect 23440 27820 23446 27832
rect 23753 27829 23765 27832
rect 23799 27829 23811 27863
rect 23753 27823 23811 27829
rect 25130 27820 25136 27872
rect 25188 27860 25194 27872
rect 25409 27863 25467 27869
rect 25409 27860 25421 27863
rect 25188 27832 25421 27860
rect 25188 27820 25194 27832
rect 25409 27829 25421 27832
rect 25455 27829 25467 27863
rect 25409 27823 25467 27829
rect 1104 27770 25852 27792
rect 1104 27718 2950 27770
rect 3002 27718 3014 27770
rect 3066 27718 3078 27770
rect 3130 27718 3142 27770
rect 3194 27718 3206 27770
rect 3258 27718 12950 27770
rect 13002 27718 13014 27770
rect 13066 27718 13078 27770
rect 13130 27718 13142 27770
rect 13194 27718 13206 27770
rect 13258 27718 22950 27770
rect 23002 27718 23014 27770
rect 23066 27718 23078 27770
rect 23130 27718 23142 27770
rect 23194 27718 23206 27770
rect 23258 27718 25852 27770
rect 1104 27696 25852 27718
rect 14642 27616 14648 27668
rect 14700 27656 14706 27668
rect 15102 27656 15108 27668
rect 14700 27628 15108 27656
rect 14700 27616 14706 27628
rect 15102 27616 15108 27628
rect 15160 27616 15166 27668
rect 20152 27659 20210 27665
rect 20152 27625 20164 27659
rect 20198 27656 20210 27659
rect 21174 27656 21180 27668
rect 20198 27628 21180 27656
rect 20198 27625 20210 27628
rect 20152 27619 20210 27625
rect 21174 27616 21180 27628
rect 21232 27616 21238 27668
rect 11974 27548 11980 27600
rect 12032 27548 12038 27600
rect 18690 27588 18696 27600
rect 17144 27560 18696 27588
rect 17144 27532 17172 27560
rect 18690 27548 18696 27560
rect 18748 27548 18754 27600
rect 21192 27560 24164 27588
rect 10505 27523 10563 27529
rect 10505 27489 10517 27523
rect 10551 27520 10563 27523
rect 13081 27523 13139 27529
rect 13081 27520 13093 27523
rect 10551 27492 13093 27520
rect 10551 27489 10563 27492
rect 10505 27483 10563 27489
rect 13081 27489 13093 27492
rect 13127 27489 13139 27523
rect 13081 27483 13139 27489
rect 15102 27480 15108 27532
rect 15160 27520 15166 27532
rect 16025 27523 16083 27529
rect 16025 27520 16037 27523
rect 15160 27492 16037 27520
rect 15160 27480 15166 27492
rect 16025 27489 16037 27492
rect 16071 27489 16083 27523
rect 17126 27520 17132 27532
rect 16025 27483 16083 27489
rect 16408 27492 17132 27520
rect 9122 27412 9128 27464
rect 9180 27452 9186 27464
rect 10229 27455 10287 27461
rect 10229 27452 10241 27455
rect 9180 27424 10241 27452
rect 9180 27412 9186 27424
rect 10229 27421 10241 27424
rect 10275 27421 10287 27455
rect 10229 27415 10287 27421
rect 10244 27316 10272 27415
rect 12066 27412 12072 27464
rect 12124 27452 12130 27464
rect 12437 27455 12495 27461
rect 12437 27452 12449 27455
rect 12124 27424 12449 27452
rect 12124 27412 12130 27424
rect 12437 27421 12449 27424
rect 12483 27421 12495 27455
rect 12437 27415 12495 27421
rect 15841 27455 15899 27461
rect 15841 27421 15853 27455
rect 15887 27452 15899 27455
rect 16206 27452 16212 27464
rect 15887 27424 16212 27452
rect 15887 27421 15899 27424
rect 15841 27415 15899 27421
rect 16206 27412 16212 27424
rect 16264 27452 16270 27464
rect 16408 27452 16436 27492
rect 17126 27480 17132 27492
rect 17184 27480 17190 27532
rect 18049 27523 18107 27529
rect 18049 27489 18061 27523
rect 18095 27520 18107 27523
rect 18414 27520 18420 27532
rect 18095 27492 18420 27520
rect 18095 27489 18107 27492
rect 18049 27483 18107 27489
rect 18414 27480 18420 27492
rect 18472 27480 18478 27532
rect 19337 27523 19395 27529
rect 19337 27489 19349 27523
rect 19383 27520 19395 27523
rect 20162 27520 20168 27532
rect 19383 27492 20168 27520
rect 19383 27489 19395 27492
rect 19337 27483 19395 27489
rect 16264 27424 16436 27452
rect 16264 27412 16270 27424
rect 16482 27412 16488 27464
rect 16540 27412 16546 27464
rect 17494 27412 17500 27464
rect 17552 27452 17558 27464
rect 17954 27452 17960 27464
rect 17552 27424 17960 27452
rect 17552 27412 17558 27424
rect 17954 27412 17960 27424
rect 18012 27412 18018 27464
rect 18877 27455 18935 27461
rect 18877 27421 18889 27455
rect 18923 27452 18935 27455
rect 19352 27452 19380 27483
rect 20162 27480 20168 27492
rect 20220 27480 20226 27532
rect 20254 27480 20260 27532
rect 20312 27520 20318 27532
rect 21192 27520 21220 27560
rect 20312 27492 21220 27520
rect 20312 27480 20318 27492
rect 22646 27480 22652 27532
rect 22704 27520 22710 27532
rect 23382 27520 23388 27532
rect 22704 27492 23388 27520
rect 22704 27480 22710 27492
rect 23382 27480 23388 27492
rect 23440 27480 23446 27532
rect 23934 27480 23940 27532
rect 23992 27480 23998 27532
rect 24136 27520 24164 27560
rect 25222 27548 25228 27600
rect 25280 27548 25286 27600
rect 26234 27520 26240 27532
rect 24136 27492 26240 27520
rect 26234 27480 26240 27492
rect 26292 27480 26298 27532
rect 18923 27424 19380 27452
rect 18923 27421 18935 27424
rect 18877 27415 18935 27421
rect 19426 27412 19432 27464
rect 19484 27452 19490 27464
rect 19886 27452 19892 27464
rect 19484 27424 19892 27452
rect 19484 27412 19490 27424
rect 19886 27412 19892 27424
rect 19944 27412 19950 27464
rect 22278 27412 22284 27464
rect 22336 27452 22342 27464
rect 22465 27455 22523 27461
rect 22465 27452 22477 27455
rect 22336 27424 22477 27452
rect 22336 27412 22342 27424
rect 22465 27421 22477 27424
rect 22511 27421 22523 27455
rect 22465 27415 22523 27421
rect 23658 27412 23664 27464
rect 23716 27412 23722 27464
rect 23753 27455 23811 27461
rect 23753 27421 23765 27455
rect 23799 27452 23811 27455
rect 24026 27452 24032 27464
rect 23799 27424 24032 27452
rect 23799 27421 23811 27424
rect 23753 27415 23811 27421
rect 24026 27412 24032 27424
rect 24084 27412 24090 27464
rect 24486 27412 24492 27464
rect 24544 27452 24550 27464
rect 24581 27455 24639 27461
rect 24581 27452 24593 27455
rect 24544 27424 24593 27452
rect 24544 27412 24550 27424
rect 24581 27421 24593 27424
rect 24627 27421 24639 27455
rect 24581 27415 24639 27421
rect 12710 27384 12716 27396
rect 11730 27356 12716 27384
rect 12710 27344 12716 27356
rect 12768 27344 12774 27396
rect 15933 27387 15991 27393
rect 15933 27353 15945 27387
rect 15979 27384 15991 27387
rect 16500 27384 16528 27412
rect 16853 27387 16911 27393
rect 16853 27384 16865 27387
rect 15979 27356 16865 27384
rect 15979 27353 15991 27356
rect 15933 27347 15991 27353
rect 16853 27353 16865 27356
rect 16899 27384 16911 27387
rect 17221 27387 17279 27393
rect 17221 27384 17233 27387
rect 16899 27356 17233 27384
rect 16899 27353 16911 27356
rect 16853 27347 16911 27353
rect 17221 27353 17233 27356
rect 17267 27384 17279 27387
rect 18598 27384 18604 27396
rect 17267 27356 18604 27384
rect 17267 27353 17279 27356
rect 17221 27347 17279 27353
rect 18598 27344 18604 27356
rect 18656 27384 18662 27396
rect 20254 27384 20260 27396
rect 18656 27356 20260 27384
rect 18656 27344 18662 27356
rect 20254 27344 20260 27356
rect 20312 27344 20318 27396
rect 21542 27384 21548 27396
rect 21390 27356 21548 27384
rect 21542 27344 21548 27356
rect 21600 27344 21606 27396
rect 22557 27387 22615 27393
rect 22557 27353 22569 27387
rect 22603 27384 22615 27387
rect 24118 27384 24124 27396
rect 22603 27356 24124 27384
rect 22603 27353 22615 27356
rect 22557 27347 22615 27353
rect 24118 27344 24124 27356
rect 24176 27344 24182 27396
rect 11330 27316 11336 27328
rect 10244 27288 11336 27316
rect 11330 27276 11336 27288
rect 11388 27276 11394 27328
rect 15470 27276 15476 27328
rect 15528 27276 15534 27328
rect 16482 27276 16488 27328
rect 16540 27276 16546 27328
rect 17037 27319 17095 27325
rect 17037 27285 17049 27319
rect 17083 27316 17095 27319
rect 17126 27316 17132 27328
rect 17083 27288 17132 27316
rect 17083 27285 17095 27288
rect 17037 27279 17095 27285
rect 17126 27276 17132 27288
rect 17184 27316 17190 27328
rect 17313 27319 17371 27325
rect 17313 27316 17325 27319
rect 17184 27288 17325 27316
rect 17184 27276 17190 27288
rect 17313 27285 17325 27288
rect 17359 27285 17371 27319
rect 17313 27279 17371 27285
rect 17402 27276 17408 27328
rect 17460 27316 17466 27328
rect 17497 27319 17555 27325
rect 17497 27316 17509 27319
rect 17460 27288 17509 27316
rect 17460 27276 17466 27288
rect 17497 27285 17509 27288
rect 17543 27285 17555 27319
rect 17497 27279 17555 27285
rect 17678 27276 17684 27328
rect 17736 27276 17742 27328
rect 18693 27319 18751 27325
rect 18693 27285 18705 27319
rect 18739 27316 18751 27319
rect 20990 27316 20996 27328
rect 18739 27288 20996 27316
rect 18739 27285 18751 27288
rect 18693 27279 18751 27285
rect 20990 27276 20996 27288
rect 21048 27276 21054 27328
rect 21174 27276 21180 27328
rect 21232 27316 21238 27328
rect 21637 27319 21695 27325
rect 21637 27316 21649 27319
rect 21232 27288 21649 27316
rect 21232 27276 21238 27288
rect 21637 27285 21649 27288
rect 21683 27285 21695 27319
rect 21637 27279 21695 27285
rect 22097 27319 22155 27325
rect 22097 27285 22109 27319
rect 22143 27316 22155 27319
rect 22278 27316 22284 27328
rect 22143 27288 22284 27316
rect 22143 27285 22155 27288
rect 22097 27279 22155 27285
rect 22278 27276 22284 27288
rect 22336 27276 22342 27328
rect 22738 27276 22744 27328
rect 22796 27316 22802 27328
rect 23293 27319 23351 27325
rect 23293 27316 23305 27319
rect 22796 27288 23305 27316
rect 22796 27276 22802 27288
rect 23293 27285 23305 27288
rect 23339 27285 23351 27319
rect 23293 27279 23351 27285
rect 1104 27226 25852 27248
rect 1104 27174 7950 27226
rect 8002 27174 8014 27226
rect 8066 27174 8078 27226
rect 8130 27174 8142 27226
rect 8194 27174 8206 27226
rect 8258 27174 17950 27226
rect 18002 27174 18014 27226
rect 18066 27174 18078 27226
rect 18130 27174 18142 27226
rect 18194 27174 18206 27226
rect 18258 27174 25852 27226
rect 1104 27152 25852 27174
rect 11517 27115 11575 27121
rect 11517 27112 11529 27115
rect 10060 27084 11529 27112
rect 10060 27044 10088 27084
rect 11517 27081 11529 27084
rect 11563 27112 11575 27115
rect 12069 27115 12127 27121
rect 12069 27112 12081 27115
rect 11563 27084 12081 27112
rect 11563 27081 11575 27084
rect 11517 27075 11575 27081
rect 12069 27081 12081 27084
rect 12115 27112 12127 27115
rect 12250 27112 12256 27124
rect 12115 27084 12256 27112
rect 12115 27081 12127 27084
rect 12069 27075 12127 27081
rect 12250 27072 12256 27084
rect 12308 27072 12314 27124
rect 14461 27115 14519 27121
rect 14461 27112 14473 27115
rect 12406 27084 14473 27112
rect 10134 27044 10140 27056
rect 10060 27016 10140 27044
rect 10134 27004 10140 27016
rect 10192 27004 10198 27056
rect 9398 26936 9404 26988
rect 9456 26936 9462 26988
rect 11514 26936 11520 26988
rect 11572 26976 11578 26988
rect 12406 26976 12434 27084
rect 14461 27081 14473 27084
rect 14507 27112 14519 27115
rect 15010 27112 15016 27124
rect 14507 27084 15016 27112
rect 14507 27081 14519 27084
rect 14461 27075 14519 27081
rect 15010 27072 15016 27084
rect 15068 27072 15074 27124
rect 18598 27072 18604 27124
rect 18656 27112 18662 27124
rect 21177 27115 21235 27121
rect 18656 27084 19564 27112
rect 18656 27072 18662 27084
rect 14642 27044 14648 27056
rect 14214 27016 14648 27044
rect 14642 27004 14648 27016
rect 14700 27004 14706 27056
rect 15194 27004 15200 27056
rect 15252 27044 15258 27056
rect 15473 27047 15531 27053
rect 15473 27044 15485 27047
rect 15252 27016 15485 27044
rect 15252 27004 15258 27016
rect 15473 27013 15485 27016
rect 15519 27044 15531 27047
rect 15930 27044 15936 27056
rect 15519 27016 15936 27044
rect 15519 27013 15531 27016
rect 15473 27007 15531 27013
rect 15930 27004 15936 27016
rect 15988 27004 15994 27056
rect 18506 27004 18512 27056
rect 18564 27044 18570 27056
rect 19536 27044 19564 27084
rect 21177 27081 21189 27115
rect 21223 27112 21235 27115
rect 23566 27112 23572 27124
rect 21223 27084 23572 27112
rect 21223 27081 21235 27084
rect 21177 27075 21235 27081
rect 23566 27072 23572 27084
rect 23624 27072 23630 27124
rect 24302 27072 24308 27124
rect 24360 27112 24366 27124
rect 25130 27112 25136 27124
rect 24360 27084 25136 27112
rect 24360 27072 24366 27084
rect 21634 27044 21640 27056
rect 18564 27016 18722 27044
rect 19536 27016 21640 27044
rect 18564 27004 18570 27016
rect 21634 27004 21640 27016
rect 21692 27004 21698 27056
rect 24780 27044 24808 27084
rect 25130 27072 25136 27084
rect 25188 27112 25194 27124
rect 25225 27115 25283 27121
rect 25225 27112 25237 27115
rect 25188 27084 25237 27112
rect 25188 27072 25194 27084
rect 25225 27081 25237 27084
rect 25271 27081 25283 27115
rect 25225 27075 25283 27081
rect 25406 27072 25412 27124
rect 25464 27112 25470 27124
rect 25501 27115 25559 27121
rect 25501 27112 25513 27115
rect 25464 27084 25513 27112
rect 25464 27072 25470 27084
rect 25501 27081 25513 27084
rect 25547 27112 25559 27115
rect 26050 27112 26056 27124
rect 25547 27084 26056 27112
rect 25547 27081 25559 27084
rect 25501 27075 25559 27081
rect 26050 27072 26056 27084
rect 26108 27072 26114 27124
rect 24702 27016 24808 27044
rect 11572 26948 12434 26976
rect 11572 26936 11578 26948
rect 14734 26936 14740 26988
rect 14792 26976 14798 26988
rect 15381 26979 15439 26985
rect 15381 26976 15393 26979
rect 14792 26948 15393 26976
rect 14792 26936 14798 26948
rect 15381 26945 15393 26948
rect 15427 26976 15439 26979
rect 16025 26979 16083 26985
rect 16025 26976 16037 26979
rect 15427 26948 16037 26976
rect 15427 26945 15439 26948
rect 15381 26939 15439 26945
rect 16025 26945 16037 26948
rect 16071 26976 16083 26979
rect 16390 26976 16396 26988
rect 16071 26948 16396 26976
rect 16071 26945 16083 26948
rect 16025 26939 16083 26945
rect 16390 26936 16396 26948
rect 16448 26936 16454 26988
rect 20441 26979 20499 26985
rect 20441 26945 20453 26979
rect 20487 26976 20499 26979
rect 21085 26979 21143 26985
rect 21085 26976 21097 26979
rect 20487 26948 21097 26976
rect 20487 26945 20499 26948
rect 20441 26939 20499 26945
rect 21085 26945 21097 26948
rect 21131 26945 21143 26979
rect 21085 26939 21143 26945
rect 9677 26911 9735 26917
rect 9677 26877 9689 26911
rect 9723 26908 9735 26911
rect 10226 26908 10232 26920
rect 9723 26880 10232 26908
rect 9723 26877 9735 26880
rect 9677 26871 9735 26877
rect 10226 26868 10232 26880
rect 10284 26868 10290 26920
rect 11330 26868 11336 26920
rect 11388 26908 11394 26920
rect 12342 26908 12348 26920
rect 11388 26880 12348 26908
rect 11388 26868 11394 26880
rect 12342 26868 12348 26880
rect 12400 26908 12406 26920
rect 12713 26911 12771 26917
rect 12713 26908 12725 26911
rect 12400 26880 12725 26908
rect 12400 26868 12406 26880
rect 12713 26877 12725 26880
rect 12759 26877 12771 26911
rect 12713 26871 12771 26877
rect 12989 26911 13047 26917
rect 12989 26877 13001 26911
rect 13035 26908 13047 26911
rect 13998 26908 14004 26920
rect 13035 26880 14004 26908
rect 13035 26877 13047 26880
rect 12989 26871 13047 26877
rect 13998 26868 14004 26880
rect 14056 26868 14062 26920
rect 15565 26911 15623 26917
rect 15565 26877 15577 26911
rect 15611 26877 15623 26911
rect 15565 26871 15623 26877
rect 17957 26911 18015 26917
rect 17957 26877 17969 26911
rect 18003 26877 18015 26911
rect 17957 26871 18015 26877
rect 18233 26911 18291 26917
rect 18233 26877 18245 26911
rect 18279 26908 18291 26911
rect 20070 26908 20076 26920
rect 18279 26880 20076 26908
rect 18279 26877 18291 26880
rect 18233 26871 18291 26877
rect 10704 26812 12848 26840
rect 9674 26732 9680 26784
rect 9732 26772 9738 26784
rect 10704 26772 10732 26812
rect 9732 26744 10732 26772
rect 9732 26732 9738 26744
rect 11146 26732 11152 26784
rect 11204 26732 11210 26784
rect 12250 26732 12256 26784
rect 12308 26772 12314 26784
rect 12710 26772 12716 26784
rect 12308 26744 12716 26772
rect 12308 26732 12314 26744
rect 12710 26732 12716 26744
rect 12768 26732 12774 26784
rect 12820 26772 12848 26812
rect 14090 26800 14096 26852
rect 14148 26840 14154 26852
rect 15102 26840 15108 26852
rect 14148 26812 15108 26840
rect 14148 26800 14154 26812
rect 15102 26800 15108 26812
rect 15160 26840 15166 26852
rect 15580 26840 15608 26871
rect 15160 26812 15608 26840
rect 15160 26800 15166 26812
rect 14274 26772 14280 26784
rect 12820 26744 14280 26772
rect 14274 26732 14280 26744
rect 14332 26732 14338 26784
rect 14366 26732 14372 26784
rect 14424 26772 14430 26784
rect 15013 26775 15071 26781
rect 15013 26772 15025 26775
rect 14424 26744 15025 26772
rect 14424 26732 14430 26744
rect 15013 26741 15025 26744
rect 15059 26741 15071 26775
rect 15013 26735 15071 26741
rect 15930 26732 15936 26784
rect 15988 26772 15994 26784
rect 16209 26775 16267 26781
rect 16209 26772 16221 26775
rect 15988 26744 16221 26772
rect 15988 26732 15994 26744
rect 16209 26741 16221 26744
rect 16255 26772 16267 26775
rect 16482 26772 16488 26784
rect 16255 26744 16488 26772
rect 16255 26741 16267 26744
rect 16209 26735 16267 26741
rect 16482 26732 16488 26744
rect 16540 26732 16546 26784
rect 17972 26772 18000 26871
rect 20070 26868 20076 26880
rect 20128 26868 20134 26920
rect 19242 26800 19248 26852
rect 19300 26840 19306 26852
rect 19705 26843 19763 26849
rect 19705 26840 19717 26843
rect 19300 26812 19717 26840
rect 19300 26800 19306 26812
rect 19705 26809 19717 26812
rect 19751 26809 19763 26843
rect 19705 26803 19763 26809
rect 19981 26843 20039 26849
rect 19981 26809 19993 26843
rect 20027 26840 20039 26843
rect 21100 26840 21128 26939
rect 21174 26936 21180 26988
rect 21232 26976 21238 26988
rect 22005 26979 22063 26985
rect 22005 26976 22017 26979
rect 21232 26948 22017 26976
rect 21232 26936 21238 26948
rect 22005 26945 22017 26948
rect 22051 26945 22063 26979
rect 22005 26939 22063 26945
rect 21266 26868 21272 26920
rect 21324 26868 21330 26920
rect 23198 26868 23204 26920
rect 23256 26868 23262 26920
rect 23477 26911 23535 26917
rect 23477 26877 23489 26911
rect 23523 26908 23535 26911
rect 25222 26908 25228 26920
rect 23523 26880 25228 26908
rect 23523 26877 23535 26880
rect 23477 26871 23535 26877
rect 25222 26868 25228 26880
rect 25280 26868 25286 26920
rect 20027 26812 21036 26840
rect 21100 26812 23336 26840
rect 20027 26809 20039 26812
rect 19981 26803 20039 26809
rect 19426 26772 19432 26784
rect 17972 26744 19432 26772
rect 19426 26732 19432 26744
rect 19484 26732 19490 26784
rect 20717 26775 20775 26781
rect 20717 26741 20729 26775
rect 20763 26772 20775 26775
rect 20898 26772 20904 26784
rect 20763 26744 20904 26772
rect 20763 26741 20775 26744
rect 20717 26735 20775 26741
rect 20898 26732 20904 26744
rect 20956 26732 20962 26784
rect 21008 26772 21036 26812
rect 21634 26772 21640 26784
rect 21008 26744 21640 26772
rect 21634 26732 21640 26744
rect 21692 26732 21698 26784
rect 22646 26732 22652 26784
rect 22704 26732 22710 26784
rect 23308 26772 23336 26812
rect 23566 26772 23572 26784
rect 23308 26744 23572 26772
rect 23566 26732 23572 26744
rect 23624 26732 23630 26784
rect 23658 26732 23664 26784
rect 23716 26772 23722 26784
rect 24486 26772 24492 26784
rect 23716 26744 24492 26772
rect 23716 26732 23722 26744
rect 24486 26732 24492 26744
rect 24544 26772 24550 26784
rect 24949 26775 25007 26781
rect 24949 26772 24961 26775
rect 24544 26744 24961 26772
rect 24544 26732 24550 26744
rect 24949 26741 24961 26744
rect 24995 26741 25007 26775
rect 24949 26735 25007 26741
rect 1104 26682 25852 26704
rect 1104 26630 2950 26682
rect 3002 26630 3014 26682
rect 3066 26630 3078 26682
rect 3130 26630 3142 26682
rect 3194 26630 3206 26682
rect 3258 26630 12950 26682
rect 13002 26630 13014 26682
rect 13066 26630 13078 26682
rect 13130 26630 13142 26682
rect 13194 26630 13206 26682
rect 13258 26630 22950 26682
rect 23002 26630 23014 26682
rect 23066 26630 23078 26682
rect 23130 26630 23142 26682
rect 23194 26630 23206 26682
rect 23258 26630 25852 26682
rect 1104 26608 25852 26630
rect 10873 26571 10931 26577
rect 10873 26537 10885 26571
rect 10919 26568 10931 26571
rect 12066 26568 12072 26580
rect 10919 26540 12072 26568
rect 10919 26537 10931 26540
rect 10873 26531 10931 26537
rect 12066 26528 12072 26540
rect 12124 26528 12130 26580
rect 13998 26528 14004 26580
rect 14056 26568 14062 26580
rect 15657 26571 15715 26577
rect 15657 26568 15669 26571
rect 14056 26540 15669 26568
rect 14056 26528 14062 26540
rect 15657 26537 15669 26540
rect 15703 26537 15715 26571
rect 15657 26531 15715 26537
rect 19692 26571 19750 26577
rect 19692 26537 19704 26571
rect 19738 26568 19750 26571
rect 22646 26568 22652 26580
rect 19738 26540 22652 26568
rect 19738 26537 19750 26540
rect 19692 26531 19750 26537
rect 22646 26528 22652 26540
rect 22704 26528 22710 26580
rect 23566 26528 23572 26580
rect 23624 26568 23630 26580
rect 25406 26568 25412 26580
rect 23624 26540 25412 26568
rect 23624 26528 23630 26540
rect 25406 26528 25412 26540
rect 25464 26528 25470 26580
rect 11793 26503 11851 26509
rect 11793 26469 11805 26503
rect 11839 26500 11851 26503
rect 12894 26500 12900 26512
rect 11839 26472 12900 26500
rect 11839 26469 11851 26472
rect 11793 26463 11851 26469
rect 12894 26460 12900 26472
rect 12952 26460 12958 26512
rect 12989 26503 13047 26509
rect 12989 26469 13001 26503
rect 13035 26500 13047 26503
rect 15102 26500 15108 26512
rect 13035 26472 15108 26500
rect 13035 26469 13047 26472
rect 12989 26463 13047 26469
rect 15102 26460 15108 26472
rect 15160 26460 15166 26512
rect 24581 26503 24639 26509
rect 16132 26472 16988 26500
rect 9122 26392 9128 26444
rect 9180 26392 9186 26444
rect 9401 26435 9459 26441
rect 9401 26401 9413 26435
rect 9447 26432 9459 26435
rect 9490 26432 9496 26444
rect 9447 26404 9496 26432
rect 9447 26401 9459 26404
rect 9401 26395 9459 26401
rect 9490 26392 9496 26404
rect 9548 26392 9554 26444
rect 10134 26392 10140 26444
rect 10192 26432 10198 26444
rect 10192 26404 11100 26432
rect 10192 26392 10198 26404
rect 11072 26364 11100 26404
rect 11146 26392 11152 26444
rect 11204 26432 11210 26444
rect 12345 26435 12403 26441
rect 12345 26432 12357 26435
rect 11204 26404 12357 26432
rect 11204 26392 11210 26404
rect 12345 26401 12357 26404
rect 12391 26401 12403 26435
rect 12345 26395 12403 26401
rect 13446 26392 13452 26444
rect 13504 26432 13510 26444
rect 13541 26435 13599 26441
rect 13541 26432 13553 26435
rect 13504 26404 13553 26432
rect 13504 26392 13510 26404
rect 13541 26401 13553 26404
rect 13587 26401 13599 26435
rect 13541 26395 13599 26401
rect 14185 26435 14243 26441
rect 14185 26401 14197 26435
rect 14231 26432 14243 26435
rect 14642 26432 14648 26444
rect 14231 26404 14648 26432
rect 14231 26401 14243 26404
rect 14185 26395 14243 26401
rect 14642 26392 14648 26404
rect 14700 26392 14706 26444
rect 15010 26392 15016 26444
rect 15068 26392 15074 26444
rect 16132 26441 16160 26472
rect 16117 26435 16175 26441
rect 16117 26401 16129 26435
rect 16163 26401 16175 26435
rect 16117 26395 16175 26401
rect 16209 26435 16267 26441
rect 16209 26401 16221 26435
rect 16255 26432 16267 26435
rect 16669 26435 16727 26441
rect 16669 26432 16681 26435
rect 16255 26404 16681 26432
rect 16255 26401 16267 26404
rect 16209 26395 16267 26401
rect 16669 26401 16681 26404
rect 16715 26401 16727 26435
rect 16669 26395 16727 26401
rect 11238 26364 11244 26376
rect 11072 26336 11244 26364
rect 11238 26324 11244 26336
rect 11296 26324 11302 26376
rect 12253 26367 12311 26373
rect 12253 26333 12265 26367
rect 12299 26364 12311 26367
rect 12802 26364 12808 26376
rect 12299 26336 12808 26364
rect 12299 26333 12311 26336
rect 12253 26327 12311 26333
rect 12802 26324 12808 26336
rect 12860 26324 12866 26376
rect 14274 26324 14280 26376
rect 14332 26364 14338 26376
rect 16224 26364 16252 26395
rect 16960 26373 16988 26472
rect 24581 26469 24593 26503
rect 24627 26500 24639 26503
rect 24670 26500 24676 26512
rect 24627 26472 24676 26500
rect 24627 26469 24639 26472
rect 24581 26463 24639 26469
rect 24670 26460 24676 26472
rect 24728 26460 24734 26512
rect 18509 26435 18567 26441
rect 18509 26401 18521 26435
rect 18555 26432 18567 26435
rect 18874 26432 18880 26444
rect 18555 26404 18880 26432
rect 18555 26401 18567 26404
rect 18509 26395 18567 26401
rect 18874 26392 18880 26404
rect 18932 26392 18938 26444
rect 19429 26435 19487 26441
rect 19429 26401 19441 26435
rect 19475 26432 19487 26435
rect 20438 26432 20444 26444
rect 19475 26404 20444 26432
rect 19475 26401 19487 26404
rect 19429 26395 19487 26401
rect 20438 26392 20444 26404
rect 20496 26392 20502 26444
rect 20714 26392 20720 26444
rect 20772 26432 20778 26444
rect 21177 26435 21235 26441
rect 21177 26432 21189 26435
rect 20772 26404 21189 26432
rect 20772 26392 20778 26404
rect 21177 26401 21189 26404
rect 21223 26432 21235 26435
rect 21266 26432 21272 26444
rect 21223 26404 21272 26432
rect 21223 26401 21235 26404
rect 21177 26395 21235 26401
rect 21266 26392 21272 26404
rect 21324 26392 21330 26444
rect 21542 26392 21548 26444
rect 21600 26432 21606 26444
rect 23201 26435 23259 26441
rect 23201 26432 23213 26435
rect 21600 26404 23213 26432
rect 21600 26392 21606 26404
rect 23201 26401 23213 26404
rect 23247 26401 23259 26435
rect 23201 26395 23259 26401
rect 25038 26392 25044 26444
rect 25096 26392 25102 26444
rect 25130 26392 25136 26444
rect 25188 26392 25194 26444
rect 14332 26336 16252 26364
rect 16945 26367 17003 26373
rect 14332 26324 14338 26336
rect 16945 26333 16957 26367
rect 16991 26364 17003 26367
rect 17954 26364 17960 26376
rect 16991 26336 17960 26364
rect 16991 26333 17003 26336
rect 16945 26327 17003 26333
rect 17954 26324 17960 26336
rect 18012 26324 18018 26376
rect 18233 26367 18291 26373
rect 18233 26333 18245 26367
rect 18279 26364 18291 26367
rect 18322 26364 18328 26376
rect 18279 26336 18328 26364
rect 18279 26333 18291 26336
rect 18233 26327 18291 26333
rect 18322 26324 18328 26336
rect 18380 26324 18386 26376
rect 20990 26324 20996 26376
rect 21048 26364 21054 26376
rect 23109 26367 23167 26373
rect 21048 26336 23060 26364
rect 21048 26324 21054 26336
rect 10134 26256 10140 26308
rect 10192 26256 10198 26308
rect 10686 26256 10692 26308
rect 10744 26296 10750 26308
rect 12161 26299 12219 26305
rect 12161 26296 12173 26299
rect 10744 26268 12173 26296
rect 10744 26256 10750 26268
rect 12161 26265 12173 26268
rect 12207 26265 12219 26299
rect 12161 26259 12219 26265
rect 12526 26256 12532 26308
rect 12584 26296 12590 26308
rect 13357 26299 13415 26305
rect 13357 26296 13369 26299
rect 12584 26268 13369 26296
rect 12584 26256 12590 26268
rect 13357 26265 13369 26268
rect 13403 26265 13415 26299
rect 13357 26259 13415 26265
rect 13449 26299 13507 26305
rect 13449 26265 13461 26299
rect 13495 26296 13507 26299
rect 13630 26296 13636 26308
rect 13495 26268 13636 26296
rect 13495 26265 13507 26268
rect 13449 26259 13507 26265
rect 13630 26256 13636 26268
rect 13688 26256 13694 26308
rect 14826 26256 14832 26308
rect 14884 26256 14890 26308
rect 14921 26299 14979 26305
rect 14921 26265 14933 26299
rect 14967 26296 14979 26299
rect 16574 26296 16580 26308
rect 14967 26268 16580 26296
rect 14967 26265 14979 26268
rect 14921 26259 14979 26265
rect 16574 26256 16580 26268
rect 16632 26256 16638 26308
rect 19978 26296 19984 26308
rect 18340 26268 19984 26296
rect 14458 26188 14464 26240
rect 14516 26188 14522 26240
rect 16022 26188 16028 26240
rect 16080 26188 16086 26240
rect 16666 26188 16672 26240
rect 16724 26228 16730 26240
rect 18340 26237 18368 26268
rect 19978 26256 19984 26268
rect 20036 26256 20042 26308
rect 20930 26268 21588 26296
rect 21560 26237 21588 26268
rect 21910 26256 21916 26308
rect 21968 26256 21974 26308
rect 22097 26299 22155 26305
rect 22097 26265 22109 26299
rect 22143 26296 22155 26299
rect 22370 26296 22376 26308
rect 22143 26268 22376 26296
rect 22143 26265 22155 26268
rect 22097 26259 22155 26265
rect 22370 26256 22376 26268
rect 22428 26256 22434 26308
rect 23032 26296 23060 26336
rect 23109 26333 23121 26367
rect 23155 26364 23167 26367
rect 25314 26364 25320 26376
rect 23155 26336 25320 26364
rect 23155 26333 23167 26336
rect 23109 26327 23167 26333
rect 25314 26324 25320 26336
rect 25372 26324 25378 26376
rect 22480 26268 22968 26296
rect 23032 26268 23796 26296
rect 17865 26231 17923 26237
rect 17865 26228 17877 26231
rect 16724 26200 17877 26228
rect 16724 26188 16730 26200
rect 17865 26197 17877 26200
rect 17911 26197 17923 26231
rect 17865 26191 17923 26197
rect 18325 26231 18383 26237
rect 18325 26197 18337 26231
rect 18371 26197 18383 26231
rect 18325 26191 18383 26197
rect 21545 26231 21603 26237
rect 21545 26197 21557 26231
rect 21591 26228 21603 26231
rect 21634 26228 21640 26240
rect 21591 26200 21640 26228
rect 21591 26197 21603 26200
rect 21545 26191 21603 26197
rect 21634 26188 21640 26200
rect 21692 26188 21698 26240
rect 22186 26188 22192 26240
rect 22244 26228 22250 26240
rect 22480 26228 22508 26268
rect 22244 26200 22508 26228
rect 22244 26188 22250 26200
rect 22554 26188 22560 26240
rect 22612 26228 22618 26240
rect 22649 26231 22707 26237
rect 22649 26228 22661 26231
rect 22612 26200 22661 26228
rect 22612 26188 22618 26200
rect 22649 26197 22661 26200
rect 22695 26197 22707 26231
rect 22940 26228 22968 26268
rect 23014 26228 23020 26240
rect 22940 26200 23020 26228
rect 22649 26191 22707 26197
rect 23014 26188 23020 26200
rect 23072 26188 23078 26240
rect 23768 26228 23796 26268
rect 23842 26256 23848 26308
rect 23900 26256 23906 26308
rect 25038 26296 25044 26308
rect 23952 26268 25044 26296
rect 23952 26228 23980 26268
rect 25038 26256 25044 26268
rect 25096 26256 25102 26308
rect 25406 26296 25412 26308
rect 25148 26268 25412 26296
rect 23768 26200 23980 26228
rect 24949 26231 25007 26237
rect 24949 26197 24961 26231
rect 24995 26228 25007 26231
rect 25148 26228 25176 26268
rect 25406 26256 25412 26268
rect 25464 26256 25470 26308
rect 24995 26200 25176 26228
rect 24995 26197 25007 26200
rect 24949 26191 25007 26197
rect 1104 26138 25852 26160
rect 1104 26086 7950 26138
rect 8002 26086 8014 26138
rect 8066 26086 8078 26138
rect 8130 26086 8142 26138
rect 8194 26086 8206 26138
rect 8258 26086 17950 26138
rect 18002 26086 18014 26138
rect 18066 26086 18078 26138
rect 18130 26086 18142 26138
rect 18194 26086 18206 26138
rect 18258 26086 25852 26138
rect 1104 26064 25852 26086
rect 12894 25984 12900 26036
rect 12952 26024 12958 26036
rect 15749 26027 15807 26033
rect 12952 25996 15056 26024
rect 12952 25984 12958 25996
rect 12710 25916 12716 25968
rect 12768 25956 12774 25968
rect 12768 25928 13110 25956
rect 12768 25916 12774 25928
rect 10505 25891 10563 25897
rect 10505 25857 10517 25891
rect 10551 25888 10563 25891
rect 11514 25888 11520 25900
rect 10551 25860 11520 25888
rect 10551 25857 10563 25860
rect 10505 25851 10563 25857
rect 11514 25848 11520 25860
rect 11572 25848 11578 25900
rect 12342 25848 12348 25900
rect 12400 25848 12406 25900
rect 14921 25891 14979 25897
rect 14921 25857 14933 25891
rect 14967 25857 14979 25891
rect 15028 25888 15056 25996
rect 15749 25993 15761 26027
rect 15795 26024 15807 26027
rect 16022 26024 16028 26036
rect 15795 25996 16028 26024
rect 15795 25993 15807 25996
rect 15749 25987 15807 25993
rect 16022 25984 16028 25996
rect 16080 25984 16086 26036
rect 16114 25984 16120 26036
rect 16172 26024 16178 26036
rect 16209 26027 16267 26033
rect 16209 26024 16221 26027
rect 16172 25996 16221 26024
rect 16172 25984 16178 25996
rect 16209 25993 16221 25996
rect 16255 25993 16267 26027
rect 16209 25987 16267 25993
rect 18233 26027 18291 26033
rect 18233 25993 18245 26027
rect 18279 26024 18291 26027
rect 18322 26024 18328 26036
rect 18279 25996 18328 26024
rect 18279 25993 18291 25996
rect 18233 25987 18291 25993
rect 18322 25984 18328 25996
rect 18380 25984 18386 26036
rect 20070 25984 20076 26036
rect 20128 26024 20134 26036
rect 20165 26027 20223 26033
rect 20165 26024 20177 26027
rect 20128 25996 20177 26024
rect 20128 25984 20134 25996
rect 20165 25993 20177 25996
rect 20211 25993 20223 26027
rect 20165 25987 20223 25993
rect 22465 26027 22523 26033
rect 22465 25993 22477 26027
rect 22511 26024 22523 26027
rect 23750 26024 23756 26036
rect 22511 25996 23756 26024
rect 22511 25993 22523 25996
rect 22465 25987 22523 25993
rect 23750 25984 23756 25996
rect 23808 25984 23814 26036
rect 24762 25984 24768 26036
rect 24820 26024 24826 26036
rect 25317 26027 25375 26033
rect 25317 26024 25329 26027
rect 24820 25996 25329 26024
rect 24820 25984 24826 25996
rect 25317 25993 25329 25996
rect 25363 25993 25375 26027
rect 25317 25987 25375 25993
rect 15102 25916 15108 25968
rect 15160 25956 15166 25968
rect 21453 25959 21511 25965
rect 15160 25928 17816 25956
rect 15160 25916 15166 25928
rect 17788 25897 17816 25928
rect 21453 25925 21465 25959
rect 21499 25956 21511 25959
rect 23845 25959 23903 25965
rect 23845 25956 23857 25959
rect 21499 25928 23857 25956
rect 21499 25925 21511 25928
rect 21453 25919 21511 25925
rect 23845 25925 23857 25928
rect 23891 25925 23903 25959
rect 23845 25919 23903 25925
rect 24118 25916 24124 25968
rect 24176 25956 24182 25968
rect 24302 25956 24308 25968
rect 24176 25928 24308 25956
rect 24176 25916 24182 25928
rect 24302 25916 24308 25928
rect 24360 25916 24366 25968
rect 17129 25891 17187 25897
rect 17129 25888 17141 25891
rect 15028 25860 17141 25888
rect 14921 25851 14979 25857
rect 17129 25857 17141 25860
rect 17175 25857 17187 25891
rect 17129 25851 17187 25857
rect 17773 25891 17831 25897
rect 17773 25857 17785 25891
rect 17819 25857 17831 25891
rect 17773 25851 17831 25857
rect 19521 25891 19579 25897
rect 19521 25857 19533 25891
rect 19567 25888 19579 25891
rect 20714 25888 20720 25900
rect 19567 25860 20720 25888
rect 19567 25857 19579 25860
rect 19521 25851 19579 25857
rect 12618 25780 12624 25832
rect 12676 25780 12682 25832
rect 12710 25780 12716 25832
rect 12768 25820 12774 25832
rect 13998 25820 14004 25832
rect 12768 25792 14004 25820
rect 12768 25780 12774 25792
rect 13998 25780 14004 25792
rect 14056 25780 14062 25832
rect 14553 25755 14611 25761
rect 14553 25752 14565 25755
rect 13648 25724 14565 25752
rect 11146 25644 11152 25696
rect 11204 25644 11210 25696
rect 11698 25644 11704 25696
rect 11756 25684 11762 25696
rect 13648 25684 13676 25724
rect 14553 25721 14565 25724
rect 14599 25721 14611 25755
rect 14936 25752 14964 25851
rect 20714 25848 20720 25860
rect 20772 25848 20778 25900
rect 20806 25848 20812 25900
rect 20864 25848 20870 25900
rect 22186 25848 22192 25900
rect 22244 25888 22250 25900
rect 22373 25891 22431 25897
rect 22373 25888 22385 25891
rect 22244 25860 22385 25888
rect 22244 25848 22250 25860
rect 22373 25857 22385 25860
rect 22419 25888 22431 25891
rect 23201 25891 23259 25897
rect 23201 25888 23213 25891
rect 22419 25860 23213 25888
rect 22419 25857 22431 25860
rect 22373 25851 22431 25857
rect 23201 25857 23213 25860
rect 23247 25857 23259 25891
rect 23201 25851 23259 25857
rect 15010 25780 15016 25832
rect 15068 25780 15074 25832
rect 15102 25780 15108 25832
rect 15160 25780 15166 25832
rect 18874 25780 18880 25832
rect 18932 25780 18938 25832
rect 22462 25780 22468 25832
rect 22520 25820 22526 25832
rect 22557 25823 22615 25829
rect 22557 25820 22569 25823
rect 22520 25792 22569 25820
rect 22520 25780 22526 25792
rect 22557 25789 22569 25792
rect 22603 25789 22615 25823
rect 22557 25783 22615 25789
rect 23014 25780 23020 25832
rect 23072 25780 23078 25832
rect 15838 25752 15844 25764
rect 14936 25724 15844 25752
rect 14553 25715 14611 25721
rect 15838 25712 15844 25724
rect 15896 25752 15902 25764
rect 16945 25755 17003 25761
rect 15896 25724 16528 25752
rect 15896 25712 15902 25724
rect 16500 25696 16528 25724
rect 16945 25721 16957 25755
rect 16991 25752 17003 25755
rect 21910 25752 21916 25764
rect 16991 25724 21916 25752
rect 16991 25721 17003 25724
rect 16945 25715 17003 25721
rect 21910 25712 21916 25724
rect 21968 25712 21974 25764
rect 11756 25656 13676 25684
rect 11756 25644 11762 25656
rect 14090 25644 14096 25696
rect 14148 25644 14154 25696
rect 15010 25644 15016 25696
rect 15068 25684 15074 25696
rect 16114 25684 16120 25696
rect 15068 25656 16120 25684
rect 15068 25644 15074 25656
rect 16114 25644 16120 25656
rect 16172 25644 16178 25696
rect 16482 25644 16488 25696
rect 16540 25644 16546 25696
rect 17589 25687 17647 25693
rect 17589 25653 17601 25687
rect 17635 25684 17647 25687
rect 18966 25684 18972 25696
rect 17635 25656 18972 25684
rect 17635 25653 17647 25656
rect 17589 25647 17647 25653
rect 18966 25644 18972 25656
rect 19024 25644 19030 25696
rect 20533 25687 20591 25693
rect 20533 25653 20545 25687
rect 20579 25684 20591 25687
rect 21634 25684 21640 25696
rect 20579 25656 21640 25684
rect 20579 25653 20591 25656
rect 20533 25647 20591 25653
rect 21634 25644 21640 25656
rect 21692 25644 21698 25696
rect 22002 25644 22008 25696
rect 22060 25644 22066 25696
rect 23032 25684 23060 25780
rect 23216 25752 23244 25851
rect 23290 25780 23296 25832
rect 23348 25820 23354 25832
rect 23566 25820 23572 25832
rect 23348 25792 23572 25820
rect 23348 25780 23354 25792
rect 23566 25780 23572 25792
rect 23624 25780 23630 25832
rect 24578 25820 24584 25832
rect 23676 25792 24584 25820
rect 23676 25752 23704 25792
rect 24578 25780 24584 25792
rect 24636 25780 24642 25832
rect 23216 25724 23704 25752
rect 23934 25684 23940 25696
rect 23032 25656 23940 25684
rect 23934 25644 23940 25656
rect 23992 25644 23998 25696
rect 1104 25594 25852 25616
rect 1104 25542 2950 25594
rect 3002 25542 3014 25594
rect 3066 25542 3078 25594
rect 3130 25542 3142 25594
rect 3194 25542 3206 25594
rect 3258 25542 12950 25594
rect 13002 25542 13014 25594
rect 13066 25542 13078 25594
rect 13130 25542 13142 25594
rect 13194 25542 13206 25594
rect 13258 25542 22950 25594
rect 23002 25542 23014 25594
rect 23066 25542 23078 25594
rect 23130 25542 23142 25594
rect 23194 25542 23206 25594
rect 23258 25542 25852 25594
rect 1104 25520 25852 25542
rect 10318 25440 10324 25492
rect 10376 25440 10382 25492
rect 12618 25440 12624 25492
rect 12676 25480 12682 25492
rect 13725 25483 13783 25489
rect 13725 25480 13737 25483
rect 12676 25452 13737 25480
rect 12676 25440 12682 25452
rect 13725 25449 13737 25452
rect 13771 25449 13783 25483
rect 13725 25443 13783 25449
rect 25222 25440 25228 25492
rect 25280 25440 25286 25492
rect 11517 25415 11575 25421
rect 11517 25381 11529 25415
rect 11563 25412 11575 25415
rect 11563 25384 18092 25412
rect 11563 25381 11575 25384
rect 11517 25375 11575 25381
rect 9582 25304 9588 25356
rect 9640 25344 9646 25356
rect 10873 25347 10931 25353
rect 10873 25344 10885 25347
rect 9640 25316 10885 25344
rect 9640 25304 9646 25316
rect 10873 25313 10885 25316
rect 10919 25313 10931 25347
rect 10873 25307 10931 25313
rect 12066 25304 12072 25356
rect 12124 25304 12130 25356
rect 12710 25344 12716 25356
rect 12176 25316 12716 25344
rect 10689 25279 10747 25285
rect 10689 25245 10701 25279
rect 10735 25276 10747 25279
rect 12176 25276 12204 25316
rect 12710 25304 12716 25316
rect 12768 25304 12774 25356
rect 14829 25347 14887 25353
rect 14829 25344 14841 25347
rect 13004 25316 14841 25344
rect 10735 25248 12204 25276
rect 10735 25245 10747 25248
rect 10689 25239 10747 25245
rect 12250 25236 12256 25288
rect 12308 25276 12314 25288
rect 13004 25276 13032 25316
rect 14829 25313 14841 25316
rect 14875 25344 14887 25347
rect 15102 25344 15108 25356
rect 14875 25316 15108 25344
rect 14875 25313 14887 25316
rect 14829 25307 14887 25313
rect 15102 25304 15108 25316
rect 15160 25304 15166 25356
rect 12308 25248 13032 25276
rect 13081 25279 13139 25285
rect 12308 25236 12314 25248
rect 13081 25245 13093 25279
rect 13127 25276 13139 25279
rect 13446 25276 13452 25288
rect 13127 25248 13452 25276
rect 13127 25245 13139 25248
rect 13081 25239 13139 25245
rect 13446 25236 13452 25248
rect 13504 25236 13510 25288
rect 17310 25236 17316 25288
rect 17368 25236 17374 25288
rect 18064 25285 18092 25384
rect 18877 25347 18935 25353
rect 18877 25313 18889 25347
rect 18923 25344 18935 25347
rect 18923 25316 22094 25344
rect 18923 25313 18935 25316
rect 18877 25307 18935 25313
rect 18049 25279 18107 25285
rect 18049 25245 18061 25279
rect 18095 25245 18107 25279
rect 18049 25239 18107 25245
rect 18156 25248 19380 25276
rect 11977 25211 12035 25217
rect 11977 25177 11989 25211
rect 12023 25208 12035 25211
rect 12158 25208 12164 25220
rect 12023 25180 12164 25208
rect 12023 25177 12035 25180
rect 11977 25171 12035 25177
rect 12158 25168 12164 25180
rect 12216 25168 12222 25220
rect 14645 25211 14703 25217
rect 13372 25180 14320 25208
rect 10318 25100 10324 25152
rect 10376 25140 10382 25152
rect 10781 25143 10839 25149
rect 10781 25140 10793 25143
rect 10376 25112 10793 25140
rect 10376 25100 10382 25112
rect 10781 25109 10793 25112
rect 10827 25109 10839 25143
rect 10781 25103 10839 25109
rect 11054 25100 11060 25152
rect 11112 25140 11118 25152
rect 11885 25143 11943 25149
rect 11885 25140 11897 25143
rect 11112 25112 11897 25140
rect 11112 25100 11118 25112
rect 11885 25109 11897 25112
rect 11931 25109 11943 25143
rect 11885 25103 11943 25109
rect 12066 25100 12072 25152
rect 12124 25140 12130 25152
rect 13372 25140 13400 25180
rect 14292 25149 14320 25180
rect 14645 25177 14657 25211
rect 14691 25208 14703 25211
rect 15657 25211 15715 25217
rect 14691 25180 15424 25208
rect 14691 25177 14703 25180
rect 14645 25171 14703 25177
rect 15396 25152 15424 25180
rect 15657 25177 15669 25211
rect 15703 25208 15715 25211
rect 18156 25208 18184 25248
rect 15703 25180 18184 25208
rect 18693 25211 18751 25217
rect 15703 25177 15715 25180
rect 15657 25171 15715 25177
rect 18693 25177 18705 25211
rect 18739 25177 18751 25211
rect 18693 25171 18751 25177
rect 12124 25112 13400 25140
rect 14277 25143 14335 25149
rect 12124 25100 12130 25112
rect 14277 25109 14289 25143
rect 14323 25109 14335 25143
rect 14277 25103 14335 25109
rect 14737 25143 14795 25149
rect 14737 25109 14749 25143
rect 14783 25140 14795 25143
rect 15286 25140 15292 25152
rect 14783 25112 15292 25140
rect 14783 25109 14795 25112
rect 14737 25103 14795 25109
rect 15286 25100 15292 25112
rect 15344 25100 15350 25152
rect 15378 25100 15384 25152
rect 15436 25100 15442 25152
rect 17865 25143 17923 25149
rect 17865 25109 17877 25143
rect 17911 25140 17923 25143
rect 18708 25140 18736 25171
rect 19352 25152 19380 25248
rect 19702 25236 19708 25288
rect 19760 25236 19766 25288
rect 20901 25279 20959 25285
rect 20901 25245 20913 25279
rect 20947 25276 20959 25279
rect 21082 25276 21088 25288
rect 20947 25248 21088 25276
rect 20947 25245 20959 25248
rect 20901 25239 20959 25245
rect 21082 25236 21088 25248
rect 21140 25276 21146 25288
rect 21450 25276 21456 25288
rect 21140 25248 21456 25276
rect 21140 25236 21146 25248
rect 21450 25236 21456 25248
rect 21508 25236 21514 25288
rect 21542 25236 21548 25288
rect 21600 25236 21606 25288
rect 22066 25276 22094 25316
rect 22649 25279 22707 25285
rect 22649 25276 22661 25279
rect 22066 25248 22661 25276
rect 22649 25245 22661 25248
rect 22695 25245 22707 25279
rect 22649 25239 22707 25245
rect 24581 25279 24639 25285
rect 24581 25245 24593 25279
rect 24627 25276 24639 25279
rect 24762 25276 24768 25288
rect 24627 25248 24768 25276
rect 24627 25245 24639 25248
rect 24581 25239 24639 25245
rect 24762 25236 24768 25248
rect 24820 25236 24826 25288
rect 23845 25211 23903 25217
rect 23845 25177 23857 25211
rect 23891 25208 23903 25211
rect 24946 25208 24952 25220
rect 23891 25180 24952 25208
rect 23891 25177 23903 25180
rect 23845 25171 23903 25177
rect 24946 25168 24952 25180
rect 25004 25168 25010 25220
rect 17911 25112 18736 25140
rect 17911 25109 17923 25112
rect 17865 25103 17923 25109
rect 19334 25100 19340 25152
rect 19392 25100 19398 25152
rect 19978 25100 19984 25152
rect 20036 25140 20042 25152
rect 20349 25143 20407 25149
rect 20349 25140 20361 25143
rect 20036 25112 20361 25140
rect 20036 25100 20042 25112
rect 20349 25109 20361 25112
rect 20395 25109 20407 25143
rect 20349 25103 20407 25109
rect 20990 25100 20996 25152
rect 21048 25100 21054 25152
rect 22186 25100 22192 25152
rect 22244 25100 22250 25152
rect 1104 25050 25852 25072
rect 1104 24998 7950 25050
rect 8002 24998 8014 25050
rect 8066 24998 8078 25050
rect 8130 24998 8142 25050
rect 8194 24998 8206 25050
rect 8258 24998 17950 25050
rect 18002 24998 18014 25050
rect 18066 24998 18078 25050
rect 18130 24998 18142 25050
rect 18194 24998 18206 25050
rect 18258 24998 25852 25050
rect 1104 24976 25852 24998
rect 10870 24896 10876 24948
rect 10928 24936 10934 24948
rect 12250 24936 12256 24948
rect 10928 24908 12256 24936
rect 10928 24896 10934 24908
rect 12250 24896 12256 24908
rect 12308 24896 12314 24948
rect 14277 24939 14335 24945
rect 14277 24905 14289 24939
rect 14323 24936 14335 24939
rect 15470 24936 15476 24948
rect 14323 24908 15476 24936
rect 14323 24905 14335 24908
rect 14277 24899 14335 24905
rect 15470 24896 15476 24908
rect 15528 24896 15534 24948
rect 15933 24939 15991 24945
rect 15933 24905 15945 24939
rect 15979 24936 15991 24939
rect 16390 24936 16396 24948
rect 15979 24908 16396 24936
rect 15979 24905 15991 24908
rect 15933 24899 15991 24905
rect 16390 24896 16396 24908
rect 16448 24936 16454 24948
rect 17402 24936 17408 24948
rect 16448 24908 17408 24936
rect 16448 24896 16454 24908
rect 17402 24896 17408 24908
rect 17460 24936 17466 24948
rect 18417 24939 18475 24945
rect 18417 24936 18429 24939
rect 17460 24908 18429 24936
rect 17460 24896 17466 24908
rect 18417 24905 18429 24908
rect 18463 24936 18475 24939
rect 19245 24939 19303 24945
rect 19245 24936 19257 24939
rect 18463 24908 19257 24936
rect 18463 24905 18475 24908
rect 18417 24899 18475 24905
rect 19245 24905 19257 24908
rect 19291 24936 19303 24939
rect 20162 24936 20168 24948
rect 19291 24908 20168 24936
rect 19291 24905 19303 24908
rect 19245 24899 19303 24905
rect 20162 24896 20168 24908
rect 20220 24896 20226 24948
rect 20806 24896 20812 24948
rect 20864 24936 20870 24948
rect 25317 24939 25375 24945
rect 25317 24936 25329 24939
rect 20864 24908 25329 24936
rect 20864 24896 20870 24908
rect 25317 24905 25329 24908
rect 25363 24936 25375 24939
rect 25406 24936 25412 24948
rect 25363 24908 25412 24936
rect 25363 24905 25375 24908
rect 25317 24899 25375 24905
rect 25406 24896 25412 24908
rect 25464 24896 25470 24948
rect 8389 24871 8447 24877
rect 8389 24837 8401 24871
rect 8435 24868 8447 24871
rect 9766 24868 9772 24880
rect 8435 24840 9772 24868
rect 8435 24837 8447 24840
rect 8389 24831 8447 24837
rect 9766 24828 9772 24840
rect 9824 24828 9830 24880
rect 11146 24828 11152 24880
rect 11204 24868 11210 24880
rect 11977 24871 12035 24877
rect 11977 24868 11989 24871
rect 11204 24840 11989 24868
rect 11204 24828 11210 24840
rect 11977 24837 11989 24840
rect 12023 24837 12035 24871
rect 11977 24831 12035 24837
rect 12710 24828 12716 24880
rect 12768 24828 12774 24880
rect 17126 24828 17132 24880
rect 17184 24868 17190 24880
rect 17221 24871 17279 24877
rect 17221 24868 17233 24871
rect 17184 24840 17233 24868
rect 17184 24828 17190 24840
rect 17221 24837 17233 24840
rect 17267 24837 17279 24871
rect 17221 24831 17279 24837
rect 11238 24800 11244 24812
rect 10626 24772 11244 24800
rect 11238 24760 11244 24772
rect 11296 24760 11302 24812
rect 14366 24760 14372 24812
rect 14424 24760 14430 24812
rect 15286 24760 15292 24812
rect 15344 24800 15350 24812
rect 17236 24800 17264 24831
rect 19978 24828 19984 24880
rect 20036 24828 20042 24880
rect 21266 24828 21272 24880
rect 21324 24868 21330 24880
rect 22465 24871 22523 24877
rect 22465 24868 22477 24871
rect 21324 24840 22477 24868
rect 21324 24828 21330 24840
rect 22465 24837 22477 24840
rect 22511 24837 22523 24871
rect 22465 24831 22523 24837
rect 24118 24828 24124 24880
rect 24176 24868 24182 24880
rect 24176 24840 24334 24868
rect 24176 24828 24182 24840
rect 18782 24800 18788 24812
rect 15344 24772 16896 24800
rect 17236 24772 18788 24800
rect 15344 24760 15350 24772
rect 16868 24744 16896 24772
rect 18782 24760 18788 24772
rect 18840 24760 18846 24812
rect 21634 24800 21640 24812
rect 21114 24772 21640 24800
rect 21634 24760 21640 24772
rect 21692 24760 21698 24812
rect 22557 24803 22615 24809
rect 22557 24769 22569 24803
rect 22603 24800 22615 24803
rect 23474 24800 23480 24812
rect 22603 24772 23480 24800
rect 22603 24769 22615 24772
rect 22557 24763 22615 24769
rect 23474 24760 23480 24772
rect 23532 24760 23538 24812
rect 8481 24735 8539 24741
rect 8481 24732 8493 24735
rect 8404 24704 8493 24732
rect 8404 24676 8432 24704
rect 8481 24701 8493 24704
rect 8527 24701 8539 24735
rect 8481 24695 8539 24701
rect 8570 24692 8576 24744
rect 8628 24692 8634 24744
rect 9217 24735 9275 24741
rect 9217 24701 9229 24735
rect 9263 24701 9275 24735
rect 9217 24695 9275 24701
rect 9493 24735 9551 24741
rect 9493 24701 9505 24735
rect 9539 24732 9551 24735
rect 10962 24732 10968 24744
rect 9539 24704 10968 24732
rect 9539 24701 9551 24704
rect 9493 24695 9551 24701
rect 8386 24624 8392 24676
rect 8444 24624 8450 24676
rect 8021 24599 8079 24605
rect 8021 24565 8033 24599
rect 8067 24596 8079 24599
rect 9122 24596 9128 24608
rect 8067 24568 9128 24596
rect 8067 24565 8079 24568
rect 8021 24559 8079 24565
rect 9122 24556 9128 24568
rect 9180 24556 9186 24608
rect 9232 24596 9260 24695
rect 10962 24692 10968 24704
rect 11020 24692 11026 24744
rect 11146 24692 11152 24744
rect 11204 24732 11210 24744
rect 11701 24735 11759 24741
rect 11701 24732 11713 24735
rect 11204 24704 11713 24732
rect 11204 24692 11210 24704
rect 11701 24701 11713 24704
rect 11747 24701 11759 24735
rect 11701 24695 11759 24701
rect 12342 24692 12348 24744
rect 12400 24732 12406 24744
rect 14461 24735 14519 24741
rect 12400 24704 13492 24732
rect 12400 24692 12406 24704
rect 11164 24664 11192 24692
rect 10520 24636 11192 24664
rect 13464 24664 13492 24704
rect 14461 24701 14473 24735
rect 14507 24701 14519 24735
rect 14461 24695 14519 24701
rect 14476 24664 14504 24695
rect 16022 24692 16028 24744
rect 16080 24692 16086 24744
rect 16117 24735 16175 24741
rect 16117 24701 16129 24735
rect 16163 24701 16175 24735
rect 16117 24695 16175 24701
rect 16132 24664 16160 24695
rect 16850 24692 16856 24744
rect 16908 24732 16914 24744
rect 17313 24735 17371 24741
rect 17313 24732 17325 24735
rect 16908 24704 17325 24732
rect 16908 24692 16914 24704
rect 13464 24636 14504 24664
rect 14568 24636 16160 24664
rect 10520 24596 10548 24636
rect 9232 24568 10548 24596
rect 10870 24556 10876 24608
rect 10928 24596 10934 24608
rect 10965 24599 11023 24605
rect 10965 24596 10977 24599
rect 10928 24568 10977 24596
rect 10928 24556 10934 24568
rect 10965 24565 10977 24568
rect 11011 24565 11023 24599
rect 10965 24559 11023 24565
rect 13446 24556 13452 24608
rect 13504 24556 13510 24608
rect 13538 24556 13544 24608
rect 13596 24596 13602 24608
rect 13909 24599 13967 24605
rect 13909 24596 13921 24599
rect 13596 24568 13921 24596
rect 13596 24556 13602 24568
rect 13909 24565 13921 24568
rect 13955 24565 13967 24599
rect 13909 24559 13967 24565
rect 13998 24556 14004 24608
rect 14056 24596 14062 24608
rect 14568 24596 14596 24636
rect 14056 24568 14596 24596
rect 14056 24556 14062 24568
rect 15378 24556 15384 24608
rect 15436 24596 15442 24608
rect 15565 24599 15623 24605
rect 15565 24596 15577 24599
rect 15436 24568 15577 24596
rect 15436 24556 15442 24568
rect 15565 24565 15577 24568
rect 15611 24565 15623 24599
rect 15565 24559 15623 24565
rect 15838 24556 15844 24608
rect 15896 24596 15902 24608
rect 16853 24599 16911 24605
rect 16853 24596 16865 24599
rect 15896 24568 16865 24596
rect 15896 24556 15902 24568
rect 16853 24565 16865 24568
rect 16899 24565 16911 24599
rect 16960 24596 16988 24704
rect 17313 24701 17325 24704
rect 17359 24701 17371 24735
rect 17313 24695 17371 24701
rect 17402 24692 17408 24744
rect 17460 24692 17466 24744
rect 18506 24692 18512 24744
rect 18564 24692 18570 24744
rect 18598 24692 18604 24744
rect 18656 24692 18662 24744
rect 19426 24692 19432 24744
rect 19484 24732 19490 24744
rect 19705 24735 19763 24741
rect 19705 24732 19717 24735
rect 19484 24704 19717 24732
rect 19484 24692 19490 24704
rect 19705 24701 19717 24704
rect 19751 24701 19763 24735
rect 19705 24695 19763 24701
rect 21453 24735 21511 24741
rect 21453 24701 21465 24735
rect 21499 24732 21511 24735
rect 21542 24732 21548 24744
rect 21499 24704 21548 24732
rect 21499 24701 21511 24704
rect 21453 24695 21511 24701
rect 21542 24692 21548 24704
rect 21600 24692 21606 24744
rect 22741 24735 22799 24741
rect 22741 24701 22753 24735
rect 22787 24701 22799 24735
rect 22741 24695 22799 24701
rect 17034 24624 17040 24676
rect 17092 24664 17098 24676
rect 17092 24636 19380 24664
rect 17092 24624 17098 24636
rect 17770 24596 17776 24608
rect 16960 24568 17776 24596
rect 16853 24559 16911 24565
rect 17770 24556 17776 24568
rect 17828 24556 17834 24608
rect 17862 24556 17868 24608
rect 17920 24596 17926 24608
rect 18049 24599 18107 24605
rect 18049 24596 18061 24599
rect 17920 24568 18061 24596
rect 17920 24556 17926 24568
rect 18049 24565 18061 24568
rect 18095 24565 18107 24599
rect 18049 24559 18107 24565
rect 18782 24556 18788 24608
rect 18840 24596 18846 24608
rect 19061 24599 19119 24605
rect 19061 24596 19073 24599
rect 18840 24568 19073 24596
rect 18840 24556 18846 24568
rect 19061 24565 19073 24568
rect 19107 24565 19119 24599
rect 19352 24596 19380 24636
rect 21634 24624 21640 24676
rect 21692 24664 21698 24676
rect 22756 24664 22784 24695
rect 23290 24692 23296 24744
rect 23348 24732 23354 24744
rect 23566 24732 23572 24744
rect 23348 24704 23572 24732
rect 23348 24692 23354 24704
rect 23566 24692 23572 24704
rect 23624 24692 23630 24744
rect 23845 24735 23903 24741
rect 23845 24701 23857 24735
rect 23891 24732 23903 24735
rect 25314 24732 25320 24744
rect 23891 24704 25320 24732
rect 23891 24701 23903 24704
rect 23845 24695 23903 24701
rect 25314 24692 25320 24704
rect 25372 24692 25378 24744
rect 21692 24636 22508 24664
rect 22756 24636 23704 24664
rect 21692 24624 21698 24636
rect 21818 24596 21824 24608
rect 19352 24568 21824 24596
rect 19061 24559 19119 24565
rect 21818 24556 21824 24568
rect 21876 24556 21882 24608
rect 22094 24556 22100 24608
rect 22152 24556 22158 24608
rect 22480 24596 22508 24636
rect 23676 24608 23704 24636
rect 23201 24599 23259 24605
rect 23201 24596 23213 24599
rect 22480 24568 23213 24596
rect 23201 24565 23213 24568
rect 23247 24596 23259 24599
rect 23474 24596 23480 24608
rect 23247 24568 23480 24596
rect 23247 24565 23259 24568
rect 23201 24559 23259 24565
rect 23474 24556 23480 24568
rect 23532 24556 23538 24608
rect 23658 24556 23664 24608
rect 23716 24556 23722 24608
rect 1104 24506 25852 24528
rect 1104 24454 2950 24506
rect 3002 24454 3014 24506
rect 3066 24454 3078 24506
rect 3130 24454 3142 24506
rect 3194 24454 3206 24506
rect 3258 24454 12950 24506
rect 13002 24454 13014 24506
rect 13066 24454 13078 24506
rect 13130 24454 13142 24506
rect 13194 24454 13206 24506
rect 13258 24454 22950 24506
rect 23002 24454 23014 24506
rect 23066 24454 23078 24506
rect 23130 24454 23142 24506
rect 23194 24454 23206 24506
rect 23258 24454 25852 24506
rect 1104 24432 25852 24454
rect 8573 24395 8631 24401
rect 8573 24361 8585 24395
rect 8619 24392 8631 24395
rect 9398 24392 9404 24404
rect 8619 24364 9404 24392
rect 8619 24361 8631 24364
rect 8573 24355 8631 24361
rect 9398 24352 9404 24364
rect 9456 24352 9462 24404
rect 12342 24392 12348 24404
rect 9508 24364 12348 24392
rect 6825 24259 6883 24265
rect 6825 24225 6837 24259
rect 6871 24256 6883 24259
rect 7742 24256 7748 24268
rect 6871 24228 7748 24256
rect 6871 24225 6883 24228
rect 6825 24219 6883 24225
rect 7742 24216 7748 24228
rect 7800 24216 7806 24268
rect 9214 24148 9220 24200
rect 9272 24188 9278 24200
rect 9508 24197 9536 24364
rect 12342 24352 12348 24364
rect 12400 24352 12406 24404
rect 12710 24352 12716 24404
rect 12768 24392 12774 24404
rect 13725 24395 13783 24401
rect 13725 24392 13737 24395
rect 12768 24364 13737 24392
rect 12768 24352 12774 24364
rect 13725 24361 13737 24364
rect 13771 24392 13783 24395
rect 15010 24392 15016 24404
rect 13771 24364 15016 24392
rect 13771 24361 13783 24364
rect 13725 24355 13783 24361
rect 15010 24352 15016 24364
rect 15068 24352 15074 24404
rect 16390 24352 16396 24404
rect 16448 24352 16454 24404
rect 16853 24395 16911 24401
rect 16853 24361 16865 24395
rect 16899 24392 16911 24395
rect 19334 24392 19340 24404
rect 16899 24364 19340 24392
rect 16899 24361 16911 24364
rect 16853 24355 16911 24361
rect 19334 24352 19340 24364
rect 19392 24352 19398 24404
rect 19702 24352 19708 24404
rect 19760 24392 19766 24404
rect 20070 24392 20076 24404
rect 19760 24364 20076 24392
rect 19760 24352 19766 24364
rect 20070 24352 20076 24364
rect 20128 24392 20134 24404
rect 21177 24395 21235 24401
rect 21177 24392 21189 24395
rect 20128 24364 21189 24392
rect 20128 24352 20134 24364
rect 21177 24361 21189 24364
rect 21223 24361 21235 24395
rect 21177 24355 21235 24361
rect 21450 24352 21456 24404
rect 21508 24352 21514 24404
rect 16022 24284 16028 24336
rect 16080 24324 16086 24336
rect 16117 24327 16175 24333
rect 16117 24324 16129 24327
rect 16080 24296 16129 24324
rect 16080 24284 16086 24296
rect 16117 24293 16129 24296
rect 16163 24324 16175 24327
rect 18506 24324 18512 24336
rect 16163 24296 18512 24324
rect 16163 24293 16175 24296
rect 16117 24287 16175 24293
rect 18506 24284 18512 24296
rect 18564 24284 18570 24336
rect 18616 24296 19380 24324
rect 18616 24265 18644 24296
rect 10873 24259 10931 24265
rect 10873 24225 10885 24259
rect 10919 24256 10931 24259
rect 18601 24259 18659 24265
rect 10919 24228 12434 24256
rect 10919 24225 10931 24228
rect 10873 24219 10931 24225
rect 9493 24191 9551 24197
rect 9493 24188 9505 24191
rect 9272 24160 9505 24188
rect 9272 24148 9278 24160
rect 9493 24157 9505 24160
rect 9539 24157 9551 24191
rect 9493 24151 9551 24157
rect 10597 24191 10655 24197
rect 10597 24157 10609 24191
rect 10643 24157 10655 24191
rect 10597 24151 10655 24157
rect 7101 24123 7159 24129
rect 7101 24089 7113 24123
rect 7147 24089 7159 24123
rect 8938 24120 8944 24132
rect 8326 24092 8944 24120
rect 7101 24083 7159 24089
rect 7116 24052 7144 24083
rect 8938 24080 8944 24092
rect 8996 24080 9002 24132
rect 10502 24120 10508 24132
rect 9692 24092 10508 24120
rect 9692 24064 9720 24092
rect 10502 24080 10508 24092
rect 10560 24080 10566 24132
rect 9217 24055 9275 24061
rect 9217 24052 9229 24055
rect 7116 24024 9229 24052
rect 9217 24021 9229 24024
rect 9263 24052 9275 24055
rect 9674 24052 9680 24064
rect 9263 24024 9680 24052
rect 9263 24021 9275 24024
rect 9217 24015 9275 24021
rect 9674 24012 9680 24024
rect 9732 24012 9738 24064
rect 10134 24012 10140 24064
rect 10192 24012 10198 24064
rect 10612 24052 10640 24151
rect 11330 24080 11336 24132
rect 11388 24080 11394 24132
rect 12406 24120 12434 24228
rect 18601 24225 18613 24259
rect 18647 24225 18659 24259
rect 18601 24219 18659 24225
rect 18785 24259 18843 24265
rect 18785 24225 18797 24259
rect 18831 24256 18843 24259
rect 19242 24256 19248 24268
rect 18831 24228 19248 24256
rect 18831 24225 18843 24228
rect 18785 24219 18843 24225
rect 19242 24216 19248 24228
rect 19300 24216 19306 24268
rect 19352 24256 19380 24296
rect 23290 24284 23296 24336
rect 23348 24284 23354 24336
rect 23934 24284 23940 24336
rect 23992 24324 23998 24336
rect 24946 24324 24952 24336
rect 23992 24296 24952 24324
rect 23992 24284 23998 24296
rect 24946 24284 24952 24296
rect 25004 24284 25010 24336
rect 20898 24256 20904 24268
rect 19352 24228 20904 24256
rect 20898 24216 20904 24228
rect 20956 24216 20962 24268
rect 21913 24259 21971 24265
rect 21913 24225 21925 24259
rect 21959 24256 21971 24259
rect 23308 24256 23336 24284
rect 21959 24228 23336 24256
rect 21959 24225 21971 24228
rect 21913 24219 21971 24225
rect 23474 24216 23480 24268
rect 23532 24256 23538 24268
rect 24118 24256 24124 24268
rect 23532 24228 24124 24256
rect 23532 24216 23538 24228
rect 24118 24216 24124 24228
rect 24176 24216 24182 24268
rect 12805 24191 12863 24197
rect 12805 24157 12817 24191
rect 12851 24188 12863 24191
rect 14090 24188 14096 24200
rect 12851 24160 14096 24188
rect 12851 24157 12863 24160
rect 12805 24151 12863 24157
rect 14090 24148 14096 24160
rect 14148 24148 14154 24200
rect 16301 24191 16359 24197
rect 16301 24157 16313 24191
rect 16347 24188 16359 24191
rect 17034 24188 17040 24200
rect 16347 24160 17040 24188
rect 16347 24157 16359 24160
rect 16301 24151 16359 24157
rect 17034 24148 17040 24160
rect 17092 24148 17098 24200
rect 17681 24191 17739 24197
rect 17681 24157 17693 24191
rect 17727 24188 17739 24191
rect 18230 24188 18236 24200
rect 17727 24160 18236 24188
rect 17727 24157 17739 24160
rect 17681 24151 17739 24157
rect 18230 24148 18236 24160
rect 18288 24148 18294 24200
rect 18509 24191 18567 24197
rect 18509 24157 18521 24191
rect 18555 24188 18567 24191
rect 18874 24188 18880 24200
rect 18555 24160 18880 24188
rect 18555 24157 18567 24160
rect 18509 24151 18567 24157
rect 18874 24148 18880 24160
rect 18932 24148 18938 24200
rect 19426 24148 19432 24200
rect 19484 24148 19490 24200
rect 23492 24188 23520 24216
rect 24581 24191 24639 24197
rect 24581 24188 24593 24191
rect 23322 24160 23520 24188
rect 23676 24160 24593 24188
rect 13449 24123 13507 24129
rect 13449 24120 13461 24123
rect 12406 24092 13461 24120
rect 13449 24089 13461 24092
rect 13495 24089 13507 24123
rect 13449 24083 13507 24089
rect 17512 24092 19656 24120
rect 11146 24052 11152 24064
rect 10612 24024 11152 24052
rect 11146 24012 11152 24024
rect 11204 24012 11210 24064
rect 17512 24061 17540 24092
rect 17497 24055 17555 24061
rect 17497 24021 17509 24055
rect 17543 24021 17555 24055
rect 17497 24015 17555 24021
rect 17678 24012 17684 24064
rect 17736 24052 17742 24064
rect 18141 24055 18199 24061
rect 18141 24052 18153 24055
rect 17736 24024 18153 24052
rect 17736 24012 17742 24024
rect 18141 24021 18153 24024
rect 18187 24021 18199 24055
rect 18141 24015 18199 24021
rect 18230 24012 18236 24064
rect 18288 24052 18294 24064
rect 19058 24052 19064 24064
rect 18288 24024 19064 24052
rect 18288 24012 18294 24024
rect 19058 24012 19064 24024
rect 19116 24012 19122 24064
rect 19628 24052 19656 24092
rect 19702 24080 19708 24132
rect 19760 24080 19766 24132
rect 21634 24120 21640 24132
rect 20930 24092 21640 24120
rect 21634 24080 21640 24092
rect 21692 24080 21698 24132
rect 22186 24080 22192 24132
rect 22244 24080 22250 24132
rect 21082 24052 21088 24064
rect 19628 24024 21088 24052
rect 21082 24012 21088 24024
rect 21140 24012 21146 24064
rect 22830 24012 22836 24064
rect 22888 24052 22894 24064
rect 23676 24061 23704 24160
rect 24581 24157 24593 24160
rect 24627 24157 24639 24191
rect 24581 24151 24639 24157
rect 23661 24055 23719 24061
rect 23661 24052 23673 24055
rect 22888 24024 23673 24052
rect 22888 24012 22894 24024
rect 23661 24021 23673 24024
rect 23707 24021 23719 24055
rect 23661 24015 23719 24021
rect 24118 24012 24124 24064
rect 24176 24012 24182 24064
rect 25222 24012 25228 24064
rect 25280 24012 25286 24064
rect 1104 23962 25852 23984
rect 1104 23910 7950 23962
rect 8002 23910 8014 23962
rect 8066 23910 8078 23962
rect 8130 23910 8142 23962
rect 8194 23910 8206 23962
rect 8258 23910 17950 23962
rect 18002 23910 18014 23962
rect 18066 23910 18078 23962
rect 18130 23910 18142 23962
rect 18194 23910 18206 23962
rect 18258 23910 25852 23962
rect 1104 23888 25852 23910
rect 10134 23848 10140 23860
rect 8864 23820 10140 23848
rect 8864 23789 8892 23820
rect 10134 23808 10140 23820
rect 10192 23808 10198 23860
rect 12529 23851 12587 23857
rect 12529 23817 12541 23851
rect 12575 23848 12587 23851
rect 12710 23848 12716 23860
rect 12575 23820 12716 23848
rect 12575 23817 12587 23820
rect 12529 23811 12587 23817
rect 12710 23808 12716 23820
rect 12768 23808 12774 23860
rect 13449 23851 13507 23857
rect 13449 23817 13461 23851
rect 13495 23817 13507 23851
rect 13449 23811 13507 23817
rect 13909 23851 13967 23857
rect 13909 23817 13921 23851
rect 13955 23848 13967 23851
rect 14458 23848 14464 23860
rect 13955 23820 14464 23848
rect 13955 23817 13967 23820
rect 13909 23811 13967 23817
rect 8849 23783 8907 23789
rect 8849 23749 8861 23783
rect 8895 23749 8907 23783
rect 8849 23743 8907 23749
rect 8938 23740 8944 23792
rect 8996 23780 9002 23792
rect 13464 23780 13492 23811
rect 14458 23808 14464 23820
rect 14516 23808 14522 23860
rect 15105 23851 15163 23857
rect 15105 23817 15117 23851
rect 15151 23848 15163 23851
rect 16393 23851 16451 23857
rect 16393 23848 16405 23851
rect 15151 23820 16405 23848
rect 15151 23817 15163 23820
rect 15105 23811 15163 23817
rect 16393 23817 16405 23820
rect 16439 23848 16451 23851
rect 17586 23848 17592 23860
rect 16439 23820 17592 23848
rect 16439 23817 16451 23820
rect 16393 23811 16451 23817
rect 17586 23808 17592 23820
rect 17644 23808 17650 23860
rect 17770 23808 17776 23860
rect 17828 23848 17834 23860
rect 18230 23848 18236 23860
rect 17828 23820 18236 23848
rect 17828 23808 17834 23820
rect 18230 23808 18236 23820
rect 18288 23848 18294 23860
rect 18877 23851 18935 23857
rect 18877 23848 18889 23851
rect 18288 23820 18889 23848
rect 18288 23808 18294 23820
rect 18877 23817 18889 23820
rect 18923 23817 18935 23851
rect 18877 23811 18935 23817
rect 19702 23808 19708 23860
rect 19760 23848 19766 23860
rect 22649 23851 22707 23857
rect 22649 23848 22661 23851
rect 19760 23820 22661 23848
rect 19760 23808 19766 23820
rect 22649 23817 22661 23820
rect 22695 23817 22707 23851
rect 25222 23848 25228 23860
rect 22649 23811 22707 23817
rect 23492 23820 25228 23848
rect 19794 23780 19800 23792
rect 8996 23752 9338 23780
rect 13464 23752 18276 23780
rect 8996 23740 9002 23752
rect 7742 23672 7748 23724
rect 7800 23712 7806 23724
rect 8573 23715 8631 23721
rect 8573 23712 8585 23715
rect 7800 23684 8585 23712
rect 7800 23672 7806 23684
rect 8573 23681 8585 23684
rect 8619 23681 8631 23715
rect 8573 23675 8631 23681
rect 12618 23672 12624 23724
rect 12676 23712 12682 23724
rect 13817 23715 13875 23721
rect 13817 23712 13829 23715
rect 12676 23684 13829 23712
rect 12676 23672 12682 23684
rect 13817 23681 13829 23684
rect 13863 23681 13875 23715
rect 13817 23675 13875 23681
rect 15013 23715 15071 23721
rect 15013 23681 15025 23715
rect 15059 23712 15071 23715
rect 15841 23715 15899 23721
rect 15841 23712 15853 23715
rect 15059 23684 15853 23712
rect 15059 23681 15071 23684
rect 15013 23675 15071 23681
rect 15841 23681 15853 23684
rect 15887 23681 15899 23715
rect 15841 23675 15899 23681
rect 16114 23672 16120 23724
rect 16172 23712 16178 23724
rect 18248 23721 18276 23752
rect 19536 23752 19800 23780
rect 17221 23715 17279 23721
rect 17221 23712 17233 23715
rect 16172 23684 17233 23712
rect 16172 23672 16178 23684
rect 17221 23681 17233 23684
rect 17267 23712 17279 23715
rect 18233 23715 18291 23721
rect 17267 23684 17540 23712
rect 17267 23681 17279 23684
rect 17221 23675 17279 23681
rect 10321 23647 10379 23653
rect 10321 23613 10333 23647
rect 10367 23644 10379 23647
rect 10594 23644 10600 23656
rect 10367 23616 10600 23644
rect 10367 23613 10379 23616
rect 10321 23607 10379 23613
rect 10594 23604 10600 23616
rect 10652 23604 10658 23656
rect 13446 23604 13452 23656
rect 13504 23644 13510 23656
rect 14001 23647 14059 23653
rect 14001 23644 14013 23647
rect 13504 23616 14013 23644
rect 13504 23604 13510 23616
rect 14001 23613 14013 23616
rect 14047 23613 14059 23647
rect 14001 23607 14059 23613
rect 15197 23647 15255 23653
rect 15197 23613 15209 23647
rect 15243 23613 15255 23647
rect 15197 23607 15255 23613
rect 11882 23536 11888 23588
rect 11940 23576 11946 23588
rect 15212 23576 15240 23607
rect 16942 23604 16948 23656
rect 17000 23644 17006 23656
rect 17126 23644 17132 23656
rect 17000 23616 17132 23644
rect 17000 23604 17006 23616
rect 17126 23604 17132 23616
rect 17184 23644 17190 23656
rect 17313 23647 17371 23653
rect 17313 23644 17325 23647
rect 17184 23616 17325 23644
rect 17184 23604 17190 23616
rect 17313 23613 17325 23616
rect 17359 23613 17371 23647
rect 17313 23607 17371 23613
rect 17405 23647 17463 23653
rect 17405 23613 17417 23647
rect 17451 23613 17463 23647
rect 17405 23607 17463 23613
rect 11940 23548 15240 23576
rect 11940 23536 11946 23548
rect 16206 23536 16212 23588
rect 16264 23576 16270 23588
rect 17420 23576 17448 23607
rect 16264 23548 17448 23576
rect 17512 23576 17540 23684
rect 18233 23681 18245 23715
rect 18279 23681 18291 23715
rect 18233 23675 18291 23681
rect 18506 23672 18512 23724
rect 18564 23672 18570 23724
rect 17770 23604 17776 23656
rect 17828 23644 17834 23656
rect 18524 23644 18552 23672
rect 18693 23647 18751 23653
rect 18693 23644 18705 23647
rect 17828 23616 18705 23644
rect 17828 23604 17834 23616
rect 18693 23613 18705 23616
rect 18739 23613 18751 23647
rect 18693 23607 18751 23613
rect 18509 23579 18567 23585
rect 18509 23576 18521 23579
rect 17512 23548 18521 23576
rect 16264 23536 16270 23548
rect 18509 23545 18521 23548
rect 18555 23576 18567 23579
rect 19536 23576 19564 23752
rect 19794 23740 19800 23752
rect 19852 23740 19858 23792
rect 20901 23783 20959 23789
rect 20901 23749 20913 23783
rect 20947 23780 20959 23783
rect 22278 23780 22284 23792
rect 20947 23752 22284 23780
rect 20947 23749 20959 23752
rect 20901 23743 20959 23749
rect 22278 23740 22284 23752
rect 22336 23740 22342 23792
rect 23382 23780 23388 23792
rect 22664 23752 23388 23780
rect 19613 23715 19671 23721
rect 19613 23681 19625 23715
rect 19659 23681 19671 23715
rect 19613 23675 19671 23681
rect 19705 23715 19763 23721
rect 19705 23681 19717 23715
rect 19751 23712 19763 23715
rect 20346 23712 20352 23724
rect 19751 23684 20352 23712
rect 19751 23681 19763 23684
rect 19705 23675 19763 23681
rect 18555 23548 19564 23576
rect 19628 23576 19656 23675
rect 20346 23672 20352 23684
rect 20404 23672 20410 23724
rect 20806 23672 20812 23724
rect 20864 23672 20870 23724
rect 22005 23715 22063 23721
rect 22005 23712 22017 23715
rect 20916 23684 22017 23712
rect 19889 23647 19947 23653
rect 19889 23613 19901 23647
rect 19935 23644 19947 23647
rect 20916 23644 20944 23684
rect 22005 23681 22017 23684
rect 22051 23712 22063 23715
rect 22462 23712 22468 23724
rect 22051 23684 22468 23712
rect 22051 23681 22063 23684
rect 22005 23675 22063 23681
rect 22462 23672 22468 23684
rect 22520 23712 22526 23724
rect 22664 23712 22692 23752
rect 23382 23740 23388 23752
rect 23440 23740 23446 23792
rect 23492 23789 23520 23820
rect 25222 23808 25228 23820
rect 25280 23808 25286 23860
rect 23477 23783 23535 23789
rect 23477 23749 23489 23783
rect 23523 23749 23535 23783
rect 23477 23743 23535 23749
rect 22520 23684 22692 23712
rect 22520 23672 22526 23684
rect 19935 23616 20944 23644
rect 19935 23613 19947 23616
rect 19889 23607 19947 23613
rect 20990 23604 20996 23656
rect 21048 23604 21054 23656
rect 21082 23604 21088 23656
rect 21140 23644 21146 23656
rect 22186 23644 22192 23656
rect 21140 23616 22192 23644
rect 21140 23604 21146 23616
rect 22186 23604 22192 23616
rect 22244 23604 22250 23656
rect 22278 23604 22284 23656
rect 22336 23644 22342 23656
rect 22646 23644 22652 23656
rect 22336 23616 22652 23644
rect 22336 23604 22342 23616
rect 22646 23604 22652 23616
rect 22704 23604 22710 23656
rect 23198 23604 23204 23656
rect 23256 23604 23262 23656
rect 23842 23644 23848 23656
rect 23308 23616 23848 23644
rect 23308 23576 23336 23616
rect 23842 23604 23848 23616
rect 23900 23604 23906 23656
rect 19628 23548 23336 23576
rect 18555 23545 18567 23548
rect 18509 23539 18567 23545
rect 10226 23468 10232 23520
rect 10284 23508 10290 23520
rect 10597 23511 10655 23517
rect 10597 23508 10609 23511
rect 10284 23480 10609 23508
rect 10284 23468 10290 23480
rect 10597 23477 10609 23480
rect 10643 23508 10655 23511
rect 11330 23508 11336 23520
rect 10643 23480 11336 23508
rect 10643 23477 10655 23480
rect 10597 23471 10655 23477
rect 11330 23468 11336 23480
rect 11388 23508 11394 23520
rect 12710 23508 12716 23520
rect 11388 23480 12716 23508
rect 11388 23468 11394 23480
rect 12710 23468 12716 23480
rect 12768 23468 12774 23520
rect 14642 23468 14648 23520
rect 14700 23468 14706 23520
rect 15102 23468 15108 23520
rect 15160 23508 15166 23520
rect 16114 23508 16120 23520
rect 15160 23480 16120 23508
rect 15160 23468 15166 23480
rect 16114 23468 16120 23480
rect 16172 23468 16178 23520
rect 16853 23511 16911 23517
rect 16853 23477 16865 23511
rect 16899 23508 16911 23511
rect 16942 23508 16948 23520
rect 16899 23480 16948 23508
rect 16899 23477 16911 23480
rect 16853 23471 16911 23477
rect 16942 23468 16948 23480
rect 17000 23468 17006 23520
rect 18049 23511 18107 23517
rect 18049 23477 18061 23511
rect 18095 23508 18107 23511
rect 18322 23508 18328 23520
rect 18095 23480 18328 23508
rect 18095 23477 18107 23480
rect 18049 23471 18107 23477
rect 18322 23468 18328 23480
rect 18380 23468 18386 23520
rect 19245 23511 19303 23517
rect 19245 23477 19257 23511
rect 19291 23508 19303 23511
rect 19886 23508 19892 23520
rect 19291 23480 19892 23508
rect 19291 23477 19303 23480
rect 19245 23471 19303 23477
rect 19886 23468 19892 23480
rect 19944 23468 19950 23520
rect 20441 23511 20499 23517
rect 20441 23477 20453 23511
rect 20487 23508 20499 23511
rect 20530 23508 20536 23520
rect 20487 23480 20536 23508
rect 20487 23477 20499 23480
rect 20441 23471 20499 23477
rect 20530 23468 20536 23480
rect 20588 23468 20594 23520
rect 20990 23468 20996 23520
rect 21048 23508 21054 23520
rect 21358 23508 21364 23520
rect 21048 23480 21364 23508
rect 21048 23468 21054 23480
rect 21358 23468 21364 23480
rect 21416 23468 21422 23520
rect 21545 23511 21603 23517
rect 21545 23477 21557 23511
rect 21591 23508 21603 23511
rect 21634 23508 21640 23520
rect 21591 23480 21640 23508
rect 21591 23477 21603 23480
rect 21545 23471 21603 23477
rect 21634 23468 21640 23480
rect 21692 23468 21698 23520
rect 22462 23468 22468 23520
rect 22520 23508 22526 23520
rect 22922 23508 22928 23520
rect 22520 23480 22928 23508
rect 22520 23468 22526 23480
rect 22922 23468 22928 23480
rect 22980 23468 22986 23520
rect 24118 23468 24124 23520
rect 24176 23508 24182 23520
rect 24596 23508 24624 23698
rect 24949 23647 25007 23653
rect 24949 23613 24961 23647
rect 24995 23644 25007 23647
rect 25130 23644 25136 23656
rect 24995 23616 25136 23644
rect 24995 23613 25007 23616
rect 24949 23607 25007 23613
rect 25130 23604 25136 23616
rect 25188 23604 25194 23656
rect 25225 23511 25283 23517
rect 25225 23508 25237 23511
rect 24176 23480 25237 23508
rect 24176 23468 24182 23480
rect 25225 23477 25237 23480
rect 25271 23508 25283 23511
rect 25409 23511 25467 23517
rect 25409 23508 25421 23511
rect 25271 23480 25421 23508
rect 25271 23477 25283 23480
rect 25225 23471 25283 23477
rect 25409 23477 25421 23480
rect 25455 23477 25467 23511
rect 25409 23471 25467 23477
rect 1104 23418 25852 23440
rect 1104 23366 2950 23418
rect 3002 23366 3014 23418
rect 3066 23366 3078 23418
rect 3130 23366 3142 23418
rect 3194 23366 3206 23418
rect 3258 23366 12950 23418
rect 13002 23366 13014 23418
rect 13066 23366 13078 23418
rect 13130 23366 13142 23418
rect 13194 23366 13206 23418
rect 13258 23366 22950 23418
rect 23002 23366 23014 23418
rect 23066 23366 23078 23418
rect 23130 23366 23142 23418
rect 23194 23366 23206 23418
rect 23258 23366 25852 23418
rect 1104 23344 25852 23366
rect 10962 23264 10968 23316
rect 11020 23304 11026 23316
rect 11241 23307 11299 23313
rect 11241 23304 11253 23307
rect 11020 23276 11253 23304
rect 11020 23264 11026 23276
rect 11241 23273 11253 23276
rect 11287 23273 11299 23307
rect 11241 23267 11299 23273
rect 14185 23307 14243 23313
rect 14185 23273 14197 23307
rect 14231 23304 14243 23307
rect 17126 23304 17132 23316
rect 14231 23276 17132 23304
rect 14231 23273 14243 23276
rect 14185 23267 14243 23273
rect 10870 23168 10876 23180
rect 9508 23140 10876 23168
rect 9508 23109 9536 23140
rect 10870 23128 10876 23140
rect 10928 23128 10934 23180
rect 13541 23171 13599 23177
rect 13541 23168 13553 23171
rect 12406 23140 13553 23168
rect 9493 23103 9551 23109
rect 9493 23069 9505 23103
rect 9539 23069 9551 23103
rect 9493 23063 9551 23069
rect 10594 23060 10600 23112
rect 10652 23060 10658 23112
rect 9122 22992 9128 23044
rect 9180 23032 9186 23044
rect 12406 23032 12434 23140
rect 13541 23137 13553 23140
rect 13587 23137 13599 23171
rect 13541 23131 13599 23137
rect 13449 23103 13507 23109
rect 13449 23069 13461 23103
rect 13495 23100 13507 23103
rect 14200 23100 14228 23267
rect 17126 23264 17132 23276
rect 17184 23264 17190 23316
rect 18969 23307 19027 23313
rect 18969 23273 18981 23307
rect 19015 23304 19027 23307
rect 19058 23304 19064 23316
rect 19015 23276 19064 23304
rect 19015 23273 19027 23276
rect 18969 23267 19027 23273
rect 19058 23264 19064 23276
rect 19116 23264 19122 23316
rect 14369 23239 14427 23245
rect 14369 23205 14381 23239
rect 14415 23236 14427 23239
rect 15102 23236 15108 23248
rect 14415 23208 15108 23236
rect 14415 23205 14427 23208
rect 14369 23199 14427 23205
rect 13495 23072 14228 23100
rect 13495 23069 13507 23072
rect 13449 23063 13507 23069
rect 9180 23004 12434 23032
rect 13357 23035 13415 23041
rect 9180 22992 9186 23004
rect 13357 23001 13369 23035
rect 13403 23032 13415 23035
rect 14384 23032 14412 23199
rect 15102 23196 15108 23208
rect 15160 23196 15166 23248
rect 17865 23239 17923 23245
rect 17865 23205 17877 23239
rect 17911 23236 17923 23239
rect 18506 23236 18512 23248
rect 17911 23208 18512 23236
rect 17911 23205 17923 23208
rect 17865 23199 17923 23205
rect 18506 23196 18512 23208
rect 18564 23196 18570 23248
rect 20809 23239 20867 23245
rect 20809 23205 20821 23239
rect 20855 23236 20867 23239
rect 22646 23236 22652 23248
rect 20855 23208 22652 23236
rect 20855 23205 20867 23208
rect 20809 23199 20867 23205
rect 22646 23196 22652 23208
rect 22704 23196 22710 23248
rect 15010 23128 15016 23180
rect 15068 23168 15074 23180
rect 15289 23171 15347 23177
rect 15289 23168 15301 23171
rect 15068 23140 15301 23168
rect 15068 23128 15074 23140
rect 15289 23137 15301 23140
rect 15335 23137 15347 23171
rect 15289 23131 15347 23137
rect 18230 23128 18236 23180
rect 18288 23168 18294 23180
rect 18325 23171 18383 23177
rect 18325 23168 18337 23171
rect 18288 23140 18337 23168
rect 18288 23128 18294 23140
rect 18325 23137 18337 23140
rect 18371 23137 18383 23171
rect 18325 23131 18383 23137
rect 18417 23171 18475 23177
rect 18417 23137 18429 23171
rect 18463 23168 18475 23171
rect 18874 23168 18880 23180
rect 18463 23140 18880 23168
rect 18463 23137 18475 23140
rect 18417 23131 18475 23137
rect 18340 23100 18368 23131
rect 18874 23128 18880 23140
rect 18932 23128 18938 23180
rect 20070 23128 20076 23180
rect 20128 23128 20134 23180
rect 23750 23128 23756 23180
rect 23808 23128 23814 23180
rect 25038 23128 25044 23180
rect 25096 23128 25102 23180
rect 25222 23128 25228 23180
rect 25280 23128 25286 23180
rect 18340 23072 19840 23100
rect 13403 23004 14412 23032
rect 18233 23035 18291 23041
rect 13403 23001 13415 23004
rect 13357 22995 13415 23001
rect 18233 23001 18245 23035
rect 18279 23032 18291 23035
rect 18782 23032 18788 23044
rect 18279 23004 18788 23032
rect 18279 23001 18291 23004
rect 18233 22995 18291 23001
rect 18782 22992 18788 23004
rect 18840 22992 18846 23044
rect 19812 23032 19840 23072
rect 19886 23060 19892 23112
rect 19944 23060 19950 23112
rect 19978 23060 19984 23112
rect 20036 23100 20042 23112
rect 20993 23103 21051 23109
rect 20993 23100 21005 23103
rect 20036 23072 21005 23100
rect 20036 23060 20042 23072
rect 20993 23069 21005 23072
rect 21039 23069 21051 23103
rect 20993 23063 21051 23069
rect 21545 23103 21603 23109
rect 21545 23069 21557 23103
rect 21591 23100 21603 23103
rect 22278 23100 22284 23112
rect 21591 23072 22284 23100
rect 21591 23069 21603 23072
rect 21545 23063 21603 23069
rect 22278 23060 22284 23072
rect 22336 23060 22342 23112
rect 22833 23103 22891 23109
rect 22833 23069 22845 23103
rect 22879 23100 22891 23103
rect 23842 23100 23848 23112
rect 22879 23072 23848 23100
rect 22879 23069 22891 23072
rect 22833 23063 22891 23069
rect 23842 23060 23848 23072
rect 23900 23060 23906 23112
rect 24949 23103 25007 23109
rect 24949 23069 24961 23103
rect 24995 23100 25007 23103
rect 26050 23100 26056 23112
rect 24995 23072 26056 23100
rect 24995 23069 25007 23072
rect 24949 23063 25007 23069
rect 25056 23044 25084 23072
rect 26050 23060 26056 23072
rect 26108 23060 26114 23112
rect 21358 23032 21364 23044
rect 19812 23004 21364 23032
rect 21358 22992 21364 23004
rect 21416 22992 21422 23044
rect 25038 22992 25044 23044
rect 25096 22992 25102 23044
rect 8478 22924 8484 22976
rect 8536 22964 8542 22976
rect 10137 22967 10195 22973
rect 10137 22964 10149 22967
rect 8536 22936 10149 22964
rect 8536 22924 8542 22936
rect 10137 22933 10149 22936
rect 10183 22933 10195 22967
rect 10137 22927 10195 22933
rect 12342 22924 12348 22976
rect 12400 22964 12406 22976
rect 12989 22967 13047 22973
rect 12989 22964 13001 22967
rect 12400 22936 13001 22964
rect 12400 22924 12406 22936
rect 12989 22933 13001 22936
rect 13035 22933 13047 22967
rect 12989 22927 13047 22933
rect 17034 22924 17040 22976
rect 17092 22964 17098 22976
rect 18598 22964 18604 22976
rect 17092 22936 18604 22964
rect 17092 22924 17098 22936
rect 18598 22924 18604 22936
rect 18656 22924 18662 22976
rect 19518 22924 19524 22976
rect 19576 22924 19582 22976
rect 19981 22967 20039 22973
rect 19981 22933 19993 22967
rect 20027 22964 20039 22967
rect 22002 22964 22008 22976
rect 20027 22936 22008 22964
rect 20027 22933 20039 22936
rect 19981 22927 20039 22933
rect 22002 22924 22008 22936
rect 22060 22924 22066 22976
rect 22189 22967 22247 22973
rect 22189 22933 22201 22967
rect 22235 22964 22247 22967
rect 23566 22964 23572 22976
rect 22235 22936 23572 22964
rect 22235 22933 22247 22936
rect 22189 22927 22247 22933
rect 23566 22924 23572 22936
rect 23624 22924 23630 22976
rect 24486 22924 24492 22976
rect 24544 22964 24550 22976
rect 24581 22967 24639 22973
rect 24581 22964 24593 22967
rect 24544 22936 24593 22964
rect 24544 22924 24550 22936
rect 24581 22933 24593 22936
rect 24627 22933 24639 22967
rect 24581 22927 24639 22933
rect 1104 22874 25852 22896
rect 1104 22822 7950 22874
rect 8002 22822 8014 22874
rect 8066 22822 8078 22874
rect 8130 22822 8142 22874
rect 8194 22822 8206 22874
rect 8258 22822 17950 22874
rect 18002 22822 18014 22874
rect 18066 22822 18078 22874
rect 18130 22822 18142 22874
rect 18194 22822 18206 22874
rect 18258 22822 25852 22874
rect 1104 22800 25852 22822
rect 9858 22760 9864 22772
rect 8864 22732 9864 22760
rect 8478 22652 8484 22704
rect 8536 22652 8542 22704
rect 8864 22692 8892 22732
rect 9858 22720 9864 22732
rect 9916 22760 9922 22772
rect 10226 22760 10232 22772
rect 9916 22732 10232 22760
rect 9916 22720 9922 22732
rect 10226 22720 10232 22732
rect 10284 22720 10290 22772
rect 11793 22763 11851 22769
rect 11793 22729 11805 22763
rect 11839 22760 11851 22763
rect 11839 22732 17080 22760
rect 11839 22729 11851 22732
rect 11793 22723 11851 22729
rect 8938 22692 8944 22704
rect 8864 22664 8944 22692
rect 8938 22652 8944 22664
rect 8996 22652 9002 22704
rect 10594 22652 10600 22704
rect 10652 22692 10658 22704
rect 15010 22692 15016 22704
rect 10652 22664 12388 22692
rect 14950 22664 15016 22692
rect 10652 22652 10658 22664
rect 7742 22584 7748 22636
rect 7800 22624 7806 22636
rect 8205 22627 8263 22633
rect 8205 22624 8217 22627
rect 7800 22596 8217 22624
rect 7800 22584 7806 22596
rect 8205 22593 8217 22596
rect 8251 22593 8263 22627
rect 8205 22587 8263 22593
rect 11790 22584 11796 22636
rect 11848 22624 11854 22636
rect 12161 22627 12219 22633
rect 12161 22624 12173 22627
rect 11848 22596 12173 22624
rect 11848 22584 11854 22596
rect 12161 22593 12173 22596
rect 12207 22593 12219 22627
rect 12161 22587 12219 22593
rect 12360 22565 12388 22664
rect 15010 22652 15016 22664
rect 15068 22652 15074 22704
rect 15749 22695 15807 22701
rect 15749 22661 15761 22695
rect 15795 22692 15807 22695
rect 16298 22692 16304 22704
rect 15795 22664 16304 22692
rect 15795 22661 15807 22664
rect 15749 22655 15807 22661
rect 16298 22652 16304 22664
rect 16356 22652 16362 22704
rect 15028 22624 15056 22652
rect 17052 22633 17080 22732
rect 17126 22720 17132 22772
rect 17184 22760 17190 22772
rect 18693 22763 18751 22769
rect 18693 22760 18705 22763
rect 17184 22732 18705 22760
rect 17184 22720 17190 22732
rect 18693 22729 18705 22732
rect 18739 22760 18751 22763
rect 19702 22760 19708 22772
rect 18739 22732 19708 22760
rect 18739 22729 18751 22732
rect 18693 22723 18751 22729
rect 19702 22720 19708 22732
rect 19760 22720 19766 22772
rect 21082 22720 21088 22772
rect 21140 22720 21146 22772
rect 18414 22652 18420 22704
rect 18472 22652 18478 22704
rect 19334 22652 19340 22704
rect 19392 22692 19398 22704
rect 21177 22695 21235 22701
rect 21177 22692 21189 22695
rect 19392 22664 21189 22692
rect 19392 22652 19398 22664
rect 21177 22661 21189 22664
rect 21223 22661 21235 22695
rect 21177 22655 21235 22661
rect 23293 22695 23351 22701
rect 23293 22661 23305 22695
rect 23339 22692 23351 22695
rect 24854 22692 24860 22704
rect 23339 22664 24860 22692
rect 23339 22661 23351 22664
rect 23293 22655 23351 22661
rect 24854 22652 24860 22664
rect 24912 22652 24918 22704
rect 17037 22627 17095 22633
rect 15028 22596 16528 22624
rect 12253 22559 12311 22565
rect 12253 22525 12265 22559
rect 12299 22525 12311 22559
rect 12253 22519 12311 22525
rect 12345 22559 12403 22565
rect 12345 22525 12357 22559
rect 12391 22525 12403 22559
rect 12345 22519 12403 22525
rect 13449 22559 13507 22565
rect 13449 22525 13461 22559
rect 13495 22525 13507 22559
rect 13449 22519 13507 22525
rect 12268 22488 12296 22519
rect 13354 22488 13360 22500
rect 12268 22460 13360 22488
rect 13354 22448 13360 22460
rect 13412 22448 13418 22500
rect 7282 22380 7288 22432
rect 7340 22420 7346 22432
rect 9950 22420 9956 22432
rect 7340 22392 9956 22420
rect 7340 22380 7346 22392
rect 9950 22380 9956 22392
rect 10008 22380 10014 22432
rect 12802 22380 12808 22432
rect 12860 22380 12866 22432
rect 13464 22420 13492 22519
rect 13722 22516 13728 22568
rect 13780 22516 13786 22568
rect 14458 22516 14464 22568
rect 14516 22556 14522 22568
rect 15933 22559 15991 22565
rect 15933 22556 15945 22559
rect 14516 22528 15945 22556
rect 14516 22516 14522 22528
rect 15933 22525 15945 22528
rect 15979 22525 15991 22559
rect 16500 22556 16528 22596
rect 17037 22593 17049 22627
rect 17083 22593 17095 22627
rect 17037 22587 17095 22593
rect 19242 22584 19248 22636
rect 19300 22624 19306 22636
rect 19981 22627 20039 22633
rect 19981 22624 19993 22627
rect 19300 22596 19993 22624
rect 19300 22584 19306 22596
rect 19981 22593 19993 22596
rect 20027 22593 20039 22627
rect 19981 22587 20039 22593
rect 20070 22584 20076 22636
rect 20128 22624 20134 22636
rect 22097 22627 22155 22633
rect 22097 22624 22109 22627
rect 20128 22596 22109 22624
rect 20128 22584 20134 22596
rect 22097 22593 22109 22596
rect 22143 22593 22155 22627
rect 22097 22587 22155 22593
rect 22370 22584 22376 22636
rect 22428 22624 22434 22636
rect 23937 22627 23995 22633
rect 23937 22624 23949 22627
rect 22428 22596 23949 22624
rect 22428 22584 22434 22596
rect 23937 22593 23949 22596
rect 23983 22593 23995 22627
rect 23937 22587 23995 22593
rect 17586 22556 17592 22568
rect 16500 22528 17592 22556
rect 15933 22519 15991 22525
rect 17586 22516 17592 22528
rect 17644 22516 17650 22568
rect 18601 22559 18659 22565
rect 18601 22525 18613 22559
rect 18647 22556 18659 22559
rect 18782 22556 18788 22568
rect 18647 22528 18788 22556
rect 18647 22525 18659 22528
rect 18601 22519 18659 22525
rect 18782 22516 18788 22528
rect 18840 22516 18846 22568
rect 19337 22559 19395 22565
rect 19337 22525 19349 22559
rect 19383 22556 19395 22559
rect 20622 22556 20628 22568
rect 19383 22528 20628 22556
rect 19383 22525 19395 22528
rect 19337 22519 19395 22525
rect 20622 22516 20628 22528
rect 20680 22516 20686 22568
rect 21269 22559 21327 22565
rect 21269 22525 21281 22559
rect 21315 22525 21327 22559
rect 21269 22519 21327 22525
rect 16114 22488 16120 22500
rect 15120 22460 16120 22488
rect 15120 22420 15148 22460
rect 16114 22448 16120 22460
rect 16172 22448 16178 22500
rect 16853 22491 16911 22497
rect 16853 22457 16865 22491
rect 16899 22488 16911 22491
rect 19978 22488 19984 22500
rect 16899 22460 19984 22488
rect 16899 22457 16911 22460
rect 16853 22451 16911 22457
rect 19978 22448 19984 22460
rect 20036 22448 20042 22500
rect 20898 22448 20904 22500
rect 20956 22488 20962 22500
rect 21284 22488 21312 22519
rect 24762 22516 24768 22568
rect 24820 22516 24826 22568
rect 20956 22460 21312 22488
rect 20956 22448 20962 22460
rect 13464 22392 15148 22420
rect 15194 22380 15200 22432
rect 15252 22420 15258 22432
rect 17402 22420 17408 22432
rect 15252 22392 17408 22420
rect 15252 22380 15258 22392
rect 17402 22380 17408 22392
rect 17460 22380 17466 22432
rect 17770 22380 17776 22432
rect 17828 22420 17834 22432
rect 18230 22420 18236 22432
rect 17828 22392 18236 22420
rect 17828 22380 17834 22392
rect 18230 22380 18236 22392
rect 18288 22380 18294 22432
rect 18414 22380 18420 22432
rect 18472 22420 18478 22432
rect 18969 22423 19027 22429
rect 18969 22420 18981 22423
rect 18472 22392 18981 22420
rect 18472 22380 18478 22392
rect 18969 22389 18981 22392
rect 19015 22420 19027 22423
rect 19058 22420 19064 22432
rect 19015 22392 19064 22420
rect 19015 22389 19027 22392
rect 18969 22383 19027 22389
rect 19058 22380 19064 22392
rect 19116 22420 19122 22432
rect 20346 22420 20352 22432
rect 19116 22392 20352 22420
rect 19116 22380 19122 22392
rect 20346 22380 20352 22392
rect 20404 22380 20410 22432
rect 20714 22380 20720 22432
rect 20772 22380 20778 22432
rect 1104 22330 25852 22352
rect 1104 22278 2950 22330
rect 3002 22278 3014 22330
rect 3066 22278 3078 22330
rect 3130 22278 3142 22330
rect 3194 22278 3206 22330
rect 3258 22278 12950 22330
rect 13002 22278 13014 22330
rect 13066 22278 13078 22330
rect 13130 22278 13142 22330
rect 13194 22278 13206 22330
rect 13258 22278 22950 22330
rect 23002 22278 23014 22330
rect 23066 22278 23078 22330
rect 23130 22278 23142 22330
rect 23194 22278 23206 22330
rect 23258 22278 25852 22330
rect 1104 22256 25852 22278
rect 7088 22219 7146 22225
rect 7088 22185 7100 22219
rect 7134 22216 7146 22219
rect 9398 22216 9404 22228
rect 7134 22188 9404 22216
rect 7134 22185 7146 22188
rect 7088 22179 7146 22185
rect 9398 22176 9404 22188
rect 9456 22176 9462 22228
rect 9950 22176 9956 22228
rect 10008 22216 10014 22228
rect 10008 22188 11836 22216
rect 10008 22176 10014 22188
rect 9490 22108 9496 22160
rect 9548 22148 9554 22160
rect 11808 22148 11836 22188
rect 12434 22176 12440 22228
rect 12492 22176 12498 22228
rect 12710 22176 12716 22228
rect 12768 22216 12774 22228
rect 12768 22188 13308 22216
rect 12768 22176 12774 22188
rect 12452 22148 12480 22176
rect 13280 22148 13308 22188
rect 13722 22176 13728 22228
rect 13780 22216 13786 22228
rect 15654 22216 15660 22228
rect 13780 22188 15660 22216
rect 13780 22176 13786 22188
rect 15654 22176 15660 22188
rect 15712 22176 15718 22228
rect 18230 22176 18236 22228
rect 18288 22216 18294 22228
rect 18288 22188 18552 22216
rect 18288 22176 18294 22188
rect 15194 22148 15200 22160
rect 9548 22120 10732 22148
rect 11808 22120 11928 22148
rect 12452 22120 13216 22148
rect 13280 22120 15200 22148
rect 9548 22108 9554 22120
rect 6825 22083 6883 22089
rect 6825 22049 6837 22083
rect 6871 22080 6883 22083
rect 7558 22080 7564 22092
rect 6871 22052 7564 22080
rect 6871 22049 6883 22052
rect 6825 22043 6883 22049
rect 7558 22040 7564 22052
rect 7616 22040 7622 22092
rect 8941 22083 8999 22089
rect 8941 22080 8953 22083
rect 8220 22052 8953 22080
rect 8220 22024 8248 22052
rect 8941 22049 8953 22052
rect 8987 22080 8999 22083
rect 9858 22080 9864 22092
rect 8987 22052 9864 22080
rect 8987 22049 8999 22052
rect 8941 22043 8999 22049
rect 9858 22040 9864 22052
rect 9916 22040 9922 22092
rect 10704 22089 10732 22120
rect 11900 22089 11928 22120
rect 10689 22083 10747 22089
rect 10689 22049 10701 22083
rect 10735 22049 10747 22083
rect 10689 22043 10747 22049
rect 11885 22083 11943 22089
rect 11885 22049 11897 22083
rect 11931 22080 11943 22083
rect 11931 22052 11965 22080
rect 11931 22049 11943 22052
rect 11885 22043 11943 22049
rect 12434 22040 12440 22092
rect 12492 22080 12498 22092
rect 12802 22080 12808 22092
rect 12492 22052 12808 22080
rect 12492 22040 12498 22052
rect 12802 22040 12808 22052
rect 12860 22080 12866 22092
rect 13188 22089 13216 22120
rect 15194 22108 15200 22120
rect 15252 22108 15258 22160
rect 18414 22108 18420 22160
rect 18472 22108 18478 22160
rect 18524 22148 18552 22188
rect 18782 22176 18788 22228
rect 18840 22216 18846 22228
rect 21174 22216 21180 22228
rect 18840 22188 21180 22216
rect 18840 22176 18846 22188
rect 21174 22176 21180 22188
rect 21232 22176 21238 22228
rect 23293 22219 23351 22225
rect 23293 22185 23305 22219
rect 23339 22216 23351 22219
rect 23382 22216 23388 22228
rect 23339 22188 23388 22216
rect 23339 22185 23351 22188
rect 23293 22179 23351 22185
rect 23382 22176 23388 22188
rect 23440 22176 23446 22228
rect 23842 22176 23848 22228
rect 23900 22176 23906 22228
rect 20438 22148 20444 22160
rect 18524 22120 19334 22148
rect 12989 22083 13047 22089
rect 12989 22080 13001 22083
rect 12860 22052 13001 22080
rect 12860 22040 12866 22052
rect 12989 22049 13001 22052
rect 13035 22049 13047 22083
rect 12989 22043 13047 22049
rect 13173 22083 13231 22089
rect 13173 22049 13185 22083
rect 13219 22080 13231 22083
rect 13219 22052 13253 22080
rect 13219 22049 13231 22052
rect 13173 22043 13231 22049
rect 15378 22040 15384 22092
rect 15436 22040 15442 22092
rect 15470 22040 15476 22092
rect 15528 22040 15534 22092
rect 16022 22040 16028 22092
rect 16080 22080 16086 22092
rect 16117 22083 16175 22089
rect 16117 22080 16129 22083
rect 16080 22052 16129 22080
rect 16080 22040 16086 22052
rect 16117 22049 16129 22052
rect 16163 22049 16175 22083
rect 16117 22043 16175 22049
rect 16393 22083 16451 22089
rect 16393 22049 16405 22083
rect 16439 22080 16451 22083
rect 17034 22080 17040 22092
rect 16439 22052 17040 22080
rect 16439 22049 16451 22052
rect 16393 22043 16451 22049
rect 17034 22040 17040 22052
rect 17092 22040 17098 22092
rect 17586 22054 17592 22106
rect 17644 22054 17650 22106
rect 19306 22080 19334 22120
rect 20364 22120 20444 22148
rect 20364 22089 20392 22120
rect 20438 22108 20444 22120
rect 20496 22108 20502 22160
rect 25406 22148 25412 22160
rect 25240 22120 25412 22148
rect 20165 22083 20223 22089
rect 20165 22080 20177 22083
rect 8202 21972 8208 22024
rect 8260 21972 8266 22024
rect 8404 21984 11652 22012
rect 6270 21836 6276 21888
rect 6328 21876 6334 21888
rect 8404 21876 8432 21984
rect 10505 21947 10563 21953
rect 10505 21913 10517 21947
rect 10551 21944 10563 21947
rect 11624 21944 11652 21984
rect 11698 21972 11704 22024
rect 11756 21972 11762 22024
rect 11793 22015 11851 22021
rect 11793 21981 11805 22015
rect 11839 22012 11851 22015
rect 11974 22012 11980 22024
rect 11839 21984 11980 22012
rect 11839 21981 11851 21984
rect 11793 21975 11851 21981
rect 11974 21972 11980 21984
rect 12032 21972 12038 22024
rect 17604 22012 17632 22054
rect 19306 22052 20177 22080
rect 20165 22049 20177 22052
rect 20211 22049 20223 22083
rect 20165 22043 20223 22049
rect 20349 22083 20407 22089
rect 20349 22049 20361 22083
rect 20395 22080 20407 22083
rect 20395 22052 20429 22080
rect 20395 22049 20407 22052
rect 20349 22043 20407 22049
rect 20806 22040 20812 22092
rect 20864 22080 20870 22092
rect 20901 22083 20959 22089
rect 20901 22080 20913 22083
rect 20864 22052 20913 22080
rect 20864 22040 20870 22052
rect 20901 22049 20913 22052
rect 20947 22049 20959 22083
rect 20901 22043 20959 22049
rect 21545 22083 21603 22089
rect 21545 22049 21557 22083
rect 21591 22080 21603 22083
rect 23290 22080 23296 22092
rect 21591 22052 23296 22080
rect 21591 22049 21603 22052
rect 21545 22043 21603 22049
rect 23290 22040 23296 22052
rect 23348 22040 23354 22092
rect 24670 22040 24676 22092
rect 24728 22080 24734 22092
rect 25240 22089 25268 22120
rect 25406 22108 25412 22120
rect 25464 22108 25470 22160
rect 25041 22083 25099 22089
rect 25041 22080 25053 22083
rect 24728 22052 25053 22080
rect 24728 22040 24734 22052
rect 25041 22049 25053 22052
rect 25087 22049 25099 22083
rect 25041 22043 25099 22049
rect 25225 22083 25283 22089
rect 25225 22049 25237 22083
rect 25271 22080 25283 22083
rect 25271 22052 25305 22080
rect 25271 22049 25283 22052
rect 25225 22043 25283 22049
rect 18693 22015 18751 22021
rect 12406 21984 15148 22012
rect 17526 21984 18552 22012
rect 12406 21944 12434 21984
rect 10551 21916 11560 21944
rect 11624 21916 12434 21944
rect 12897 21947 12955 21953
rect 10551 21913 10563 21916
rect 10505 21907 10563 21913
rect 6328 21848 8432 21876
rect 6328 21836 6334 21848
rect 8478 21836 8484 21888
rect 8536 21876 8542 21888
rect 8573 21879 8631 21885
rect 8573 21876 8585 21879
rect 8536 21848 8585 21876
rect 8536 21836 8542 21848
rect 8573 21845 8585 21848
rect 8619 21845 8631 21879
rect 8573 21839 8631 21845
rect 9490 21836 9496 21888
rect 9548 21836 9554 21888
rect 10042 21836 10048 21888
rect 10100 21876 10106 21888
rect 10137 21879 10195 21885
rect 10137 21876 10149 21879
rect 10100 21848 10149 21876
rect 10100 21836 10106 21848
rect 10137 21845 10149 21848
rect 10183 21845 10195 21879
rect 10137 21839 10195 21845
rect 10594 21836 10600 21888
rect 10652 21836 10658 21888
rect 11238 21836 11244 21888
rect 11296 21876 11302 21888
rect 11333 21879 11391 21885
rect 11333 21876 11345 21879
rect 11296 21848 11345 21876
rect 11296 21836 11302 21848
rect 11333 21845 11345 21848
rect 11379 21845 11391 21879
rect 11532 21876 11560 21916
rect 12897 21913 12909 21947
rect 12943 21944 12955 21947
rect 13354 21944 13360 21956
rect 12943 21916 13360 21944
rect 12943 21913 12955 21916
rect 12897 21907 12955 21913
rect 13354 21904 13360 21916
rect 13412 21904 13418 21956
rect 15120 21944 15148 21984
rect 18414 21944 18420 21956
rect 15120 21916 15424 21944
rect 11606 21876 11612 21888
rect 11532 21848 11612 21876
rect 11333 21839 11391 21845
rect 11606 21836 11612 21848
rect 11664 21836 11670 21888
rect 12526 21836 12532 21888
rect 12584 21836 12590 21888
rect 14918 21836 14924 21888
rect 14976 21836 14982 21888
rect 15286 21836 15292 21888
rect 15344 21836 15350 21888
rect 15396 21876 15424 21916
rect 17696 21916 18420 21944
rect 17696 21876 17724 21916
rect 18414 21904 18420 21916
rect 18472 21904 18478 21956
rect 15396 21848 17724 21876
rect 17770 21836 17776 21888
rect 17828 21876 17834 21888
rect 17865 21879 17923 21885
rect 17865 21876 17877 21879
rect 17828 21848 17877 21876
rect 17828 21836 17834 21848
rect 17865 21845 17877 21848
rect 17911 21845 17923 21879
rect 17865 21839 17923 21845
rect 18233 21879 18291 21885
rect 18233 21845 18245 21879
rect 18279 21876 18291 21879
rect 18524 21876 18552 21984
rect 18693 21981 18705 22015
rect 18739 22012 18751 22015
rect 21266 22012 21272 22024
rect 18739 21984 21272 22012
rect 18739 21981 18751 21984
rect 18693 21975 18751 21981
rect 21266 21972 21272 21984
rect 21324 21972 21330 22024
rect 23106 21972 23112 22024
rect 23164 22012 23170 22024
rect 24029 22015 24087 22021
rect 24029 22012 24041 22015
rect 23164 21984 24041 22012
rect 23164 21972 23170 21984
rect 24029 21981 24041 21984
rect 24075 21981 24087 22015
rect 24029 21975 24087 21981
rect 20346 21944 20352 21956
rect 19720 21916 20352 21944
rect 18598 21876 18604 21888
rect 18279 21848 18604 21876
rect 18279 21845 18291 21848
rect 18233 21839 18291 21845
rect 18598 21836 18604 21848
rect 18656 21836 18662 21888
rect 19334 21836 19340 21888
rect 19392 21836 19398 21888
rect 19720 21885 19748 21916
rect 20346 21904 20352 21916
rect 20404 21904 20410 21956
rect 21818 21904 21824 21956
rect 21876 21904 21882 21956
rect 23198 21944 23204 21956
rect 23046 21916 23204 21944
rect 23198 21904 23204 21916
rect 23256 21904 23262 21956
rect 24949 21947 25007 21953
rect 24949 21944 24961 21947
rect 23492 21916 24961 21944
rect 19705 21879 19763 21885
rect 19705 21845 19717 21879
rect 19751 21845 19763 21879
rect 19705 21839 19763 21845
rect 20073 21879 20131 21885
rect 20073 21845 20085 21879
rect 20119 21876 20131 21879
rect 20162 21876 20168 21888
rect 20119 21848 20168 21876
rect 20119 21845 20131 21848
rect 20073 21839 20131 21845
rect 20162 21836 20168 21848
rect 20220 21836 20226 21888
rect 20622 21836 20628 21888
rect 20680 21876 20686 21888
rect 23492 21876 23520 21916
rect 24949 21913 24961 21916
rect 24995 21913 25007 21947
rect 24949 21907 25007 21913
rect 20680 21848 23520 21876
rect 20680 21836 20686 21848
rect 24578 21836 24584 21888
rect 24636 21836 24642 21888
rect 1104 21786 25852 21808
rect 1104 21734 7950 21786
rect 8002 21734 8014 21786
rect 8066 21734 8078 21786
rect 8130 21734 8142 21786
rect 8194 21734 8206 21786
rect 8258 21734 17950 21786
rect 18002 21734 18014 21786
rect 18066 21734 18078 21786
rect 18130 21734 18142 21786
rect 18194 21734 18206 21786
rect 18258 21734 25852 21786
rect 1104 21712 25852 21734
rect 9766 21632 9772 21684
rect 9824 21672 9830 21684
rect 10321 21675 10379 21681
rect 10321 21672 10333 21675
rect 9824 21644 10333 21672
rect 9824 21632 9830 21644
rect 10321 21641 10333 21644
rect 10367 21641 10379 21675
rect 10321 21635 10379 21641
rect 10689 21675 10747 21681
rect 10689 21641 10701 21675
rect 10735 21672 10747 21675
rect 14642 21672 14648 21684
rect 10735 21644 14648 21672
rect 10735 21641 10747 21644
rect 10689 21635 10747 21641
rect 14642 21632 14648 21644
rect 14700 21632 14706 21684
rect 15654 21632 15660 21684
rect 15712 21632 15718 21684
rect 19242 21632 19248 21684
rect 19300 21632 19306 21684
rect 20162 21632 20168 21684
rect 20220 21672 20226 21684
rect 20530 21672 20536 21684
rect 20220 21644 20536 21672
rect 20220 21632 20226 21644
rect 20530 21632 20536 21644
rect 20588 21632 20594 21684
rect 22465 21675 22523 21681
rect 22465 21641 22477 21675
rect 22511 21672 22523 21675
rect 22554 21672 22560 21684
rect 22511 21644 22560 21672
rect 22511 21641 22523 21644
rect 22465 21635 22523 21641
rect 22554 21632 22560 21644
rect 22612 21632 22618 21684
rect 22738 21632 22744 21684
rect 22796 21672 22802 21684
rect 25041 21675 25099 21681
rect 25041 21672 25053 21675
rect 22796 21644 25053 21672
rect 22796 21632 22802 21644
rect 25041 21641 25053 21644
rect 25087 21641 25099 21675
rect 25041 21635 25099 21641
rect 8294 21564 8300 21616
rect 8352 21564 8358 21616
rect 9858 21564 9864 21616
rect 9916 21564 9922 21616
rect 13630 21564 13636 21616
rect 13688 21564 13694 21616
rect 14918 21564 14924 21616
rect 14976 21604 14982 21616
rect 14976 21576 18460 21604
rect 14976 21564 14982 21576
rect 11701 21539 11759 21545
rect 11701 21505 11713 21539
rect 11747 21536 11759 21539
rect 12710 21536 12716 21548
rect 11747 21508 12716 21536
rect 11747 21505 11759 21508
rect 11701 21499 11759 21505
rect 12710 21496 12716 21508
rect 12768 21496 12774 21548
rect 15013 21539 15071 21545
rect 15013 21536 15025 21539
rect 14568 21508 15025 21536
rect 7558 21428 7564 21480
rect 7616 21428 7622 21480
rect 7837 21471 7895 21477
rect 7837 21437 7849 21471
rect 7883 21468 7895 21471
rect 8570 21468 8576 21480
rect 7883 21440 8576 21468
rect 7883 21437 7895 21440
rect 7837 21431 7895 21437
rect 8570 21428 8576 21440
rect 8628 21428 8634 21480
rect 9582 21428 9588 21480
rect 9640 21428 9646 21480
rect 10410 21428 10416 21480
rect 10468 21468 10474 21480
rect 10781 21471 10839 21477
rect 10781 21468 10793 21471
rect 10468 21440 10793 21468
rect 10468 21428 10474 21440
rect 10781 21437 10793 21440
rect 10827 21437 10839 21471
rect 10781 21431 10839 21437
rect 10873 21471 10931 21477
rect 10873 21437 10885 21471
rect 10919 21437 10931 21471
rect 10873 21431 10931 21437
rect 9398 21360 9404 21412
rect 9456 21400 9462 21412
rect 10888 21400 10916 21431
rect 11146 21428 11152 21480
rect 11204 21468 11210 21480
rect 12618 21468 12624 21480
rect 11204 21440 12624 21468
rect 11204 21428 11210 21440
rect 12618 21428 12624 21440
rect 12676 21468 12682 21480
rect 12805 21471 12863 21477
rect 12805 21468 12817 21471
rect 12676 21440 12817 21468
rect 12676 21428 12682 21440
rect 12805 21437 12817 21440
rect 12851 21437 12863 21471
rect 12805 21431 12863 21437
rect 13081 21471 13139 21477
rect 13081 21437 13093 21471
rect 13127 21468 13139 21471
rect 13814 21468 13820 21480
rect 13127 21440 13820 21468
rect 13127 21437 13139 21440
rect 13081 21431 13139 21437
rect 13814 21428 13820 21440
rect 13872 21468 13878 21480
rect 14090 21468 14096 21480
rect 13872 21440 14096 21468
rect 13872 21428 13878 21440
rect 14090 21428 14096 21440
rect 14148 21428 14154 21480
rect 14568 21477 14596 21508
rect 15013 21505 15025 21508
rect 15059 21536 15071 21539
rect 15470 21536 15476 21548
rect 15059 21508 15476 21536
rect 15059 21505 15071 21508
rect 15013 21499 15071 21505
rect 15470 21496 15476 21508
rect 15528 21496 15534 21548
rect 16574 21496 16580 21548
rect 16632 21536 16638 21548
rect 18432 21545 18460 21576
rect 19058 21564 19064 21616
rect 19116 21604 19122 21616
rect 19337 21607 19395 21613
rect 19337 21604 19349 21607
rect 19116 21576 19349 21604
rect 19116 21564 19122 21576
rect 19337 21573 19349 21576
rect 19383 21573 19395 21607
rect 23106 21604 23112 21616
rect 19337 21567 19395 21573
rect 19444 21576 23112 21604
rect 16853 21539 16911 21545
rect 16853 21536 16865 21539
rect 16632 21508 16865 21536
rect 16632 21496 16638 21508
rect 16853 21505 16865 21508
rect 16899 21505 16911 21539
rect 16853 21499 16911 21505
rect 18417 21539 18475 21545
rect 18417 21505 18429 21539
rect 18463 21505 18475 21539
rect 18417 21499 18475 21505
rect 18966 21496 18972 21548
rect 19024 21536 19030 21548
rect 19444 21536 19472 21576
rect 23106 21564 23112 21576
rect 23164 21564 23170 21616
rect 23198 21564 23204 21616
rect 23256 21604 23262 21616
rect 24026 21604 24032 21616
rect 23256 21576 24032 21604
rect 23256 21564 23262 21576
rect 24026 21564 24032 21576
rect 24084 21564 24090 21616
rect 24118 21564 24124 21616
rect 24176 21564 24182 21616
rect 19024 21508 19472 21536
rect 20257 21539 20315 21545
rect 19024 21496 19030 21508
rect 20257 21505 20269 21539
rect 20303 21536 20315 21539
rect 22002 21536 22008 21548
rect 20303 21508 22008 21536
rect 20303 21505 20315 21508
rect 20257 21499 20315 21505
rect 22002 21496 22008 21508
rect 22060 21496 22066 21548
rect 22373 21539 22431 21545
rect 22373 21505 22385 21539
rect 22419 21536 22431 21539
rect 22554 21536 22560 21548
rect 22419 21508 22560 21536
rect 22419 21505 22431 21508
rect 22373 21499 22431 21505
rect 22554 21496 22560 21508
rect 22612 21496 22618 21548
rect 23290 21496 23296 21548
rect 23348 21496 23354 21548
rect 14553 21471 14611 21477
rect 14553 21437 14565 21471
rect 14599 21437 14611 21471
rect 14553 21431 14611 21437
rect 15102 21428 15108 21480
rect 15160 21468 15166 21480
rect 19334 21468 19340 21480
rect 15160 21440 19340 21468
rect 15160 21428 15166 21440
rect 19334 21428 19340 21440
rect 19392 21428 19398 21480
rect 19521 21471 19579 21477
rect 19521 21437 19533 21471
rect 19567 21468 19579 21471
rect 20898 21468 20904 21480
rect 19567 21440 20904 21468
rect 19567 21437 19579 21440
rect 19521 21431 19579 21437
rect 20898 21428 20904 21440
rect 20956 21428 20962 21480
rect 21269 21471 21327 21477
rect 21269 21437 21281 21471
rect 21315 21468 21327 21471
rect 22649 21471 22707 21477
rect 21315 21440 22094 21468
rect 21315 21437 21327 21440
rect 21269 21431 21327 21437
rect 9456 21372 10916 21400
rect 9456 21360 9462 21372
rect 11790 21360 11796 21412
rect 11848 21400 11854 21412
rect 11848 21372 12940 21400
rect 11848 21360 11854 21372
rect 12345 21335 12403 21341
rect 12345 21301 12357 21335
rect 12391 21332 12403 21335
rect 12710 21332 12716 21344
rect 12391 21304 12716 21332
rect 12391 21301 12403 21304
rect 12345 21295 12403 21301
rect 12710 21292 12716 21304
rect 12768 21292 12774 21344
rect 12912 21332 12940 21372
rect 15378 21360 15384 21412
rect 15436 21400 15442 21412
rect 17865 21403 17923 21409
rect 15436 21372 17632 21400
rect 15436 21360 15442 21372
rect 14734 21332 14740 21344
rect 12912 21304 14740 21332
rect 14734 21292 14740 21304
rect 14792 21292 14798 21344
rect 15470 21292 15476 21344
rect 15528 21332 15534 21344
rect 17497 21335 17555 21341
rect 17497 21332 17509 21335
rect 15528 21304 17509 21332
rect 15528 21292 15534 21304
rect 17497 21301 17509 21304
rect 17543 21301 17555 21335
rect 17604 21332 17632 21372
rect 17865 21369 17877 21403
rect 17911 21400 17923 21403
rect 18598 21400 18604 21412
rect 17911 21372 18604 21400
rect 17911 21369 17923 21372
rect 17865 21363 17923 21369
rect 18598 21360 18604 21372
rect 18656 21360 18662 21412
rect 19352 21400 19380 21428
rect 21082 21400 21088 21412
rect 19352 21372 21088 21400
rect 21082 21360 21088 21372
rect 21140 21360 21146 21412
rect 22066 21400 22094 21440
rect 22649 21437 22661 21471
rect 22695 21468 22707 21471
rect 22922 21468 22928 21480
rect 22695 21440 22928 21468
rect 22695 21437 22707 21440
rect 22649 21431 22707 21437
rect 22922 21428 22928 21440
rect 22980 21428 22986 21480
rect 23569 21471 23627 21477
rect 23569 21437 23581 21471
rect 23615 21468 23627 21471
rect 25406 21468 25412 21480
rect 23615 21440 25412 21468
rect 23615 21437 23627 21440
rect 23569 21431 23627 21437
rect 25406 21428 25412 21440
rect 25464 21428 25470 21480
rect 22066 21372 23428 21400
rect 23400 21344 23428 21372
rect 18233 21335 18291 21341
rect 18233 21332 18245 21335
rect 17604 21304 18245 21332
rect 17497 21295 17555 21301
rect 18233 21301 18245 21304
rect 18279 21301 18291 21335
rect 18233 21295 18291 21301
rect 18877 21335 18935 21341
rect 18877 21301 18889 21335
rect 18923 21332 18935 21335
rect 20438 21332 20444 21344
rect 18923 21304 20444 21332
rect 18923 21301 18935 21304
rect 18877 21295 18935 21301
rect 20438 21292 20444 21304
rect 20496 21292 20502 21344
rect 21726 21292 21732 21344
rect 21784 21332 21790 21344
rect 22005 21335 22063 21341
rect 22005 21332 22017 21335
rect 21784 21304 22017 21332
rect 21784 21292 21790 21304
rect 22005 21301 22017 21304
rect 22051 21301 22063 21335
rect 22005 21295 22063 21301
rect 23382 21292 23388 21344
rect 23440 21292 23446 21344
rect 24118 21292 24124 21344
rect 24176 21332 24182 21344
rect 25317 21335 25375 21341
rect 25317 21332 25329 21335
rect 24176 21304 25329 21332
rect 24176 21292 24182 21304
rect 25317 21301 25329 21304
rect 25363 21301 25375 21335
rect 25317 21295 25375 21301
rect 1104 21242 25852 21264
rect 1104 21190 2950 21242
rect 3002 21190 3014 21242
rect 3066 21190 3078 21242
rect 3130 21190 3142 21242
rect 3194 21190 3206 21242
rect 3258 21190 12950 21242
rect 13002 21190 13014 21242
rect 13066 21190 13078 21242
rect 13130 21190 13142 21242
rect 13194 21190 13206 21242
rect 13258 21190 22950 21242
rect 23002 21190 23014 21242
rect 23066 21190 23078 21242
rect 23130 21190 23142 21242
rect 23194 21190 23206 21242
rect 23258 21190 25852 21242
rect 1104 21168 25852 21190
rect 8570 21088 8576 21140
rect 8628 21088 8634 21140
rect 9677 21131 9735 21137
rect 9677 21097 9689 21131
rect 9723 21128 9735 21131
rect 10686 21128 10692 21140
rect 9723 21100 10692 21128
rect 9723 21097 9735 21100
rect 9677 21091 9735 21097
rect 10686 21088 10692 21100
rect 10744 21088 10750 21140
rect 10796 21100 12756 21128
rect 5258 21020 5264 21072
rect 5316 21060 5322 21072
rect 10796 21060 10824 21100
rect 5316 21032 10824 21060
rect 12728 21060 12756 21100
rect 12802 21088 12808 21140
rect 12860 21128 12866 21140
rect 13538 21128 13544 21140
rect 12860 21100 13544 21128
rect 12860 21088 12866 21100
rect 13538 21088 13544 21100
rect 13596 21088 13602 21140
rect 15194 21088 15200 21140
rect 15252 21128 15258 21140
rect 16114 21128 16120 21140
rect 15252 21100 16120 21128
rect 15252 21088 15258 21100
rect 16114 21088 16120 21100
rect 16172 21088 16178 21140
rect 16482 21088 16488 21140
rect 16540 21128 16546 21140
rect 16945 21131 17003 21137
rect 16945 21128 16957 21131
rect 16540 21100 16957 21128
rect 16540 21088 16546 21100
rect 16945 21097 16957 21100
rect 16991 21128 17003 21131
rect 17034 21128 17040 21140
rect 16991 21100 17040 21128
rect 16991 21097 17003 21100
rect 16945 21091 17003 21097
rect 17034 21088 17040 21100
rect 17092 21088 17098 21140
rect 17635 21131 17693 21137
rect 17635 21097 17647 21131
rect 17681 21128 17693 21131
rect 19978 21128 19984 21140
rect 17681 21100 19984 21128
rect 17681 21097 17693 21100
rect 17635 21091 17693 21097
rect 19978 21088 19984 21100
rect 20036 21088 20042 21140
rect 20254 21088 20260 21140
rect 20312 21128 20318 21140
rect 21637 21131 21695 21137
rect 21637 21128 21649 21131
rect 20312 21100 21649 21128
rect 20312 21088 20318 21100
rect 21637 21097 21649 21100
rect 21683 21097 21695 21131
rect 21637 21091 21695 21097
rect 22002 21088 22008 21140
rect 22060 21088 22066 21140
rect 15102 21060 15108 21072
rect 12728 21032 15108 21060
rect 5316 21020 5322 21032
rect 15102 21020 15108 21032
rect 15160 21020 15166 21072
rect 16500 21032 21220 21060
rect 10226 20952 10232 21004
rect 10284 20952 10290 21004
rect 11146 20952 11152 21004
rect 11204 20952 11210 21004
rect 13354 20952 13360 21004
rect 13412 20952 13418 21004
rect 15470 20952 15476 21004
rect 15528 20952 15534 21004
rect 16022 20952 16028 21004
rect 16080 20992 16086 21004
rect 16500 20992 16528 21032
rect 16080 20964 16528 20992
rect 17405 20995 17463 21001
rect 16080 20952 16086 20964
rect 17405 20961 17417 20995
rect 17451 20992 17463 20995
rect 18322 20992 18328 21004
rect 17451 20964 18328 20992
rect 17451 20961 17463 20964
rect 17405 20955 17463 20961
rect 18322 20952 18328 20964
rect 18380 20952 18386 21004
rect 19978 20952 19984 21004
rect 20036 20952 20042 21004
rect 7929 20927 7987 20933
rect 7929 20893 7941 20927
rect 7975 20924 7987 20927
rect 8478 20924 8484 20936
rect 7975 20896 8484 20924
rect 7975 20893 7987 20896
rect 7929 20887 7987 20893
rect 8478 20884 8484 20896
rect 8536 20884 8542 20936
rect 9490 20884 9496 20936
rect 9548 20924 9554 20936
rect 10045 20927 10103 20933
rect 10045 20924 10057 20927
rect 9548 20896 10057 20924
rect 9548 20884 9554 20896
rect 10045 20893 10057 20896
rect 10091 20893 10103 20927
rect 10045 20887 10103 20893
rect 15194 20884 15200 20936
rect 15252 20884 15258 20936
rect 18414 20884 18420 20936
rect 18472 20924 18478 20936
rect 18877 20927 18935 20933
rect 18877 20924 18889 20927
rect 18472 20896 18889 20924
rect 18472 20884 18478 20896
rect 18877 20893 18889 20896
rect 18923 20893 18935 20927
rect 18877 20887 18935 20893
rect 19797 20927 19855 20933
rect 19797 20893 19809 20927
rect 19843 20924 19855 20927
rect 19886 20924 19892 20936
rect 19843 20896 19892 20924
rect 19843 20893 19855 20896
rect 19797 20887 19855 20893
rect 19886 20884 19892 20896
rect 19944 20884 19950 20936
rect 20993 20927 21051 20933
rect 20993 20893 21005 20927
rect 21039 20924 21051 20927
rect 21082 20924 21088 20936
rect 21039 20896 21088 20924
rect 21039 20893 21051 20896
rect 20993 20887 21051 20893
rect 21082 20884 21088 20896
rect 21140 20884 21146 20936
rect 21192 20924 21220 21032
rect 22186 21020 22192 21072
rect 22244 21060 22250 21072
rect 22244 21032 25084 21060
rect 22244 21020 22250 21032
rect 21269 20995 21327 21001
rect 21269 20961 21281 20995
rect 21315 20992 21327 20995
rect 23845 20995 23903 21001
rect 21315 20964 22600 20992
rect 21315 20961 21327 20964
rect 21269 20955 21327 20961
rect 22189 20927 22247 20933
rect 22189 20924 22201 20927
rect 21192 20896 22201 20924
rect 22189 20893 22201 20896
rect 22235 20893 22247 20927
rect 22189 20887 22247 20893
rect 11422 20816 11428 20868
rect 11480 20816 11486 20868
rect 11808 20828 11914 20856
rect 8294 20748 8300 20800
rect 8352 20788 8358 20800
rect 8478 20788 8484 20800
rect 8352 20760 8484 20788
rect 8352 20748 8358 20760
rect 8478 20748 8484 20760
rect 8536 20748 8542 20800
rect 9401 20791 9459 20797
rect 9401 20757 9413 20791
rect 9447 20788 9459 20791
rect 10137 20791 10195 20797
rect 10137 20788 10149 20791
rect 9447 20760 10149 20788
rect 9447 20757 9459 20760
rect 9401 20751 9459 20757
rect 10137 20757 10149 20760
rect 10183 20788 10195 20791
rect 10226 20788 10232 20800
rect 10183 20760 10232 20788
rect 10183 20757 10195 20760
rect 10137 20751 10195 20757
rect 10226 20748 10232 20760
rect 10284 20748 10290 20800
rect 10962 20748 10968 20800
rect 11020 20788 11026 20800
rect 11808 20788 11836 20828
rect 13354 20816 13360 20868
rect 13412 20856 13418 20868
rect 13630 20856 13636 20868
rect 13412 20828 13636 20856
rect 13412 20816 13418 20828
rect 13630 20816 13636 20828
rect 13688 20856 13694 20868
rect 13817 20859 13875 20865
rect 13817 20856 13829 20859
rect 13688 20828 13829 20856
rect 13688 20816 13694 20828
rect 13817 20825 13829 20828
rect 13863 20856 13875 20859
rect 14645 20859 14703 20865
rect 14645 20856 14657 20859
rect 13863 20828 14657 20856
rect 13863 20825 13875 20828
rect 13817 20819 13875 20825
rect 14645 20825 14657 20828
rect 14691 20856 14703 20859
rect 14829 20859 14887 20865
rect 14829 20856 14841 20859
rect 14691 20828 14841 20856
rect 14691 20825 14703 20828
rect 14645 20819 14703 20825
rect 14829 20825 14841 20828
rect 14875 20856 14887 20859
rect 14875 20828 15962 20856
rect 14875 20825 14887 20828
rect 14829 20819 14887 20825
rect 19702 20816 19708 20868
rect 19760 20856 19766 20868
rect 22002 20856 22008 20868
rect 19760 20828 22008 20856
rect 19760 20816 19766 20828
rect 11020 20760 11836 20788
rect 12897 20791 12955 20797
rect 11020 20748 11026 20760
rect 12897 20757 12909 20791
rect 12943 20788 12955 20791
rect 14090 20788 14096 20800
rect 12943 20760 14096 20788
rect 12943 20757 12955 20760
rect 12897 20751 12955 20757
rect 14090 20748 14096 20760
rect 14148 20788 14154 20800
rect 14734 20788 14740 20800
rect 14148 20760 14740 20788
rect 14148 20748 14154 20760
rect 14734 20748 14740 20760
rect 14792 20748 14798 20800
rect 18693 20791 18751 20797
rect 18693 20757 18705 20791
rect 18739 20788 18751 20791
rect 19334 20788 19340 20800
rect 18739 20760 19340 20788
rect 18739 20757 18751 20760
rect 18693 20751 18751 20757
rect 19334 20748 19340 20760
rect 19392 20748 19398 20800
rect 19429 20791 19487 20797
rect 19429 20757 19441 20791
rect 19475 20788 19487 20791
rect 19794 20788 19800 20800
rect 19475 20760 19800 20788
rect 19475 20757 19487 20760
rect 19429 20751 19487 20757
rect 19794 20748 19800 20760
rect 19852 20748 19858 20800
rect 19904 20797 19932 20828
rect 22002 20816 22008 20828
rect 22060 20816 22066 20868
rect 19889 20791 19947 20797
rect 19889 20757 19901 20791
rect 19935 20757 19947 20791
rect 19889 20751 19947 20757
rect 20625 20791 20683 20797
rect 20625 20757 20637 20791
rect 20671 20788 20683 20791
rect 20898 20788 20904 20800
rect 20671 20760 20904 20788
rect 20671 20757 20683 20760
rect 20625 20751 20683 20757
rect 20898 20748 20904 20760
rect 20956 20748 20962 20800
rect 21082 20748 21088 20800
rect 21140 20788 21146 20800
rect 21358 20788 21364 20800
rect 21140 20760 21364 20788
rect 21140 20748 21146 20760
rect 21358 20748 21364 20760
rect 21416 20748 21422 20800
rect 22572 20788 22600 20964
rect 23845 20961 23857 20995
rect 23891 20992 23903 20995
rect 24854 20992 24860 21004
rect 23891 20964 24860 20992
rect 23891 20961 23903 20964
rect 23845 20955 23903 20961
rect 24854 20952 24860 20964
rect 24912 20952 24918 21004
rect 25056 21001 25084 21032
rect 25041 20995 25099 21001
rect 25041 20961 25053 20995
rect 25087 20961 25099 20995
rect 25041 20955 25099 20961
rect 25133 20995 25191 21001
rect 25133 20961 25145 20995
rect 25179 20961 25191 20995
rect 25133 20955 25191 20961
rect 22646 20884 22652 20936
rect 22704 20884 22710 20936
rect 23934 20884 23940 20936
rect 23992 20924 23998 20936
rect 25148 20924 25176 20955
rect 23992 20896 25176 20924
rect 23992 20884 23998 20896
rect 23750 20816 23756 20868
rect 23808 20856 23814 20868
rect 25498 20856 25504 20868
rect 23808 20828 25504 20856
rect 23808 20816 23814 20828
rect 25498 20816 25504 20828
rect 25556 20816 25562 20868
rect 22646 20788 22652 20800
rect 22572 20760 22652 20788
rect 22646 20748 22652 20760
rect 22704 20748 22710 20800
rect 24581 20791 24639 20797
rect 24581 20757 24593 20791
rect 24627 20788 24639 20791
rect 24854 20788 24860 20800
rect 24627 20760 24860 20788
rect 24627 20757 24639 20760
rect 24581 20751 24639 20757
rect 24854 20748 24860 20760
rect 24912 20748 24918 20800
rect 24946 20748 24952 20800
rect 25004 20788 25010 20800
rect 25866 20788 25872 20800
rect 25004 20760 25872 20788
rect 25004 20748 25010 20760
rect 25866 20748 25872 20760
rect 25924 20748 25930 20800
rect 1104 20698 25852 20720
rect 1104 20646 7950 20698
rect 8002 20646 8014 20698
rect 8066 20646 8078 20698
rect 8130 20646 8142 20698
rect 8194 20646 8206 20698
rect 8258 20646 17950 20698
rect 18002 20646 18014 20698
rect 18066 20646 18078 20698
rect 18130 20646 18142 20698
rect 18194 20646 18206 20698
rect 18258 20646 25852 20698
rect 1104 20624 25852 20646
rect 8021 20587 8079 20593
rect 8021 20553 8033 20587
rect 8067 20584 8079 20587
rect 9306 20584 9312 20596
rect 8067 20556 9312 20584
rect 8067 20553 8079 20556
rect 8021 20547 8079 20553
rect 9306 20544 9312 20556
rect 9364 20544 9370 20596
rect 11422 20544 11428 20596
rect 11480 20584 11486 20596
rect 12345 20587 12403 20593
rect 12345 20584 12357 20587
rect 11480 20556 12357 20584
rect 11480 20544 11486 20556
rect 12345 20553 12357 20556
rect 12391 20553 12403 20587
rect 12345 20547 12403 20553
rect 15013 20587 15071 20593
rect 15013 20553 15025 20587
rect 15059 20553 15071 20587
rect 15013 20547 15071 20553
rect 15473 20587 15531 20593
rect 15473 20553 15485 20587
rect 15519 20584 15531 20587
rect 15838 20584 15844 20596
rect 15519 20556 15844 20584
rect 15519 20553 15531 20556
rect 15473 20547 15531 20553
rect 8481 20519 8539 20525
rect 8481 20485 8493 20519
rect 8527 20516 8539 20519
rect 10134 20516 10140 20528
rect 8527 20488 10140 20516
rect 8527 20485 8539 20488
rect 8481 20479 8539 20485
rect 10134 20476 10140 20488
rect 10192 20476 10198 20528
rect 12710 20476 12716 20528
rect 12768 20516 12774 20528
rect 13081 20519 13139 20525
rect 13081 20516 13093 20519
rect 12768 20488 13093 20516
rect 12768 20476 12774 20488
rect 13081 20485 13093 20488
rect 13127 20485 13139 20519
rect 13081 20479 13139 20485
rect 13354 20476 13360 20528
rect 13412 20516 13418 20528
rect 15028 20516 15056 20547
rect 15838 20544 15844 20556
rect 15896 20544 15902 20596
rect 19242 20584 19248 20596
rect 17512 20556 19248 20584
rect 17512 20516 17540 20556
rect 19242 20544 19248 20556
rect 19300 20544 19306 20596
rect 19797 20587 19855 20593
rect 19797 20553 19809 20587
rect 19843 20584 19855 20587
rect 19886 20584 19892 20596
rect 19843 20556 19892 20584
rect 19843 20553 19855 20556
rect 19797 20547 19855 20553
rect 19886 20544 19892 20556
rect 19944 20544 19950 20596
rect 21818 20544 21824 20596
rect 21876 20584 21882 20596
rect 23109 20587 23167 20593
rect 23109 20584 23121 20587
rect 21876 20556 23121 20584
rect 21876 20544 21882 20556
rect 23109 20553 23121 20556
rect 23155 20553 23167 20587
rect 23109 20547 23167 20553
rect 25222 20544 25228 20596
rect 25280 20584 25286 20596
rect 25317 20587 25375 20593
rect 25317 20584 25329 20587
rect 25280 20556 25329 20584
rect 25280 20544 25286 20556
rect 25317 20553 25329 20556
rect 25363 20553 25375 20587
rect 25317 20547 25375 20553
rect 19610 20516 19616 20528
rect 13412 20488 13570 20516
rect 15028 20488 17540 20516
rect 19260 20488 19616 20516
rect 13412 20476 13418 20488
rect 6733 20451 6791 20457
rect 6733 20417 6745 20451
rect 6779 20448 6791 20451
rect 8294 20448 8300 20460
rect 6779 20420 8300 20448
rect 6779 20417 6791 20420
rect 6733 20411 6791 20417
rect 8294 20408 8300 20420
rect 8352 20408 8358 20460
rect 8389 20451 8447 20457
rect 8389 20417 8401 20451
rect 8435 20448 8447 20451
rect 9030 20448 9036 20460
rect 8435 20420 9036 20448
rect 8435 20417 8447 20420
rect 8389 20411 8447 20417
rect 9030 20408 9036 20420
rect 9088 20408 9094 20460
rect 11698 20408 11704 20460
rect 11756 20408 11762 20460
rect 15381 20451 15439 20457
rect 15381 20448 15393 20451
rect 14292 20420 15393 20448
rect 8573 20383 8631 20389
rect 8573 20349 8585 20383
rect 8619 20349 8631 20383
rect 8573 20343 8631 20349
rect 7650 20272 7656 20324
rect 7708 20312 7714 20324
rect 8588 20312 8616 20343
rect 12618 20340 12624 20392
rect 12676 20380 12682 20392
rect 12805 20383 12863 20389
rect 12805 20380 12817 20383
rect 12676 20352 12817 20380
rect 12676 20340 12682 20352
rect 12805 20349 12817 20352
rect 12851 20349 12863 20383
rect 12805 20343 12863 20349
rect 13538 20340 13544 20392
rect 13596 20380 13602 20392
rect 14292 20380 14320 20420
rect 15381 20417 15393 20420
rect 15427 20417 15439 20451
rect 18598 20448 18604 20460
rect 18262 20420 18604 20448
rect 15381 20411 15439 20417
rect 18598 20408 18604 20420
rect 18656 20448 18662 20460
rect 19260 20457 19288 20488
rect 19610 20476 19616 20488
rect 19668 20476 19674 20528
rect 22002 20476 22008 20528
rect 22060 20476 22066 20528
rect 24118 20476 24124 20528
rect 24176 20516 24182 20528
rect 24176 20488 24334 20516
rect 24176 20476 24182 20488
rect 19245 20451 19303 20457
rect 18656 20420 18920 20448
rect 18656 20408 18662 20420
rect 13596 20352 14320 20380
rect 14553 20383 14611 20389
rect 13596 20340 13602 20352
rect 14553 20349 14565 20383
rect 14599 20380 14611 20383
rect 14642 20380 14648 20392
rect 14599 20352 14648 20380
rect 14599 20349 14611 20352
rect 14553 20343 14611 20349
rect 14642 20340 14648 20352
rect 14700 20380 14706 20392
rect 15565 20383 15623 20389
rect 15565 20380 15577 20383
rect 14700 20352 15577 20380
rect 14700 20340 14706 20352
rect 15565 20349 15577 20352
rect 15611 20349 15623 20383
rect 15565 20343 15623 20349
rect 16853 20383 16911 20389
rect 16853 20349 16865 20383
rect 16899 20349 16911 20383
rect 16853 20343 16911 20349
rect 17129 20383 17187 20389
rect 17129 20349 17141 20383
rect 17175 20380 17187 20383
rect 18782 20380 18788 20392
rect 17175 20352 18788 20380
rect 17175 20349 17187 20352
rect 17129 20343 17187 20349
rect 7708 20284 8616 20312
rect 7708 20272 7714 20284
rect 7190 20204 7196 20256
rect 7248 20244 7254 20256
rect 7377 20247 7435 20253
rect 7377 20244 7389 20247
rect 7248 20216 7389 20244
rect 7248 20204 7254 20216
rect 7377 20213 7389 20216
rect 7423 20213 7435 20247
rect 16868 20244 16896 20343
rect 18782 20340 18788 20352
rect 18840 20340 18846 20392
rect 18892 20380 18920 20420
rect 19245 20417 19257 20451
rect 19291 20417 19303 20451
rect 19245 20411 19303 20417
rect 19334 20408 19340 20460
rect 19392 20448 19398 20460
rect 20073 20451 20131 20457
rect 20073 20448 20085 20451
rect 19392 20420 20085 20448
rect 19392 20408 19398 20420
rect 20073 20417 20085 20420
rect 20119 20417 20131 20451
rect 20073 20411 20131 20417
rect 21174 20408 21180 20460
rect 21232 20448 21238 20460
rect 21821 20451 21879 20457
rect 21821 20448 21833 20451
rect 21232 20420 21833 20448
rect 21232 20408 21238 20420
rect 21821 20417 21833 20420
rect 21867 20417 21879 20451
rect 21821 20411 21879 20417
rect 22465 20451 22523 20457
rect 22465 20417 22477 20451
rect 22511 20448 22523 20451
rect 22738 20448 22744 20460
rect 22511 20420 22744 20448
rect 22511 20417 22523 20420
rect 22465 20411 22523 20417
rect 22738 20408 22744 20420
rect 22796 20408 22802 20460
rect 19610 20380 19616 20392
rect 18892 20352 19616 20380
rect 19610 20340 19616 20352
rect 19668 20340 19674 20392
rect 21269 20383 21327 20389
rect 21269 20349 21281 20383
rect 21315 20380 21327 20383
rect 23198 20380 23204 20392
rect 21315 20352 23204 20380
rect 21315 20349 21327 20352
rect 21269 20343 21327 20349
rect 23198 20340 23204 20352
rect 23256 20340 23262 20392
rect 23290 20340 23296 20392
rect 23348 20380 23354 20392
rect 23569 20383 23627 20389
rect 23569 20380 23581 20383
rect 23348 20352 23581 20380
rect 23348 20340 23354 20352
rect 23569 20349 23581 20352
rect 23615 20349 23627 20383
rect 23569 20343 23627 20349
rect 23845 20383 23903 20389
rect 23845 20349 23857 20383
rect 23891 20380 23903 20383
rect 23891 20352 25084 20380
rect 23891 20349 23903 20352
rect 23845 20343 23903 20349
rect 19426 20312 19432 20324
rect 18524 20284 19432 20312
rect 18524 20244 18552 20284
rect 19426 20272 19432 20284
rect 19484 20312 19490 20324
rect 19886 20312 19892 20324
rect 19484 20284 19892 20312
rect 19484 20272 19490 20284
rect 19886 20272 19892 20284
rect 19944 20272 19950 20324
rect 25056 20256 25084 20352
rect 16868 20216 18552 20244
rect 18601 20247 18659 20253
rect 7377 20207 7435 20213
rect 18601 20213 18613 20247
rect 18647 20244 18659 20247
rect 18690 20244 18696 20256
rect 18647 20216 18696 20244
rect 18647 20213 18659 20216
rect 18601 20207 18659 20213
rect 18690 20204 18696 20216
rect 18748 20244 18754 20256
rect 18966 20244 18972 20256
rect 18748 20216 18972 20244
rect 18748 20204 18754 20216
rect 18966 20204 18972 20216
rect 19024 20204 19030 20256
rect 19058 20204 19064 20256
rect 19116 20204 19122 20256
rect 19610 20204 19616 20256
rect 19668 20204 19674 20256
rect 25038 20204 25044 20256
rect 25096 20204 25102 20256
rect 1104 20154 25852 20176
rect 1104 20102 2950 20154
rect 3002 20102 3014 20154
rect 3066 20102 3078 20154
rect 3130 20102 3142 20154
rect 3194 20102 3206 20154
rect 3258 20102 12950 20154
rect 13002 20102 13014 20154
rect 13066 20102 13078 20154
rect 13130 20102 13142 20154
rect 13194 20102 13206 20154
rect 13258 20102 22950 20154
rect 23002 20102 23014 20154
rect 23066 20102 23078 20154
rect 23130 20102 23142 20154
rect 23194 20102 23206 20154
rect 23258 20102 25852 20154
rect 1104 20080 25852 20102
rect 8478 20000 8484 20052
rect 8536 20000 8542 20052
rect 9858 20000 9864 20052
rect 9916 20040 9922 20052
rect 10962 20040 10968 20052
rect 9916 20012 10968 20040
rect 9916 20000 9922 20012
rect 10962 20000 10968 20012
rect 11020 20040 11026 20052
rect 11149 20043 11207 20049
rect 11149 20040 11161 20043
rect 11020 20012 11161 20040
rect 11020 20000 11026 20012
rect 11149 20009 11161 20012
rect 11195 20009 11207 20043
rect 11149 20003 11207 20009
rect 11885 20043 11943 20049
rect 11885 20009 11897 20043
rect 11931 20040 11943 20043
rect 18693 20043 18751 20049
rect 18693 20040 18705 20043
rect 11931 20012 15792 20040
rect 11931 20009 11943 20012
rect 11885 20003 11943 20009
rect 6365 19907 6423 19913
rect 6365 19873 6377 19907
rect 6411 19904 6423 19907
rect 6730 19904 6736 19916
rect 6411 19876 6736 19904
rect 6411 19873 6423 19876
rect 6365 19867 6423 19873
rect 6730 19864 6736 19876
rect 6788 19864 6794 19916
rect 8496 19836 8524 20000
rect 9122 19972 9128 19984
rect 7774 19808 8524 19836
rect 9048 19944 9128 19972
rect 6641 19771 6699 19777
rect 6641 19737 6653 19771
rect 6687 19768 6699 19771
rect 6687 19740 7052 19768
rect 6687 19737 6699 19740
rect 6641 19731 6699 19737
rect 7024 19712 7052 19740
rect 8404 19712 8432 19808
rect 8478 19728 8484 19780
rect 8536 19768 8542 19780
rect 9048 19768 9076 19944
rect 9122 19932 9128 19944
rect 9180 19932 9186 19984
rect 10873 19907 10931 19913
rect 10873 19873 10885 19907
rect 10919 19904 10931 19907
rect 11698 19904 11704 19916
rect 10919 19876 11704 19904
rect 10919 19873 10931 19876
rect 10873 19867 10931 19873
rect 11698 19864 11704 19876
rect 11756 19904 11762 19916
rect 12437 19907 12495 19913
rect 12437 19904 12449 19907
rect 11756 19876 12449 19904
rect 11756 19864 11762 19876
rect 12437 19873 12449 19876
rect 12483 19873 12495 19907
rect 12437 19867 12495 19873
rect 9122 19796 9128 19848
rect 9180 19796 9186 19848
rect 12342 19796 12348 19848
rect 12400 19796 12406 19848
rect 12618 19796 12624 19848
rect 12676 19836 12682 19848
rect 14277 19839 14335 19845
rect 14277 19836 14289 19839
rect 12676 19808 14289 19836
rect 12676 19796 12682 19808
rect 14277 19805 14289 19808
rect 14323 19805 14335 19839
rect 15764 19836 15792 20012
rect 16960 20012 18705 20040
rect 15930 19932 15936 19984
rect 15988 19972 15994 19984
rect 16960 19972 16988 20012
rect 18693 20009 18705 20012
rect 18739 20009 18751 20043
rect 18693 20003 18751 20009
rect 22186 20000 22192 20052
rect 22244 20040 22250 20052
rect 24213 20043 24271 20049
rect 24213 20040 24225 20043
rect 22244 20012 24225 20040
rect 22244 20000 22250 20012
rect 24213 20009 24225 20012
rect 24259 20040 24271 20043
rect 24946 20040 24952 20052
rect 24259 20012 24952 20040
rect 24259 20009 24271 20012
rect 24213 20003 24271 20009
rect 24946 20000 24952 20012
rect 25004 20000 25010 20052
rect 25225 20043 25283 20049
rect 25225 20009 25237 20043
rect 25271 20040 25283 20043
rect 25314 20040 25320 20052
rect 25271 20012 25320 20040
rect 25271 20009 25283 20012
rect 25225 20003 25283 20009
rect 25314 20000 25320 20012
rect 25372 20000 25378 20052
rect 15988 19944 16988 19972
rect 15988 19932 15994 19944
rect 17402 19932 17408 19984
rect 17460 19972 17466 19984
rect 17497 19975 17555 19981
rect 17497 19972 17509 19975
rect 17460 19944 17509 19972
rect 17460 19932 17466 19944
rect 17497 19941 17509 19944
rect 17543 19941 17555 19975
rect 17497 19935 17555 19941
rect 17770 19932 17776 19984
rect 17828 19972 17834 19984
rect 17828 19944 18092 19972
rect 17828 19932 17834 19944
rect 16025 19907 16083 19913
rect 16025 19873 16037 19907
rect 16071 19904 16083 19907
rect 16574 19904 16580 19916
rect 16071 19876 16580 19904
rect 16071 19873 16083 19876
rect 16025 19867 16083 19873
rect 16574 19864 16580 19876
rect 16632 19864 16638 19916
rect 17862 19864 17868 19916
rect 17920 19904 17926 19916
rect 18064 19913 18092 19944
rect 17957 19907 18015 19913
rect 17957 19904 17969 19907
rect 17920 19876 17969 19904
rect 17920 19864 17926 19876
rect 17957 19873 17969 19876
rect 18003 19873 18015 19907
rect 17957 19867 18015 19873
rect 18049 19907 18107 19913
rect 18049 19873 18061 19907
rect 18095 19873 18107 19907
rect 18049 19867 18107 19873
rect 19886 19864 19892 19916
rect 19944 19864 19950 19916
rect 16853 19839 16911 19845
rect 16853 19836 16865 19839
rect 15764 19808 16865 19836
rect 14277 19799 14335 19805
rect 16853 19805 16865 19808
rect 16899 19805 16911 19839
rect 16853 19799 16911 19805
rect 18877 19839 18935 19845
rect 18877 19805 18889 19839
rect 18923 19836 18935 19839
rect 19150 19836 19156 19848
rect 18923 19808 19156 19836
rect 18923 19805 18935 19808
rect 18877 19799 18935 19805
rect 19150 19796 19156 19808
rect 19208 19796 19214 19848
rect 22097 19839 22155 19845
rect 22097 19805 22109 19839
rect 22143 19805 22155 19839
rect 22097 19799 22155 19805
rect 24581 19839 24639 19845
rect 24581 19805 24593 19839
rect 24627 19836 24639 19839
rect 25130 19836 25136 19848
rect 24627 19808 25136 19836
rect 24627 19805 24639 19808
rect 24581 19799 24639 19805
rect 9401 19771 9459 19777
rect 9401 19768 9413 19771
rect 8536 19740 9413 19768
rect 8536 19728 8542 19740
rect 9401 19737 9413 19740
rect 9447 19737 9459 19771
rect 9858 19768 9864 19780
rect 9401 19731 9459 19737
rect 9508 19740 9864 19768
rect 9508 19712 9536 19740
rect 9858 19728 9864 19740
rect 9916 19728 9922 19780
rect 12253 19771 12311 19777
rect 12253 19768 12265 19771
rect 10704 19740 12265 19768
rect 7006 19660 7012 19712
rect 7064 19700 7070 19712
rect 7282 19700 7288 19712
rect 7064 19672 7288 19700
rect 7064 19660 7070 19672
rect 7282 19660 7288 19672
rect 7340 19660 7346 19712
rect 8113 19703 8171 19709
rect 8113 19669 8125 19703
rect 8159 19700 8171 19703
rect 8294 19700 8300 19712
rect 8159 19672 8300 19700
rect 8159 19669 8171 19672
rect 8113 19663 8171 19669
rect 8294 19660 8300 19672
rect 8352 19660 8358 19712
rect 8386 19660 8392 19712
rect 8444 19700 8450 19712
rect 9490 19700 9496 19712
rect 8444 19672 9496 19700
rect 8444 19660 8450 19672
rect 9490 19660 9496 19672
rect 9548 19660 9554 19712
rect 9674 19660 9680 19712
rect 9732 19700 9738 19712
rect 10704 19700 10732 19740
rect 12253 19737 12265 19740
rect 12299 19737 12311 19771
rect 12253 19731 12311 19737
rect 14550 19728 14556 19780
rect 14608 19728 14614 19780
rect 18414 19768 18420 19780
rect 14660 19740 15042 19768
rect 16684 19740 18420 19768
rect 9732 19672 10732 19700
rect 9732 19660 9738 19672
rect 10962 19660 10968 19712
rect 11020 19700 11026 19712
rect 13078 19700 13084 19712
rect 11020 19672 13084 19700
rect 11020 19660 11026 19672
rect 13078 19660 13084 19672
rect 13136 19700 13142 19712
rect 13354 19700 13360 19712
rect 13136 19672 13360 19700
rect 13136 19660 13142 19672
rect 13354 19660 13360 19672
rect 13412 19700 13418 19712
rect 14660 19700 14688 19740
rect 13412 19672 14688 19700
rect 14936 19700 14964 19740
rect 16684 19709 16712 19740
rect 18414 19728 18420 19740
rect 18472 19728 18478 19780
rect 20162 19728 20168 19780
rect 20220 19728 20226 19780
rect 22112 19768 22140 19799
rect 25130 19796 25136 19808
rect 25188 19796 25194 19848
rect 22278 19768 22284 19780
rect 20272 19740 20654 19768
rect 22112 19740 22284 19768
rect 16301 19703 16359 19709
rect 16301 19700 16313 19703
rect 14936 19672 16313 19700
rect 13412 19660 13418 19672
rect 16301 19669 16313 19672
rect 16347 19669 16359 19703
rect 16301 19663 16359 19669
rect 16669 19703 16727 19709
rect 16669 19669 16681 19703
rect 16715 19669 16727 19703
rect 16669 19663 16727 19669
rect 16758 19660 16764 19712
rect 16816 19700 16822 19712
rect 17865 19703 17923 19709
rect 17865 19700 17877 19703
rect 16816 19672 17877 19700
rect 16816 19660 16822 19672
rect 17865 19669 17877 19672
rect 17911 19669 17923 19703
rect 17865 19663 17923 19669
rect 19429 19703 19487 19709
rect 19429 19669 19441 19703
rect 19475 19700 19487 19703
rect 19610 19700 19616 19712
rect 19475 19672 19616 19700
rect 19475 19669 19487 19672
rect 19429 19663 19487 19669
rect 19610 19660 19616 19672
rect 19668 19700 19674 19712
rect 20272 19700 20300 19740
rect 22278 19728 22284 19740
rect 22336 19728 22342 19780
rect 22370 19728 22376 19780
rect 22428 19728 22434 19780
rect 24118 19768 24124 19780
rect 23598 19740 24124 19768
rect 24118 19728 24124 19740
rect 24176 19728 24182 19780
rect 19668 19672 20300 19700
rect 21637 19703 21695 19709
rect 19668 19660 19674 19672
rect 21637 19669 21649 19703
rect 21683 19700 21695 19703
rect 22002 19700 22008 19712
rect 21683 19672 22008 19700
rect 21683 19669 21695 19672
rect 21637 19663 21695 19669
rect 22002 19660 22008 19672
rect 22060 19660 22066 19712
rect 23845 19703 23903 19709
rect 23845 19669 23857 19703
rect 23891 19700 23903 19703
rect 23934 19700 23940 19712
rect 23891 19672 23940 19700
rect 23891 19669 23903 19672
rect 23845 19663 23903 19669
rect 23934 19660 23940 19672
rect 23992 19660 23998 19712
rect 1104 19610 25852 19632
rect 1104 19558 7950 19610
rect 8002 19558 8014 19610
rect 8066 19558 8078 19610
rect 8130 19558 8142 19610
rect 8194 19558 8206 19610
rect 8258 19558 17950 19610
rect 18002 19558 18014 19610
rect 18066 19558 18078 19610
rect 18130 19558 18142 19610
rect 18194 19558 18206 19610
rect 18258 19558 25852 19610
rect 1104 19536 25852 19558
rect 7558 19496 7564 19508
rect 7484 19468 7564 19496
rect 6822 19320 6828 19372
rect 6880 19360 6886 19372
rect 7484 19369 7512 19468
rect 7558 19456 7564 19468
rect 7616 19496 7622 19508
rect 9122 19496 9128 19508
rect 7616 19468 9128 19496
rect 7616 19456 7622 19468
rect 9122 19456 9128 19468
rect 9180 19456 9186 19508
rect 9217 19499 9275 19505
rect 9217 19465 9229 19499
rect 9263 19496 9275 19499
rect 9306 19496 9312 19508
rect 9263 19468 9312 19496
rect 9263 19465 9275 19468
rect 9217 19459 9275 19465
rect 9306 19456 9312 19468
rect 9364 19456 9370 19508
rect 9490 19456 9496 19508
rect 9548 19456 9554 19508
rect 10137 19499 10195 19505
rect 10137 19465 10149 19499
rect 10183 19496 10195 19499
rect 10318 19496 10324 19508
rect 10183 19468 10324 19496
rect 10183 19465 10195 19468
rect 10137 19459 10195 19465
rect 10318 19456 10324 19468
rect 10376 19456 10382 19508
rect 10597 19499 10655 19505
rect 10597 19465 10609 19499
rect 10643 19496 10655 19499
rect 12710 19496 12716 19508
rect 10643 19468 12716 19496
rect 10643 19465 10655 19468
rect 10597 19459 10655 19465
rect 12710 19456 12716 19468
rect 12768 19456 12774 19508
rect 12802 19456 12808 19508
rect 12860 19496 12866 19508
rect 14093 19499 14151 19505
rect 14093 19496 14105 19499
rect 12860 19468 14105 19496
rect 12860 19456 12866 19468
rect 14093 19465 14105 19468
rect 14139 19465 14151 19499
rect 15657 19499 15715 19505
rect 14093 19459 14151 19465
rect 14200 19468 14780 19496
rect 9508 19428 9536 19456
rect 12618 19428 12624 19440
rect 8970 19400 9536 19428
rect 12360 19400 12624 19428
rect 7469 19363 7527 19369
rect 7469 19360 7481 19363
rect 6880 19332 7481 19360
rect 6880 19320 6886 19332
rect 7469 19329 7481 19332
rect 7515 19329 7527 19363
rect 7469 19323 7527 19329
rect 9861 19363 9919 19369
rect 9861 19329 9873 19363
rect 9907 19360 9919 19363
rect 10318 19360 10324 19372
rect 9907 19332 10324 19360
rect 9907 19329 9919 19332
rect 9861 19323 9919 19329
rect 10318 19320 10324 19332
rect 10376 19360 10382 19372
rect 12360 19369 12388 19400
rect 12618 19388 12624 19400
rect 12676 19388 12682 19440
rect 13078 19388 13084 19440
rect 13136 19388 13142 19440
rect 13906 19388 13912 19440
rect 13964 19428 13970 19440
rect 14200 19428 14228 19468
rect 14642 19428 14648 19440
rect 13964 19400 14228 19428
rect 14568 19400 14648 19428
rect 13964 19388 13970 19400
rect 14568 19369 14596 19400
rect 14642 19388 14648 19400
rect 14700 19388 14706 19440
rect 14752 19428 14780 19468
rect 15657 19465 15669 19499
rect 15703 19496 15715 19499
rect 16022 19496 16028 19508
rect 15703 19468 16028 19496
rect 15703 19465 15715 19468
rect 15657 19459 15715 19465
rect 16022 19456 16028 19468
rect 16080 19456 16086 19508
rect 16390 19456 16396 19508
rect 16448 19496 16454 19508
rect 16758 19496 16764 19508
rect 16448 19468 16764 19496
rect 16448 19456 16454 19468
rect 16758 19456 16764 19468
rect 16816 19456 16822 19508
rect 16853 19499 16911 19505
rect 16853 19465 16865 19499
rect 16899 19465 16911 19499
rect 16853 19459 16911 19465
rect 16868 19428 16896 19459
rect 16942 19456 16948 19508
rect 17000 19496 17006 19508
rect 17313 19499 17371 19505
rect 17313 19496 17325 19499
rect 17000 19468 17325 19496
rect 17000 19456 17006 19468
rect 17313 19465 17325 19468
rect 17359 19465 17371 19499
rect 17313 19459 17371 19465
rect 18782 19456 18788 19508
rect 18840 19456 18846 19508
rect 18966 19456 18972 19508
rect 19024 19496 19030 19508
rect 20073 19499 20131 19505
rect 20073 19496 20085 19499
rect 19024 19468 20085 19496
rect 19024 19456 19030 19468
rect 20073 19465 20085 19468
rect 20119 19465 20131 19499
rect 20073 19459 20131 19465
rect 20438 19456 20444 19508
rect 20496 19456 20502 19508
rect 20533 19499 20591 19505
rect 20533 19465 20545 19499
rect 20579 19496 20591 19499
rect 20714 19496 20720 19508
rect 20579 19468 20720 19496
rect 20579 19465 20591 19468
rect 20533 19459 20591 19465
rect 20714 19456 20720 19468
rect 20772 19456 20778 19508
rect 21450 19456 21456 19508
rect 21508 19496 21514 19508
rect 22189 19499 22247 19505
rect 22189 19496 22201 19499
rect 21508 19468 22201 19496
rect 21508 19456 21514 19468
rect 22189 19465 22201 19468
rect 22235 19465 22247 19499
rect 22189 19459 22247 19465
rect 22649 19499 22707 19505
rect 22649 19465 22661 19499
rect 22695 19496 22707 19499
rect 24486 19496 24492 19508
rect 22695 19468 24492 19496
rect 22695 19465 22707 19468
rect 22649 19459 22707 19465
rect 24486 19456 24492 19468
rect 24544 19456 24550 19508
rect 20254 19428 20260 19440
rect 14752 19400 15976 19428
rect 16868 19400 20260 19428
rect 10505 19363 10563 19369
rect 10505 19360 10517 19363
rect 10376 19332 10517 19360
rect 10376 19320 10382 19332
rect 10505 19329 10517 19332
rect 10551 19329 10563 19363
rect 10505 19323 10563 19329
rect 12345 19363 12403 19369
rect 12345 19329 12357 19363
rect 12391 19329 12403 19363
rect 12345 19323 12403 19329
rect 14553 19363 14611 19369
rect 14553 19329 14565 19363
rect 14599 19329 14611 19363
rect 15197 19363 15255 19369
rect 15197 19360 15209 19363
rect 14553 19323 14611 19329
rect 14660 19332 15209 19360
rect 7745 19295 7803 19301
rect 7745 19261 7757 19295
rect 7791 19292 7803 19295
rect 9766 19292 9772 19304
rect 7791 19264 9772 19292
rect 7791 19261 7803 19264
rect 7745 19255 7803 19261
rect 9766 19252 9772 19264
rect 9824 19252 9830 19304
rect 10689 19295 10747 19301
rect 10689 19261 10701 19295
rect 10735 19292 10747 19295
rect 11146 19292 11152 19304
rect 10735 19264 11152 19292
rect 10735 19261 10747 19264
rect 10689 19255 10747 19261
rect 8772 19196 9628 19224
rect 3510 19116 3516 19168
rect 3568 19156 3574 19168
rect 8772 19156 8800 19196
rect 3568 19128 8800 19156
rect 9600 19156 9628 19196
rect 10502 19184 10508 19236
rect 10560 19224 10566 19236
rect 10704 19224 10732 19255
rect 11146 19252 11152 19264
rect 11204 19252 11210 19304
rect 12621 19295 12679 19301
rect 12621 19261 12633 19295
rect 12667 19292 12679 19295
rect 14660 19292 14688 19332
rect 15197 19329 15209 19332
rect 15243 19329 15255 19363
rect 15197 19323 15255 19329
rect 15841 19363 15899 19369
rect 15841 19329 15853 19363
rect 15887 19329 15899 19363
rect 15948 19360 15976 19400
rect 20254 19388 20260 19400
rect 20312 19388 20318 19440
rect 24118 19388 24124 19440
rect 24176 19388 24182 19440
rect 17221 19363 17279 19369
rect 17221 19360 17233 19363
rect 15948 19332 17233 19360
rect 15841 19323 15899 19329
rect 17221 19329 17233 19332
rect 17267 19329 17279 19363
rect 17221 19323 17279 19329
rect 12667 19264 14688 19292
rect 12667 19261 12679 19264
rect 12621 19255 12679 19261
rect 10560 19196 10732 19224
rect 10560 19184 10566 19196
rect 10962 19184 10968 19236
rect 11020 19224 11026 19236
rect 11517 19227 11575 19233
rect 11517 19224 11529 19227
rect 11020 19196 11529 19224
rect 11020 19184 11026 19196
rect 11517 19193 11529 19196
rect 11563 19193 11575 19227
rect 11517 19187 11575 19193
rect 14090 19184 14096 19236
rect 14148 19224 14154 19236
rect 15856 19224 15884 19323
rect 17770 19320 17776 19372
rect 17828 19360 17834 19372
rect 18141 19363 18199 19369
rect 18141 19360 18153 19363
rect 17828 19332 18153 19360
rect 17828 19320 17834 19332
rect 18141 19329 18153 19332
rect 18187 19329 18199 19363
rect 18141 19323 18199 19329
rect 19242 19320 19248 19372
rect 19300 19360 19306 19372
rect 19429 19363 19487 19369
rect 19429 19360 19441 19363
rect 19300 19332 19441 19360
rect 19300 19320 19306 19332
rect 19429 19329 19441 19332
rect 19475 19329 19487 19363
rect 19429 19323 19487 19329
rect 21453 19363 21511 19369
rect 21453 19329 21465 19363
rect 21499 19360 21511 19363
rect 22462 19360 22468 19372
rect 21499 19332 22468 19360
rect 21499 19329 21511 19332
rect 21453 19323 21511 19329
rect 22462 19320 22468 19332
rect 22520 19320 22526 19372
rect 22554 19320 22560 19372
rect 22612 19320 22618 19372
rect 16574 19252 16580 19304
rect 16632 19292 16638 19304
rect 17405 19295 17463 19301
rect 17405 19292 17417 19295
rect 16632 19264 17417 19292
rect 16632 19252 16638 19264
rect 17405 19261 17417 19264
rect 17451 19261 17463 19295
rect 17405 19255 17463 19261
rect 20717 19295 20775 19301
rect 20717 19261 20729 19295
rect 20763 19292 20775 19295
rect 22002 19292 22008 19304
rect 20763 19264 22008 19292
rect 20763 19261 20775 19264
rect 20717 19255 20775 19261
rect 22002 19252 22008 19264
rect 22060 19252 22066 19304
rect 22738 19252 22744 19304
rect 22796 19252 22802 19304
rect 23290 19252 23296 19304
rect 23348 19292 23354 19304
rect 23385 19295 23443 19301
rect 23385 19292 23397 19295
rect 23348 19264 23397 19292
rect 23348 19252 23354 19264
rect 23385 19261 23397 19264
rect 23431 19261 23443 19295
rect 23385 19255 23443 19261
rect 23661 19295 23719 19301
rect 23661 19261 23673 19295
rect 23707 19292 23719 19295
rect 25222 19292 25228 19304
rect 23707 19264 25228 19292
rect 23707 19261 23719 19264
rect 23661 19255 23719 19261
rect 25222 19252 25228 19264
rect 25280 19252 25286 19304
rect 14148 19196 15884 19224
rect 14148 19184 14154 19196
rect 21082 19184 21088 19236
rect 21140 19224 21146 19236
rect 21821 19227 21879 19233
rect 21821 19224 21833 19227
rect 21140 19196 21833 19224
rect 21140 19184 21146 19196
rect 21821 19193 21833 19196
rect 21867 19193 21879 19227
rect 25409 19227 25467 19233
rect 25409 19224 25421 19227
rect 21821 19187 21879 19193
rect 24688 19196 25421 19224
rect 11330 19156 11336 19168
rect 9600 19128 11336 19156
rect 3568 19116 3574 19128
rect 11330 19116 11336 19128
rect 11388 19116 11394 19168
rect 14366 19116 14372 19168
rect 14424 19156 14430 19168
rect 18782 19156 18788 19168
rect 14424 19128 18788 19156
rect 14424 19116 14430 19128
rect 18782 19116 18788 19128
rect 18840 19116 18846 19168
rect 19242 19116 19248 19168
rect 19300 19116 19306 19168
rect 19702 19116 19708 19168
rect 19760 19116 19766 19168
rect 21266 19116 21272 19168
rect 21324 19116 21330 19168
rect 22738 19116 22744 19168
rect 22796 19156 22802 19168
rect 23750 19156 23756 19168
rect 22796 19128 23756 19156
rect 22796 19116 22802 19128
rect 23750 19116 23756 19128
rect 23808 19116 23814 19168
rect 24118 19116 24124 19168
rect 24176 19156 24182 19168
rect 24688 19156 24716 19196
rect 25409 19193 25421 19196
rect 25455 19193 25467 19227
rect 25409 19187 25467 19193
rect 24176 19128 24716 19156
rect 24176 19116 24182 19128
rect 25130 19116 25136 19168
rect 25188 19116 25194 19168
rect 1104 19066 25852 19088
rect 1104 19014 2950 19066
rect 3002 19014 3014 19066
rect 3066 19014 3078 19066
rect 3130 19014 3142 19066
rect 3194 19014 3206 19066
rect 3258 19014 12950 19066
rect 13002 19014 13014 19066
rect 13066 19014 13078 19066
rect 13130 19014 13142 19066
rect 13194 19014 13206 19066
rect 13258 19014 22950 19066
rect 23002 19014 23014 19066
rect 23066 19014 23078 19066
rect 23130 19014 23142 19066
rect 23194 19014 23206 19066
rect 23258 19014 25852 19066
rect 1104 18992 25852 19014
rect 9769 18955 9827 18961
rect 9769 18921 9781 18955
rect 9815 18952 9827 18955
rect 9815 18924 11100 18952
rect 9815 18921 9827 18924
rect 9769 18915 9827 18921
rect 10965 18887 11023 18893
rect 10965 18853 10977 18887
rect 11011 18853 11023 18887
rect 11072 18884 11100 18924
rect 11330 18912 11336 18964
rect 11388 18952 11394 18964
rect 22186 18952 22192 18964
rect 11388 18924 22192 18952
rect 11388 18912 11394 18924
rect 22186 18912 22192 18924
rect 22244 18912 22250 18964
rect 25317 18955 25375 18961
rect 25317 18921 25329 18955
rect 25363 18952 25375 18955
rect 25406 18952 25412 18964
rect 25363 18924 25412 18952
rect 25363 18921 25375 18924
rect 25317 18915 25375 18921
rect 25406 18912 25412 18924
rect 25464 18912 25470 18964
rect 14090 18884 14096 18896
rect 11072 18856 14096 18884
rect 10965 18847 11023 18853
rect 6822 18776 6828 18828
rect 6880 18776 6886 18828
rect 7101 18819 7159 18825
rect 7101 18785 7113 18819
rect 7147 18816 7159 18819
rect 7190 18816 7196 18828
rect 7147 18788 7196 18816
rect 7147 18785 7159 18788
rect 7101 18779 7159 18785
rect 7190 18776 7196 18788
rect 7248 18776 7254 18828
rect 8294 18776 8300 18828
rect 8352 18816 8358 18828
rect 10321 18819 10379 18825
rect 10321 18816 10333 18819
rect 8352 18788 10333 18816
rect 8352 18776 8358 18788
rect 10321 18785 10333 18788
rect 10367 18785 10379 18819
rect 10980 18816 11008 18847
rect 14090 18844 14096 18856
rect 14148 18844 14154 18896
rect 14277 18887 14335 18893
rect 14277 18853 14289 18887
rect 14323 18853 14335 18887
rect 14277 18847 14335 18853
rect 17957 18887 18015 18893
rect 17957 18853 17969 18887
rect 18003 18884 18015 18887
rect 19058 18884 19064 18896
rect 18003 18856 19064 18884
rect 18003 18853 18015 18856
rect 17957 18847 18015 18853
rect 10980 18788 11468 18816
rect 10321 18779 10379 18785
rect 8386 18748 8392 18760
rect 8234 18720 8392 18748
rect 8386 18708 8392 18720
rect 8444 18748 8450 18760
rect 8754 18748 8760 18760
rect 8444 18720 8760 18748
rect 8444 18708 8450 18720
rect 8754 18708 8760 18720
rect 8812 18708 8818 18760
rect 10778 18708 10784 18760
rect 10836 18748 10842 18760
rect 10962 18748 10968 18760
rect 10836 18720 10968 18748
rect 10836 18708 10842 18720
rect 10962 18708 10968 18720
rect 11020 18748 11026 18760
rect 11440 18748 11468 18788
rect 11514 18776 11520 18828
rect 11572 18776 11578 18828
rect 12526 18748 12532 18760
rect 11020 18720 11376 18748
rect 11440 18720 12532 18748
rect 11020 18708 11026 18720
rect 10137 18683 10195 18689
rect 10137 18680 10149 18683
rect 8404 18652 10149 18680
rect 7374 18572 7380 18624
rect 7432 18612 7438 18624
rect 8404 18612 8432 18652
rect 10137 18649 10149 18652
rect 10183 18649 10195 18683
rect 10137 18643 10195 18649
rect 10229 18683 10287 18689
rect 10229 18649 10241 18683
rect 10275 18680 10287 18683
rect 11238 18680 11244 18692
rect 10275 18652 11244 18680
rect 10275 18649 10287 18652
rect 10229 18643 10287 18649
rect 11238 18640 11244 18652
rect 11296 18640 11302 18692
rect 11348 18680 11376 18720
rect 12526 18708 12532 18720
rect 12584 18708 12590 18760
rect 14292 18748 14320 18847
rect 19058 18844 19064 18856
rect 19116 18844 19122 18896
rect 20162 18844 20168 18896
rect 20220 18884 20226 18896
rect 21361 18887 21419 18893
rect 21361 18884 21373 18887
rect 20220 18856 21373 18884
rect 20220 18844 20226 18856
rect 21361 18853 21373 18856
rect 21407 18853 21419 18887
rect 21361 18847 21419 18853
rect 14734 18776 14740 18828
rect 14792 18816 14798 18828
rect 14829 18819 14887 18825
rect 14829 18816 14841 18819
rect 14792 18788 14841 18816
rect 14792 18776 14798 18788
rect 14829 18785 14841 18788
rect 14875 18785 14887 18819
rect 14829 18779 14887 18785
rect 16298 18776 16304 18828
rect 16356 18816 16362 18828
rect 17126 18816 17132 18828
rect 16356 18788 17132 18816
rect 16356 18776 16362 18788
rect 17126 18776 17132 18788
rect 17184 18776 17190 18828
rect 17218 18776 17224 18828
rect 17276 18776 17282 18828
rect 17405 18819 17463 18825
rect 17405 18785 17417 18819
rect 17451 18816 17463 18819
rect 17770 18816 17776 18828
rect 17451 18788 17776 18816
rect 17451 18785 17463 18788
rect 17405 18779 17463 18785
rect 17770 18776 17776 18788
rect 17828 18776 17834 18828
rect 18509 18819 18567 18825
rect 18509 18816 18521 18819
rect 17880 18788 18521 18816
rect 15286 18748 15292 18760
rect 14292 18720 15292 18748
rect 15286 18708 15292 18720
rect 15344 18708 15350 18760
rect 16209 18751 16267 18757
rect 16209 18717 16221 18751
rect 16255 18748 16267 18751
rect 17494 18748 17500 18760
rect 16255 18720 17500 18748
rect 16255 18717 16267 18720
rect 16209 18711 16267 18717
rect 17494 18708 17500 18720
rect 17552 18708 17558 18760
rect 17586 18708 17592 18760
rect 17644 18748 17650 18760
rect 17880 18748 17908 18788
rect 18509 18785 18521 18788
rect 18555 18785 18567 18819
rect 18509 18779 18567 18785
rect 18782 18776 18788 18828
rect 18840 18816 18846 18828
rect 21821 18819 21879 18825
rect 18840 18788 21312 18816
rect 18840 18776 18846 18788
rect 17644 18720 17908 18748
rect 18417 18751 18475 18757
rect 17644 18708 17650 18720
rect 18417 18717 18429 18751
rect 18463 18748 18475 18751
rect 18598 18748 18604 18760
rect 18463 18720 18604 18748
rect 18463 18717 18475 18720
rect 18417 18711 18475 18717
rect 18598 18708 18604 18720
rect 18656 18708 18662 18760
rect 18690 18708 18696 18760
rect 18748 18748 18754 18760
rect 19429 18751 19487 18757
rect 19429 18748 19441 18751
rect 18748 18720 19441 18748
rect 18748 18708 18754 18720
rect 19429 18717 19441 18720
rect 19475 18717 19487 18751
rect 19429 18711 19487 18717
rect 20714 18708 20720 18760
rect 20772 18748 20778 18760
rect 21174 18748 21180 18760
rect 20772 18720 21180 18748
rect 20772 18708 20778 18720
rect 21174 18708 21180 18720
rect 21232 18708 21238 18760
rect 21284 18748 21312 18788
rect 21821 18785 21833 18819
rect 21867 18816 21879 18819
rect 22554 18816 22560 18828
rect 21867 18788 22560 18816
rect 21867 18785 21879 18788
rect 21821 18779 21879 18785
rect 22554 18776 22560 18788
rect 22612 18776 22618 18828
rect 23382 18776 23388 18828
rect 23440 18816 23446 18828
rect 23477 18819 23535 18825
rect 23477 18816 23489 18819
rect 23440 18788 23489 18816
rect 23440 18776 23446 18788
rect 23477 18785 23489 18788
rect 23523 18785 23535 18819
rect 23477 18779 23535 18785
rect 22649 18751 22707 18757
rect 22649 18748 22661 18751
rect 21284 18720 22661 18748
rect 22649 18717 22661 18720
rect 22695 18717 22707 18751
rect 22649 18711 22707 18717
rect 24673 18751 24731 18757
rect 24673 18717 24685 18751
rect 24719 18748 24731 18751
rect 25314 18748 25320 18760
rect 24719 18720 25320 18748
rect 24719 18717 24731 18720
rect 24673 18711 24731 18717
rect 25314 18708 25320 18720
rect 25372 18708 25378 18760
rect 11425 18683 11483 18689
rect 11425 18680 11437 18683
rect 11348 18652 11437 18680
rect 11425 18649 11437 18652
rect 11471 18649 11483 18683
rect 11425 18643 11483 18649
rect 12161 18683 12219 18689
rect 12161 18649 12173 18683
rect 12207 18680 12219 18683
rect 12207 18652 12434 18680
rect 12207 18649 12219 18652
rect 12161 18643 12219 18649
rect 7432 18584 8432 18612
rect 7432 18572 7438 18584
rect 8478 18572 8484 18624
rect 8536 18612 8542 18624
rect 8573 18615 8631 18621
rect 8573 18612 8585 18615
rect 8536 18584 8585 18612
rect 8536 18572 8542 18584
rect 8573 18581 8585 18584
rect 8619 18581 8631 18615
rect 8573 18575 8631 18581
rect 9125 18615 9183 18621
rect 9125 18581 9137 18615
rect 9171 18612 9183 18615
rect 9490 18612 9496 18624
rect 9171 18584 9496 18612
rect 9171 18581 9183 18584
rect 9125 18575 9183 18581
rect 9490 18572 9496 18584
rect 9548 18572 9554 18624
rect 11333 18615 11391 18621
rect 11333 18581 11345 18615
rect 11379 18612 11391 18615
rect 11698 18612 11704 18624
rect 11379 18584 11704 18612
rect 11379 18581 11391 18584
rect 11333 18575 11391 18581
rect 11698 18572 11704 18584
rect 11756 18572 11762 18624
rect 12406 18612 12434 18652
rect 12618 18640 12624 18692
rect 12676 18680 12682 18692
rect 12897 18683 12955 18689
rect 12897 18680 12909 18683
rect 12676 18652 12909 18680
rect 12676 18640 12682 18652
rect 12897 18649 12909 18652
rect 12943 18649 12955 18683
rect 14737 18683 14795 18689
rect 14737 18680 14749 18683
rect 12897 18643 12955 18649
rect 13648 18652 14749 18680
rect 13648 18624 13676 18652
rect 14737 18649 14749 18652
rect 14783 18649 14795 18683
rect 14737 18643 14795 18649
rect 15746 18640 15752 18692
rect 15804 18680 15810 18692
rect 20806 18680 20812 18692
rect 15804 18652 20812 18680
rect 15804 18640 15810 18652
rect 20806 18640 20812 18652
rect 20864 18640 20870 18692
rect 21910 18640 21916 18692
rect 21968 18680 21974 18692
rect 22738 18680 22744 18692
rect 21968 18652 22744 18680
rect 21968 18640 21974 18652
rect 22738 18640 22744 18652
rect 22796 18640 22802 18692
rect 13446 18612 13452 18624
rect 12406 18584 13452 18612
rect 13446 18572 13452 18584
rect 13504 18572 13510 18624
rect 13630 18572 13636 18624
rect 13688 18572 13694 18624
rect 13909 18615 13967 18621
rect 13909 18581 13921 18615
rect 13955 18612 13967 18615
rect 13998 18612 14004 18624
rect 13955 18584 14004 18612
rect 13955 18581 13967 18584
rect 13909 18575 13967 18581
rect 13998 18572 14004 18584
rect 14056 18572 14062 18624
rect 14642 18572 14648 18624
rect 14700 18572 14706 18624
rect 16025 18615 16083 18621
rect 16025 18581 16037 18615
rect 16071 18612 16083 18615
rect 16114 18612 16120 18624
rect 16071 18584 16120 18612
rect 16071 18581 16083 18584
rect 16025 18575 16083 18581
rect 16114 18572 16120 18584
rect 16172 18572 16178 18624
rect 16761 18615 16819 18621
rect 16761 18581 16773 18615
rect 16807 18612 16819 18615
rect 17034 18612 17040 18624
rect 16807 18584 17040 18612
rect 16807 18581 16819 18584
rect 16761 18575 16819 18581
rect 17034 18572 17040 18584
rect 17092 18572 17098 18624
rect 17126 18572 17132 18624
rect 17184 18612 17190 18624
rect 18325 18615 18383 18621
rect 18325 18612 18337 18615
rect 17184 18584 18337 18612
rect 17184 18572 17190 18584
rect 18325 18581 18337 18584
rect 18371 18612 18383 18615
rect 18969 18615 19027 18621
rect 18969 18612 18981 18615
rect 18371 18584 18981 18612
rect 18371 18581 18383 18584
rect 18325 18575 18383 18581
rect 18969 18581 18981 18584
rect 19015 18612 19027 18615
rect 19702 18612 19708 18624
rect 19015 18584 19708 18612
rect 19015 18581 19027 18584
rect 18969 18575 19027 18581
rect 19702 18572 19708 18584
rect 19760 18572 19766 18624
rect 20070 18572 20076 18624
rect 20128 18572 20134 18624
rect 20438 18572 20444 18624
rect 20496 18572 20502 18624
rect 22186 18572 22192 18624
rect 22244 18612 22250 18624
rect 22281 18615 22339 18621
rect 22281 18612 22293 18615
rect 22244 18584 22293 18612
rect 22244 18572 22250 18584
rect 22281 18581 22293 18584
rect 22327 18581 22339 18615
rect 22281 18575 22339 18581
rect 1104 18522 25852 18544
rect 1104 18470 7950 18522
rect 8002 18470 8014 18522
rect 8066 18470 8078 18522
rect 8130 18470 8142 18522
rect 8194 18470 8206 18522
rect 8258 18470 17950 18522
rect 18002 18470 18014 18522
rect 18066 18470 18078 18522
rect 18130 18470 18142 18522
rect 18194 18470 18206 18522
rect 18258 18470 25852 18522
rect 1104 18448 25852 18470
rect 7929 18411 7987 18417
rect 7929 18377 7941 18411
rect 7975 18408 7987 18411
rect 8662 18408 8668 18420
rect 7975 18380 8668 18408
rect 7975 18377 7987 18380
rect 7929 18371 7987 18377
rect 8662 18368 8668 18380
rect 8720 18368 8726 18420
rect 9582 18368 9588 18420
rect 9640 18408 9646 18420
rect 11514 18408 11520 18420
rect 9640 18380 11520 18408
rect 9640 18368 9646 18380
rect 11514 18368 11520 18380
rect 11572 18368 11578 18420
rect 11698 18368 11704 18420
rect 11756 18368 11762 18420
rect 12710 18368 12716 18420
rect 12768 18408 12774 18420
rect 13173 18411 13231 18417
rect 13173 18408 13185 18411
rect 12768 18380 13185 18408
rect 12768 18368 12774 18380
rect 13173 18377 13185 18380
rect 13219 18377 13231 18411
rect 13173 18371 13231 18377
rect 13630 18368 13636 18420
rect 13688 18368 13694 18420
rect 14550 18368 14556 18420
rect 14608 18408 14614 18420
rect 15013 18411 15071 18417
rect 15013 18408 15025 18411
rect 14608 18380 15025 18408
rect 14608 18368 14614 18380
rect 15013 18377 15025 18380
rect 15059 18377 15071 18411
rect 15013 18371 15071 18377
rect 15194 18368 15200 18420
rect 15252 18408 15258 18420
rect 20070 18408 20076 18420
rect 15252 18380 16896 18408
rect 15252 18368 15258 18380
rect 9401 18343 9459 18349
rect 9401 18309 9413 18343
rect 9447 18340 9459 18343
rect 9600 18340 9628 18368
rect 9447 18312 9628 18340
rect 9447 18309 9459 18312
rect 9401 18303 9459 18309
rect 9858 18300 9864 18352
rect 9916 18300 9922 18352
rect 11146 18300 11152 18352
rect 11204 18300 11210 18352
rect 13648 18340 13676 18368
rect 16206 18340 16212 18352
rect 12820 18312 13676 18340
rect 14384 18312 16212 18340
rect 8294 18232 8300 18284
rect 8352 18232 8358 18284
rect 8386 18164 8392 18216
rect 8444 18164 8450 18216
rect 8481 18207 8539 18213
rect 8481 18173 8493 18207
rect 8527 18173 8539 18207
rect 8481 18167 8539 18173
rect 7742 18096 7748 18148
rect 7800 18136 7806 18148
rect 8496 18136 8524 18167
rect 9122 18164 9128 18216
rect 9180 18204 9186 18216
rect 9398 18204 9404 18216
rect 9180 18176 9404 18204
rect 9180 18164 9186 18176
rect 9398 18164 9404 18176
rect 9456 18164 9462 18216
rect 12820 18145 12848 18312
rect 13541 18275 13599 18281
rect 13541 18241 13553 18275
rect 13587 18241 13599 18275
rect 13541 18235 13599 18241
rect 12805 18139 12863 18145
rect 12805 18136 12817 18139
rect 7800 18108 8524 18136
rect 11440 18108 12817 18136
rect 7800 18096 7806 18108
rect 5166 18028 5172 18080
rect 5224 18068 5230 18080
rect 11440 18068 11468 18108
rect 12805 18105 12817 18108
rect 12851 18105 12863 18139
rect 13556 18136 13584 18235
rect 13630 18232 13636 18284
rect 13688 18272 13694 18284
rect 13906 18272 13912 18284
rect 13688 18244 13912 18272
rect 13688 18232 13694 18244
rect 13906 18232 13912 18244
rect 13964 18232 13970 18284
rect 14384 18281 14412 18312
rect 16206 18300 16212 18312
rect 16264 18300 16270 18352
rect 16868 18284 16896 18380
rect 17144 18380 20076 18408
rect 17144 18349 17172 18380
rect 20070 18368 20076 18380
rect 20128 18368 20134 18420
rect 22370 18368 22376 18420
rect 22428 18408 22434 18420
rect 22649 18411 22707 18417
rect 22649 18408 22661 18411
rect 22428 18380 22661 18408
rect 22428 18368 22434 18380
rect 22649 18377 22661 18380
rect 22695 18377 22707 18411
rect 25682 18408 25688 18420
rect 22649 18371 22707 18377
rect 23492 18380 25688 18408
rect 17129 18343 17187 18349
rect 17129 18309 17141 18343
rect 17175 18309 17187 18343
rect 17129 18303 17187 18309
rect 17862 18300 17868 18352
rect 17920 18300 17926 18352
rect 18598 18300 18604 18352
rect 18656 18340 18662 18352
rect 18877 18343 18935 18349
rect 18877 18340 18889 18343
rect 18656 18312 18889 18340
rect 18656 18300 18662 18312
rect 18877 18309 18889 18312
rect 18923 18309 18935 18343
rect 20990 18340 20996 18352
rect 18877 18303 18935 18309
rect 19628 18312 20996 18340
rect 14369 18275 14427 18281
rect 14369 18241 14381 18275
rect 14415 18241 14427 18275
rect 14369 18235 14427 18241
rect 15473 18275 15531 18281
rect 15473 18241 15485 18275
rect 15519 18272 15531 18275
rect 15519 18244 16804 18272
rect 15519 18241 15531 18244
rect 15473 18235 15531 18241
rect 13725 18207 13783 18213
rect 13725 18173 13737 18207
rect 13771 18204 13783 18207
rect 13771 18176 13952 18204
rect 13771 18173 13783 18176
rect 13725 18167 13783 18173
rect 13814 18136 13820 18148
rect 13556 18108 13820 18136
rect 12805 18099 12863 18105
rect 13814 18096 13820 18108
rect 13872 18096 13878 18148
rect 5224 18040 11468 18068
rect 5224 18028 5230 18040
rect 11514 18028 11520 18080
rect 11572 18068 11578 18080
rect 12526 18068 12532 18080
rect 11572 18040 12532 18068
rect 11572 18028 11578 18040
rect 12526 18028 12532 18040
rect 12584 18068 12590 18080
rect 13924 18068 13952 18176
rect 15746 18164 15752 18216
rect 15804 18164 15810 18216
rect 16776 18204 16804 18244
rect 16850 18232 16856 18284
rect 16908 18232 16914 18284
rect 19628 18281 19656 18312
rect 20990 18300 20996 18312
rect 21048 18300 21054 18352
rect 21269 18343 21327 18349
rect 21269 18309 21281 18343
rect 21315 18340 21327 18343
rect 21634 18340 21640 18352
rect 21315 18312 21640 18340
rect 21315 18309 21327 18312
rect 21269 18303 21327 18309
rect 21634 18300 21640 18312
rect 21692 18340 21698 18352
rect 23492 18340 23520 18380
rect 25682 18368 25688 18380
rect 25740 18368 25746 18420
rect 21692 18312 23520 18340
rect 21692 18300 21698 18312
rect 23566 18300 23572 18352
rect 23624 18300 23630 18352
rect 19613 18275 19671 18281
rect 19613 18241 19625 18275
rect 19659 18241 19671 18275
rect 19613 18235 19671 18241
rect 20254 18232 20260 18284
rect 20312 18232 20318 18284
rect 22002 18232 22008 18284
rect 22060 18232 22066 18284
rect 19242 18204 19248 18216
rect 16776 18176 19248 18204
rect 19242 18164 19248 18176
rect 19300 18164 19306 18216
rect 20438 18164 20444 18216
rect 20496 18204 20502 18216
rect 20990 18204 20996 18216
rect 20496 18176 20996 18204
rect 20496 18164 20502 18176
rect 20990 18164 20996 18176
rect 21048 18204 21054 18216
rect 22186 18204 22192 18216
rect 21048 18176 22192 18204
rect 21048 18164 21054 18176
rect 22186 18164 22192 18176
rect 22244 18164 22250 18216
rect 22278 18164 22284 18216
rect 22336 18204 22342 18216
rect 23290 18204 23296 18216
rect 22336 18176 23296 18204
rect 22336 18164 22342 18176
rect 23290 18164 23296 18176
rect 23348 18164 23354 18216
rect 24118 18204 24124 18216
rect 23400 18176 24124 18204
rect 20717 18139 20775 18145
rect 18156 18108 18920 18136
rect 12584 18040 13952 18068
rect 12584 18028 12590 18040
rect 17218 18028 17224 18080
rect 17276 18068 17282 18080
rect 18156 18068 18184 18108
rect 18892 18080 18920 18108
rect 20717 18105 20729 18139
rect 20763 18136 20775 18139
rect 21910 18136 21916 18148
rect 20763 18108 21916 18136
rect 20763 18105 20775 18108
rect 20717 18099 20775 18105
rect 21910 18096 21916 18108
rect 21968 18096 21974 18148
rect 22204 18136 22232 18164
rect 22925 18139 22983 18145
rect 22925 18136 22937 18139
rect 22204 18108 22937 18136
rect 22925 18105 22937 18108
rect 22971 18136 22983 18139
rect 23400 18136 23428 18176
rect 24118 18164 24124 18176
rect 24176 18204 24182 18216
rect 24688 18204 24716 18258
rect 24176 18176 24716 18204
rect 25317 18207 25375 18213
rect 24176 18164 24182 18176
rect 25317 18173 25329 18207
rect 25363 18173 25375 18207
rect 25317 18167 25375 18173
rect 22971 18108 23428 18136
rect 22971 18105 22983 18108
rect 22925 18099 22983 18105
rect 17276 18040 18184 18068
rect 17276 18028 17282 18040
rect 18598 18028 18604 18080
rect 18656 18028 18662 18080
rect 18874 18028 18880 18080
rect 18932 18068 18938 18080
rect 19061 18071 19119 18077
rect 19061 18068 19073 18071
rect 18932 18040 19073 18068
rect 18932 18028 18938 18040
rect 19061 18037 19073 18040
rect 19107 18037 19119 18071
rect 19061 18031 19119 18037
rect 19429 18071 19487 18077
rect 19429 18037 19441 18071
rect 19475 18068 19487 18071
rect 19610 18068 19616 18080
rect 19475 18040 19616 18068
rect 19475 18037 19487 18040
rect 19429 18031 19487 18037
rect 19610 18028 19616 18040
rect 19668 18028 19674 18080
rect 20070 18028 20076 18080
rect 20128 18028 20134 18080
rect 20901 18071 20959 18077
rect 20901 18037 20913 18071
rect 20947 18068 20959 18071
rect 20990 18068 20996 18080
rect 20947 18040 20996 18068
rect 20947 18037 20959 18040
rect 20901 18031 20959 18037
rect 20990 18028 20996 18040
rect 21048 18028 21054 18080
rect 21358 18028 21364 18080
rect 21416 18028 21422 18080
rect 23382 18028 23388 18080
rect 23440 18068 23446 18080
rect 25332 18068 25360 18167
rect 23440 18040 25360 18068
rect 23440 18028 23446 18040
rect 1104 17978 25852 18000
rect 1104 17926 2950 17978
rect 3002 17926 3014 17978
rect 3066 17926 3078 17978
rect 3130 17926 3142 17978
rect 3194 17926 3206 17978
rect 3258 17926 12950 17978
rect 13002 17926 13014 17978
rect 13066 17926 13078 17978
rect 13130 17926 13142 17978
rect 13194 17926 13206 17978
rect 13258 17926 22950 17978
rect 23002 17926 23014 17978
rect 23066 17926 23078 17978
rect 23130 17926 23142 17978
rect 23194 17926 23206 17978
rect 23258 17926 25852 17978
rect 1104 17904 25852 17926
rect 8754 17824 8760 17876
rect 8812 17824 8818 17876
rect 9033 17867 9091 17873
rect 9033 17864 9045 17867
rect 8956 17836 9045 17864
rect 7653 17799 7711 17805
rect 7653 17765 7665 17799
rect 7699 17796 7711 17799
rect 7699 17768 8248 17796
rect 7699 17765 7711 17768
rect 7653 17759 7711 17765
rect 8220 17660 8248 17768
rect 8297 17731 8355 17737
rect 8297 17697 8309 17731
rect 8343 17728 8355 17731
rect 8956 17728 8984 17836
rect 9033 17833 9045 17836
rect 9079 17864 9091 17867
rect 10686 17864 10692 17876
rect 9079 17836 10692 17864
rect 9079 17833 9091 17836
rect 9033 17827 9091 17833
rect 10686 17824 10692 17836
rect 10744 17824 10750 17876
rect 10870 17824 10876 17876
rect 10928 17864 10934 17876
rect 10928 17836 11192 17864
rect 10928 17824 10934 17836
rect 11054 17796 11060 17808
rect 8343 17700 8984 17728
rect 9324 17768 11060 17796
rect 8343 17697 8355 17700
rect 8297 17691 8355 17697
rect 9324 17660 9352 17768
rect 11054 17756 11060 17768
rect 11112 17756 11118 17808
rect 11164 17796 11192 17836
rect 11238 17824 11244 17876
rect 11296 17864 11302 17876
rect 11793 17867 11851 17873
rect 11793 17864 11805 17867
rect 11296 17836 11805 17864
rect 11296 17824 11302 17836
rect 11793 17833 11805 17836
rect 11839 17833 11851 17867
rect 11793 17827 11851 17833
rect 13446 17824 13452 17876
rect 13504 17864 13510 17876
rect 17310 17864 17316 17876
rect 13504 17836 17316 17864
rect 13504 17824 13510 17836
rect 17310 17824 17316 17836
rect 17368 17824 17374 17876
rect 19426 17864 19432 17876
rect 17420 17836 19432 17864
rect 11330 17796 11336 17808
rect 11164 17768 11336 17796
rect 11330 17756 11336 17768
rect 11388 17796 11394 17808
rect 11609 17799 11667 17805
rect 11609 17796 11621 17799
rect 11388 17768 11621 17796
rect 11388 17756 11394 17768
rect 11609 17765 11621 17768
rect 11655 17796 11667 17799
rect 12158 17796 12164 17808
rect 11655 17768 12164 17796
rect 11655 17765 11667 17768
rect 11609 17759 11667 17765
rect 12158 17756 12164 17768
rect 12216 17756 12222 17808
rect 12434 17796 12440 17808
rect 12406 17756 12440 17796
rect 12492 17756 12498 17808
rect 9398 17688 9404 17740
rect 9456 17728 9462 17740
rect 10965 17731 11023 17737
rect 10965 17728 10977 17731
rect 9456 17700 10977 17728
rect 9456 17688 9462 17700
rect 10965 17697 10977 17700
rect 11011 17697 11023 17731
rect 12406 17728 12434 17756
rect 10965 17691 11023 17697
rect 11072 17700 12434 17728
rect 11072 17672 11100 17700
rect 8220 17632 9352 17660
rect 10229 17663 10287 17669
rect 10229 17629 10241 17663
rect 10275 17660 10287 17663
rect 10870 17660 10876 17672
rect 10275 17632 10876 17660
rect 10275 17629 10287 17632
rect 10229 17623 10287 17629
rect 10870 17620 10876 17632
rect 10928 17620 10934 17672
rect 11054 17620 11060 17672
rect 11112 17620 11118 17672
rect 12802 17620 12808 17672
rect 12860 17620 12866 17672
rect 8113 17595 8171 17601
rect 8113 17592 8125 17595
rect 7300 17564 8125 17592
rect 3786 17484 3792 17536
rect 3844 17524 3850 17536
rect 7300 17533 7328 17564
rect 8113 17561 8125 17564
rect 8159 17561 8171 17595
rect 8113 17555 8171 17561
rect 11238 17552 11244 17604
rect 11296 17592 11302 17604
rect 12066 17592 12072 17604
rect 11296 17564 12072 17592
rect 11296 17552 11302 17564
rect 12066 17552 12072 17564
rect 12124 17552 12130 17604
rect 12158 17552 12164 17604
rect 12216 17592 12222 17604
rect 13464 17592 13492 17824
rect 13814 17756 13820 17808
rect 13872 17796 13878 17808
rect 13909 17799 13967 17805
rect 13909 17796 13921 17799
rect 13872 17768 13921 17796
rect 13872 17756 13878 17768
rect 13909 17765 13921 17768
rect 13955 17796 13967 17799
rect 17420 17796 17448 17836
rect 19426 17824 19432 17836
rect 19484 17824 19490 17876
rect 21174 17824 21180 17876
rect 21232 17824 21238 17876
rect 21634 17824 21640 17876
rect 21692 17824 21698 17876
rect 21818 17824 21824 17876
rect 21876 17864 21882 17876
rect 26142 17864 26148 17876
rect 21876 17836 26148 17864
rect 21876 17824 21882 17836
rect 26142 17824 26148 17836
rect 26200 17824 26206 17876
rect 17862 17796 17868 17808
rect 13955 17768 17448 17796
rect 17788 17768 17868 17796
rect 13955 17765 13967 17768
rect 13909 17759 13967 17765
rect 14369 17731 14427 17737
rect 14369 17697 14381 17731
rect 14415 17728 14427 17731
rect 14642 17728 14648 17740
rect 14415 17700 14648 17728
rect 14415 17697 14427 17700
rect 14369 17691 14427 17697
rect 14642 17688 14648 17700
rect 14700 17688 14706 17740
rect 16666 17688 16672 17740
rect 16724 17728 16730 17740
rect 17788 17728 17816 17768
rect 17862 17756 17868 17768
rect 17920 17756 17926 17808
rect 17957 17799 18015 17805
rect 17957 17765 17969 17799
rect 18003 17796 18015 17799
rect 19150 17796 19156 17808
rect 18003 17768 19156 17796
rect 18003 17765 18015 17768
rect 17957 17759 18015 17765
rect 19150 17756 19156 17768
rect 19208 17756 19214 17808
rect 16724 17700 17816 17728
rect 18417 17731 18475 17737
rect 16724 17688 16730 17700
rect 18417 17697 18429 17731
rect 18463 17728 18475 17731
rect 18506 17728 18512 17740
rect 18463 17700 18512 17728
rect 18463 17697 18475 17700
rect 18417 17691 18475 17697
rect 18506 17688 18512 17700
rect 18564 17688 18570 17740
rect 18598 17688 18604 17740
rect 18656 17688 18662 17740
rect 18782 17688 18788 17740
rect 18840 17728 18846 17740
rect 18969 17731 19027 17737
rect 18969 17728 18981 17731
rect 18840 17700 18981 17728
rect 18840 17688 18846 17700
rect 18969 17697 18981 17700
rect 19015 17697 19027 17731
rect 18969 17691 19027 17697
rect 23845 17731 23903 17737
rect 23845 17697 23857 17731
rect 23891 17728 23903 17731
rect 24854 17728 24860 17740
rect 23891 17700 24860 17728
rect 23891 17697 23903 17700
rect 23845 17691 23903 17697
rect 24854 17688 24860 17700
rect 24912 17688 24918 17740
rect 24946 17688 24952 17740
rect 25004 17728 25010 17740
rect 25041 17731 25099 17737
rect 25041 17728 25053 17731
rect 25004 17700 25053 17728
rect 25004 17688 25010 17700
rect 25041 17697 25053 17700
rect 25087 17697 25099 17731
rect 25041 17691 25099 17697
rect 25130 17688 25136 17740
rect 25188 17688 25194 17740
rect 16758 17620 16764 17672
rect 16816 17660 16822 17672
rect 16853 17663 16911 17669
rect 16853 17660 16865 17663
rect 16816 17632 16865 17660
rect 16816 17620 16822 17632
rect 16853 17629 16865 17632
rect 16899 17629 16911 17663
rect 16853 17623 16911 17629
rect 18322 17620 18328 17672
rect 18380 17660 18386 17672
rect 19429 17663 19487 17669
rect 19429 17660 19441 17663
rect 18380 17632 19441 17660
rect 18380 17620 18386 17632
rect 19429 17629 19441 17632
rect 19475 17629 19487 17663
rect 19429 17623 19487 17629
rect 21910 17620 21916 17672
rect 21968 17660 21974 17672
rect 22005 17663 22063 17669
rect 22005 17660 22017 17663
rect 21968 17632 22017 17660
rect 21968 17620 21974 17632
rect 22005 17629 22017 17632
rect 22051 17629 22063 17663
rect 22005 17623 22063 17629
rect 22646 17620 22652 17672
rect 22704 17620 22710 17672
rect 12216 17564 13492 17592
rect 12216 17552 12222 17564
rect 13998 17552 14004 17604
rect 14056 17592 14062 17604
rect 15194 17592 15200 17604
rect 14056 17564 15200 17592
rect 14056 17552 14062 17564
rect 15194 17552 15200 17564
rect 15252 17552 15258 17604
rect 15562 17552 15568 17604
rect 15620 17592 15626 17604
rect 17313 17595 17371 17601
rect 15620 17564 16896 17592
rect 15620 17552 15626 17564
rect 7285 17527 7343 17533
rect 7285 17524 7297 17527
rect 3844 17496 7297 17524
rect 3844 17484 3850 17496
rect 7285 17493 7297 17496
rect 7331 17493 7343 17527
rect 7285 17487 7343 17493
rect 7834 17484 7840 17536
rect 7892 17524 7898 17536
rect 8021 17527 8079 17533
rect 8021 17524 8033 17527
rect 7892 17496 8033 17524
rect 7892 17484 7898 17496
rect 8021 17493 8033 17496
rect 8067 17493 8079 17527
rect 8021 17487 8079 17493
rect 9766 17484 9772 17536
rect 9824 17524 9830 17536
rect 11256 17524 11284 17552
rect 9824 17496 11284 17524
rect 9824 17484 9830 17496
rect 11514 17484 11520 17536
rect 11572 17484 11578 17536
rect 13446 17484 13452 17536
rect 13504 17484 13510 17536
rect 13906 17484 13912 17536
rect 13964 17524 13970 17536
rect 15013 17527 15071 17533
rect 15013 17524 15025 17527
rect 13964 17496 15025 17524
rect 13964 17484 13970 17496
rect 15013 17493 15025 17496
rect 15059 17493 15071 17527
rect 15013 17487 15071 17493
rect 15654 17484 15660 17536
rect 15712 17484 15718 17536
rect 16669 17527 16727 17533
rect 16669 17493 16681 17527
rect 16715 17524 16727 17527
rect 16758 17524 16764 17536
rect 16715 17496 16764 17524
rect 16715 17493 16727 17496
rect 16669 17487 16727 17493
rect 16758 17484 16764 17496
rect 16816 17484 16822 17536
rect 16868 17524 16896 17564
rect 17313 17561 17325 17595
rect 17359 17592 17371 17595
rect 19242 17592 19248 17604
rect 17359 17564 19248 17592
rect 17359 17561 17371 17564
rect 17313 17555 17371 17561
rect 19242 17552 19248 17564
rect 19300 17552 19306 17604
rect 19334 17552 19340 17604
rect 19392 17592 19398 17604
rect 19705 17595 19763 17601
rect 19705 17592 19717 17595
rect 19392 17564 19717 17592
rect 19392 17552 19398 17564
rect 19705 17561 19717 17564
rect 19751 17561 19763 17595
rect 20990 17592 20996 17604
rect 20930 17564 20996 17592
rect 19705 17555 19763 17561
rect 20990 17552 20996 17564
rect 21048 17592 21054 17604
rect 21358 17592 21364 17604
rect 21048 17564 21364 17592
rect 21048 17552 21054 17564
rect 21358 17552 21364 17564
rect 21416 17552 21422 17604
rect 18325 17527 18383 17533
rect 18325 17524 18337 17527
rect 16868 17496 18337 17524
rect 18325 17493 18337 17496
rect 18371 17493 18383 17527
rect 18325 17487 18383 17493
rect 18782 17484 18788 17536
rect 18840 17524 18846 17536
rect 21008 17524 21036 17552
rect 18840 17496 21036 17524
rect 18840 17484 18846 17496
rect 22094 17484 22100 17536
rect 22152 17484 22158 17536
rect 24578 17484 24584 17536
rect 24636 17484 24642 17536
rect 24946 17484 24952 17536
rect 25004 17484 25010 17536
rect 1104 17434 25852 17456
rect 1104 17382 7950 17434
rect 8002 17382 8014 17434
rect 8066 17382 8078 17434
rect 8130 17382 8142 17434
rect 8194 17382 8206 17434
rect 8258 17382 17950 17434
rect 18002 17382 18014 17434
rect 18066 17382 18078 17434
rect 18130 17382 18142 17434
rect 18194 17382 18206 17434
rect 18258 17382 25852 17434
rect 1104 17360 25852 17382
rect 7834 17280 7840 17332
rect 7892 17320 7898 17332
rect 8021 17323 8079 17329
rect 8021 17320 8033 17323
rect 7892 17292 8033 17320
rect 7892 17280 7898 17292
rect 8021 17289 8033 17292
rect 8067 17289 8079 17323
rect 8021 17283 8079 17289
rect 9490 17280 9496 17332
rect 9548 17280 9554 17332
rect 10321 17323 10379 17329
rect 10321 17289 10333 17323
rect 10367 17289 10379 17323
rect 10321 17283 10379 17289
rect 8570 17212 8576 17264
rect 8628 17252 8634 17264
rect 10336 17252 10364 17283
rect 11606 17280 11612 17332
rect 11664 17320 11670 17332
rect 11701 17323 11759 17329
rect 11701 17320 11713 17323
rect 11664 17292 11713 17320
rect 11664 17280 11670 17292
rect 11701 17289 11713 17292
rect 11747 17289 11759 17323
rect 11701 17283 11759 17289
rect 12897 17323 12955 17329
rect 12897 17289 12909 17323
rect 12943 17289 12955 17323
rect 12897 17283 12955 17289
rect 13265 17323 13323 17329
rect 13265 17289 13277 17323
rect 13311 17320 13323 17323
rect 13906 17320 13912 17332
rect 13311 17292 13912 17320
rect 13311 17289 13323 17292
rect 13265 17283 13323 17289
rect 8628 17224 10364 17252
rect 10781 17255 10839 17261
rect 8628 17212 8634 17224
rect 10781 17221 10793 17255
rect 10827 17252 10839 17255
rect 12250 17252 12256 17264
rect 10827 17224 12256 17252
rect 10827 17221 10839 17224
rect 10781 17215 10839 17221
rect 12250 17212 12256 17224
rect 12308 17212 12314 17264
rect 12912 17252 12940 17283
rect 13906 17280 13912 17292
rect 13964 17280 13970 17332
rect 15102 17320 15108 17332
rect 14384 17292 15108 17320
rect 13538 17252 13544 17264
rect 12912 17224 13544 17252
rect 13538 17212 13544 17224
rect 13596 17212 13602 17264
rect 6917 17187 6975 17193
rect 6917 17153 6929 17187
rect 6963 17184 6975 17187
rect 7650 17184 7656 17196
rect 6963 17156 7656 17184
rect 6963 17153 6975 17156
rect 6917 17147 6975 17153
rect 7650 17144 7656 17156
rect 7708 17144 7714 17196
rect 9214 17144 9220 17196
rect 9272 17184 9278 17196
rect 10689 17187 10747 17193
rect 9272 17156 9720 17184
rect 9272 17144 9278 17156
rect 9692 17125 9720 17156
rect 10689 17153 10701 17187
rect 10735 17184 10747 17187
rect 11698 17184 11704 17196
rect 10735 17156 11704 17184
rect 10735 17153 10747 17156
rect 10689 17147 10747 17153
rect 11698 17144 11704 17156
rect 11756 17144 11762 17196
rect 12066 17144 12072 17196
rect 12124 17144 12130 17196
rect 14384 17184 14412 17292
rect 15102 17280 15108 17292
rect 15160 17280 15166 17332
rect 19242 17280 19248 17332
rect 19300 17320 19306 17332
rect 21085 17323 21143 17329
rect 21085 17320 21097 17323
rect 19300 17292 21097 17320
rect 19300 17280 19306 17292
rect 21085 17289 21097 17292
rect 21131 17289 21143 17323
rect 21085 17283 21143 17289
rect 21174 17280 21180 17332
rect 21232 17280 21238 17332
rect 15194 17212 15200 17264
rect 15252 17212 15258 17264
rect 17037 17255 17095 17261
rect 17037 17221 17049 17255
rect 17083 17252 17095 17255
rect 17310 17252 17316 17264
rect 17083 17224 17316 17252
rect 17083 17221 17095 17224
rect 17037 17215 17095 17221
rect 17310 17212 17316 17224
rect 17368 17212 17374 17264
rect 19518 17212 19524 17264
rect 19576 17252 19582 17264
rect 19889 17255 19947 17261
rect 19889 17252 19901 17255
rect 19576 17224 19901 17252
rect 19576 17212 19582 17224
rect 19889 17221 19901 17224
rect 19935 17221 19947 17255
rect 19889 17215 19947 17221
rect 20806 17212 20812 17264
rect 20864 17252 20870 17264
rect 23293 17255 23351 17261
rect 20864 17224 23060 17252
rect 20864 17212 20870 17224
rect 14461 17187 14519 17193
rect 14461 17184 14473 17187
rect 14384 17156 14473 17184
rect 14461 17153 14473 17156
rect 14507 17153 14519 17187
rect 14461 17147 14519 17153
rect 16850 17144 16856 17196
rect 16908 17184 16914 17196
rect 18049 17187 18107 17193
rect 18049 17184 18061 17187
rect 16908 17156 18061 17184
rect 16908 17144 16914 17156
rect 18049 17153 18061 17156
rect 18095 17184 18107 17187
rect 18322 17184 18328 17196
rect 18095 17156 18328 17184
rect 18095 17153 18107 17156
rect 18049 17147 18107 17153
rect 18322 17144 18328 17156
rect 18380 17144 18386 17196
rect 18598 17144 18604 17196
rect 18656 17184 18662 17196
rect 18693 17187 18751 17193
rect 18693 17184 18705 17187
rect 18656 17156 18705 17184
rect 18656 17144 18662 17156
rect 18693 17153 18705 17156
rect 18739 17153 18751 17187
rect 18693 17147 18751 17153
rect 19242 17144 19248 17196
rect 19300 17184 19306 17196
rect 20349 17187 20407 17193
rect 20349 17184 20361 17187
rect 19300 17156 20361 17184
rect 19300 17144 19306 17156
rect 20349 17153 20361 17156
rect 20395 17184 20407 17187
rect 20395 17156 21312 17184
rect 20395 17153 20407 17156
rect 20349 17147 20407 17153
rect 9585 17119 9643 17125
rect 9585 17116 9597 17119
rect 8864 17088 9597 17116
rect 8864 16992 8892 17088
rect 9585 17085 9597 17088
rect 9631 17085 9643 17119
rect 9585 17079 9643 17085
rect 9677 17119 9735 17125
rect 9677 17085 9689 17119
rect 9723 17085 9735 17119
rect 9677 17079 9735 17085
rect 10873 17119 10931 17125
rect 10873 17085 10885 17119
rect 10919 17085 10931 17119
rect 10873 17079 10931 17085
rect 9306 17008 9312 17060
rect 9364 17048 9370 17060
rect 10888 17048 10916 17079
rect 12158 17076 12164 17128
rect 12216 17076 12222 17128
rect 12253 17119 12311 17125
rect 12253 17085 12265 17119
rect 12299 17085 12311 17119
rect 12253 17079 12311 17085
rect 9364 17020 10916 17048
rect 9364 17008 9370 17020
rect 11146 17008 11152 17060
rect 11204 17048 11210 17060
rect 12268 17048 12296 17079
rect 13354 17076 13360 17128
rect 13412 17076 13418 17128
rect 13541 17119 13599 17125
rect 13541 17085 13553 17119
rect 13587 17116 13599 17119
rect 13722 17116 13728 17128
rect 13587 17088 13728 17116
rect 13587 17085 13599 17088
rect 13541 17079 13599 17085
rect 13722 17076 13728 17088
rect 13780 17076 13786 17128
rect 14737 17119 14795 17125
rect 14737 17085 14749 17119
rect 14783 17116 14795 17119
rect 15470 17116 15476 17128
rect 14783 17088 15476 17116
rect 14783 17085 14795 17088
rect 14737 17079 14795 17085
rect 15470 17076 15476 17088
rect 15528 17076 15534 17128
rect 16298 17076 16304 17128
rect 16356 17116 16362 17128
rect 21284 17125 21312 17156
rect 22186 17144 22192 17196
rect 22244 17144 22250 17196
rect 23032 17184 23060 17224
rect 23293 17221 23305 17255
rect 23339 17252 23351 17255
rect 24854 17252 24860 17264
rect 23339 17224 24860 17252
rect 23339 17221 23351 17224
rect 23293 17215 23351 17221
rect 24854 17212 24860 17224
rect 24912 17212 24918 17264
rect 23937 17187 23995 17193
rect 23937 17184 23949 17187
rect 23032 17156 23949 17184
rect 23937 17153 23949 17156
rect 23983 17153 23995 17187
rect 23937 17147 23995 17153
rect 21269 17119 21327 17125
rect 16356 17088 19472 17116
rect 16356 17076 16362 17088
rect 12342 17048 12348 17060
rect 11204 17020 12348 17048
rect 11204 17008 11210 17020
rect 12342 17008 12348 17020
rect 12400 17008 12406 17060
rect 13372 17048 13400 17076
rect 13909 17051 13967 17057
rect 13909 17048 13921 17051
rect 13372 17020 13921 17048
rect 13909 17017 13921 17020
rect 13955 17017 13967 17051
rect 13909 17011 13967 17017
rect 16206 17008 16212 17060
rect 16264 17008 16270 17060
rect 16574 17008 16580 17060
rect 16632 17048 16638 17060
rect 19337 17051 19395 17057
rect 19337 17048 19349 17051
rect 16632 17020 19349 17048
rect 16632 17008 16638 17020
rect 19337 17017 19349 17020
rect 19383 17017 19395 17051
rect 19444 17048 19472 17088
rect 21269 17085 21281 17119
rect 21315 17116 21327 17119
rect 23382 17116 23388 17128
rect 21315 17088 23388 17116
rect 21315 17085 21327 17088
rect 21269 17079 21327 17085
rect 23382 17076 23388 17088
rect 23440 17076 23446 17128
rect 24762 17076 24768 17128
rect 24820 17076 24826 17128
rect 24578 17048 24584 17060
rect 19444 17020 24584 17048
rect 19337 17011 19395 17017
rect 24578 17008 24584 17020
rect 24636 17008 24642 17060
rect 7561 16983 7619 16989
rect 7561 16949 7573 16983
rect 7607 16980 7619 16983
rect 7834 16980 7840 16992
rect 7607 16952 7840 16980
rect 7607 16949 7619 16952
rect 7561 16943 7619 16949
rect 7834 16940 7840 16952
rect 7892 16940 7898 16992
rect 8846 16940 8852 16992
rect 8904 16940 8910 16992
rect 9125 16983 9183 16989
rect 9125 16949 9137 16983
rect 9171 16980 9183 16983
rect 11974 16980 11980 16992
rect 9171 16952 11980 16980
rect 9171 16949 9183 16952
rect 9125 16943 9183 16949
rect 11974 16940 11980 16952
rect 12032 16940 12038 16992
rect 15194 16940 15200 16992
rect 15252 16980 15258 16992
rect 16666 16980 16672 16992
rect 15252 16952 16672 16980
rect 15252 16940 15258 16952
rect 16666 16940 16672 16952
rect 16724 16940 16730 16992
rect 16850 16940 16856 16992
rect 16908 16980 16914 16992
rect 19981 16983 20039 16989
rect 19981 16980 19993 16983
rect 16908 16952 19993 16980
rect 16908 16940 16914 16952
rect 19981 16949 19993 16952
rect 20027 16949 20039 16983
rect 19981 16943 20039 16949
rect 20717 16983 20775 16989
rect 20717 16949 20729 16983
rect 20763 16980 20775 16983
rect 22370 16980 22376 16992
rect 20763 16952 22376 16980
rect 20763 16949 20775 16952
rect 20717 16943 20775 16949
rect 22370 16940 22376 16952
rect 22428 16940 22434 16992
rect 1104 16890 25852 16912
rect 1104 16838 2950 16890
rect 3002 16838 3014 16890
rect 3066 16838 3078 16890
rect 3130 16838 3142 16890
rect 3194 16838 3206 16890
rect 3258 16838 12950 16890
rect 13002 16838 13014 16890
rect 13066 16838 13078 16890
rect 13130 16838 13142 16890
rect 13194 16838 13206 16890
rect 13258 16838 22950 16890
rect 23002 16838 23014 16890
rect 23066 16838 23078 16890
rect 23130 16838 23142 16890
rect 23194 16838 23206 16890
rect 23258 16838 25852 16890
rect 1104 16816 25852 16838
rect 7650 16736 7656 16788
rect 7708 16736 7714 16788
rect 8021 16779 8079 16785
rect 8021 16745 8033 16779
rect 8067 16776 8079 16779
rect 8754 16776 8760 16788
rect 8067 16748 8760 16776
rect 8067 16745 8079 16748
rect 8021 16739 8079 16745
rect 8036 16708 8064 16739
rect 8754 16736 8760 16748
rect 8812 16776 8818 16788
rect 9582 16776 9588 16788
rect 8812 16748 9588 16776
rect 8812 16736 8818 16748
rect 9582 16736 9588 16748
rect 9640 16736 9646 16788
rect 11146 16736 11152 16788
rect 11204 16776 11210 16788
rect 11425 16779 11483 16785
rect 11425 16776 11437 16779
rect 11204 16748 11437 16776
rect 11204 16736 11210 16748
rect 11425 16745 11437 16748
rect 11471 16745 11483 16779
rect 11425 16739 11483 16745
rect 12434 16736 12440 16788
rect 12492 16776 12498 16788
rect 13998 16776 14004 16788
rect 12492 16748 14004 16776
rect 12492 16736 12498 16748
rect 13998 16736 14004 16748
rect 14056 16736 14062 16788
rect 16666 16736 16672 16788
rect 16724 16776 16730 16788
rect 17037 16779 17095 16785
rect 17037 16776 17049 16779
rect 16724 16748 17049 16776
rect 16724 16736 16730 16748
rect 17037 16745 17049 16748
rect 17083 16745 17095 16779
rect 17037 16739 17095 16745
rect 17310 16736 17316 16788
rect 17368 16776 17374 16788
rect 18322 16776 18328 16788
rect 17368 16748 18328 16776
rect 17368 16736 17374 16748
rect 18322 16736 18328 16748
rect 18380 16776 18386 16788
rect 18969 16779 19027 16785
rect 18969 16776 18981 16779
rect 18380 16748 18981 16776
rect 18380 16736 18386 16748
rect 18969 16745 18981 16748
rect 19015 16745 19027 16779
rect 18969 16739 19027 16745
rect 12989 16711 13047 16717
rect 12989 16708 13001 16711
rect 7300 16680 8064 16708
rect 10704 16680 13001 16708
rect 5905 16643 5963 16649
rect 5905 16609 5917 16643
rect 5951 16640 5963 16643
rect 6822 16640 6828 16652
rect 5951 16612 6828 16640
rect 5951 16609 5963 16612
rect 5905 16603 5963 16609
rect 6822 16600 6828 16612
rect 6880 16600 6886 16652
rect 7300 16558 7328 16680
rect 7466 16600 7472 16652
rect 7524 16640 7530 16652
rect 9674 16640 9680 16652
rect 7524 16612 9680 16640
rect 7524 16600 7530 16612
rect 9674 16600 9680 16612
rect 9732 16600 9738 16652
rect 10704 16649 10732 16680
rect 12989 16677 13001 16680
rect 13035 16677 13047 16711
rect 14277 16711 14335 16717
rect 14277 16708 14289 16711
rect 12989 16671 13047 16677
rect 13464 16680 14289 16708
rect 10689 16643 10747 16649
rect 10689 16609 10701 16643
rect 10735 16609 10747 16643
rect 10689 16603 10747 16609
rect 10873 16643 10931 16649
rect 10873 16609 10885 16643
rect 10919 16640 10931 16643
rect 11238 16640 11244 16652
rect 10919 16612 11244 16640
rect 10919 16609 10931 16612
rect 10873 16603 10931 16609
rect 11238 16600 11244 16612
rect 11296 16600 11302 16652
rect 12342 16600 12348 16652
rect 12400 16600 12406 16652
rect 13354 16640 13360 16652
rect 12452 16612 13360 16640
rect 10594 16532 10600 16584
rect 10652 16532 10658 16584
rect 11054 16532 11060 16584
rect 11112 16572 11118 16584
rect 12452 16572 12480 16612
rect 13354 16600 13360 16612
rect 13412 16640 13418 16652
rect 13464 16649 13492 16680
rect 14277 16677 14289 16680
rect 14323 16677 14335 16711
rect 14277 16671 14335 16677
rect 18141 16711 18199 16717
rect 18141 16677 18153 16711
rect 18187 16708 18199 16711
rect 18414 16708 18420 16720
rect 18187 16680 18420 16708
rect 18187 16677 18199 16680
rect 18141 16671 18199 16677
rect 13449 16643 13507 16649
rect 13449 16640 13461 16643
rect 13412 16612 13461 16640
rect 13412 16600 13418 16612
rect 13449 16609 13461 16612
rect 13495 16609 13507 16643
rect 13449 16603 13507 16609
rect 13538 16600 13544 16652
rect 13596 16600 13602 16652
rect 14090 16600 14096 16652
rect 14148 16600 14154 16652
rect 15013 16643 15071 16649
rect 15013 16609 15025 16643
rect 15059 16640 15071 16643
rect 15746 16640 15752 16652
rect 15059 16612 15752 16640
rect 15059 16609 15071 16612
rect 15013 16603 15071 16609
rect 15746 16600 15752 16612
rect 15804 16600 15810 16652
rect 15933 16643 15991 16649
rect 15933 16609 15945 16643
rect 15979 16640 15991 16643
rect 16482 16640 16488 16652
rect 15979 16612 16488 16640
rect 15979 16609 15991 16612
rect 15933 16603 15991 16609
rect 16482 16600 16488 16612
rect 16540 16600 16546 16652
rect 11112 16544 12480 16572
rect 11112 16532 11118 16544
rect 15654 16532 15660 16584
rect 15712 16532 15718 16584
rect 17678 16532 17684 16584
rect 17736 16572 17742 16584
rect 17773 16575 17831 16581
rect 17773 16572 17785 16575
rect 17736 16544 17785 16572
rect 17736 16532 17742 16544
rect 17773 16541 17785 16544
rect 17819 16541 17831 16575
rect 17773 16535 17831 16541
rect 6178 16464 6184 16516
rect 6236 16464 6242 16516
rect 9953 16507 10011 16513
rect 9953 16473 9965 16507
rect 9999 16504 10011 16507
rect 10612 16504 10640 16532
rect 12161 16507 12219 16513
rect 9999 16476 10548 16504
rect 10612 16476 11836 16504
rect 9999 16473 10011 16476
rect 9953 16467 10011 16473
rect 10229 16439 10287 16445
rect 10229 16405 10241 16439
rect 10275 16436 10287 16439
rect 10410 16436 10416 16448
rect 10275 16408 10416 16436
rect 10275 16405 10287 16408
rect 10229 16399 10287 16405
rect 10410 16396 10416 16408
rect 10468 16396 10474 16448
rect 10520 16436 10548 16476
rect 10597 16439 10655 16445
rect 10597 16436 10609 16439
rect 10520 16408 10609 16436
rect 10597 16405 10609 16408
rect 10643 16436 10655 16439
rect 10686 16436 10692 16448
rect 10643 16408 10692 16436
rect 10643 16405 10655 16408
rect 10597 16399 10655 16405
rect 10686 16396 10692 16408
rect 10744 16436 10750 16448
rect 10962 16436 10968 16448
rect 10744 16408 10968 16436
rect 10744 16396 10750 16408
rect 10962 16396 10968 16408
rect 11020 16396 11026 16448
rect 11808 16445 11836 16476
rect 12161 16473 12173 16507
rect 12207 16504 12219 16507
rect 13630 16504 13636 16516
rect 12207 16476 13636 16504
rect 12207 16473 12219 16476
rect 12161 16467 12219 16473
rect 13630 16464 13636 16476
rect 13688 16464 13694 16516
rect 16945 16507 17003 16513
rect 16945 16473 16957 16507
rect 16991 16504 17003 16507
rect 18156 16504 18184 16671
rect 18414 16668 18420 16680
rect 18472 16668 18478 16720
rect 18598 16532 18604 16584
rect 18656 16532 18662 16584
rect 18984 16572 19012 16739
rect 19426 16736 19432 16788
rect 19484 16776 19490 16788
rect 25774 16776 25780 16788
rect 19484 16748 25780 16776
rect 19484 16736 19490 16748
rect 25774 16736 25780 16748
rect 25832 16736 25838 16788
rect 19429 16575 19487 16581
rect 19429 16572 19441 16575
rect 18984 16544 19441 16572
rect 19429 16541 19441 16544
rect 19475 16541 19487 16575
rect 20714 16572 20720 16584
rect 19429 16535 19487 16541
rect 19628 16544 20720 16572
rect 19628 16504 19656 16544
rect 20714 16532 20720 16544
rect 20772 16532 20778 16584
rect 20809 16575 20867 16581
rect 20809 16541 20821 16575
rect 20855 16572 20867 16575
rect 20990 16572 20996 16584
rect 20855 16544 20996 16572
rect 20855 16541 20867 16544
rect 20809 16535 20867 16541
rect 20990 16532 20996 16544
rect 21048 16532 21054 16584
rect 21913 16575 21971 16581
rect 21913 16541 21925 16575
rect 21959 16572 21971 16575
rect 22554 16572 22560 16584
rect 21959 16544 22560 16572
rect 21959 16541 21971 16544
rect 21913 16535 21971 16541
rect 22554 16532 22560 16544
rect 22612 16532 22618 16584
rect 22738 16532 22744 16584
rect 22796 16532 22802 16584
rect 23934 16532 23940 16584
rect 23992 16572 23998 16584
rect 24581 16575 24639 16581
rect 24581 16572 24593 16575
rect 23992 16544 24593 16572
rect 23992 16532 23998 16544
rect 24581 16541 24593 16544
rect 24627 16541 24639 16575
rect 24581 16535 24639 16541
rect 25222 16532 25228 16584
rect 25280 16532 25286 16584
rect 16991 16476 18184 16504
rect 18432 16476 19656 16504
rect 16991 16473 17003 16476
rect 16945 16467 17003 16473
rect 11793 16439 11851 16445
rect 11793 16405 11805 16439
rect 11839 16405 11851 16439
rect 11793 16399 11851 16405
rect 12253 16439 12311 16445
rect 12253 16405 12265 16439
rect 12299 16436 12311 16439
rect 12434 16436 12440 16448
rect 12299 16408 12440 16436
rect 12299 16405 12311 16408
rect 12253 16399 12311 16405
rect 12434 16396 12440 16408
rect 12492 16396 12498 16448
rect 13357 16439 13415 16445
rect 13357 16405 13369 16439
rect 13403 16436 13415 16439
rect 14090 16436 14096 16448
rect 13403 16408 14096 16436
rect 13403 16405 13415 16408
rect 13357 16399 13415 16405
rect 14090 16396 14096 16408
rect 14148 16396 14154 16448
rect 15289 16439 15347 16445
rect 15289 16405 15301 16439
rect 15335 16436 15347 16439
rect 16390 16436 16396 16448
rect 15335 16408 16396 16436
rect 15335 16405 15347 16408
rect 15289 16399 15347 16405
rect 16390 16396 16396 16408
rect 16448 16396 16454 16448
rect 17402 16396 17408 16448
rect 17460 16436 17466 16448
rect 18432 16445 18460 16476
rect 19702 16464 19708 16516
rect 19760 16504 19766 16516
rect 20165 16507 20223 16513
rect 20165 16504 20177 16507
rect 19760 16476 20177 16504
rect 19760 16464 19766 16476
rect 20165 16473 20177 16476
rect 20211 16504 20223 16507
rect 20622 16504 20628 16516
rect 20211 16476 20628 16504
rect 20211 16473 20223 16476
rect 20165 16467 20223 16473
rect 20622 16464 20628 16476
rect 20680 16464 20686 16516
rect 23845 16507 23903 16513
rect 23845 16473 23857 16507
rect 23891 16504 23903 16507
rect 24946 16504 24952 16516
rect 23891 16476 24952 16504
rect 23891 16473 23903 16476
rect 23845 16467 23903 16473
rect 24946 16464 24952 16476
rect 25004 16464 25010 16516
rect 17589 16439 17647 16445
rect 17589 16436 17601 16439
rect 17460 16408 17601 16436
rect 17460 16396 17466 16408
rect 17589 16405 17601 16408
rect 17635 16405 17647 16439
rect 17589 16399 17647 16405
rect 18417 16439 18475 16445
rect 18417 16405 18429 16439
rect 18463 16405 18475 16439
rect 18417 16399 18475 16405
rect 18874 16396 18880 16448
rect 18932 16436 18938 16448
rect 19242 16436 19248 16448
rect 18932 16408 19248 16436
rect 18932 16396 18938 16408
rect 19242 16396 19248 16408
rect 19300 16396 19306 16448
rect 19978 16396 19984 16448
rect 20036 16436 20042 16448
rect 21453 16439 21511 16445
rect 21453 16436 21465 16439
rect 20036 16408 21465 16436
rect 20036 16396 20042 16408
rect 21453 16405 21465 16408
rect 21499 16405 21511 16439
rect 21453 16399 21511 16405
rect 21542 16396 21548 16448
rect 21600 16436 21606 16448
rect 24854 16436 24860 16448
rect 21600 16408 24860 16436
rect 21600 16396 21606 16408
rect 24854 16396 24860 16408
rect 24912 16396 24918 16448
rect 1104 16346 25852 16368
rect 1104 16294 7950 16346
rect 8002 16294 8014 16346
rect 8066 16294 8078 16346
rect 8130 16294 8142 16346
rect 8194 16294 8206 16346
rect 8258 16294 17950 16346
rect 18002 16294 18014 16346
rect 18066 16294 18078 16346
rect 18130 16294 18142 16346
rect 18194 16294 18206 16346
rect 18258 16294 25852 16346
rect 1104 16272 25852 16294
rect 5442 16192 5448 16244
rect 5500 16232 5506 16244
rect 11054 16232 11060 16244
rect 5500 16204 11060 16232
rect 5500 16192 5506 16204
rect 11054 16192 11060 16204
rect 11112 16192 11118 16244
rect 11606 16192 11612 16244
rect 11664 16232 11670 16244
rect 12618 16232 12624 16244
rect 11664 16204 12624 16232
rect 11664 16192 11670 16204
rect 12618 16192 12624 16204
rect 12676 16192 12682 16244
rect 14093 16235 14151 16241
rect 14093 16201 14105 16235
rect 14139 16201 14151 16235
rect 14093 16195 14151 16201
rect 7834 16124 7840 16176
rect 7892 16124 7898 16176
rect 9582 16164 9588 16176
rect 9062 16136 9588 16164
rect 9582 16124 9588 16136
rect 9640 16164 9646 16176
rect 9861 16167 9919 16173
rect 9861 16164 9873 16167
rect 9640 16136 9873 16164
rect 9640 16124 9646 16136
rect 9861 16133 9873 16136
rect 9907 16164 9919 16167
rect 11514 16164 11520 16176
rect 9907 16136 11520 16164
rect 9907 16133 9919 16136
rect 9861 16127 9919 16133
rect 11514 16124 11520 16136
rect 11572 16164 11578 16176
rect 12434 16164 12440 16176
rect 11572 16136 12440 16164
rect 11572 16124 11578 16136
rect 12434 16124 12440 16136
rect 12492 16124 12498 16176
rect 14108 16164 14136 16195
rect 15470 16192 15476 16244
rect 15528 16232 15534 16244
rect 16301 16235 16359 16241
rect 16301 16232 16313 16235
rect 15528 16204 16313 16232
rect 15528 16192 15534 16204
rect 16301 16201 16313 16204
rect 16347 16201 16359 16235
rect 18598 16232 18604 16244
rect 16301 16195 16359 16201
rect 16408 16204 18604 16232
rect 16408 16164 16436 16204
rect 18598 16192 18604 16204
rect 18656 16192 18662 16244
rect 19245 16235 19303 16241
rect 19245 16201 19257 16235
rect 19291 16232 19303 16235
rect 19334 16232 19340 16244
rect 19291 16204 19340 16232
rect 19291 16201 19303 16204
rect 19245 16195 19303 16201
rect 19334 16192 19340 16204
rect 19392 16192 19398 16244
rect 21542 16232 21548 16244
rect 19904 16204 21548 16232
rect 14108 16136 16436 16164
rect 16853 16167 16911 16173
rect 16853 16133 16865 16167
rect 16899 16164 16911 16167
rect 17218 16164 17224 16176
rect 16899 16136 17224 16164
rect 16899 16133 16911 16136
rect 16853 16127 16911 16133
rect 17218 16124 17224 16136
rect 17276 16124 17282 16176
rect 17957 16167 18015 16173
rect 17957 16133 17969 16167
rect 18003 16164 18015 16167
rect 19904 16164 19932 16204
rect 21542 16192 21548 16204
rect 21600 16192 21606 16244
rect 21634 16192 21640 16244
rect 21692 16232 21698 16244
rect 21692 16204 24348 16232
rect 21692 16192 21698 16204
rect 18003 16136 19932 16164
rect 18003 16133 18015 16136
rect 17957 16127 18015 16133
rect 19978 16124 19984 16176
rect 20036 16124 20042 16176
rect 21358 16164 21364 16176
rect 21206 16136 21364 16164
rect 21358 16124 21364 16136
rect 21416 16164 21422 16176
rect 21910 16164 21916 16176
rect 21416 16136 21916 16164
rect 21416 16124 21422 16136
rect 21910 16124 21916 16136
rect 21968 16124 21974 16176
rect 24320 16164 24348 16204
rect 25038 16192 25044 16244
rect 25096 16232 25102 16244
rect 25133 16235 25191 16241
rect 25133 16232 25145 16235
rect 25096 16204 25145 16232
rect 25096 16192 25102 16204
rect 25133 16201 25145 16204
rect 25179 16201 25191 16235
rect 25133 16195 25191 16201
rect 25409 16167 25467 16173
rect 25409 16164 25421 16167
rect 24320 16136 25421 16164
rect 25409 16133 25421 16136
rect 25455 16164 25467 16167
rect 25866 16164 25872 16176
rect 25455 16136 25872 16164
rect 25455 16133 25467 16136
rect 25409 16127 25467 16133
rect 25866 16124 25872 16136
rect 25924 16124 25930 16176
rect 6914 16056 6920 16108
rect 6972 16096 6978 16108
rect 7561 16099 7619 16105
rect 7561 16096 7573 16099
rect 6972 16068 7573 16096
rect 6972 16056 6978 16068
rect 7561 16065 7573 16068
rect 7607 16065 7619 16099
rect 7561 16059 7619 16065
rect 11606 16056 11612 16108
rect 11664 16096 11670 16108
rect 11701 16099 11759 16105
rect 11701 16096 11713 16099
rect 11664 16068 11713 16096
rect 11664 16056 11670 16068
rect 11701 16065 11713 16068
rect 11747 16065 11759 16099
rect 11701 16059 11759 16065
rect 14461 16099 14519 16105
rect 14461 16065 14473 16099
rect 14507 16096 14519 16099
rect 15286 16096 15292 16108
rect 14507 16068 15292 16096
rect 14507 16065 14519 16068
rect 14461 16059 14519 16065
rect 15286 16056 15292 16068
rect 15344 16056 15350 16108
rect 15657 16099 15715 16105
rect 15657 16065 15669 16099
rect 15703 16096 15715 16099
rect 15838 16096 15844 16108
rect 15703 16068 15844 16096
rect 15703 16065 15715 16068
rect 15657 16059 15715 16065
rect 15838 16056 15844 16068
rect 15896 16056 15902 16108
rect 18598 16056 18604 16108
rect 18656 16056 18662 16108
rect 24489 16099 24547 16105
rect 23414 16068 23612 16096
rect 9582 15988 9588 16040
rect 9640 15988 9646 16040
rect 11977 16031 12035 16037
rect 11977 15997 11989 16031
rect 12023 16028 12035 16031
rect 13446 16028 13452 16040
rect 12023 16000 13452 16028
rect 12023 15997 12035 16000
rect 11977 15991 12035 15997
rect 13446 15988 13452 16000
rect 13504 15988 13510 16040
rect 14550 15988 14556 16040
rect 14608 15988 14614 16040
rect 14645 16031 14703 16037
rect 14645 15997 14657 16031
rect 14691 15997 14703 16031
rect 14645 15991 14703 15997
rect 13725 15963 13783 15969
rect 13725 15960 13737 15963
rect 13372 15932 13737 15960
rect 12434 15852 12440 15904
rect 12492 15892 12498 15904
rect 13372 15892 13400 15932
rect 13725 15929 13737 15932
rect 13771 15960 13783 15963
rect 13906 15960 13912 15972
rect 13771 15932 13912 15960
rect 13771 15929 13783 15932
rect 13725 15923 13783 15929
rect 13906 15920 13912 15932
rect 13964 15920 13970 15972
rect 14660 15960 14688 15991
rect 19702 15988 19708 16040
rect 19760 15988 19766 16040
rect 20438 16028 20444 16040
rect 19812 16000 20444 16028
rect 14568 15932 14688 15960
rect 12492 15864 13400 15892
rect 12492 15852 12498 15864
rect 13446 15852 13452 15904
rect 13504 15892 13510 15904
rect 14568 15892 14596 15932
rect 17494 15920 17500 15972
rect 17552 15960 17558 15972
rect 19812 15960 19840 16000
rect 20438 15988 20444 16000
rect 20496 15988 20502 16040
rect 20622 15988 20628 16040
rect 20680 16028 20686 16040
rect 22005 16031 22063 16037
rect 22005 16028 22017 16031
rect 20680 16000 22017 16028
rect 20680 15988 20686 16000
rect 22005 15997 22017 16000
rect 22051 16028 22063 16031
rect 22278 16028 22284 16040
rect 22051 16000 22284 16028
rect 22051 15997 22063 16000
rect 22005 15991 22063 15997
rect 22278 15988 22284 16000
rect 22336 15988 22342 16040
rect 23584 15972 23612 16068
rect 24489 16065 24501 16099
rect 24535 16096 24547 16099
rect 25130 16096 25136 16108
rect 24535 16068 25136 16096
rect 24535 16065 24547 16068
rect 24489 16059 24547 16065
rect 25130 16056 25136 16068
rect 25188 16056 25194 16108
rect 17552 15932 19840 15960
rect 21453 15963 21511 15969
rect 17552 15920 17558 15932
rect 21453 15929 21465 15963
rect 21499 15929 21511 15963
rect 21453 15923 21511 15929
rect 13504 15864 14596 15892
rect 13504 15852 13510 15864
rect 17310 15852 17316 15904
rect 17368 15852 17374 15904
rect 19334 15852 19340 15904
rect 19392 15892 19398 15904
rect 20162 15892 20168 15904
rect 19392 15864 20168 15892
rect 19392 15852 19398 15864
rect 20162 15852 20168 15864
rect 20220 15852 20226 15904
rect 20530 15852 20536 15904
rect 20588 15892 20594 15904
rect 21468 15892 21496 15923
rect 23566 15920 23572 15972
rect 23624 15960 23630 15972
rect 24121 15963 24179 15969
rect 24121 15960 24133 15963
rect 23624 15932 24133 15960
rect 23624 15920 23630 15932
rect 24121 15929 24133 15932
rect 24167 15929 24179 15963
rect 24121 15923 24179 15929
rect 22262 15895 22320 15901
rect 22262 15892 22274 15895
rect 20588 15864 22274 15892
rect 20588 15852 20594 15864
rect 22262 15861 22274 15864
rect 22308 15861 22320 15895
rect 22262 15855 22320 15861
rect 23750 15852 23756 15904
rect 23808 15852 23814 15904
rect 1104 15802 25852 15824
rect 1104 15750 2950 15802
rect 3002 15750 3014 15802
rect 3066 15750 3078 15802
rect 3130 15750 3142 15802
rect 3194 15750 3206 15802
rect 3258 15750 12950 15802
rect 13002 15750 13014 15802
rect 13066 15750 13078 15802
rect 13130 15750 13142 15802
rect 13194 15750 13206 15802
rect 13258 15750 22950 15802
rect 23002 15750 23014 15802
rect 23066 15750 23078 15802
rect 23130 15750 23142 15802
rect 23194 15750 23206 15802
rect 23258 15750 25852 15802
rect 1104 15728 25852 15750
rect 7742 15648 7748 15700
rect 7800 15688 7806 15700
rect 8113 15691 8171 15697
rect 8113 15688 8125 15691
rect 7800 15660 8125 15688
rect 7800 15648 7806 15660
rect 8113 15657 8125 15660
rect 8159 15657 8171 15691
rect 8113 15651 8171 15657
rect 8481 15691 8539 15697
rect 8481 15657 8493 15691
rect 8527 15688 8539 15691
rect 8754 15688 8760 15700
rect 8527 15660 8760 15688
rect 8527 15657 8539 15660
rect 8481 15651 8539 15657
rect 8754 15648 8760 15660
rect 8812 15648 8818 15700
rect 9306 15648 9312 15700
rect 9364 15688 9370 15700
rect 12989 15691 13047 15697
rect 9364 15660 12434 15688
rect 9364 15648 9370 15660
rect 8772 15620 8800 15648
rect 9585 15623 9643 15629
rect 9585 15620 9597 15623
rect 8772 15592 9597 15620
rect 9585 15589 9597 15592
rect 9631 15589 9643 15623
rect 12406 15620 12434 15660
rect 12989 15657 13001 15691
rect 13035 15688 13047 15691
rect 14550 15688 14556 15700
rect 13035 15660 14556 15688
rect 13035 15657 13047 15660
rect 12989 15651 13047 15657
rect 14550 15648 14556 15660
rect 14608 15648 14614 15700
rect 16316 15660 17540 15688
rect 16316 15620 16344 15660
rect 12406 15592 16344 15620
rect 17512 15620 17540 15660
rect 17770 15648 17776 15700
rect 17828 15688 17834 15700
rect 17957 15691 18015 15697
rect 17957 15688 17969 15691
rect 17828 15660 17969 15688
rect 17828 15648 17834 15660
rect 17957 15657 17969 15660
rect 18003 15657 18015 15691
rect 21634 15688 21640 15700
rect 17957 15651 18015 15657
rect 18064 15660 21640 15688
rect 18064 15620 18092 15660
rect 21634 15648 21640 15660
rect 21692 15648 21698 15700
rect 17512 15592 18092 15620
rect 9585 15583 9643 15589
rect 6641 15555 6699 15561
rect 6641 15521 6653 15555
rect 6687 15552 6699 15555
rect 9398 15552 9404 15564
rect 6687 15524 9404 15552
rect 6687 15521 6699 15524
rect 6641 15515 6699 15521
rect 9398 15512 9404 15524
rect 9456 15512 9462 15564
rect 6362 15444 6368 15496
rect 6420 15444 6426 15496
rect 8754 15416 8760 15428
rect 7866 15388 8760 15416
rect 8754 15376 8760 15388
rect 8812 15376 8818 15428
rect 9600 15348 9628 15583
rect 11238 15512 11244 15564
rect 11296 15552 11302 15564
rect 11974 15552 11980 15564
rect 11296 15524 11980 15552
rect 11296 15512 11302 15524
rect 11974 15512 11980 15524
rect 12032 15512 12038 15564
rect 12345 15555 12403 15561
rect 12345 15521 12357 15555
rect 12391 15552 12403 15555
rect 12434 15552 12440 15564
rect 12391 15524 12440 15552
rect 12391 15521 12403 15524
rect 12345 15515 12403 15521
rect 12434 15512 12440 15524
rect 12492 15512 12498 15564
rect 12802 15512 12808 15564
rect 12860 15552 12866 15564
rect 13541 15555 13599 15561
rect 13541 15552 13553 15555
rect 12860 15524 13553 15552
rect 12860 15512 12866 15524
rect 13541 15521 13553 15524
rect 13587 15521 13599 15555
rect 13541 15515 13599 15521
rect 15286 15512 15292 15564
rect 15344 15512 15350 15564
rect 16209 15555 16267 15561
rect 16209 15521 16221 15555
rect 16255 15552 16267 15555
rect 19429 15555 19487 15561
rect 19429 15552 19441 15555
rect 16255 15524 19441 15552
rect 16255 15521 16267 15524
rect 16209 15515 16267 15521
rect 19429 15521 19441 15524
rect 19475 15552 19487 15555
rect 19702 15552 19708 15564
rect 19475 15524 19708 15552
rect 19475 15521 19487 15524
rect 19429 15515 19487 15521
rect 19702 15512 19708 15524
rect 19760 15512 19766 15564
rect 20438 15512 20444 15564
rect 20496 15552 20502 15564
rect 20496 15524 21864 15552
rect 20496 15512 20502 15524
rect 9950 15444 9956 15496
rect 10008 15444 10014 15496
rect 18693 15487 18751 15493
rect 18693 15453 18705 15487
rect 18739 15484 18751 15487
rect 19334 15484 19340 15496
rect 18739 15456 19340 15484
rect 18739 15453 18751 15456
rect 18693 15447 18751 15453
rect 19334 15444 19340 15456
rect 19392 15444 19398 15496
rect 21836 15493 21864 15524
rect 22278 15512 22284 15564
rect 22336 15512 22342 15564
rect 22557 15555 22615 15561
rect 22557 15521 22569 15555
rect 22603 15552 22615 15555
rect 25225 15555 25283 15561
rect 25225 15552 25237 15555
rect 22603 15524 25237 15552
rect 22603 15521 22615 15524
rect 22557 15515 22615 15521
rect 25225 15521 25237 15524
rect 25271 15521 25283 15555
rect 25225 15515 25283 15521
rect 21821 15487 21879 15493
rect 21821 15453 21833 15487
rect 21867 15453 21879 15487
rect 21821 15447 21879 15453
rect 23842 15444 23848 15496
rect 23900 15484 23906 15496
rect 24581 15487 24639 15493
rect 24581 15484 24593 15487
rect 23900 15456 24593 15484
rect 23900 15444 23906 15456
rect 24581 15453 24593 15456
rect 24627 15453 24639 15487
rect 24581 15447 24639 15453
rect 10226 15376 10232 15428
rect 10284 15376 10290 15428
rect 13449 15419 13507 15425
rect 10336 15388 10718 15416
rect 10336 15348 10364 15388
rect 13449 15385 13461 15419
rect 13495 15416 13507 15419
rect 14829 15419 14887 15425
rect 14829 15416 14841 15419
rect 13495 15388 14841 15416
rect 13495 15385 13507 15388
rect 13449 15379 13507 15385
rect 14829 15385 14841 15388
rect 14875 15416 14887 15419
rect 16485 15419 16543 15425
rect 14875 15388 16436 15416
rect 14875 15385 14887 15388
rect 14829 15379 14887 15385
rect 9600 15320 10364 15348
rect 12710 15308 12716 15360
rect 12768 15348 12774 15360
rect 13354 15348 13360 15360
rect 12768 15320 13360 15348
rect 12768 15308 12774 15320
rect 13354 15308 13360 15320
rect 13412 15308 13418 15360
rect 14274 15308 14280 15360
rect 14332 15308 14338 15360
rect 15841 15351 15899 15357
rect 15841 15317 15853 15351
rect 15887 15348 15899 15351
rect 16022 15348 16028 15360
rect 15887 15320 16028 15348
rect 15887 15317 15899 15320
rect 15841 15311 15899 15317
rect 16022 15308 16028 15320
rect 16080 15308 16086 15360
rect 16408 15348 16436 15388
rect 16485 15385 16497 15419
rect 16531 15416 16543 15419
rect 16574 15416 16580 15428
rect 16531 15388 16580 15416
rect 16531 15385 16543 15388
rect 16485 15379 16543 15385
rect 16574 15376 16580 15388
rect 16632 15376 16638 15428
rect 16942 15376 16948 15428
rect 17000 15376 17006 15428
rect 19705 15419 19763 15425
rect 19705 15385 19717 15419
rect 19751 15416 19763 15419
rect 21910 15416 21916 15428
rect 19751 15388 19932 15416
rect 20930 15388 21916 15416
rect 19751 15385 19763 15388
rect 19705 15379 19763 15385
rect 19904 15360 19932 15388
rect 21910 15376 21916 15388
rect 21968 15376 21974 15428
rect 23566 15376 23572 15428
rect 23624 15376 23630 15428
rect 17218 15348 17224 15360
rect 16408 15320 17224 15348
rect 17218 15308 17224 15320
rect 17276 15308 17282 15360
rect 18509 15351 18567 15357
rect 18509 15317 18521 15351
rect 18555 15348 18567 15351
rect 18782 15348 18788 15360
rect 18555 15320 18788 15348
rect 18555 15317 18567 15320
rect 18509 15311 18567 15317
rect 18782 15308 18788 15320
rect 18840 15308 18846 15360
rect 19518 15308 19524 15360
rect 19576 15348 19582 15360
rect 19886 15348 19892 15360
rect 19576 15320 19892 15348
rect 19576 15308 19582 15320
rect 19886 15308 19892 15320
rect 19944 15308 19950 15360
rect 20990 15308 20996 15360
rect 21048 15348 21054 15360
rect 21177 15351 21235 15357
rect 21177 15348 21189 15351
rect 21048 15320 21189 15348
rect 21048 15308 21054 15320
rect 21177 15317 21189 15320
rect 21223 15317 21235 15351
rect 21177 15311 21235 15317
rect 21634 15308 21640 15360
rect 21692 15308 21698 15360
rect 22462 15308 22468 15360
rect 22520 15348 22526 15360
rect 24029 15351 24087 15357
rect 24029 15348 24041 15351
rect 22520 15320 24041 15348
rect 22520 15308 22526 15320
rect 24029 15317 24041 15320
rect 24075 15317 24087 15351
rect 24029 15311 24087 15317
rect 1104 15258 25852 15280
rect 1104 15206 7950 15258
rect 8002 15206 8014 15258
rect 8066 15206 8078 15258
rect 8130 15206 8142 15258
rect 8194 15206 8206 15258
rect 8258 15206 17950 15258
rect 18002 15206 18014 15258
rect 18066 15206 18078 15258
rect 18130 15206 18142 15258
rect 18194 15206 18206 15258
rect 18258 15206 25852 15258
rect 1104 15184 25852 15206
rect 6178 15104 6184 15156
rect 6236 15144 6242 15156
rect 7285 15147 7343 15153
rect 7285 15144 7297 15147
rect 6236 15116 7297 15144
rect 6236 15104 6242 15116
rect 7285 15113 7297 15116
rect 7331 15113 7343 15147
rect 7285 15107 7343 15113
rect 10597 15147 10655 15153
rect 10597 15113 10609 15147
rect 10643 15144 10655 15147
rect 10643 15116 11284 15144
rect 10643 15113 10655 15116
rect 10597 15107 10655 15113
rect 8754 15036 8760 15088
rect 8812 15036 8818 15088
rect 9769 15079 9827 15085
rect 9769 15045 9781 15079
rect 9815 15076 9827 15079
rect 10226 15076 10232 15088
rect 9815 15048 10232 15076
rect 9815 15045 9827 15048
rect 9769 15039 9827 15045
rect 10226 15036 10232 15048
rect 10284 15036 10290 15088
rect 11256 15076 11284 15116
rect 11330 15104 11336 15156
rect 11388 15104 11394 15156
rect 12710 15144 12716 15156
rect 11624 15116 12716 15144
rect 11514 15076 11520 15088
rect 11256 15048 11520 15076
rect 11514 15036 11520 15048
rect 11572 15036 11578 15088
rect 3418 14968 3424 15020
rect 3476 15008 3482 15020
rect 5258 15008 5264 15020
rect 3476 14980 5264 15008
rect 3476 14968 3482 14980
rect 5258 14968 5264 14980
rect 5316 14968 5322 15020
rect 6641 15011 6699 15017
rect 6641 14977 6653 15011
rect 6687 15008 6699 15011
rect 7558 15008 7564 15020
rect 6687 14980 7564 15008
rect 6687 14977 6699 14980
rect 6641 14971 6699 14977
rect 7558 14968 7564 14980
rect 7616 14968 7622 15020
rect 9674 14968 9680 15020
rect 9732 15008 9738 15020
rect 9732 14980 10824 15008
rect 9732 14968 9738 14980
rect 6362 14900 6368 14952
rect 6420 14940 6426 14952
rect 7745 14943 7803 14949
rect 7745 14940 7757 14943
rect 6420 14912 7757 14940
rect 6420 14900 6426 14912
rect 7745 14909 7757 14912
rect 7791 14909 7803 14943
rect 7745 14903 7803 14909
rect 8021 14943 8079 14949
rect 8021 14909 8033 14943
rect 8067 14940 8079 14943
rect 8570 14940 8576 14952
rect 8067 14912 8576 14940
rect 8067 14909 8079 14912
rect 8021 14903 8079 14909
rect 7760 14804 7788 14903
rect 8570 14900 8576 14912
rect 8628 14900 8634 14952
rect 10796 14949 10824 14980
rect 10962 14968 10968 15020
rect 11020 15008 11026 15020
rect 11624 15008 11652 15116
rect 12710 15104 12716 15116
rect 12768 15104 12774 15156
rect 13633 15147 13691 15153
rect 13633 15113 13645 15147
rect 13679 15144 13691 15147
rect 13722 15144 13728 15156
rect 13679 15116 13728 15144
rect 13679 15113 13691 15116
rect 13633 15107 13691 15113
rect 13722 15104 13728 15116
rect 13780 15104 13786 15156
rect 14001 15147 14059 15153
rect 14001 15113 14013 15147
rect 14047 15144 14059 15147
rect 14274 15144 14280 15156
rect 14047 15116 14280 15144
rect 14047 15113 14059 15116
rect 14001 15107 14059 15113
rect 14274 15104 14280 15116
rect 14332 15104 14338 15156
rect 15286 15104 15292 15156
rect 15344 15144 15350 15156
rect 19521 15147 19579 15153
rect 19521 15144 19533 15147
rect 15344 15116 19533 15144
rect 15344 15104 15350 15116
rect 19521 15113 19533 15116
rect 19567 15113 19579 15147
rect 19521 15107 19579 15113
rect 19794 15104 19800 15156
rect 19852 15144 19858 15156
rect 19981 15147 20039 15153
rect 19981 15144 19993 15147
rect 19852 15116 19993 15144
rect 19852 15104 19858 15116
rect 19981 15113 19993 15116
rect 20027 15113 20039 15147
rect 19981 15107 20039 15113
rect 20346 15104 20352 15156
rect 20404 15144 20410 15156
rect 21177 15147 21235 15153
rect 21177 15144 21189 15147
rect 20404 15116 21189 15144
rect 20404 15104 20410 15116
rect 21177 15113 21189 15116
rect 21223 15113 21235 15147
rect 21177 15107 21235 15113
rect 21910 15104 21916 15156
rect 21968 15144 21974 15156
rect 22097 15147 22155 15153
rect 22097 15144 22109 15147
rect 21968 15116 22109 15144
rect 21968 15104 21974 15116
rect 22097 15113 22109 15116
rect 22143 15144 22155 15147
rect 23566 15144 23572 15156
rect 22143 15116 23572 15144
rect 22143 15113 22155 15116
rect 22097 15107 22155 15113
rect 23566 15104 23572 15116
rect 23624 15104 23630 15156
rect 12618 15036 12624 15088
rect 12676 15076 12682 15088
rect 14182 15076 14188 15088
rect 12676 15048 14188 15076
rect 12676 15036 12682 15048
rect 14182 15036 14188 15048
rect 14240 15076 14246 15088
rect 14458 15076 14464 15088
rect 14240 15048 14464 15076
rect 14240 15036 14246 15048
rect 14458 15036 14464 15048
rect 14516 15036 14522 15088
rect 16206 15076 16212 15088
rect 14844 15048 16212 15076
rect 11020 14980 11652 15008
rect 11701 15011 11759 15017
rect 11020 14968 11026 14980
rect 11701 14977 11713 15011
rect 11747 15008 11759 15011
rect 13446 15008 13452 15020
rect 11747 14980 13452 15008
rect 11747 14977 11759 14980
rect 11701 14971 11759 14977
rect 13446 14968 13452 14980
rect 13504 14968 13510 15020
rect 14093 15011 14151 15017
rect 14093 14977 14105 15011
rect 14139 15008 14151 15011
rect 14550 15008 14556 15020
rect 14139 14980 14556 15008
rect 14139 14977 14151 14980
rect 14093 14971 14151 14977
rect 10689 14943 10747 14949
rect 10689 14909 10701 14943
rect 10735 14909 10747 14943
rect 10689 14903 10747 14909
rect 10781 14943 10839 14949
rect 10781 14909 10793 14943
rect 10827 14909 10839 14943
rect 10781 14903 10839 14909
rect 13357 14943 13415 14949
rect 13357 14909 13369 14943
rect 13403 14940 13415 14943
rect 14108 14940 14136 14971
rect 14550 14968 14556 14980
rect 14608 14968 14614 15020
rect 13403 14912 14136 14940
rect 14277 14943 14335 14949
rect 13403 14909 13415 14912
rect 13357 14903 13415 14909
rect 14277 14909 14289 14943
rect 14323 14940 14335 14943
rect 14844 14940 14872 15048
rect 16206 15036 16212 15048
rect 16264 15036 16270 15088
rect 16942 15036 16948 15088
rect 17000 15076 17006 15088
rect 18049 15079 18107 15085
rect 18049 15076 18061 15079
rect 17000 15048 18061 15076
rect 17000 15036 17006 15048
rect 18049 15045 18061 15048
rect 18095 15045 18107 15079
rect 18049 15039 18107 15045
rect 18601 15079 18659 15085
rect 18601 15045 18613 15079
rect 18647 15076 18659 15079
rect 18966 15076 18972 15088
rect 18647 15048 18972 15076
rect 18647 15045 18659 15048
rect 18601 15039 18659 15045
rect 18966 15036 18972 15048
rect 19024 15036 19030 15088
rect 20806 15036 20812 15088
rect 20864 15076 20870 15088
rect 20864 15048 21404 15076
rect 20864 15036 20870 15048
rect 14921 15011 14979 15017
rect 14921 14977 14933 15011
rect 14967 15008 14979 15011
rect 15933 15011 15991 15017
rect 15933 15008 15945 15011
rect 14967 14980 15945 15008
rect 14967 14977 14979 14980
rect 14921 14971 14979 14977
rect 15933 14977 15945 14980
rect 15979 14977 15991 15011
rect 18690 15008 18696 15020
rect 15933 14971 15991 14977
rect 16224 14980 18696 15008
rect 14323 14912 14872 14940
rect 14323 14909 14335 14912
rect 14277 14903 14335 14909
rect 10134 14832 10140 14884
rect 10192 14872 10198 14884
rect 10229 14875 10287 14881
rect 10229 14872 10241 14875
rect 10192 14844 10241 14872
rect 10192 14832 10198 14844
rect 10229 14841 10241 14844
rect 10275 14841 10287 14875
rect 10704 14872 10732 14903
rect 16022 14900 16028 14952
rect 16080 14900 16086 14952
rect 16224 14949 16252 14980
rect 18690 14968 18696 14980
rect 18748 14968 18754 15020
rect 18874 14968 18880 15020
rect 18932 15008 18938 15020
rect 19889 15011 19947 15017
rect 19889 15008 19901 15011
rect 18932 14980 19901 15008
rect 18932 14968 18938 14980
rect 19889 14977 19901 14980
rect 19935 14977 19947 15011
rect 19889 14971 19947 14977
rect 21082 14968 21088 15020
rect 21140 14968 21146 15020
rect 21376 15008 21404 15048
rect 21450 15036 21456 15088
rect 21508 15076 21514 15088
rect 21508 15048 23980 15076
rect 21508 15036 21514 15048
rect 22462 15008 22468 15020
rect 21376 14980 22468 15008
rect 22462 14968 22468 14980
rect 22520 14968 22526 15020
rect 23952 15017 23980 15048
rect 23937 15011 23995 15017
rect 23937 14977 23949 15011
rect 23983 14977 23995 15011
rect 23937 14971 23995 14977
rect 16209 14943 16267 14949
rect 16209 14909 16221 14943
rect 16255 14909 16267 14943
rect 16209 14903 16267 14909
rect 16853 14943 16911 14949
rect 16853 14909 16865 14943
rect 16899 14909 16911 14943
rect 16853 14903 16911 14909
rect 17129 14943 17187 14949
rect 17129 14909 17141 14943
rect 17175 14940 17187 14943
rect 19794 14940 19800 14952
rect 17175 14912 19800 14940
rect 17175 14909 17187 14912
rect 17129 14903 17187 14909
rect 11422 14872 11428 14884
rect 10704 14844 11428 14872
rect 10229 14835 10287 14841
rect 11422 14832 11428 14844
rect 11480 14832 11486 14884
rect 12897 14875 12955 14881
rect 12897 14841 12909 14875
rect 12943 14872 12955 14875
rect 13446 14872 13452 14884
rect 12943 14844 13452 14872
rect 12943 14841 12955 14844
rect 12897 14835 12955 14841
rect 13446 14832 13452 14844
rect 13504 14832 13510 14884
rect 15562 14832 15568 14884
rect 15620 14832 15626 14884
rect 16868 14872 16896 14903
rect 19794 14900 19800 14912
rect 19852 14900 19858 14952
rect 20165 14943 20223 14949
rect 20165 14909 20177 14943
rect 20211 14940 20223 14943
rect 20990 14940 20996 14952
rect 20211 14912 20996 14940
rect 20211 14909 20223 14912
rect 20165 14903 20223 14909
rect 20990 14900 20996 14912
rect 21048 14900 21054 14952
rect 21361 14943 21419 14949
rect 21361 14909 21373 14943
rect 21407 14940 21419 14943
rect 23750 14940 23756 14952
rect 21407 14912 23756 14940
rect 21407 14909 21419 14912
rect 21361 14903 21419 14909
rect 23750 14900 23756 14912
rect 23808 14900 23814 14952
rect 24762 14900 24768 14952
rect 24820 14900 24826 14952
rect 19426 14872 19432 14884
rect 16868 14844 19432 14872
rect 19426 14832 19432 14844
rect 19484 14832 19490 14884
rect 19702 14832 19708 14884
rect 19760 14872 19766 14884
rect 25590 14872 25596 14884
rect 19760 14844 25596 14872
rect 19760 14832 19766 14844
rect 25590 14832 25596 14844
rect 25648 14832 25654 14884
rect 9950 14804 9956 14816
rect 7760 14776 9956 14804
rect 9950 14764 9956 14776
rect 10008 14764 10014 14816
rect 10318 14764 10324 14816
rect 10376 14804 10382 14816
rect 12345 14807 12403 14813
rect 12345 14804 12357 14807
rect 10376 14776 12357 14804
rect 10376 14764 10382 14776
rect 12345 14773 12357 14776
rect 12391 14773 12403 14807
rect 12345 14767 12403 14773
rect 13173 14807 13231 14813
rect 13173 14773 13185 14807
rect 13219 14804 13231 14807
rect 13538 14804 13544 14816
rect 13219 14776 13544 14804
rect 13219 14773 13231 14776
rect 13173 14767 13231 14773
rect 13538 14764 13544 14776
rect 13596 14764 13602 14816
rect 18690 14764 18696 14816
rect 18748 14764 18754 14816
rect 19058 14764 19064 14816
rect 19116 14804 19122 14816
rect 20717 14807 20775 14813
rect 20717 14804 20729 14807
rect 19116 14776 20729 14804
rect 19116 14764 19122 14776
rect 20717 14773 20729 14776
rect 20763 14773 20775 14807
rect 20717 14767 20775 14773
rect 22554 14764 22560 14816
rect 22612 14804 22618 14816
rect 23109 14807 23167 14813
rect 23109 14804 23121 14807
rect 22612 14776 23121 14804
rect 22612 14764 22618 14776
rect 23109 14773 23121 14776
rect 23155 14773 23167 14807
rect 23109 14767 23167 14773
rect 23477 14807 23535 14813
rect 23477 14773 23489 14807
rect 23523 14804 23535 14807
rect 23566 14804 23572 14816
rect 23523 14776 23572 14804
rect 23523 14773 23535 14776
rect 23477 14767 23535 14773
rect 23566 14764 23572 14776
rect 23624 14804 23630 14816
rect 23661 14807 23719 14813
rect 23661 14804 23673 14807
rect 23624 14776 23673 14804
rect 23624 14764 23630 14776
rect 23661 14773 23673 14776
rect 23707 14804 23719 14807
rect 23842 14804 23848 14816
rect 23707 14776 23848 14804
rect 23707 14773 23719 14776
rect 23661 14767 23719 14773
rect 23842 14764 23848 14776
rect 23900 14764 23906 14816
rect 1104 14714 25852 14736
rect 1104 14662 2950 14714
rect 3002 14662 3014 14714
rect 3066 14662 3078 14714
rect 3130 14662 3142 14714
rect 3194 14662 3206 14714
rect 3258 14662 12950 14714
rect 13002 14662 13014 14714
rect 13066 14662 13078 14714
rect 13130 14662 13142 14714
rect 13194 14662 13206 14714
rect 13258 14662 22950 14714
rect 23002 14662 23014 14714
rect 23066 14662 23078 14714
rect 23130 14662 23142 14714
rect 23194 14662 23206 14714
rect 23258 14662 25852 14714
rect 1104 14640 25852 14662
rect 8570 14560 8576 14612
rect 8628 14560 8634 14612
rect 9030 14560 9036 14612
rect 9088 14600 9094 14612
rect 9125 14603 9183 14609
rect 9125 14600 9137 14603
rect 9088 14572 9137 14600
rect 9088 14560 9094 14572
rect 9125 14569 9137 14572
rect 9171 14569 9183 14603
rect 9125 14563 9183 14569
rect 11698 14560 11704 14612
rect 11756 14560 11762 14612
rect 14366 14560 14372 14612
rect 14424 14560 14430 14612
rect 14734 14560 14740 14612
rect 14792 14600 14798 14612
rect 16850 14600 16856 14612
rect 14792 14572 16856 14600
rect 14792 14560 14798 14572
rect 16850 14560 16856 14572
rect 16908 14560 16914 14612
rect 18322 14560 18328 14612
rect 18380 14560 18386 14612
rect 19426 14560 19432 14612
rect 19484 14600 19490 14612
rect 19521 14603 19579 14609
rect 19521 14600 19533 14603
rect 19484 14572 19533 14600
rect 19484 14560 19490 14572
rect 19521 14569 19533 14572
rect 19567 14569 19579 14603
rect 19521 14563 19579 14569
rect 20901 14603 20959 14609
rect 20901 14569 20913 14603
rect 20947 14600 20959 14603
rect 22646 14600 22652 14612
rect 20947 14572 22652 14600
rect 20947 14569 20959 14572
rect 20901 14563 20959 14569
rect 22646 14560 22652 14572
rect 22704 14560 22710 14612
rect 12342 14492 12348 14544
rect 12400 14532 12406 14544
rect 15013 14535 15071 14541
rect 15013 14532 15025 14535
rect 12400 14504 15025 14532
rect 12400 14492 12406 14504
rect 15013 14501 15025 14504
rect 15059 14501 15071 14535
rect 15013 14495 15071 14501
rect 15102 14492 15108 14544
rect 15160 14532 15166 14544
rect 19058 14532 19064 14544
rect 15160 14504 19064 14532
rect 15160 14492 15166 14504
rect 19058 14492 19064 14504
rect 19116 14492 19122 14544
rect 19334 14492 19340 14544
rect 19392 14532 19398 14544
rect 20070 14532 20076 14544
rect 19392 14504 20076 14532
rect 19392 14492 19398 14504
rect 20070 14492 20076 14504
rect 20128 14492 20134 14544
rect 21821 14535 21879 14541
rect 21821 14501 21833 14535
rect 21867 14532 21879 14535
rect 22278 14532 22284 14544
rect 21867 14504 22284 14532
rect 21867 14501 21879 14504
rect 21821 14495 21879 14501
rect 22278 14492 22284 14504
rect 22336 14492 22342 14544
rect 7558 14424 7564 14476
rect 7616 14464 7622 14476
rect 9674 14464 9680 14476
rect 7616 14436 9680 14464
rect 7616 14424 7622 14436
rect 9674 14424 9680 14436
rect 9732 14424 9738 14476
rect 9950 14424 9956 14476
rect 10008 14464 10014 14476
rect 11057 14467 11115 14473
rect 11057 14464 11069 14467
rect 10008 14436 11069 14464
rect 10008 14424 10014 14436
rect 11057 14433 11069 14436
rect 11103 14433 11115 14467
rect 11057 14427 11115 14433
rect 11974 14424 11980 14476
rect 12032 14464 12038 14476
rect 12253 14467 12311 14473
rect 12253 14464 12265 14467
rect 12032 14436 12265 14464
rect 12032 14424 12038 14436
rect 12253 14433 12265 14436
rect 12299 14433 12311 14467
rect 12253 14427 12311 14433
rect 13446 14424 13452 14476
rect 13504 14424 13510 14476
rect 13633 14467 13691 14473
rect 13633 14433 13645 14467
rect 13679 14464 13691 14467
rect 15378 14464 15384 14476
rect 13679 14436 15384 14464
rect 13679 14433 13691 14436
rect 13633 14427 13691 14433
rect 7742 14356 7748 14408
rect 7800 14396 7806 14408
rect 7929 14399 7987 14405
rect 7929 14396 7941 14399
rect 7800 14368 7941 14396
rect 7800 14356 7806 14368
rect 7929 14365 7941 14368
rect 7975 14365 7987 14399
rect 7929 14359 7987 14365
rect 8938 14356 8944 14408
rect 8996 14396 9002 14408
rect 9582 14396 9588 14408
rect 8996 14368 9588 14396
rect 8996 14356 9002 14368
rect 9582 14356 9588 14368
rect 9640 14356 9646 14408
rect 10321 14399 10379 14405
rect 10321 14365 10333 14399
rect 10367 14396 10379 14399
rect 11330 14396 11336 14408
rect 10367 14368 11336 14396
rect 10367 14365 10379 14368
rect 10321 14359 10379 14365
rect 11330 14356 11336 14368
rect 11388 14356 11394 14408
rect 13648 14396 13676 14427
rect 15378 14424 15384 14436
rect 15436 14424 15442 14476
rect 15562 14424 15568 14476
rect 15620 14424 15626 14476
rect 17221 14467 17279 14473
rect 17221 14433 17233 14467
rect 17267 14464 17279 14467
rect 18322 14464 18328 14476
rect 17267 14436 18328 14464
rect 17267 14433 17279 14436
rect 17221 14427 17279 14433
rect 18322 14424 18328 14436
rect 18380 14424 18386 14476
rect 19150 14424 19156 14476
rect 19208 14464 19214 14476
rect 19208 14436 19748 14464
rect 19208 14424 19214 14436
rect 11440 14368 13676 14396
rect 14553 14399 14611 14405
rect 9600 14328 9628 14356
rect 11440 14328 11468 14368
rect 14553 14365 14565 14399
rect 14599 14396 14611 14399
rect 15194 14396 15200 14408
rect 14599 14368 15200 14396
rect 14599 14365 14611 14368
rect 14553 14359 14611 14365
rect 15194 14356 15200 14368
rect 15252 14356 15258 14408
rect 17497 14399 17555 14405
rect 17497 14365 17509 14399
rect 17543 14365 17555 14399
rect 17497 14359 17555 14365
rect 18877 14399 18935 14405
rect 18877 14365 18889 14399
rect 18923 14396 18935 14399
rect 19334 14396 19340 14408
rect 18923 14368 19340 14396
rect 18923 14365 18935 14368
rect 18877 14359 18935 14365
rect 9600 14300 11468 14328
rect 12069 14331 12127 14337
rect 12069 14297 12081 14331
rect 12115 14328 12127 14331
rect 12526 14328 12532 14340
rect 12115 14300 12532 14328
rect 12115 14297 12127 14300
rect 12069 14291 12127 14297
rect 12526 14288 12532 14300
rect 12584 14288 12590 14340
rect 13357 14331 13415 14337
rect 13357 14297 13369 14331
rect 13403 14328 13415 14331
rect 13538 14328 13544 14340
rect 13403 14300 13544 14328
rect 13403 14297 13415 14300
rect 13357 14291 13415 14297
rect 13538 14288 13544 14300
rect 13596 14288 13602 14340
rect 17512 14328 17540 14359
rect 19334 14356 19340 14368
rect 19392 14356 19398 14408
rect 19720 14405 19748 14436
rect 19794 14424 19800 14476
rect 19852 14464 19858 14476
rect 22186 14464 22192 14476
rect 19852 14436 22192 14464
rect 19852 14424 19858 14436
rect 22186 14424 22192 14436
rect 22244 14424 22250 14476
rect 22554 14424 22560 14476
rect 22612 14424 22618 14476
rect 19705 14399 19763 14405
rect 19705 14365 19717 14399
rect 19751 14365 19763 14399
rect 19705 14359 19763 14365
rect 20349 14399 20407 14405
rect 20349 14365 20361 14399
rect 20395 14365 20407 14399
rect 20349 14359 20407 14365
rect 19794 14328 19800 14340
rect 15396 14300 16344 14328
rect 17512 14300 19800 14328
rect 9490 14220 9496 14272
rect 9548 14220 9554 14272
rect 9582 14220 9588 14272
rect 9640 14220 9646 14272
rect 10226 14220 10232 14272
rect 10284 14260 10290 14272
rect 10962 14260 10968 14272
rect 10284 14232 10968 14260
rect 10284 14220 10290 14232
rect 10962 14220 10968 14232
rect 11020 14220 11026 14272
rect 12161 14263 12219 14269
rect 12161 14229 12173 14263
rect 12207 14260 12219 14263
rect 12710 14260 12716 14272
rect 12207 14232 12716 14260
rect 12207 14229 12219 14232
rect 12161 14223 12219 14229
rect 12710 14220 12716 14232
rect 12768 14220 12774 14272
rect 12802 14220 12808 14272
rect 12860 14260 12866 14272
rect 15396 14269 15424 14300
rect 16316 14272 16344 14300
rect 19794 14288 19800 14300
rect 19852 14288 19858 14340
rect 20364 14328 20392 14359
rect 20714 14356 20720 14408
rect 20772 14396 20778 14408
rect 21085 14399 21143 14405
rect 21085 14396 21097 14399
rect 20772 14368 21097 14396
rect 20772 14356 20778 14368
rect 21085 14365 21097 14368
rect 21131 14365 21143 14399
rect 21726 14396 21732 14408
rect 21085 14359 21143 14365
rect 21192 14368 21732 14396
rect 21192 14328 21220 14368
rect 21726 14356 21732 14368
rect 21784 14356 21790 14408
rect 22278 14356 22284 14408
rect 22336 14356 22342 14408
rect 24670 14356 24676 14408
rect 24728 14396 24734 14408
rect 24765 14399 24823 14405
rect 24765 14396 24777 14399
rect 24728 14368 24777 14396
rect 24728 14356 24734 14368
rect 24765 14365 24777 14368
rect 24811 14365 24823 14399
rect 24765 14359 24823 14365
rect 21637 14331 21695 14337
rect 21637 14328 21649 14331
rect 20364 14300 21220 14328
rect 21284 14300 21649 14328
rect 12989 14263 13047 14269
rect 12989 14260 13001 14263
rect 12860 14232 13001 14260
rect 12860 14220 12866 14232
rect 12989 14229 13001 14232
rect 13035 14229 13047 14263
rect 12989 14223 13047 14229
rect 15381 14263 15439 14269
rect 15381 14229 15393 14263
rect 15427 14229 15439 14263
rect 15381 14223 15439 14229
rect 15473 14263 15531 14269
rect 15473 14229 15485 14263
rect 15519 14260 15531 14263
rect 16022 14260 16028 14272
rect 15519 14232 16028 14260
rect 15519 14229 15531 14232
rect 15473 14223 15531 14229
rect 16022 14220 16028 14232
rect 16080 14220 16086 14272
rect 16298 14220 16304 14272
rect 16356 14220 16362 14272
rect 16574 14220 16580 14272
rect 16632 14220 16638 14272
rect 18693 14263 18751 14269
rect 18693 14229 18705 14263
rect 18739 14260 18751 14263
rect 19426 14260 19432 14272
rect 18739 14232 19432 14260
rect 18739 14229 18751 14232
rect 18693 14223 18751 14229
rect 19426 14220 19432 14232
rect 19484 14220 19490 14272
rect 19886 14220 19892 14272
rect 19944 14260 19950 14272
rect 20165 14263 20223 14269
rect 20165 14260 20177 14263
rect 19944 14232 20177 14260
rect 19944 14220 19950 14232
rect 20165 14229 20177 14232
rect 20211 14229 20223 14263
rect 20165 14223 20223 14229
rect 20346 14220 20352 14272
rect 20404 14260 20410 14272
rect 21284 14260 21312 14300
rect 21637 14297 21649 14300
rect 21683 14297 21695 14331
rect 23842 14328 23848 14340
rect 23782 14300 23848 14328
rect 21637 14291 21695 14297
rect 23842 14288 23848 14300
rect 23900 14328 23906 14340
rect 23900 14300 25084 14328
rect 23900 14288 23906 14300
rect 25056 14272 25084 14300
rect 20404 14232 21312 14260
rect 20404 14220 20410 14232
rect 21358 14220 21364 14272
rect 21416 14260 21422 14272
rect 22094 14260 22100 14272
rect 21416 14232 22100 14260
rect 21416 14220 21422 14232
rect 22094 14220 22100 14232
rect 22152 14220 22158 14272
rect 24026 14220 24032 14272
rect 24084 14220 24090 14272
rect 24486 14220 24492 14272
rect 24544 14260 24550 14272
rect 24581 14263 24639 14269
rect 24581 14260 24593 14263
rect 24544 14232 24593 14260
rect 24544 14220 24550 14232
rect 24581 14229 24593 14232
rect 24627 14229 24639 14263
rect 24581 14223 24639 14229
rect 25038 14220 25044 14272
rect 25096 14220 25102 14272
rect 1104 14170 25852 14192
rect 1104 14118 7950 14170
rect 8002 14118 8014 14170
rect 8066 14118 8078 14170
rect 8130 14118 8142 14170
rect 8194 14118 8206 14170
rect 8258 14118 17950 14170
rect 18002 14118 18014 14170
rect 18066 14118 18078 14170
rect 18130 14118 18142 14170
rect 18194 14118 18206 14170
rect 18258 14118 25852 14170
rect 1104 14096 25852 14118
rect 8294 14016 8300 14068
rect 8352 14056 8358 14068
rect 9125 14059 9183 14065
rect 9125 14056 9137 14059
rect 8352 14028 9137 14056
rect 8352 14016 8358 14028
rect 9125 14025 9137 14028
rect 9171 14025 9183 14059
rect 9125 14019 9183 14025
rect 9490 14016 9496 14068
rect 9548 14056 9554 14068
rect 10413 14059 10471 14065
rect 10413 14056 10425 14059
rect 9548 14028 10425 14056
rect 9548 14016 9554 14028
rect 10413 14025 10425 14028
rect 10459 14025 10471 14059
rect 10413 14019 10471 14025
rect 12250 14016 12256 14068
rect 12308 14056 12314 14068
rect 12345 14059 12403 14065
rect 12345 14056 12357 14059
rect 12308 14028 12357 14056
rect 12308 14016 12314 14028
rect 12345 14025 12357 14028
rect 12391 14025 12403 14059
rect 12345 14019 12403 14025
rect 12713 14059 12771 14065
rect 12713 14025 12725 14059
rect 12759 14056 12771 14059
rect 14642 14056 14648 14068
rect 12759 14028 14648 14056
rect 12759 14025 12771 14028
rect 12713 14019 12771 14025
rect 14642 14016 14648 14028
rect 14700 14016 14706 14068
rect 15841 14059 15899 14065
rect 15841 14025 15853 14059
rect 15887 14056 15899 14059
rect 16482 14056 16488 14068
rect 15887 14028 16488 14056
rect 15887 14025 15899 14028
rect 15841 14019 15899 14025
rect 7098 13988 7104 14000
rect 6564 13960 7104 13988
rect 6362 13880 6368 13932
rect 6420 13920 6426 13932
rect 6564 13929 6592 13960
rect 7098 13948 7104 13960
rect 7156 13948 7162 14000
rect 8665 13991 8723 13997
rect 8665 13988 8677 13991
rect 8050 13960 8677 13988
rect 8665 13957 8677 13960
rect 8711 13988 8723 13991
rect 8754 13988 8760 14000
rect 8711 13960 8760 13988
rect 8711 13957 8723 13960
rect 8665 13951 8723 13957
rect 8754 13948 8760 13960
rect 8812 13948 8818 14000
rect 10134 13988 10140 14000
rect 9508 13960 10140 13988
rect 9508 13929 9536 13960
rect 10134 13948 10140 13960
rect 10192 13948 10198 14000
rect 10873 13991 10931 13997
rect 10873 13957 10885 13991
rect 10919 13988 10931 13991
rect 12618 13988 12624 14000
rect 10919 13960 12624 13988
rect 10919 13957 10931 13960
rect 10873 13951 10931 13957
rect 12618 13948 12624 13960
rect 12676 13948 12682 14000
rect 6549 13923 6607 13929
rect 6549 13920 6561 13923
rect 6420 13892 6561 13920
rect 6420 13880 6426 13892
rect 6549 13889 6561 13892
rect 6595 13889 6607 13923
rect 6549 13883 6607 13889
rect 9493 13923 9551 13929
rect 9493 13889 9505 13923
rect 9539 13889 9551 13923
rect 9493 13883 9551 13889
rect 9585 13923 9643 13929
rect 9585 13889 9597 13923
rect 9631 13920 9643 13923
rect 9766 13920 9772 13932
rect 9631 13892 9772 13920
rect 9631 13889 9643 13892
rect 9585 13883 9643 13889
rect 9766 13880 9772 13892
rect 9824 13880 9830 13932
rect 10781 13923 10839 13929
rect 10781 13889 10793 13923
rect 10827 13920 10839 13923
rect 11701 13923 11759 13929
rect 11701 13920 11713 13923
rect 10827 13892 11713 13920
rect 10827 13889 10839 13892
rect 10781 13883 10839 13889
rect 11701 13889 11713 13892
rect 11747 13889 11759 13923
rect 11701 13883 11759 13889
rect 12805 13923 12863 13929
rect 12805 13889 12817 13923
rect 12851 13920 12863 13923
rect 13446 13920 13452 13932
rect 12851 13892 13452 13920
rect 12851 13889 12863 13892
rect 12805 13883 12863 13889
rect 13446 13880 13452 13892
rect 13504 13880 13510 13932
rect 14918 13880 14924 13932
rect 14976 13880 14982 13932
rect 15562 13920 15568 13932
rect 15120 13892 15568 13920
rect 7558 13812 7564 13864
rect 7616 13852 7622 13864
rect 8297 13855 8355 13861
rect 8297 13852 8309 13855
rect 7616 13824 8309 13852
rect 7616 13812 7622 13824
rect 8297 13821 8309 13824
rect 8343 13821 8355 13855
rect 8297 13815 8355 13821
rect 9398 13812 9404 13864
rect 9456 13852 9462 13864
rect 9677 13855 9735 13861
rect 9677 13852 9689 13855
rect 9456 13824 9689 13852
rect 9456 13812 9462 13824
rect 9677 13821 9689 13824
rect 9723 13821 9735 13855
rect 9677 13815 9735 13821
rect 11057 13855 11115 13861
rect 11057 13821 11069 13855
rect 11103 13821 11115 13855
rect 11057 13815 11115 13821
rect 12897 13855 12955 13861
rect 12897 13821 12909 13855
rect 12943 13821 12955 13855
rect 12897 13815 12955 13821
rect 6812 13719 6870 13725
rect 6812 13685 6824 13719
rect 6858 13716 6870 13719
rect 9490 13716 9496 13728
rect 6858 13688 9496 13716
rect 6858 13685 6870 13688
rect 6812 13679 6870 13685
rect 9490 13676 9496 13688
rect 9548 13716 9554 13728
rect 11072 13716 11100 13815
rect 11974 13744 11980 13796
rect 12032 13784 12038 13796
rect 12912 13784 12940 13815
rect 13538 13812 13544 13864
rect 13596 13812 13602 13864
rect 14366 13812 14372 13864
rect 14424 13852 14430 13864
rect 15120 13852 15148 13892
rect 15562 13880 15568 13892
rect 15620 13880 15626 13932
rect 14424 13824 15148 13852
rect 15289 13855 15347 13861
rect 14424 13812 14430 13824
rect 15289 13821 15301 13855
rect 15335 13852 15347 13855
rect 15838 13852 15844 13864
rect 15335 13824 15844 13852
rect 15335 13821 15347 13824
rect 15289 13815 15347 13821
rect 15838 13812 15844 13824
rect 15896 13812 15902 13864
rect 12032 13756 12940 13784
rect 12032 13744 12038 13756
rect 14918 13744 14924 13796
rect 14976 13784 14982 13796
rect 15948 13784 15976 14028
rect 16482 14016 16488 14028
rect 16540 14056 16546 14068
rect 16942 14056 16948 14068
rect 16540 14028 16948 14056
rect 16540 14016 16546 14028
rect 16942 14016 16948 14028
rect 17000 14056 17006 14068
rect 17000 14028 17264 14056
rect 17000 14016 17006 14028
rect 16117 13991 16175 13997
rect 16117 13957 16129 13991
rect 16163 13988 16175 13991
rect 17126 13988 17132 14000
rect 16163 13960 17132 13988
rect 16163 13957 16175 13960
rect 16117 13951 16175 13957
rect 17126 13948 17132 13960
rect 17184 13948 17190 14000
rect 17236 13988 17264 14028
rect 17512 14028 18276 14056
rect 17512 13988 17540 14028
rect 17236 13960 17618 13988
rect 18248 13920 18276 14028
rect 18598 14016 18604 14068
rect 18656 14016 18662 14068
rect 19794 14016 19800 14068
rect 19852 14056 19858 14068
rect 19852 14028 23060 14056
rect 19852 14016 19858 14028
rect 18414 13948 18420 14000
rect 18472 13988 18478 14000
rect 19061 13991 19119 13997
rect 19061 13988 19073 13991
rect 18472 13960 19073 13988
rect 18472 13948 18478 13960
rect 19061 13957 19073 13960
rect 19107 13957 19119 13991
rect 19061 13951 19119 13957
rect 19426 13948 19432 14000
rect 19484 13988 19490 14000
rect 19484 13960 22140 13988
rect 19484 13948 19490 13960
rect 20349 13923 20407 13929
rect 20349 13920 20361 13923
rect 18248 13906 20361 13920
rect 18262 13892 20361 13906
rect 20349 13889 20361 13892
rect 20395 13889 20407 13923
rect 20349 13883 20407 13889
rect 20809 13923 20867 13929
rect 20809 13889 20821 13923
rect 20855 13920 20867 13923
rect 21358 13920 21364 13932
rect 20855 13892 21364 13920
rect 20855 13889 20867 13892
rect 20809 13883 20867 13889
rect 21358 13880 21364 13892
rect 21416 13880 21422 13932
rect 22112 13929 22140 13960
rect 21453 13923 21511 13929
rect 21453 13889 21465 13923
rect 21499 13889 21511 13923
rect 21453 13883 21511 13889
rect 22097 13923 22155 13929
rect 22097 13889 22109 13923
rect 22143 13889 22155 13923
rect 23032 13920 23060 14028
rect 23293 13991 23351 13997
rect 23293 13957 23305 13991
rect 23339 13988 23351 13991
rect 24854 13988 24860 14000
rect 23339 13960 24860 13988
rect 23339 13957 23351 13960
rect 23293 13951 23351 13957
rect 24854 13948 24860 13960
rect 24912 13948 24918 14000
rect 25130 13948 25136 14000
rect 25188 13948 25194 14000
rect 23937 13923 23995 13929
rect 23937 13920 23949 13923
rect 23032 13892 23949 13920
rect 22097 13883 22155 13889
rect 23937 13889 23949 13892
rect 23983 13889 23995 13923
rect 23937 13883 23995 13889
rect 16853 13855 16911 13861
rect 16853 13821 16865 13855
rect 16899 13852 16911 13855
rect 17862 13852 17868 13864
rect 16899 13824 17868 13852
rect 16899 13821 16911 13824
rect 16853 13815 16911 13821
rect 17862 13812 17868 13824
rect 17920 13812 17926 13864
rect 19889 13855 19947 13861
rect 19889 13821 19901 13855
rect 19935 13852 19947 13855
rect 20254 13852 20260 13864
rect 19935 13824 20260 13852
rect 19935 13821 19947 13824
rect 19889 13815 19947 13821
rect 20254 13812 20260 13824
rect 20312 13812 20318 13864
rect 21468 13852 21496 13883
rect 22830 13852 22836 13864
rect 21468 13824 22836 13852
rect 22830 13812 22836 13824
rect 22888 13812 22894 13864
rect 21910 13784 21916 13796
rect 14976 13756 15976 13784
rect 18156 13756 21916 13784
rect 14976 13744 14982 13756
rect 11882 13716 11888 13728
rect 9548 13688 11888 13716
rect 9548 13676 9554 13688
rect 11882 13676 11888 13688
rect 11940 13676 11946 13728
rect 13804 13719 13862 13725
rect 13804 13685 13816 13719
rect 13850 13716 13862 13719
rect 15194 13716 15200 13728
rect 13850 13688 15200 13716
rect 13850 13685 13862 13688
rect 13804 13679 13862 13685
rect 15194 13676 15200 13688
rect 15252 13676 15258 13728
rect 15930 13676 15936 13728
rect 15988 13716 15994 13728
rect 16298 13716 16304 13728
rect 15988 13688 16304 13716
rect 15988 13676 15994 13688
rect 16298 13676 16304 13688
rect 16356 13676 16362 13728
rect 17116 13719 17174 13725
rect 17116 13685 17128 13719
rect 17162 13716 17174 13719
rect 17218 13716 17224 13728
rect 17162 13688 17224 13716
rect 17162 13685 17174 13688
rect 17116 13679 17174 13685
rect 17218 13676 17224 13688
rect 17276 13716 17282 13728
rect 17586 13716 17592 13728
rect 17276 13688 17592 13716
rect 17276 13676 17282 13688
rect 17586 13676 17592 13688
rect 17644 13676 17650 13728
rect 17678 13676 17684 13728
rect 17736 13716 17742 13728
rect 18156 13716 18184 13756
rect 21910 13744 21916 13756
rect 21968 13784 21974 13796
rect 26602 13784 26608 13796
rect 21968 13756 26608 13784
rect 21968 13744 21974 13756
rect 26602 13744 26608 13756
rect 26660 13744 26666 13796
rect 17736 13688 18184 13716
rect 17736 13676 17742 13688
rect 19334 13676 19340 13728
rect 19392 13716 19398 13728
rect 20530 13716 20536 13728
rect 19392 13688 20536 13716
rect 19392 13676 19398 13688
rect 20530 13676 20536 13688
rect 20588 13676 20594 13728
rect 20622 13676 20628 13728
rect 20680 13676 20686 13728
rect 21266 13676 21272 13728
rect 21324 13676 21330 13728
rect 1104 13626 25852 13648
rect 1104 13574 2950 13626
rect 3002 13574 3014 13626
rect 3066 13574 3078 13626
rect 3130 13574 3142 13626
rect 3194 13574 3206 13626
rect 3258 13574 12950 13626
rect 13002 13574 13014 13626
rect 13066 13574 13078 13626
rect 13130 13574 13142 13626
rect 13194 13574 13206 13626
rect 13258 13574 22950 13626
rect 23002 13574 23014 13626
rect 23066 13574 23078 13626
rect 23130 13574 23142 13626
rect 23194 13574 23206 13626
rect 23258 13574 25852 13626
rect 1104 13552 25852 13574
rect 7009 13515 7067 13521
rect 7009 13481 7021 13515
rect 7055 13512 7067 13515
rect 7374 13512 7380 13524
rect 7055 13484 7380 13512
rect 7055 13481 7067 13484
rect 7009 13475 7067 13481
rect 7374 13472 7380 13484
rect 7432 13472 7438 13524
rect 13906 13472 13912 13524
rect 13964 13512 13970 13524
rect 14182 13512 14188 13524
rect 13964 13484 14188 13512
rect 13964 13472 13970 13484
rect 14182 13472 14188 13484
rect 14240 13472 14246 13524
rect 15010 13472 15016 13524
rect 15068 13512 15074 13524
rect 20530 13512 20536 13524
rect 15068 13484 20536 13512
rect 15068 13472 15074 13484
rect 20530 13472 20536 13484
rect 20588 13472 20594 13524
rect 16393 13447 16451 13453
rect 16393 13413 16405 13447
rect 16439 13444 16451 13447
rect 24762 13444 24768 13456
rect 16439 13416 18920 13444
rect 16439 13413 16451 13416
rect 16393 13407 16451 13413
rect 7006 13336 7012 13388
rect 7064 13376 7070 13388
rect 7561 13379 7619 13385
rect 7561 13376 7573 13379
rect 7064 13348 7573 13376
rect 7064 13336 7070 13348
rect 7561 13345 7573 13348
rect 7607 13345 7619 13379
rect 11698 13376 11704 13388
rect 7561 13339 7619 13345
rect 9784 13348 11704 13376
rect 9214 13268 9220 13320
rect 9272 13308 9278 13320
rect 9784 13317 9812 13348
rect 11698 13336 11704 13348
rect 11756 13376 11762 13388
rect 12805 13379 12863 13385
rect 12805 13376 12817 13379
rect 11756 13348 12817 13376
rect 11756 13336 11762 13348
rect 12805 13345 12817 13348
rect 12851 13376 12863 13379
rect 13538 13376 13544 13388
rect 12851 13348 13544 13376
rect 12851 13345 12863 13348
rect 12805 13339 12863 13345
rect 13538 13336 13544 13348
rect 13596 13336 13602 13388
rect 14185 13379 14243 13385
rect 14185 13345 14197 13379
rect 14231 13376 14243 13379
rect 14918 13376 14924 13388
rect 14231 13348 14924 13376
rect 14231 13345 14243 13348
rect 14185 13339 14243 13345
rect 14918 13336 14924 13348
rect 14976 13336 14982 13388
rect 15378 13336 15384 13388
rect 15436 13376 15442 13388
rect 15749 13379 15807 13385
rect 15749 13376 15761 13379
rect 15436 13348 15761 13376
rect 15436 13336 15442 13348
rect 15749 13345 15761 13348
rect 15795 13345 15807 13379
rect 15749 13339 15807 13345
rect 9769 13311 9827 13317
rect 9769 13308 9781 13311
rect 9272 13280 9781 13308
rect 9272 13268 9278 13280
rect 9769 13277 9781 13280
rect 9815 13277 9827 13311
rect 9769 13271 9827 13277
rect 11330 13268 11336 13320
rect 11388 13308 11394 13320
rect 11977 13311 12035 13317
rect 11977 13308 11989 13311
rect 11388 13280 11989 13308
rect 11388 13268 11394 13280
rect 11977 13277 11989 13280
rect 12023 13308 12035 13311
rect 13173 13311 13231 13317
rect 13173 13308 13185 13311
rect 12023 13280 13185 13308
rect 12023 13277 12035 13280
rect 11977 13271 12035 13277
rect 13173 13277 13185 13280
rect 13219 13277 13231 13311
rect 13173 13271 13231 13277
rect 13725 13311 13783 13317
rect 13725 13277 13737 13311
rect 13771 13308 13783 13311
rect 15286 13308 15292 13320
rect 13771 13280 15292 13308
rect 13771 13277 13783 13280
rect 13725 13271 13783 13277
rect 15286 13268 15292 13280
rect 15344 13268 15350 13320
rect 15764 13308 15792 13339
rect 15838 13336 15844 13388
rect 15896 13376 15902 13388
rect 16945 13379 17003 13385
rect 16945 13376 16957 13379
rect 15896 13348 16957 13376
rect 15896 13336 15902 13348
rect 16945 13345 16957 13348
rect 16991 13345 17003 13379
rect 16945 13339 17003 13345
rect 16390 13308 16396 13320
rect 15764 13280 16396 13308
rect 16390 13268 16396 13280
rect 16448 13268 16454 13320
rect 16574 13268 16580 13320
rect 16632 13308 16638 13320
rect 16761 13311 16819 13317
rect 16761 13308 16773 13311
rect 16632 13280 16773 13308
rect 16632 13268 16638 13280
rect 16761 13277 16773 13280
rect 16807 13277 16819 13311
rect 16761 13271 16819 13277
rect 17586 13268 17592 13320
rect 17644 13308 17650 13320
rect 17770 13308 17776 13320
rect 17644 13280 17776 13308
rect 17644 13268 17650 13280
rect 17770 13268 17776 13280
rect 17828 13268 17834 13320
rect 18322 13268 18328 13320
rect 18380 13268 18386 13320
rect 18892 13317 18920 13416
rect 20732 13416 24768 13444
rect 19242 13336 19248 13388
rect 19300 13376 19306 13388
rect 20732 13385 20760 13416
rect 24762 13404 24768 13416
rect 24820 13404 24826 13456
rect 20717 13379 20775 13385
rect 19300 13348 20668 13376
rect 19300 13336 19306 13348
rect 18877 13311 18935 13317
rect 18877 13277 18889 13311
rect 18923 13277 18935 13311
rect 18877 13271 18935 13277
rect 6178 13200 6184 13252
rect 6236 13240 6242 13252
rect 7469 13243 7527 13249
rect 7469 13240 7481 13243
rect 6236 13212 7481 13240
rect 6236 13200 6242 13212
rect 7469 13209 7481 13212
rect 7515 13209 7527 13243
rect 7469 13203 7527 13209
rect 8754 13200 8760 13252
rect 8812 13240 8818 13252
rect 10045 13243 10103 13249
rect 8812 13212 9674 13240
rect 8812 13200 8818 13212
rect 7374 13132 7380 13184
rect 7432 13132 7438 13184
rect 9122 13132 9128 13184
rect 9180 13132 9186 13184
rect 9646 13172 9674 13212
rect 10045 13209 10057 13243
rect 10091 13240 10103 13243
rect 10318 13240 10324 13252
rect 10091 13212 10324 13240
rect 10091 13209 10103 13212
rect 10045 13203 10103 13209
rect 10318 13200 10324 13212
rect 10376 13200 10382 13252
rect 10502 13240 10508 13252
rect 10428 13212 10508 13240
rect 10428 13172 10456 13212
rect 10502 13200 10508 13212
rect 10560 13200 10566 13252
rect 14553 13243 14611 13249
rect 14553 13209 14565 13243
rect 14599 13240 14611 13243
rect 17494 13240 17500 13252
rect 14599 13212 17500 13240
rect 14599 13209 14611 13212
rect 14553 13203 14611 13209
rect 17494 13200 17500 13212
rect 17552 13200 17558 13252
rect 18340 13240 18368 13268
rect 18340 13212 18736 13240
rect 9646 13144 10456 13172
rect 11054 13132 11060 13184
rect 11112 13172 11118 13184
rect 11517 13175 11575 13181
rect 11517 13172 11529 13175
rect 11112 13144 11529 13172
rect 11112 13132 11118 13144
rect 11517 13141 11529 13144
rect 11563 13141 11575 13175
rect 11517 13135 11575 13141
rect 13446 13132 13452 13184
rect 13504 13172 13510 13184
rect 13541 13175 13599 13181
rect 13541 13172 13553 13175
rect 13504 13144 13553 13172
rect 13504 13132 13510 13144
rect 13541 13141 13553 13144
rect 13587 13141 13599 13175
rect 13541 13135 13599 13141
rect 15197 13175 15255 13181
rect 15197 13141 15209 13175
rect 15243 13172 15255 13175
rect 15378 13172 15384 13184
rect 15243 13144 15384 13172
rect 15243 13141 15255 13144
rect 15197 13135 15255 13141
rect 15378 13132 15384 13144
rect 15436 13132 15442 13184
rect 15562 13132 15568 13184
rect 15620 13132 15626 13184
rect 15654 13132 15660 13184
rect 15712 13132 15718 13184
rect 15746 13132 15752 13184
rect 15804 13172 15810 13184
rect 16853 13175 16911 13181
rect 16853 13172 16865 13175
rect 15804 13144 16865 13172
rect 15804 13132 15810 13144
rect 16853 13141 16865 13144
rect 16899 13141 16911 13175
rect 16853 13135 16911 13141
rect 18233 13175 18291 13181
rect 18233 13141 18245 13175
rect 18279 13172 18291 13175
rect 18322 13172 18328 13184
rect 18279 13144 18328 13172
rect 18279 13141 18291 13144
rect 18233 13135 18291 13141
rect 18322 13132 18328 13144
rect 18380 13132 18386 13184
rect 18708 13181 18736 13212
rect 19518 13200 19524 13252
rect 19576 13240 19582 13252
rect 19576 13212 19748 13240
rect 19576 13200 19582 13212
rect 18693 13175 18751 13181
rect 18693 13141 18705 13175
rect 18739 13141 18751 13175
rect 18693 13135 18751 13141
rect 19334 13132 19340 13184
rect 19392 13172 19398 13184
rect 19613 13175 19671 13181
rect 19613 13172 19625 13175
rect 19392 13144 19625 13172
rect 19392 13132 19398 13144
rect 19613 13141 19625 13144
rect 19659 13141 19671 13175
rect 19720 13172 19748 13212
rect 20070 13172 20076 13184
rect 19720 13144 20076 13172
rect 19613 13135 19671 13141
rect 20070 13132 20076 13144
rect 20128 13132 20134 13184
rect 20162 13132 20168 13184
rect 20220 13132 20226 13184
rect 20530 13132 20536 13184
rect 20588 13132 20594 13184
rect 20640 13181 20668 13348
rect 20717 13345 20729 13379
rect 20763 13345 20775 13379
rect 20717 13339 20775 13345
rect 22097 13379 22155 13385
rect 22097 13345 22109 13379
rect 22143 13376 22155 13379
rect 24026 13376 24032 13388
rect 22143 13348 24032 13376
rect 22143 13345 22155 13348
rect 22097 13339 22155 13345
rect 24026 13336 24032 13348
rect 24084 13376 24090 13388
rect 24084 13348 24624 13376
rect 24084 13336 24090 13348
rect 20898 13268 20904 13320
rect 20956 13308 20962 13320
rect 22833 13311 22891 13317
rect 20956 13280 21956 13308
rect 20956 13268 20962 13280
rect 20714 13200 20720 13252
rect 20772 13240 20778 13252
rect 21928 13249 21956 13280
rect 22833 13277 22845 13311
rect 22879 13308 22891 13311
rect 23750 13308 23756 13320
rect 22879 13280 23756 13308
rect 22879 13277 22891 13280
rect 22833 13271 22891 13277
rect 23750 13268 23756 13280
rect 23808 13268 23814 13320
rect 24596 13317 24624 13348
rect 24581 13311 24639 13317
rect 24581 13277 24593 13311
rect 24627 13277 24639 13311
rect 24581 13271 24639 13277
rect 21821 13243 21879 13249
rect 21821 13240 21833 13243
rect 20772 13212 21833 13240
rect 20772 13200 20778 13212
rect 21821 13209 21833 13212
rect 21867 13209 21879 13243
rect 21821 13203 21879 13209
rect 21913 13243 21971 13249
rect 21913 13209 21925 13243
rect 21959 13209 21971 13243
rect 21913 13203 21971 13209
rect 23845 13243 23903 13249
rect 23845 13209 23857 13243
rect 23891 13240 23903 13243
rect 24946 13240 24952 13252
rect 23891 13212 24952 13240
rect 23891 13209 23903 13212
rect 23845 13203 23903 13209
rect 24946 13200 24952 13212
rect 25004 13200 25010 13252
rect 20625 13175 20683 13181
rect 20625 13141 20637 13175
rect 20671 13172 20683 13175
rect 20990 13172 20996 13184
rect 20671 13144 20996 13172
rect 20671 13141 20683 13144
rect 20625 13135 20683 13141
rect 20990 13132 20996 13144
rect 21048 13132 21054 13184
rect 21453 13175 21511 13181
rect 21453 13141 21465 13175
rect 21499 13172 21511 13175
rect 21726 13172 21732 13184
rect 21499 13144 21732 13172
rect 21499 13141 21511 13144
rect 21453 13135 21511 13141
rect 21726 13132 21732 13144
rect 21784 13132 21790 13184
rect 23290 13132 23296 13184
rect 23348 13172 23354 13184
rect 25225 13175 25283 13181
rect 25225 13172 25237 13175
rect 23348 13144 25237 13172
rect 23348 13132 23354 13144
rect 25225 13141 25237 13144
rect 25271 13141 25283 13175
rect 25225 13135 25283 13141
rect 1104 13082 25852 13104
rect 1104 13030 7950 13082
rect 8002 13030 8014 13082
rect 8066 13030 8078 13082
rect 8130 13030 8142 13082
rect 8194 13030 8206 13082
rect 8258 13030 17950 13082
rect 18002 13030 18014 13082
rect 18066 13030 18078 13082
rect 18130 13030 18142 13082
rect 18194 13030 18206 13082
rect 18258 13030 25852 13082
rect 1104 13008 25852 13030
rect 6549 12971 6607 12977
rect 6549 12937 6561 12971
rect 6595 12968 6607 12971
rect 7374 12968 7380 12980
rect 6595 12940 7380 12968
rect 6595 12937 6607 12940
rect 6549 12931 6607 12937
rect 7374 12928 7380 12940
rect 7432 12928 7438 12980
rect 8386 12928 8392 12980
rect 8444 12968 8450 12980
rect 10321 12971 10379 12977
rect 10321 12968 10333 12971
rect 8444 12940 10333 12968
rect 8444 12928 8450 12940
rect 10321 12937 10333 12940
rect 10367 12937 10379 12971
rect 13998 12968 14004 12980
rect 10321 12931 10379 12937
rect 10428 12940 14004 12968
rect 8754 12900 8760 12912
rect 8694 12872 8760 12900
rect 8754 12860 8760 12872
rect 8812 12900 8818 12912
rect 9217 12903 9275 12909
rect 9217 12900 9229 12903
rect 8812 12872 9229 12900
rect 8812 12860 8818 12872
rect 9217 12869 9229 12872
rect 9263 12869 9275 12903
rect 10428 12900 10456 12940
rect 13998 12928 14004 12940
rect 14056 12928 14062 12980
rect 14093 12971 14151 12977
rect 14093 12937 14105 12971
rect 14139 12968 14151 12971
rect 15746 12968 15752 12980
rect 14139 12940 15752 12968
rect 14139 12937 14151 12940
rect 14093 12931 14151 12937
rect 15746 12928 15752 12940
rect 15804 12928 15810 12980
rect 16117 12971 16175 12977
rect 16117 12937 16129 12971
rect 16163 12968 16175 12971
rect 20898 12968 20904 12980
rect 16163 12940 18184 12968
rect 16163 12937 16175 12940
rect 16117 12931 16175 12937
rect 9217 12863 9275 12869
rect 9324 12872 10456 12900
rect 10689 12903 10747 12909
rect 7098 12792 7104 12844
rect 7156 12832 7162 12844
rect 7193 12835 7251 12841
rect 7193 12832 7205 12835
rect 7156 12804 7205 12832
rect 7156 12792 7162 12804
rect 7193 12801 7205 12804
rect 7239 12801 7251 12835
rect 7193 12795 7251 12801
rect 7469 12767 7527 12773
rect 7469 12733 7481 12767
rect 7515 12764 7527 12767
rect 9324 12764 9352 12872
rect 10689 12869 10701 12903
rect 10735 12900 10747 12903
rect 12618 12900 12624 12912
rect 10735 12872 12624 12900
rect 10735 12869 10747 12872
rect 10689 12863 10747 12869
rect 12618 12860 12624 12872
rect 12676 12860 12682 12912
rect 15102 12900 15108 12912
rect 12912 12872 15108 12900
rect 9398 12792 9404 12844
rect 9456 12832 9462 12844
rect 10781 12835 10839 12841
rect 9456 12804 10548 12832
rect 9456 12792 9462 12804
rect 7515 12736 8616 12764
rect 7515 12733 7527 12736
rect 7469 12727 7527 12733
rect 8588 12708 8616 12736
rect 8680 12736 9352 12764
rect 10520 12764 10548 12804
rect 10781 12801 10793 12835
rect 10827 12832 10839 12835
rect 11974 12832 11980 12844
rect 10827 12804 11980 12832
rect 10827 12801 10839 12804
rect 10781 12795 10839 12801
rect 11974 12792 11980 12804
rect 12032 12792 12038 12844
rect 12161 12835 12219 12841
rect 12161 12801 12173 12835
rect 12207 12832 12219 12835
rect 12912 12832 12940 12872
rect 15102 12860 15108 12872
rect 15160 12860 15166 12912
rect 16206 12900 16212 12912
rect 15672 12872 16212 12900
rect 12207 12804 12940 12832
rect 12207 12801 12219 12804
rect 12161 12795 12219 12801
rect 12986 12792 12992 12844
rect 13044 12792 13050 12844
rect 13081 12835 13139 12841
rect 13081 12801 13093 12835
rect 13127 12832 13139 12835
rect 13354 12832 13360 12844
rect 13127 12804 13360 12832
rect 13127 12801 13139 12804
rect 13081 12795 13139 12801
rect 13354 12792 13360 12804
rect 13412 12792 13418 12844
rect 14274 12792 14280 12844
rect 14332 12832 14338 12844
rect 15672 12841 15700 12872
rect 16206 12860 16212 12872
rect 16264 12860 16270 12912
rect 18156 12900 18184 12940
rect 19996 12940 20904 12968
rect 19996 12909 20024 12940
rect 20898 12928 20904 12940
rect 20956 12928 20962 12980
rect 20990 12928 20996 12980
rect 21048 12968 21054 12980
rect 22465 12971 22523 12977
rect 22465 12968 22477 12971
rect 21048 12940 22477 12968
rect 21048 12928 21054 12940
rect 22465 12937 22477 12940
rect 22511 12937 22523 12971
rect 22465 12931 22523 12937
rect 24762 12928 24768 12980
rect 24820 12928 24826 12980
rect 19981 12903 20039 12909
rect 18156 12872 19196 12900
rect 14461 12835 14519 12841
rect 14461 12832 14473 12835
rect 14332 12804 14473 12832
rect 14332 12792 14338 12804
rect 14461 12801 14473 12804
rect 14507 12801 14519 12835
rect 14461 12795 14519 12801
rect 14553 12835 14611 12841
rect 14553 12801 14565 12835
rect 14599 12832 14611 12835
rect 15657 12835 15715 12841
rect 14599 12804 15516 12832
rect 14599 12801 14611 12804
rect 14553 12795 14611 12801
rect 10873 12767 10931 12773
rect 10873 12764 10885 12767
rect 10520 12736 10885 12764
rect 8570 12656 8576 12708
rect 8628 12656 8634 12708
rect 7650 12588 7656 12640
rect 7708 12628 7714 12640
rect 8680 12628 8708 12736
rect 10873 12733 10885 12736
rect 10919 12733 10931 12767
rect 10873 12727 10931 12733
rect 11606 12724 11612 12776
rect 11664 12764 11670 12776
rect 13173 12767 13231 12773
rect 13173 12764 13185 12767
rect 11664 12736 13185 12764
rect 11664 12724 11670 12736
rect 13173 12733 13185 12736
rect 13219 12764 13231 12767
rect 14366 12764 14372 12776
rect 13219 12736 14372 12764
rect 13219 12733 13231 12736
rect 13173 12727 13231 12733
rect 14366 12724 14372 12736
rect 14424 12724 14430 12776
rect 14737 12767 14795 12773
rect 14737 12733 14749 12767
rect 14783 12764 14795 12767
rect 15102 12764 15108 12776
rect 14783 12736 15108 12764
rect 14783 12733 14795 12736
rect 14737 12727 14795 12733
rect 15102 12724 15108 12736
rect 15160 12724 15166 12776
rect 8941 12699 8999 12705
rect 8941 12665 8953 12699
rect 8987 12696 8999 12699
rect 9398 12696 9404 12708
rect 8987 12668 9404 12696
rect 8987 12665 8999 12668
rect 8941 12659 8999 12665
rect 9398 12656 9404 12668
rect 9456 12656 9462 12708
rect 9674 12656 9680 12708
rect 9732 12696 9738 12708
rect 12621 12699 12679 12705
rect 12621 12696 12633 12699
rect 9732 12668 12633 12696
rect 9732 12656 9738 12668
rect 12621 12665 12633 12668
rect 12667 12665 12679 12699
rect 12621 12659 12679 12665
rect 13998 12656 14004 12708
rect 14056 12696 14062 12708
rect 15197 12699 15255 12705
rect 15197 12696 15209 12699
rect 14056 12668 15209 12696
rect 14056 12656 14062 12668
rect 15197 12665 15209 12668
rect 15243 12696 15255 12699
rect 15286 12696 15292 12708
rect 15243 12668 15292 12696
rect 15243 12665 15255 12668
rect 15197 12659 15255 12665
rect 15286 12656 15292 12668
rect 15344 12656 15350 12708
rect 15488 12696 15516 12804
rect 15657 12801 15669 12835
rect 15703 12801 15715 12835
rect 15657 12795 15715 12801
rect 15746 12792 15752 12844
rect 15804 12832 15810 12844
rect 16301 12835 16359 12841
rect 16301 12832 16313 12835
rect 15804 12804 16313 12832
rect 15804 12792 15810 12804
rect 16301 12801 16313 12804
rect 16347 12801 16359 12835
rect 16301 12795 16359 12801
rect 16761 12835 16819 12841
rect 16761 12801 16773 12835
rect 16807 12832 16819 12835
rect 16942 12832 16948 12844
rect 16807 12804 16948 12832
rect 16807 12801 16819 12804
rect 16761 12795 16819 12801
rect 15562 12724 15568 12776
rect 15620 12764 15626 12776
rect 15930 12764 15936 12776
rect 15620 12736 15936 12764
rect 15620 12724 15626 12736
rect 15930 12724 15936 12736
rect 15988 12724 15994 12776
rect 16776 12696 16804 12795
rect 16942 12792 16948 12804
rect 17000 12792 17006 12844
rect 17221 12835 17279 12841
rect 17221 12801 17233 12835
rect 17267 12832 17279 12835
rect 18414 12832 18420 12844
rect 17267 12804 18420 12832
rect 17267 12801 17279 12804
rect 17221 12795 17279 12801
rect 18414 12792 18420 12804
rect 18472 12792 18478 12844
rect 19058 12792 19064 12844
rect 19116 12792 19122 12844
rect 19168 12832 19196 12872
rect 19981 12869 19993 12903
rect 20027 12869 20039 12903
rect 19981 12863 20039 12869
rect 20070 12860 20076 12912
rect 20128 12900 20134 12912
rect 20441 12903 20499 12909
rect 20441 12900 20453 12903
rect 20128 12872 20453 12900
rect 20128 12860 20134 12872
rect 20441 12869 20453 12872
rect 20487 12869 20499 12903
rect 20441 12863 20499 12869
rect 20530 12860 20536 12912
rect 20588 12900 20594 12912
rect 20625 12903 20683 12909
rect 20625 12900 20637 12903
rect 20588 12872 20637 12900
rect 20588 12860 20594 12872
rect 20625 12869 20637 12872
rect 20671 12869 20683 12903
rect 20625 12863 20683 12869
rect 21450 12860 21456 12912
rect 21508 12860 21514 12912
rect 22370 12900 22376 12912
rect 22204 12872 22376 12900
rect 20346 12832 20352 12844
rect 19168 12804 20352 12832
rect 20346 12792 20352 12804
rect 20404 12792 20410 12844
rect 21269 12835 21327 12841
rect 21269 12801 21281 12835
rect 21315 12832 21327 12835
rect 21542 12832 21548 12844
rect 21315 12804 21548 12832
rect 21315 12801 21327 12804
rect 21269 12795 21327 12801
rect 21542 12792 21548 12804
rect 21600 12792 21606 12844
rect 22204 12841 22232 12872
rect 22370 12860 22376 12872
rect 22428 12860 22434 12912
rect 23290 12860 23296 12912
rect 23348 12860 23354 12912
rect 25130 12900 25136 12912
rect 24518 12872 25136 12900
rect 25130 12860 25136 12872
rect 25188 12860 25194 12912
rect 22189 12835 22247 12841
rect 22189 12801 22201 12835
rect 22235 12801 22247 12835
rect 22189 12795 22247 12801
rect 22278 12792 22284 12844
rect 22336 12832 22342 12844
rect 22830 12832 22836 12844
rect 22336 12804 22836 12832
rect 22336 12792 22342 12804
rect 22830 12792 22836 12804
rect 22888 12832 22894 12844
rect 23017 12835 23075 12841
rect 23017 12832 23029 12835
rect 22888 12804 23029 12832
rect 22888 12792 22894 12804
rect 23017 12801 23029 12804
rect 23063 12801 23075 12835
rect 23017 12795 23075 12801
rect 17862 12724 17868 12776
rect 17920 12764 17926 12776
rect 17957 12767 18015 12773
rect 17957 12764 17969 12767
rect 17920 12736 17969 12764
rect 17920 12724 17926 12736
rect 17957 12733 17969 12736
rect 18003 12733 18015 12767
rect 17957 12727 18015 12733
rect 18506 12724 18512 12776
rect 18564 12764 18570 12776
rect 19153 12767 19211 12773
rect 19153 12764 19165 12767
rect 18564 12736 19165 12764
rect 18564 12724 18570 12736
rect 19153 12733 19165 12736
rect 19199 12733 19211 12767
rect 19153 12727 19211 12733
rect 19242 12724 19248 12776
rect 19300 12724 19306 12776
rect 19352 12736 22048 12764
rect 19352 12696 19380 12736
rect 21082 12696 21088 12708
rect 15488 12668 16804 12696
rect 18064 12668 19380 12696
rect 19904 12668 21088 12696
rect 7708 12600 8708 12628
rect 7708 12588 7714 12600
rect 11606 12588 11612 12640
rect 11664 12588 11670 12640
rect 11977 12631 12035 12637
rect 11977 12597 11989 12631
rect 12023 12628 12035 12631
rect 12342 12628 12348 12640
rect 12023 12600 12348 12628
rect 12023 12597 12035 12600
rect 11977 12591 12035 12597
rect 12342 12588 12348 12600
rect 12400 12588 12406 12640
rect 12986 12588 12992 12640
rect 13044 12628 13050 12640
rect 13722 12628 13728 12640
rect 13044 12600 13728 12628
rect 13044 12588 13050 12600
rect 13722 12588 13728 12600
rect 13780 12588 13786 12640
rect 15473 12631 15531 12637
rect 15473 12597 15485 12631
rect 15519 12628 15531 12631
rect 15838 12628 15844 12640
rect 15519 12600 15844 12628
rect 15519 12597 15531 12600
rect 15473 12591 15531 12597
rect 15838 12588 15844 12600
rect 15896 12588 15902 12640
rect 15930 12588 15936 12640
rect 15988 12628 15994 12640
rect 16945 12631 17003 12637
rect 16945 12628 16957 12631
rect 15988 12600 16957 12628
rect 15988 12588 15994 12600
rect 16945 12597 16957 12600
rect 16991 12628 17003 12631
rect 17678 12628 17684 12640
rect 16991 12600 17684 12628
rect 16991 12597 17003 12600
rect 16945 12591 17003 12597
rect 17678 12588 17684 12600
rect 17736 12588 17742 12640
rect 17770 12588 17776 12640
rect 17828 12628 17834 12640
rect 18064 12628 18092 12668
rect 17828 12600 18092 12628
rect 18693 12631 18751 12637
rect 17828 12588 17834 12600
rect 18693 12597 18705 12631
rect 18739 12628 18751 12631
rect 19904 12628 19932 12668
rect 21082 12656 21088 12668
rect 21140 12656 21146 12708
rect 22020 12705 22048 12736
rect 22005 12699 22063 12705
rect 22005 12665 22017 12699
rect 22051 12665 22063 12699
rect 22005 12659 22063 12665
rect 18739 12600 19932 12628
rect 18739 12597 18751 12600
rect 18693 12591 18751 12597
rect 20070 12588 20076 12640
rect 20128 12588 20134 12640
rect 22278 12588 22284 12640
rect 22336 12628 22342 12640
rect 22649 12631 22707 12637
rect 22649 12628 22661 12631
rect 22336 12600 22661 12628
rect 22336 12588 22342 12600
rect 22649 12597 22661 12600
rect 22695 12597 22707 12631
rect 22649 12591 22707 12597
rect 25130 12588 25136 12640
rect 25188 12588 25194 12640
rect 1104 12538 25852 12560
rect 1104 12486 2950 12538
rect 3002 12486 3014 12538
rect 3066 12486 3078 12538
rect 3130 12486 3142 12538
rect 3194 12486 3206 12538
rect 3258 12486 12950 12538
rect 13002 12486 13014 12538
rect 13066 12486 13078 12538
rect 13130 12486 13142 12538
rect 13194 12486 13206 12538
rect 13258 12486 22950 12538
rect 23002 12486 23014 12538
rect 23066 12486 23078 12538
rect 23130 12486 23142 12538
rect 23194 12486 23206 12538
rect 23258 12486 25852 12538
rect 1104 12464 25852 12486
rect 7466 12384 7472 12436
rect 7524 12424 7530 12436
rect 7837 12427 7895 12433
rect 7837 12424 7849 12427
rect 7524 12396 7849 12424
rect 7524 12384 7530 12396
rect 7837 12393 7849 12396
rect 7883 12393 7895 12427
rect 7837 12387 7895 12393
rect 9766 12384 9772 12436
rect 9824 12384 9830 12436
rect 11422 12384 11428 12436
rect 11480 12384 11486 12436
rect 12066 12384 12072 12436
rect 12124 12424 12130 12436
rect 12621 12427 12679 12433
rect 12621 12424 12633 12427
rect 12124 12396 12633 12424
rect 12124 12384 12130 12396
rect 12621 12393 12633 12396
rect 12667 12393 12679 12427
rect 12621 12387 12679 12393
rect 13630 12384 13636 12436
rect 13688 12424 13694 12436
rect 14369 12427 14427 12433
rect 14369 12424 14381 12427
rect 13688 12396 14381 12424
rect 13688 12384 13694 12396
rect 14369 12393 14381 12396
rect 14415 12393 14427 12427
rect 14369 12387 14427 12393
rect 17957 12427 18015 12433
rect 17957 12393 17969 12427
rect 18003 12424 18015 12427
rect 18414 12424 18420 12436
rect 18003 12396 18420 12424
rect 18003 12393 18015 12396
rect 17957 12387 18015 12393
rect 18414 12384 18420 12396
rect 18472 12384 18478 12436
rect 20073 12427 20131 12433
rect 20073 12393 20085 12427
rect 20119 12424 20131 12427
rect 20346 12424 20352 12436
rect 20119 12396 20352 12424
rect 20119 12393 20131 12396
rect 20073 12387 20131 12393
rect 15654 12356 15660 12368
rect 11900 12328 15660 12356
rect 8478 12248 8484 12300
rect 8536 12248 8542 12300
rect 10413 12291 10471 12297
rect 10413 12257 10425 12291
rect 10459 12288 10471 12291
rect 10778 12288 10784 12300
rect 10459 12260 10784 12288
rect 10459 12257 10471 12260
rect 10413 12251 10471 12257
rect 10778 12248 10784 12260
rect 10836 12248 10842 12300
rect 11900 12297 11928 12328
rect 15654 12316 15660 12328
rect 15712 12316 15718 12368
rect 16853 12359 16911 12365
rect 16853 12325 16865 12359
rect 16899 12325 16911 12359
rect 16853 12319 16911 12325
rect 11885 12291 11943 12297
rect 11885 12257 11897 12291
rect 11931 12257 11943 12291
rect 11885 12251 11943 12257
rect 12066 12248 12072 12300
rect 12124 12248 12130 12300
rect 12434 12248 12440 12300
rect 12492 12288 12498 12300
rect 13173 12291 13231 12297
rect 13173 12288 13185 12291
rect 12492 12260 13185 12288
rect 12492 12248 12498 12260
rect 13173 12257 13185 12260
rect 13219 12288 13231 12291
rect 14182 12288 14188 12300
rect 13219 12260 14188 12288
rect 13219 12257 13231 12260
rect 13173 12251 13231 12257
rect 14182 12248 14188 12260
rect 14240 12288 14246 12300
rect 14921 12291 14979 12297
rect 14921 12288 14933 12291
rect 14240 12260 14933 12288
rect 14240 12248 14246 12260
rect 14921 12257 14933 12260
rect 14967 12257 14979 12291
rect 14921 12251 14979 12257
rect 15010 12248 15016 12300
rect 15068 12248 15074 12300
rect 15286 12248 15292 12300
rect 15344 12288 15350 12300
rect 16758 12288 16764 12300
rect 15344 12260 16764 12288
rect 15344 12248 15350 12260
rect 16758 12248 16764 12260
rect 16816 12248 16822 12300
rect 8205 12223 8263 12229
rect 8205 12189 8217 12223
rect 8251 12220 8263 12223
rect 9122 12220 9128 12232
rect 8251 12192 9128 12220
rect 8251 12189 8263 12192
rect 8205 12183 8263 12189
rect 9122 12180 9128 12192
rect 9180 12180 9186 12232
rect 10229 12223 10287 12229
rect 10229 12189 10241 12223
rect 10275 12220 10287 12223
rect 12802 12220 12808 12232
rect 10275 12192 12808 12220
rect 10275 12189 10287 12192
rect 10229 12183 10287 12189
rect 12802 12180 12808 12192
rect 12860 12180 12866 12232
rect 13081 12223 13139 12229
rect 13081 12189 13093 12223
rect 13127 12220 13139 12223
rect 14274 12220 14280 12232
rect 13127 12192 14280 12220
rect 13127 12189 13139 12192
rect 13081 12183 13139 12189
rect 5074 12112 5080 12164
rect 5132 12152 5138 12164
rect 9401 12155 9459 12161
rect 9401 12152 9413 12155
rect 5132 12124 9413 12152
rect 5132 12112 5138 12124
rect 9401 12121 9413 12124
rect 9447 12152 9459 12155
rect 10137 12155 10195 12161
rect 10137 12152 10149 12155
rect 9447 12124 10149 12152
rect 9447 12121 9459 12124
rect 9401 12115 9459 12121
rect 10137 12121 10149 12124
rect 10183 12152 10195 12155
rect 10870 12152 10876 12164
rect 10183 12124 10876 12152
rect 10183 12121 10195 12124
rect 10137 12115 10195 12121
rect 10870 12112 10876 12124
rect 10928 12112 10934 12164
rect 11793 12155 11851 12161
rect 11793 12121 11805 12155
rect 11839 12152 11851 12155
rect 12434 12152 12440 12164
rect 11839 12124 12440 12152
rect 11839 12121 11851 12124
rect 11793 12115 11851 12121
rect 12434 12112 12440 12124
rect 12492 12112 12498 12164
rect 13096 12152 13124 12183
rect 14274 12180 14280 12192
rect 14332 12180 14338 12232
rect 14366 12180 14372 12232
rect 14424 12220 14430 12232
rect 14829 12223 14887 12229
rect 14829 12220 14841 12223
rect 14424 12192 14841 12220
rect 14424 12180 14430 12192
rect 14829 12189 14841 12192
rect 14875 12220 14887 12223
rect 15028 12220 15056 12248
rect 16298 12220 16304 12232
rect 14875 12192 15056 12220
rect 15120 12192 16304 12220
rect 14875 12189 14887 12192
rect 14829 12183 14887 12189
rect 15120 12152 15148 12192
rect 16298 12180 16304 12192
rect 16356 12180 16362 12232
rect 16393 12223 16451 12229
rect 16393 12189 16405 12223
rect 16439 12220 16451 12223
rect 16868 12220 16896 12319
rect 17678 12316 17684 12368
rect 17736 12356 17742 12368
rect 18782 12356 18788 12368
rect 17736 12328 18788 12356
rect 17736 12316 17742 12328
rect 18782 12316 18788 12328
rect 18840 12316 18846 12368
rect 17497 12291 17555 12297
rect 17497 12257 17509 12291
rect 17543 12288 17555 12291
rect 18598 12288 18604 12300
rect 17543 12260 18604 12288
rect 17543 12257 17555 12260
rect 17497 12251 17555 12257
rect 18598 12248 18604 12260
rect 18656 12248 18662 12300
rect 16439 12192 16896 12220
rect 17313 12223 17371 12229
rect 16439 12189 16451 12192
rect 16393 12183 16451 12189
rect 17313 12189 17325 12223
rect 17359 12220 17371 12223
rect 18966 12220 18972 12232
rect 17359 12192 18972 12220
rect 17359 12189 17371 12192
rect 17313 12183 17371 12189
rect 18966 12180 18972 12192
rect 19024 12180 19030 12232
rect 19521 12223 19579 12229
rect 19521 12189 19533 12223
rect 19567 12220 19579 12223
rect 20088 12220 20116 12387
rect 20346 12384 20352 12396
rect 20404 12384 20410 12436
rect 21726 12316 21732 12368
rect 21784 12356 21790 12368
rect 21910 12356 21916 12368
rect 21784 12328 21916 12356
rect 21784 12316 21790 12328
rect 21910 12316 21916 12328
rect 21968 12316 21974 12368
rect 20254 12248 20260 12300
rect 20312 12288 20318 12300
rect 20349 12291 20407 12297
rect 20349 12288 20361 12291
rect 20312 12260 20361 12288
rect 20312 12248 20318 12260
rect 20349 12257 20361 12260
rect 20395 12257 20407 12291
rect 20349 12251 20407 12257
rect 19567 12192 20116 12220
rect 19567 12189 19579 12192
rect 19521 12183 19579 12189
rect 22186 12180 22192 12232
rect 22244 12220 22250 12232
rect 22649 12223 22707 12229
rect 22649 12220 22661 12223
rect 22244 12192 22661 12220
rect 22244 12180 22250 12192
rect 22649 12189 22661 12192
rect 22695 12189 22707 12223
rect 22649 12183 22707 12189
rect 24673 12223 24731 12229
rect 24673 12189 24685 12223
rect 24719 12220 24731 12223
rect 24762 12220 24768 12232
rect 24719 12192 24768 12220
rect 24719 12189 24731 12192
rect 24673 12183 24731 12189
rect 24762 12180 24768 12192
rect 24820 12180 24826 12232
rect 18322 12152 18328 12164
rect 12912 12124 13124 12152
rect 13280 12124 15148 12152
rect 15488 12124 18328 12152
rect 6914 12044 6920 12096
rect 6972 12084 6978 12096
rect 8297 12087 8355 12093
rect 8297 12084 8309 12087
rect 6972 12056 8309 12084
rect 6972 12044 6978 12056
rect 8297 12053 8309 12056
rect 8343 12053 8355 12087
rect 8297 12047 8355 12053
rect 8754 12044 8760 12096
rect 8812 12084 8818 12096
rect 8941 12087 8999 12093
rect 8941 12084 8953 12087
rect 8812 12056 8953 12084
rect 8812 12044 8818 12056
rect 8941 12053 8953 12056
rect 8987 12084 8999 12087
rect 9030 12084 9036 12096
rect 8987 12056 9036 12084
rect 8987 12053 8999 12056
rect 8941 12047 8999 12053
rect 9030 12044 9036 12056
rect 9088 12044 9094 12096
rect 9122 12044 9128 12096
rect 9180 12084 9186 12096
rect 12912 12084 12940 12124
rect 9180 12056 12940 12084
rect 12989 12087 13047 12093
rect 9180 12044 9186 12056
rect 12989 12053 13001 12087
rect 13035 12084 13047 12087
rect 13280 12084 13308 12124
rect 13035 12056 13308 12084
rect 13035 12053 13047 12056
rect 12989 12047 13047 12053
rect 13354 12044 13360 12096
rect 13412 12084 13418 12096
rect 13630 12084 13636 12096
rect 13412 12056 13636 12084
rect 13412 12044 13418 12056
rect 13630 12044 13636 12056
rect 13688 12044 13694 12096
rect 13909 12087 13967 12093
rect 13909 12053 13921 12087
rect 13955 12084 13967 12087
rect 14366 12084 14372 12096
rect 13955 12056 14372 12084
rect 13955 12053 13967 12056
rect 13909 12047 13967 12053
rect 14366 12044 14372 12056
rect 14424 12044 14430 12096
rect 14734 12044 14740 12096
rect 14792 12044 14798 12096
rect 14918 12044 14924 12096
rect 14976 12084 14982 12096
rect 15488 12084 15516 12124
rect 18322 12112 18328 12124
rect 18380 12112 18386 12164
rect 18414 12112 18420 12164
rect 18472 12152 18478 12164
rect 18601 12155 18659 12161
rect 18601 12152 18613 12155
rect 18472 12124 18613 12152
rect 18472 12112 18478 12124
rect 18601 12121 18613 12124
rect 18647 12152 18659 12155
rect 19150 12152 19156 12164
rect 18647 12124 19156 12152
rect 18647 12121 18659 12124
rect 18601 12115 18659 12121
rect 19150 12112 19156 12124
rect 19208 12112 19214 12164
rect 19705 12155 19763 12161
rect 19705 12121 19717 12155
rect 19751 12152 19763 12155
rect 20346 12152 20352 12164
rect 19751 12124 20352 12152
rect 19751 12121 19763 12124
rect 19705 12115 19763 12121
rect 20346 12112 20352 12124
rect 20404 12112 20410 12164
rect 20622 12112 20628 12164
rect 20680 12112 20686 12164
rect 21910 12152 21916 12164
rect 21850 12124 21916 12152
rect 21910 12112 21916 12124
rect 21968 12152 21974 12164
rect 22278 12152 22284 12164
rect 21968 12124 22284 12152
rect 21968 12112 21974 12124
rect 22278 12112 22284 12124
rect 22336 12112 22342 12164
rect 23845 12155 23903 12161
rect 23845 12121 23857 12155
rect 23891 12152 23903 12155
rect 24946 12152 24952 12164
rect 23891 12124 24952 12152
rect 23891 12121 23903 12124
rect 23845 12115 23903 12121
rect 24946 12112 24952 12124
rect 25004 12112 25010 12164
rect 14976 12056 15516 12084
rect 15565 12087 15623 12093
rect 14976 12044 14982 12056
rect 15565 12053 15577 12087
rect 15611 12084 15623 12087
rect 16114 12084 16120 12096
rect 15611 12056 16120 12084
rect 15611 12053 15623 12056
rect 15565 12047 15623 12053
rect 16114 12044 16120 12056
rect 16172 12044 16178 12096
rect 16206 12044 16212 12096
rect 16264 12044 16270 12096
rect 16758 12044 16764 12096
rect 16816 12084 16822 12096
rect 17221 12087 17279 12093
rect 17221 12084 17233 12087
rect 16816 12056 17233 12084
rect 16816 12044 16822 12056
rect 17221 12053 17233 12056
rect 17267 12053 17279 12087
rect 17221 12047 17279 12053
rect 18233 12087 18291 12093
rect 18233 12053 18245 12087
rect 18279 12084 18291 12087
rect 18506 12084 18512 12096
rect 18279 12056 18512 12084
rect 18279 12053 18291 12056
rect 18233 12047 18291 12053
rect 18506 12044 18512 12056
rect 18564 12044 18570 12096
rect 18693 12087 18751 12093
rect 18693 12053 18705 12087
rect 18739 12084 18751 12087
rect 18966 12084 18972 12096
rect 18739 12056 18972 12084
rect 18739 12053 18751 12056
rect 18693 12047 18751 12053
rect 18966 12044 18972 12056
rect 19024 12044 19030 12096
rect 19426 12044 19432 12096
rect 19484 12084 19490 12096
rect 22097 12087 22155 12093
rect 22097 12084 22109 12087
rect 19484 12056 22109 12084
rect 19484 12044 19490 12056
rect 22097 12053 22109 12056
rect 22143 12053 22155 12087
rect 22097 12047 22155 12053
rect 23382 12044 23388 12096
rect 23440 12084 23446 12096
rect 25317 12087 25375 12093
rect 25317 12084 25329 12087
rect 23440 12056 25329 12084
rect 23440 12044 23446 12056
rect 25317 12053 25329 12056
rect 25363 12053 25375 12087
rect 25317 12047 25375 12053
rect 1104 11994 25852 12016
rect 1104 11942 7950 11994
rect 8002 11942 8014 11994
rect 8066 11942 8078 11994
rect 8130 11942 8142 11994
rect 8194 11942 8206 11994
rect 8258 11942 17950 11994
rect 18002 11942 18014 11994
rect 18066 11942 18078 11994
rect 18130 11942 18142 11994
rect 18194 11942 18206 11994
rect 18258 11942 25852 11994
rect 1104 11920 25852 11942
rect 8941 11883 8999 11889
rect 8941 11849 8953 11883
rect 8987 11849 8999 11883
rect 8941 11843 8999 11849
rect 9401 11883 9459 11889
rect 9401 11849 9413 11883
rect 9447 11880 9459 11883
rect 9674 11880 9680 11892
rect 9447 11852 9680 11880
rect 9447 11849 9459 11852
rect 9401 11843 9459 11849
rect 8956 11812 8984 11843
rect 9674 11840 9680 11852
rect 9732 11840 9738 11892
rect 10134 11840 10140 11892
rect 10192 11840 10198 11892
rect 11054 11880 11060 11892
rect 10428 11852 11060 11880
rect 9582 11812 9588 11824
rect 8956 11784 9588 11812
rect 9582 11772 9588 11784
rect 9640 11772 9646 11824
rect 7837 11747 7895 11753
rect 7837 11713 7849 11747
rect 7883 11713 7895 11747
rect 7837 11707 7895 11713
rect 7852 11676 7880 11707
rect 8754 11704 8760 11756
rect 8812 11744 8818 11756
rect 9309 11747 9367 11753
rect 9309 11744 9321 11747
rect 8812 11716 9321 11744
rect 8812 11704 8818 11716
rect 9309 11713 9321 11716
rect 9355 11713 9367 11747
rect 10428 11744 10456 11852
rect 11054 11840 11060 11852
rect 11112 11840 11118 11892
rect 11514 11840 11520 11892
rect 11572 11880 11578 11892
rect 11977 11883 12035 11889
rect 11977 11880 11989 11883
rect 11572 11852 11989 11880
rect 11572 11840 11578 11852
rect 11977 11849 11989 11852
rect 12023 11849 12035 11883
rect 11977 11843 12035 11849
rect 12158 11840 12164 11892
rect 12216 11880 12222 11892
rect 13173 11883 13231 11889
rect 13173 11880 13185 11883
rect 12216 11852 13185 11880
rect 12216 11840 12222 11852
rect 13173 11849 13185 11852
rect 13219 11849 13231 11883
rect 13173 11843 13231 11849
rect 13262 11840 13268 11892
rect 13320 11880 13326 11892
rect 13633 11883 13691 11889
rect 13633 11880 13645 11883
rect 13320 11852 13645 11880
rect 13320 11840 13326 11852
rect 13633 11849 13645 11852
rect 13679 11849 13691 11883
rect 13633 11843 13691 11849
rect 13814 11840 13820 11892
rect 13872 11880 13878 11892
rect 14369 11883 14427 11889
rect 14369 11880 14381 11883
rect 13872 11852 14381 11880
rect 13872 11840 13878 11852
rect 14369 11849 14381 11852
rect 14415 11849 14427 11883
rect 14369 11843 14427 11849
rect 14458 11840 14464 11892
rect 14516 11880 14522 11892
rect 14737 11883 14795 11889
rect 14737 11880 14749 11883
rect 14516 11852 14749 11880
rect 14516 11840 14522 11852
rect 14737 11849 14749 11852
rect 14783 11880 14795 11883
rect 14826 11880 14832 11892
rect 14783 11852 14832 11880
rect 14783 11849 14795 11852
rect 14737 11843 14795 11849
rect 14826 11840 14832 11852
rect 14884 11840 14890 11892
rect 15194 11840 15200 11892
rect 15252 11880 15258 11892
rect 16209 11883 16267 11889
rect 16209 11880 16221 11883
rect 15252 11852 16221 11880
rect 15252 11840 15258 11852
rect 16209 11849 16221 11852
rect 16255 11849 16267 11883
rect 16209 11843 16267 11849
rect 17034 11840 17040 11892
rect 17092 11880 17098 11892
rect 17313 11883 17371 11889
rect 17313 11880 17325 11883
rect 17092 11852 17325 11880
rect 17092 11840 17098 11852
rect 17313 11849 17325 11852
rect 17359 11849 17371 11883
rect 17313 11843 17371 11849
rect 18049 11883 18107 11889
rect 18049 11849 18061 11883
rect 18095 11880 18107 11883
rect 18874 11880 18880 11892
rect 18095 11852 18880 11880
rect 18095 11849 18107 11852
rect 18049 11843 18107 11849
rect 18874 11840 18880 11852
rect 18932 11840 18938 11892
rect 19150 11840 19156 11892
rect 19208 11880 19214 11892
rect 19245 11883 19303 11889
rect 19245 11880 19257 11883
rect 19208 11852 19257 11880
rect 19208 11840 19214 11852
rect 19245 11849 19257 11852
rect 19291 11849 19303 11883
rect 19245 11843 19303 11849
rect 19613 11883 19671 11889
rect 19613 11849 19625 11883
rect 19659 11880 19671 11883
rect 19659 11852 20576 11880
rect 19659 11849 19671 11852
rect 19613 11843 19671 11849
rect 13541 11815 13599 11821
rect 13541 11781 13553 11815
rect 13587 11781 13599 11815
rect 13541 11775 13599 11781
rect 9309 11707 9367 11713
rect 9416 11716 10456 11744
rect 10505 11747 10563 11753
rect 9416 11676 9444 11716
rect 10505 11713 10517 11747
rect 10551 11744 10563 11747
rect 11422 11744 11428 11756
rect 10551 11716 11428 11744
rect 10551 11713 10563 11716
rect 10505 11707 10563 11713
rect 11422 11704 11428 11716
rect 11480 11704 11486 11756
rect 12250 11704 12256 11756
rect 12308 11744 12314 11756
rect 12345 11747 12403 11753
rect 12345 11744 12357 11747
rect 12308 11716 12357 11744
rect 12308 11704 12314 11716
rect 12345 11713 12357 11716
rect 12391 11713 12403 11747
rect 12345 11707 12403 11713
rect 12434 11704 12440 11756
rect 12492 11704 12498 11756
rect 7852 11648 9444 11676
rect 9490 11636 9496 11688
rect 9548 11676 9554 11688
rect 9585 11679 9643 11685
rect 9585 11676 9597 11679
rect 9548 11648 9597 11676
rect 9548 11636 9554 11648
rect 9585 11645 9597 11648
rect 9631 11676 9643 11679
rect 9950 11676 9956 11688
rect 9631 11648 9956 11676
rect 9631 11645 9643 11648
rect 9585 11639 9643 11645
rect 9950 11636 9956 11648
rect 10008 11636 10014 11688
rect 10597 11679 10655 11685
rect 10597 11645 10609 11679
rect 10643 11645 10655 11679
rect 10597 11639 10655 11645
rect 8481 11611 8539 11617
rect 8481 11577 8493 11611
rect 8527 11608 8539 11611
rect 9398 11608 9404 11620
rect 8527 11580 9404 11608
rect 8527 11577 8539 11580
rect 8481 11571 8539 11577
rect 9398 11568 9404 11580
rect 9456 11568 9462 11620
rect 7190 11500 7196 11552
rect 7248 11540 7254 11552
rect 9122 11540 9128 11552
rect 7248 11512 9128 11540
rect 7248 11500 7254 11512
rect 9122 11500 9128 11512
rect 9180 11500 9186 11552
rect 10612 11540 10640 11639
rect 10778 11636 10784 11688
rect 10836 11636 10842 11688
rect 11054 11636 11060 11688
rect 11112 11676 11118 11688
rect 11882 11676 11888 11688
rect 11112 11648 11888 11676
rect 11112 11636 11118 11648
rect 11882 11636 11888 11648
rect 11940 11636 11946 11688
rect 12066 11636 12072 11688
rect 12124 11676 12130 11688
rect 12529 11679 12587 11685
rect 12529 11676 12541 11679
rect 12124 11648 12541 11676
rect 12124 11636 12130 11648
rect 12529 11645 12541 11648
rect 12575 11645 12587 11679
rect 13556 11676 13584 11775
rect 13998 11772 14004 11824
rect 14056 11812 14062 11824
rect 14056 11784 15700 11812
rect 14056 11772 14062 11784
rect 14826 11704 14832 11756
rect 14884 11704 14890 11756
rect 15102 11704 15108 11756
rect 15160 11744 15166 11756
rect 15565 11747 15623 11753
rect 15565 11744 15577 11747
rect 15160 11716 15577 11744
rect 15160 11704 15166 11716
rect 15565 11713 15577 11716
rect 15611 11713 15623 11747
rect 15672 11744 15700 11784
rect 16114 11772 16120 11824
rect 16172 11812 16178 11824
rect 19981 11815 20039 11821
rect 19981 11812 19993 11815
rect 16172 11784 19993 11812
rect 16172 11772 16178 11784
rect 19981 11781 19993 11784
rect 20027 11781 20039 11815
rect 20548 11812 20576 11852
rect 20622 11840 20628 11892
rect 20680 11880 20686 11892
rect 22649 11883 22707 11889
rect 22649 11880 22661 11883
rect 20680 11852 22661 11880
rect 20680 11840 20686 11852
rect 22649 11849 22661 11852
rect 22695 11849 22707 11883
rect 22649 11843 22707 11849
rect 20714 11812 20720 11824
rect 20548 11784 20720 11812
rect 19981 11775 20039 11781
rect 20714 11772 20720 11784
rect 20772 11772 20778 11824
rect 20901 11815 20959 11821
rect 20901 11781 20913 11815
rect 20947 11812 20959 11815
rect 21637 11815 21695 11821
rect 21637 11812 21649 11815
rect 20947 11784 21649 11812
rect 20947 11781 20959 11784
rect 20901 11775 20959 11781
rect 21637 11781 21649 11784
rect 21683 11812 21695 11815
rect 21726 11812 21732 11824
rect 21683 11784 21732 11812
rect 21683 11781 21695 11784
rect 21637 11775 21695 11781
rect 21726 11772 21732 11784
rect 21784 11772 21790 11824
rect 23382 11772 23388 11824
rect 23440 11772 23446 11824
rect 25130 11812 25136 11824
rect 24610 11784 25136 11812
rect 25130 11772 25136 11784
rect 25188 11772 25194 11824
rect 17221 11747 17279 11753
rect 17221 11744 17233 11747
rect 15672 11716 17233 11744
rect 15565 11707 15623 11713
rect 17221 11713 17233 11716
rect 17267 11713 17279 11747
rect 17221 11707 17279 11713
rect 18417 11747 18475 11753
rect 18417 11713 18429 11747
rect 18463 11713 18475 11747
rect 18417 11707 18475 11713
rect 13817 11679 13875 11685
rect 13556 11648 13676 11676
rect 12529 11639 12587 11645
rect 11238 11540 11244 11552
rect 10612 11512 11244 11540
rect 11238 11500 11244 11512
rect 11296 11500 11302 11552
rect 12802 11500 12808 11552
rect 12860 11540 12866 11552
rect 13262 11540 13268 11552
rect 12860 11512 13268 11540
rect 12860 11500 12866 11512
rect 13262 11500 13268 11512
rect 13320 11500 13326 11552
rect 13648 11540 13676 11648
rect 13817 11645 13829 11679
rect 13863 11676 13875 11679
rect 14182 11676 14188 11688
rect 13863 11648 14188 11676
rect 13863 11645 13875 11648
rect 13817 11639 13875 11645
rect 14182 11636 14188 11648
rect 14240 11676 14246 11688
rect 14921 11679 14979 11685
rect 14921 11676 14933 11679
rect 14240 11648 14933 11676
rect 14240 11636 14246 11648
rect 14921 11645 14933 11648
rect 14967 11645 14979 11679
rect 14921 11639 14979 11645
rect 17402 11636 17408 11688
rect 17460 11636 17466 11688
rect 14090 11568 14096 11620
rect 14148 11608 14154 11620
rect 18432 11608 18460 11707
rect 19058 11704 19064 11756
rect 19116 11744 19122 11756
rect 20073 11747 20131 11753
rect 20073 11744 20085 11747
rect 19116 11716 20085 11744
rect 19116 11704 19122 11716
rect 20073 11713 20085 11716
rect 20119 11713 20131 11747
rect 20073 11707 20131 11713
rect 20438 11704 20444 11756
rect 20496 11744 20502 11756
rect 21361 11747 21419 11753
rect 21361 11744 21373 11747
rect 20496 11716 21373 11744
rect 20496 11704 20502 11716
rect 21361 11713 21373 11716
rect 21407 11713 21419 11747
rect 21361 11707 21419 11713
rect 21450 11704 21456 11756
rect 21508 11744 21514 11756
rect 21993 11747 22051 11753
rect 21993 11744 22005 11747
rect 21508 11716 22005 11744
rect 21508 11704 21514 11716
rect 21993 11713 22005 11716
rect 22039 11713 22051 11747
rect 21993 11707 22051 11713
rect 22278 11704 22284 11756
rect 22336 11744 22342 11756
rect 22830 11744 22836 11756
rect 22336 11716 22836 11744
rect 22336 11704 22342 11716
rect 22830 11704 22836 11716
rect 22888 11744 22894 11756
rect 23109 11747 23167 11753
rect 23109 11744 23121 11747
rect 22888 11716 23121 11744
rect 22888 11704 22894 11716
rect 23109 11713 23121 11716
rect 23155 11713 23167 11747
rect 23109 11707 23167 11713
rect 18506 11636 18512 11688
rect 18564 11636 18570 11688
rect 18693 11679 18751 11685
rect 18693 11645 18705 11679
rect 18739 11676 18751 11679
rect 19426 11676 19432 11688
rect 18739 11648 19432 11676
rect 18739 11645 18751 11648
rect 18693 11639 18751 11645
rect 19426 11636 19432 11648
rect 19484 11636 19490 11688
rect 20257 11679 20315 11685
rect 20257 11645 20269 11679
rect 20303 11676 20315 11679
rect 20806 11676 20812 11688
rect 20303 11648 20812 11676
rect 20303 11645 20315 11648
rect 20257 11639 20315 11645
rect 20806 11636 20812 11648
rect 20864 11636 20870 11688
rect 14148 11580 18460 11608
rect 18524 11608 18552 11636
rect 19061 11611 19119 11617
rect 19061 11608 19073 11611
rect 18524 11580 19073 11608
rect 14148 11568 14154 11580
rect 19061 11577 19073 11580
rect 19107 11577 19119 11611
rect 19061 11571 19119 11577
rect 19150 11568 19156 11620
rect 19208 11608 19214 11620
rect 19702 11608 19708 11620
rect 19208 11580 19708 11608
rect 19208 11568 19214 11580
rect 19702 11568 19708 11580
rect 19760 11568 19766 11620
rect 14182 11540 14188 11552
rect 13648 11512 14188 11540
rect 14182 11500 14188 11512
rect 14240 11540 14246 11552
rect 15286 11540 15292 11552
rect 14240 11512 15292 11540
rect 14240 11500 14246 11512
rect 15286 11500 15292 11512
rect 15344 11500 15350 11552
rect 16853 11543 16911 11549
rect 16853 11509 16865 11543
rect 16899 11540 16911 11543
rect 18598 11540 18604 11552
rect 16899 11512 18604 11540
rect 16899 11509 16911 11512
rect 16853 11503 16911 11509
rect 18598 11500 18604 11512
rect 18656 11500 18662 11552
rect 20714 11500 20720 11552
rect 20772 11540 20778 11552
rect 20993 11543 21051 11549
rect 20993 11540 21005 11543
rect 20772 11512 21005 11540
rect 20772 11500 20778 11512
rect 20993 11509 21005 11512
rect 21039 11509 21051 11543
rect 20993 11503 21051 11509
rect 24578 11500 24584 11552
rect 24636 11540 24642 11552
rect 24857 11543 24915 11549
rect 24857 11540 24869 11543
rect 24636 11512 24869 11540
rect 24636 11500 24642 11512
rect 24857 11509 24869 11512
rect 24903 11509 24915 11543
rect 24857 11503 24915 11509
rect 25130 11500 25136 11552
rect 25188 11500 25194 11552
rect 1104 11450 25852 11472
rect 1104 11398 2950 11450
rect 3002 11398 3014 11450
rect 3066 11398 3078 11450
rect 3130 11398 3142 11450
rect 3194 11398 3206 11450
rect 3258 11398 12950 11450
rect 13002 11398 13014 11450
rect 13066 11398 13078 11450
rect 13130 11398 13142 11450
rect 13194 11398 13206 11450
rect 13258 11398 22950 11450
rect 23002 11398 23014 11450
rect 23066 11398 23078 11450
rect 23130 11398 23142 11450
rect 23194 11398 23206 11450
rect 23258 11398 25852 11450
rect 1104 11376 25852 11398
rect 8570 11296 8576 11348
rect 8628 11296 8634 11348
rect 10778 11296 10784 11348
rect 10836 11336 10842 11348
rect 10836 11308 12434 11336
rect 10836 11296 10842 11308
rect 10336 11240 11376 11268
rect 9125 11203 9183 11209
rect 9125 11169 9137 11203
rect 9171 11200 9183 11203
rect 9490 11200 9496 11212
rect 9171 11172 9496 11200
rect 9171 11169 9183 11172
rect 9125 11163 9183 11169
rect 9490 11160 9496 11172
rect 9548 11160 9554 11212
rect 10042 11160 10048 11212
rect 10100 11200 10106 11212
rect 10336 11209 10364 11240
rect 10321 11203 10379 11209
rect 10321 11200 10333 11203
rect 10100 11172 10333 11200
rect 10100 11160 10106 11172
rect 10321 11169 10333 11172
rect 10367 11169 10379 11203
rect 10321 11163 10379 11169
rect 7929 11135 7987 11141
rect 7929 11101 7941 11135
rect 7975 11101 7987 11135
rect 7929 11095 7987 11101
rect 9401 11135 9459 11141
rect 9401 11101 9413 11135
rect 9447 11132 9459 11135
rect 10870 11132 10876 11144
rect 9447 11104 10876 11132
rect 9447 11101 9459 11104
rect 9401 11095 9459 11101
rect 7944 11064 7972 11095
rect 10870 11092 10876 11104
rect 10928 11092 10934 11144
rect 11348 11132 11376 11240
rect 11790 11160 11796 11212
rect 11848 11160 11854 11212
rect 11882 11160 11888 11212
rect 11940 11160 11946 11212
rect 12406 11200 12434 11308
rect 12618 11296 12624 11348
rect 12676 11296 12682 11348
rect 12986 11296 12992 11348
rect 13044 11336 13050 11348
rect 15378 11336 15384 11348
rect 13044 11308 15384 11336
rect 13044 11296 13050 11308
rect 15378 11296 15384 11308
rect 15436 11296 15442 11348
rect 16393 11339 16451 11345
rect 16393 11305 16405 11339
rect 16439 11336 16451 11339
rect 17218 11336 17224 11348
rect 16439 11308 17224 11336
rect 16439 11305 16451 11308
rect 16393 11299 16451 11305
rect 17218 11296 17224 11308
rect 17276 11336 17282 11348
rect 17402 11336 17408 11348
rect 17276 11308 17408 11336
rect 17276 11296 17282 11308
rect 17402 11296 17408 11308
rect 17460 11296 17466 11348
rect 17773 11339 17831 11345
rect 17773 11305 17785 11339
rect 17819 11336 17831 11339
rect 18322 11336 18328 11348
rect 17819 11308 18328 11336
rect 17819 11305 17831 11308
rect 17773 11299 17831 11305
rect 18322 11296 18328 11308
rect 18380 11296 18386 11348
rect 18414 11296 18420 11348
rect 18472 11336 18478 11348
rect 18690 11336 18696 11348
rect 18472 11308 18696 11336
rect 18472 11296 18478 11308
rect 18690 11296 18696 11308
rect 18748 11336 18754 11348
rect 18785 11339 18843 11345
rect 18785 11336 18797 11339
rect 18748 11308 18797 11336
rect 18748 11296 18754 11308
rect 18785 11305 18797 11308
rect 18831 11305 18843 11339
rect 18785 11299 18843 11305
rect 19058 11296 19064 11348
rect 19116 11296 19122 11348
rect 19426 11296 19432 11348
rect 19484 11336 19490 11348
rect 19613 11339 19671 11345
rect 19613 11336 19625 11339
rect 19484 11308 19625 11336
rect 19484 11296 19490 11308
rect 19613 11305 19625 11308
rect 19659 11305 19671 11339
rect 19613 11299 19671 11305
rect 21542 11296 21548 11348
rect 21600 11296 21606 11348
rect 12894 11228 12900 11280
rect 12952 11268 12958 11280
rect 13633 11271 13691 11277
rect 13633 11268 13645 11271
rect 12952 11240 13645 11268
rect 12952 11228 12958 11240
rect 13633 11237 13645 11240
rect 13679 11237 13691 11271
rect 13633 11231 13691 11237
rect 13265 11203 13323 11209
rect 13265 11200 13277 11203
rect 12406 11172 13277 11200
rect 13265 11169 13277 11172
rect 13311 11200 13323 11203
rect 13446 11200 13452 11212
rect 13311 11172 13452 11200
rect 13311 11169 13323 11172
rect 13265 11163 13323 11169
rect 13446 11160 13452 11172
rect 13504 11160 13510 11212
rect 13648 11200 13676 11231
rect 13814 11228 13820 11280
rect 13872 11268 13878 11280
rect 13909 11271 13967 11277
rect 13909 11268 13921 11271
rect 13872 11240 13921 11268
rect 13872 11228 13878 11240
rect 13909 11237 13921 11240
rect 13955 11268 13967 11271
rect 14550 11268 14556 11280
rect 13955 11240 14556 11268
rect 13955 11237 13967 11240
rect 13909 11231 13967 11237
rect 14550 11228 14556 11240
rect 14608 11228 14614 11280
rect 16868 11240 17540 11268
rect 14366 11200 14372 11212
rect 13648 11172 14372 11200
rect 14366 11160 14372 11172
rect 14424 11160 14430 11212
rect 14645 11203 14703 11209
rect 14645 11169 14657 11203
rect 14691 11200 14703 11203
rect 15010 11200 15016 11212
rect 14691 11172 15016 11200
rect 14691 11169 14703 11172
rect 14645 11163 14703 11169
rect 15010 11160 15016 11172
rect 15068 11200 15074 11212
rect 16868 11200 16896 11240
rect 15068 11172 16896 11200
rect 15068 11160 15074 11172
rect 11701 11135 11759 11141
rect 11701 11132 11713 11135
rect 11348 11104 11713 11132
rect 11701 11101 11713 11104
rect 11747 11132 11759 11135
rect 13630 11132 13636 11144
rect 11747 11104 13636 11132
rect 11747 11101 11759 11104
rect 11701 11095 11759 11101
rect 13630 11092 13636 11104
rect 13688 11092 13694 11144
rect 14182 11092 14188 11144
rect 14240 11092 14246 11144
rect 17037 11135 17095 11141
rect 17037 11101 17049 11135
rect 17083 11101 17095 11135
rect 17037 11095 17095 11101
rect 10778 11064 10784 11076
rect 7944 11036 10784 11064
rect 10778 11024 10784 11036
rect 10836 11024 10842 11076
rect 11256 11036 12572 11064
rect 10689 10999 10747 11005
rect 10689 10965 10701 10999
rect 10735 10996 10747 10999
rect 11256 10996 11284 11036
rect 10735 10968 11284 10996
rect 10735 10965 10747 10968
rect 10689 10959 10747 10965
rect 11330 10956 11336 11008
rect 11388 10956 11394 11008
rect 12544 10996 12572 11036
rect 12618 11024 12624 11076
rect 12676 11064 12682 11076
rect 12894 11064 12900 11076
rect 12676 11036 12900 11064
rect 12676 11024 12682 11036
rect 12894 11024 12900 11036
rect 12952 11024 12958 11076
rect 12986 11024 12992 11076
rect 13044 11024 13050 11076
rect 13081 11067 13139 11073
rect 13081 11033 13093 11067
rect 13127 11064 13139 11067
rect 14274 11064 14280 11076
rect 13127 11036 14280 11064
rect 13127 11033 13139 11036
rect 13081 11027 13139 11033
rect 14274 11024 14280 11036
rect 14332 11024 14338 11076
rect 14369 11067 14427 11073
rect 14369 11033 14381 11067
rect 14415 11064 14427 11067
rect 14458 11064 14464 11076
rect 14415 11036 14464 11064
rect 14415 11033 14427 11036
rect 14369 11027 14427 11033
rect 14458 11024 14464 11036
rect 14516 11024 14522 11076
rect 14918 11024 14924 11076
rect 14976 11024 14982 11076
rect 16482 11064 16488 11076
rect 16146 11036 16488 11064
rect 16482 11024 16488 11036
rect 16540 11024 16546 11076
rect 14090 10996 14096 11008
rect 12544 10968 14096 10996
rect 14090 10956 14096 10968
rect 14148 10956 14154 11008
rect 16666 10956 16672 11008
rect 16724 10996 16730 11008
rect 16853 10999 16911 11005
rect 16853 10996 16865 10999
rect 16724 10968 16865 10996
rect 16724 10956 16730 10968
rect 16853 10965 16865 10968
rect 16899 10965 16911 10999
rect 16853 10959 16911 10965
rect 16942 10956 16948 11008
rect 17000 10996 17006 11008
rect 17052 10996 17080 11095
rect 17402 11092 17408 11144
rect 17460 11092 17466 11144
rect 17512 11132 17540 11240
rect 18506 11228 18512 11280
rect 18564 11268 18570 11280
rect 18966 11268 18972 11280
rect 18564 11240 18972 11268
rect 18564 11228 18570 11240
rect 18966 11228 18972 11240
rect 19024 11228 19030 11280
rect 19702 11268 19708 11280
rect 19444 11240 19708 11268
rect 18138 11160 18144 11212
rect 18196 11200 18202 11212
rect 18325 11203 18383 11209
rect 18325 11200 18337 11203
rect 18196 11172 18337 11200
rect 18196 11160 18202 11172
rect 18325 11169 18337 11172
rect 18371 11169 18383 11203
rect 18325 11163 18383 11169
rect 19150 11160 19156 11212
rect 19208 11200 19214 11212
rect 19334 11200 19340 11212
rect 19208 11172 19340 11200
rect 19208 11160 19214 11172
rect 19334 11160 19340 11172
rect 19392 11160 19398 11212
rect 17862 11132 17868 11144
rect 17512 11104 17868 11132
rect 17862 11092 17868 11104
rect 17920 11132 17926 11144
rect 19444 11132 19472 11240
rect 19702 11228 19708 11240
rect 19760 11228 19766 11280
rect 20806 11228 20812 11280
rect 20864 11268 20870 11280
rect 22741 11271 22799 11277
rect 22741 11268 22753 11271
rect 20864 11240 22753 11268
rect 20864 11228 20870 11240
rect 22741 11237 22753 11240
rect 22787 11237 22799 11271
rect 22741 11231 22799 11237
rect 19978 11200 19984 11212
rect 19536 11172 19984 11200
rect 19536 11141 19564 11172
rect 19978 11160 19984 11172
rect 20036 11160 20042 11212
rect 20162 11160 20168 11212
rect 20220 11200 20226 11212
rect 23201 11203 23259 11209
rect 23201 11200 23213 11203
rect 20220 11172 23213 11200
rect 20220 11160 20226 11172
rect 23201 11169 23213 11172
rect 23247 11169 23259 11203
rect 23201 11163 23259 11169
rect 23385 11203 23443 11209
rect 23385 11169 23397 11203
rect 23431 11169 23443 11203
rect 23385 11163 23443 11169
rect 17920 11104 19472 11132
rect 19521 11135 19579 11141
rect 17920 11092 17926 11104
rect 19521 11101 19533 11135
rect 19567 11101 19579 11135
rect 20441 11135 20499 11141
rect 19521 11095 19579 11101
rect 20180 11104 20392 11132
rect 18233 11067 18291 11073
rect 18233 11033 18245 11067
rect 18279 11064 18291 11067
rect 18414 11064 18420 11076
rect 18279 11036 18420 11064
rect 18279 11033 18291 11036
rect 18233 11027 18291 11033
rect 18414 11024 18420 11036
rect 18472 11024 18478 11076
rect 18690 11024 18696 11076
rect 18748 11064 18754 11076
rect 20180 11064 20208 11104
rect 18748 11036 20208 11064
rect 20257 11067 20315 11073
rect 18748 11024 18754 11036
rect 20257 11033 20269 11067
rect 20303 11033 20315 11067
rect 20364 11064 20392 11104
rect 20441 11101 20453 11135
rect 20487 11132 20499 11135
rect 20990 11132 20996 11144
rect 20487 11104 20996 11132
rect 20487 11101 20499 11104
rect 20441 11095 20499 11101
rect 20990 11092 20996 11104
rect 21048 11092 21054 11144
rect 21085 11135 21143 11141
rect 21085 11101 21097 11135
rect 21131 11132 21143 11135
rect 21358 11132 21364 11144
rect 21131 11104 21364 11132
rect 21131 11101 21143 11104
rect 21085 11095 21143 11101
rect 21358 11092 21364 11104
rect 21416 11092 21422 11144
rect 21726 11092 21732 11144
rect 21784 11092 21790 11144
rect 23400 11132 23428 11163
rect 24578 11132 24584 11144
rect 22066 11104 23244 11132
rect 23400 11104 24584 11132
rect 22066 11064 22094 11104
rect 20364 11036 22094 11064
rect 22465 11067 22523 11073
rect 20257 11027 20315 11033
rect 22465 11033 22477 11067
rect 22511 11064 22523 11067
rect 23109 11067 23167 11073
rect 23109 11064 23121 11067
rect 22511 11036 23121 11064
rect 22511 11033 22523 11036
rect 22465 11027 22523 11033
rect 23109 11033 23121 11036
rect 23155 11033 23167 11067
rect 23216 11064 23244 11104
rect 24578 11092 24584 11104
rect 24636 11092 24642 11144
rect 23474 11064 23480 11076
rect 23216 11036 23480 11064
rect 23109 11027 23167 11033
rect 17000 10968 17080 10996
rect 17000 10956 17006 10968
rect 17862 10956 17868 11008
rect 17920 10996 17926 11008
rect 18141 10999 18199 11005
rect 18141 10996 18153 10999
rect 17920 10968 18153 10996
rect 17920 10956 17926 10968
rect 18141 10965 18153 10968
rect 18187 10965 18199 10999
rect 18141 10959 18199 10965
rect 19334 10956 19340 11008
rect 19392 10996 19398 11008
rect 19794 10996 19800 11008
rect 19392 10968 19800 10996
rect 19392 10956 19398 10968
rect 19794 10956 19800 10968
rect 19852 10956 19858 11008
rect 20272 10996 20300 11027
rect 20438 10996 20444 11008
rect 20272 10968 20444 10996
rect 20438 10956 20444 10968
rect 20496 10956 20502 11008
rect 20898 10956 20904 11008
rect 20956 10956 20962 11008
rect 21358 10956 21364 11008
rect 21416 10996 21422 11008
rect 22480 10996 22508 11027
rect 23474 11024 23480 11036
rect 23532 11024 23538 11076
rect 21416 10968 22508 10996
rect 21416 10956 21422 10968
rect 25222 10956 25228 11008
rect 25280 10956 25286 11008
rect 1104 10906 25852 10928
rect 1104 10854 7950 10906
rect 8002 10854 8014 10906
rect 8066 10854 8078 10906
rect 8130 10854 8142 10906
rect 8194 10854 8206 10906
rect 8258 10854 17950 10906
rect 18002 10854 18014 10906
rect 18066 10854 18078 10906
rect 18130 10854 18142 10906
rect 18194 10854 18206 10906
rect 18258 10854 25852 10906
rect 1104 10832 25852 10854
rect 10778 10752 10784 10804
rect 10836 10792 10842 10804
rect 10965 10795 11023 10801
rect 10965 10792 10977 10795
rect 10836 10764 10977 10792
rect 10836 10752 10842 10764
rect 10965 10761 10977 10764
rect 11011 10761 11023 10795
rect 10965 10755 11023 10761
rect 11422 10752 11428 10804
rect 11480 10792 11486 10804
rect 11701 10795 11759 10801
rect 11701 10792 11713 10795
rect 11480 10764 11713 10792
rect 11480 10752 11486 10764
rect 11701 10761 11713 10764
rect 11747 10761 11759 10795
rect 11701 10755 11759 10761
rect 11790 10752 11796 10804
rect 11848 10792 11854 10804
rect 12161 10795 12219 10801
rect 12161 10792 12173 10795
rect 11848 10764 12173 10792
rect 11848 10752 11854 10764
rect 12161 10761 12173 10764
rect 12207 10792 12219 10795
rect 12250 10792 12256 10804
rect 12207 10764 12256 10792
rect 12207 10761 12219 10764
rect 12161 10755 12219 10761
rect 12250 10752 12256 10764
rect 12308 10752 12314 10804
rect 12526 10752 12532 10804
rect 12584 10752 12590 10804
rect 13722 10752 13728 10804
rect 13780 10792 13786 10804
rect 13909 10795 13967 10801
rect 13909 10792 13921 10795
rect 13780 10764 13921 10792
rect 13780 10752 13786 10764
rect 13909 10761 13921 10764
rect 13955 10761 13967 10795
rect 13909 10755 13967 10761
rect 14366 10752 14372 10804
rect 14424 10752 14430 10804
rect 15197 10795 15255 10801
rect 15197 10761 15209 10795
rect 15243 10792 15255 10795
rect 15562 10792 15568 10804
rect 15243 10764 15568 10792
rect 15243 10761 15255 10764
rect 15197 10755 15255 10761
rect 15562 10752 15568 10764
rect 15620 10792 15626 10804
rect 15930 10792 15936 10804
rect 15620 10764 15936 10792
rect 15620 10752 15626 10764
rect 15930 10752 15936 10764
rect 15988 10752 15994 10804
rect 16114 10752 16120 10804
rect 16172 10792 16178 10804
rect 20622 10792 20628 10804
rect 16172 10764 20628 10792
rect 16172 10752 16178 10764
rect 20622 10752 20628 10764
rect 20680 10752 20686 10804
rect 20898 10752 20904 10804
rect 20956 10792 20962 10804
rect 20956 10764 21312 10792
rect 20956 10752 20962 10764
rect 8938 10684 8944 10736
rect 8996 10724 9002 10736
rect 9493 10727 9551 10733
rect 9493 10724 9505 10727
rect 8996 10696 9505 10724
rect 8996 10684 9002 10696
rect 9493 10693 9505 10696
rect 9539 10693 9551 10727
rect 9493 10687 9551 10693
rect 10502 10684 10508 10736
rect 10560 10684 10566 10736
rect 12989 10727 13047 10733
rect 12989 10724 13001 10727
rect 12406 10696 13001 10724
rect 9214 10616 9220 10668
rect 9272 10616 9278 10668
rect 8938 10548 8944 10600
rect 8996 10588 9002 10600
rect 12406 10588 12434 10696
rect 12989 10693 13001 10696
rect 13035 10724 13047 10727
rect 13814 10724 13820 10736
rect 13035 10696 13820 10724
rect 13035 10693 13047 10696
rect 12989 10687 13047 10693
rect 13814 10684 13820 10696
rect 13872 10684 13878 10736
rect 13924 10696 16160 10724
rect 12897 10659 12955 10665
rect 12897 10625 12909 10659
rect 12943 10656 12955 10659
rect 13722 10656 13728 10668
rect 12943 10628 13728 10656
rect 12943 10625 12955 10628
rect 12897 10619 12955 10625
rect 13722 10616 13728 10628
rect 13780 10616 13786 10668
rect 8996 10560 12434 10588
rect 13173 10591 13231 10597
rect 8996 10548 9002 10560
rect 13173 10557 13185 10591
rect 13219 10588 13231 10591
rect 13354 10588 13360 10600
rect 13219 10560 13360 10588
rect 13219 10557 13231 10560
rect 13173 10551 13231 10557
rect 13354 10548 13360 10560
rect 13412 10588 13418 10600
rect 13924 10588 13952 10696
rect 14277 10659 14335 10665
rect 14277 10625 14289 10659
rect 14323 10656 14335 10659
rect 14734 10656 14740 10668
rect 14323 10628 14740 10656
rect 14323 10625 14335 10628
rect 14277 10619 14335 10625
rect 14734 10616 14740 10628
rect 14792 10616 14798 10668
rect 15841 10659 15899 10665
rect 15841 10656 15853 10659
rect 15304 10628 15853 10656
rect 13412 10560 13952 10588
rect 14461 10591 14519 10597
rect 13412 10548 13418 10560
rect 14461 10557 14473 10591
rect 14507 10557 14519 10591
rect 14461 10551 14519 10557
rect 14476 10520 14504 10551
rect 13556 10492 14504 10520
rect 14752 10520 14780 10616
rect 14921 10591 14979 10597
rect 14921 10557 14933 10591
rect 14967 10588 14979 10591
rect 15304 10588 15332 10628
rect 15841 10625 15853 10628
rect 15887 10625 15899 10659
rect 15841 10619 15899 10625
rect 14967 10560 15332 10588
rect 14967 10557 14979 10560
rect 14921 10551 14979 10557
rect 15378 10520 15384 10532
rect 14752 10492 15384 10520
rect 13556 10464 13584 10492
rect 15378 10480 15384 10492
rect 15436 10480 15442 10532
rect 15473 10523 15531 10529
rect 15473 10489 15485 10523
rect 15519 10520 15531 10523
rect 15562 10520 15568 10532
rect 15519 10492 15568 10520
rect 15519 10489 15531 10492
rect 15473 10483 15531 10489
rect 15562 10480 15568 10492
rect 15620 10480 15626 10532
rect 15856 10520 15884 10619
rect 16132 10597 16160 10696
rect 16666 10684 16672 10736
rect 16724 10724 16730 10736
rect 18049 10727 18107 10733
rect 16724 10696 18000 10724
rect 16724 10684 16730 10696
rect 16853 10659 16911 10665
rect 16853 10625 16865 10659
rect 16899 10656 16911 10659
rect 17218 10656 17224 10668
rect 16899 10628 17224 10656
rect 16899 10625 16911 10628
rect 16853 10619 16911 10625
rect 17218 10616 17224 10628
rect 17276 10616 17282 10668
rect 17310 10616 17316 10668
rect 17368 10656 17374 10668
rect 17972 10656 18000 10696
rect 18049 10693 18061 10727
rect 18095 10724 18107 10727
rect 19610 10724 19616 10736
rect 18095 10696 19616 10724
rect 18095 10693 18107 10696
rect 18049 10687 18107 10693
rect 19610 10684 19616 10696
rect 19668 10684 19674 10736
rect 21284 10724 21312 10764
rect 21450 10752 21456 10804
rect 21508 10752 21514 10804
rect 22738 10752 22744 10804
rect 22796 10792 22802 10804
rect 23293 10795 23351 10801
rect 23293 10792 23305 10795
rect 22796 10764 23305 10792
rect 22796 10752 22802 10764
rect 23293 10761 23305 10764
rect 23339 10761 23351 10795
rect 23293 10755 23351 10761
rect 23382 10724 23388 10736
rect 21284 10696 23388 10724
rect 23382 10684 23388 10696
rect 23440 10684 23446 10736
rect 18690 10656 18696 10668
rect 17368 10628 17540 10656
rect 17972 10628 18696 10656
rect 17368 10616 17374 10628
rect 16117 10591 16175 10597
rect 16117 10557 16129 10591
rect 16163 10588 16175 10591
rect 17402 10588 17408 10600
rect 16163 10560 17408 10588
rect 16163 10557 16175 10560
rect 16117 10551 16175 10557
rect 17402 10548 17408 10560
rect 17460 10548 17466 10600
rect 17512 10588 17540 10628
rect 18690 10616 18696 10628
rect 18748 10616 18754 10668
rect 19058 10616 19064 10668
rect 19116 10616 19122 10668
rect 19702 10616 19708 10668
rect 19760 10616 19766 10668
rect 21910 10656 21916 10668
rect 21114 10628 21916 10656
rect 21910 10616 21916 10628
rect 21968 10616 21974 10668
rect 23474 10616 23480 10668
rect 23532 10616 23538 10668
rect 23934 10616 23940 10668
rect 23992 10616 23998 10668
rect 19981 10591 20039 10597
rect 17512 10560 19748 10588
rect 19720 10532 19748 10560
rect 19981 10557 19993 10591
rect 20027 10588 20039 10591
rect 20070 10588 20076 10600
rect 20027 10560 20076 10588
rect 20027 10557 20039 10560
rect 19981 10551 20039 10557
rect 20070 10548 20076 10560
rect 20128 10548 20134 10600
rect 22002 10548 22008 10600
rect 22060 10548 22066 10600
rect 22281 10591 22339 10597
rect 22281 10557 22293 10591
rect 22327 10588 22339 10591
rect 23658 10588 23664 10600
rect 22327 10560 23664 10588
rect 22327 10557 22339 10560
rect 22281 10551 22339 10557
rect 23658 10548 23664 10560
rect 23716 10548 23722 10600
rect 24762 10548 24768 10600
rect 24820 10548 24826 10600
rect 15856 10492 19334 10520
rect 13538 10412 13544 10464
rect 13596 10412 13602 10464
rect 14182 10412 14188 10464
rect 14240 10452 14246 10464
rect 14826 10452 14832 10464
rect 14240 10424 14832 10452
rect 14240 10412 14246 10424
rect 14826 10412 14832 10424
rect 14884 10452 14890 10464
rect 16482 10452 16488 10464
rect 14884 10424 16488 10452
rect 14884 10412 14890 10424
rect 16482 10412 16488 10424
rect 16540 10412 16546 10464
rect 16666 10412 16672 10464
rect 16724 10452 16730 10464
rect 17497 10455 17555 10461
rect 17497 10452 17509 10455
rect 16724 10424 17509 10452
rect 16724 10412 16730 10424
rect 17497 10421 17509 10424
rect 17543 10421 17555 10455
rect 17497 10415 17555 10421
rect 18141 10455 18199 10461
rect 18141 10421 18153 10455
rect 18187 10452 18199 10455
rect 18322 10452 18328 10464
rect 18187 10424 18328 10452
rect 18187 10421 18199 10424
rect 18141 10415 18199 10421
rect 18322 10412 18328 10424
rect 18380 10412 18386 10464
rect 18690 10412 18696 10464
rect 18748 10412 18754 10464
rect 19150 10412 19156 10464
rect 19208 10412 19214 10464
rect 19306 10452 19334 10492
rect 19702 10480 19708 10532
rect 19760 10480 19766 10532
rect 20162 10452 20168 10464
rect 19306 10424 20168 10452
rect 20162 10412 20168 10424
rect 20220 10412 20226 10464
rect 1104 10362 25852 10384
rect 1104 10310 2950 10362
rect 3002 10310 3014 10362
rect 3066 10310 3078 10362
rect 3130 10310 3142 10362
rect 3194 10310 3206 10362
rect 3258 10310 12950 10362
rect 13002 10310 13014 10362
rect 13066 10310 13078 10362
rect 13130 10310 13142 10362
rect 13194 10310 13206 10362
rect 13258 10310 22950 10362
rect 23002 10310 23014 10362
rect 23066 10310 23078 10362
rect 23130 10310 23142 10362
rect 23194 10310 23206 10362
rect 23258 10310 25852 10362
rect 1104 10288 25852 10310
rect 12710 10208 12716 10260
rect 12768 10208 12774 10260
rect 13722 10208 13728 10260
rect 13780 10248 13786 10260
rect 15562 10248 15568 10260
rect 13780 10220 15568 10248
rect 13780 10208 13786 10220
rect 15562 10208 15568 10220
rect 15620 10208 15626 10260
rect 15654 10208 15660 10260
rect 15712 10208 15718 10260
rect 16574 10208 16580 10260
rect 16632 10248 16638 10260
rect 16853 10251 16911 10257
rect 16853 10248 16865 10251
rect 16632 10220 16865 10248
rect 16632 10208 16638 10220
rect 16853 10217 16865 10220
rect 16899 10217 16911 10251
rect 16853 10211 16911 10217
rect 17310 10208 17316 10260
rect 17368 10248 17374 10260
rect 19610 10248 19616 10260
rect 17368 10220 19616 10248
rect 17368 10208 17374 10220
rect 19610 10208 19616 10220
rect 19668 10208 19674 10260
rect 19794 10208 19800 10260
rect 19852 10248 19858 10260
rect 19852 10220 19932 10248
rect 19852 10208 19858 10220
rect 12434 10140 12440 10192
rect 12492 10180 12498 10192
rect 14461 10183 14519 10189
rect 14461 10180 14473 10183
rect 12492 10152 14473 10180
rect 12492 10140 12498 10152
rect 14461 10149 14473 10152
rect 14507 10149 14519 10183
rect 15580 10180 15608 10208
rect 16022 10180 16028 10192
rect 14461 10143 14519 10149
rect 14752 10152 15148 10180
rect 15580 10152 16028 10180
rect 9122 10072 9128 10124
rect 9180 10072 9186 10124
rect 9398 10072 9404 10124
rect 9456 10072 9462 10124
rect 11054 10112 11060 10124
rect 10520 10084 11060 10112
rect 10520 10056 10548 10084
rect 11054 10072 11060 10084
rect 11112 10112 11118 10124
rect 11149 10115 11207 10121
rect 11149 10112 11161 10115
rect 11112 10084 11161 10112
rect 11112 10072 11118 10084
rect 11149 10081 11161 10084
rect 11195 10081 11207 10115
rect 11149 10075 11207 10081
rect 11330 10072 11336 10124
rect 11388 10112 11394 10124
rect 11977 10115 12035 10121
rect 11977 10112 11989 10115
rect 11388 10084 11989 10112
rect 11388 10072 11394 10084
rect 11977 10081 11989 10084
rect 12023 10081 12035 10115
rect 11977 10075 12035 10081
rect 12069 10115 12127 10121
rect 12069 10081 12081 10115
rect 12115 10081 12127 10115
rect 12069 10075 12127 10081
rect 8573 10047 8631 10053
rect 8573 10013 8585 10047
rect 8619 10013 8631 10047
rect 8573 10007 8631 10013
rect 8588 9976 8616 10007
rect 10502 10004 10508 10056
rect 10560 10004 10566 10056
rect 12084 10044 12112 10075
rect 13354 10072 13360 10124
rect 13412 10072 13418 10124
rect 14752 10112 14780 10152
rect 14918 10112 14924 10124
rect 14108 10084 14780 10112
rect 14844 10084 14924 10112
rect 10888 10016 12112 10044
rect 9674 9976 9680 9988
rect 8588 9948 9680 9976
rect 9674 9936 9680 9948
rect 9732 9936 9738 9988
rect 8386 9868 8392 9920
rect 8444 9868 8450 9920
rect 10410 9868 10416 9920
rect 10468 9908 10474 9920
rect 10888 9917 10916 10016
rect 12618 10004 12624 10056
rect 12676 10044 12682 10056
rect 13173 10047 13231 10053
rect 13173 10044 13185 10047
rect 12676 10016 13185 10044
rect 12676 10004 12682 10016
rect 13173 10013 13185 10016
rect 13219 10013 13231 10047
rect 13173 10007 13231 10013
rect 13538 10004 13544 10056
rect 13596 10044 13602 10056
rect 14108 10053 14136 10084
rect 14844 10053 14872 10084
rect 14918 10072 14924 10084
rect 14976 10072 14982 10124
rect 15120 10121 15148 10152
rect 16022 10140 16028 10152
rect 16080 10140 16086 10192
rect 16482 10180 16488 10192
rect 16132 10152 16488 10180
rect 16132 10121 16160 10152
rect 16482 10140 16488 10152
rect 16540 10180 16546 10192
rect 16540 10152 17540 10180
rect 16540 10140 16546 10152
rect 15105 10115 15163 10121
rect 15105 10081 15117 10115
rect 15151 10112 15163 10115
rect 16117 10115 16175 10121
rect 15151 10084 15608 10112
rect 15151 10081 15163 10084
rect 15105 10075 15163 10081
rect 15580 10056 15608 10084
rect 16117 10081 16129 10115
rect 16163 10081 16175 10115
rect 16117 10075 16175 10081
rect 16209 10115 16267 10121
rect 16209 10081 16221 10115
rect 16255 10081 16267 10115
rect 16209 10075 16267 10081
rect 14093 10047 14151 10053
rect 14093 10044 14105 10047
rect 13596 10016 14105 10044
rect 13596 10004 13602 10016
rect 14093 10013 14105 10016
rect 14139 10013 14151 10047
rect 14093 10007 14151 10013
rect 14829 10047 14887 10053
rect 14829 10013 14841 10047
rect 14875 10013 14887 10047
rect 14829 10007 14887 10013
rect 15562 10004 15568 10056
rect 15620 10044 15626 10056
rect 16224 10044 16252 10075
rect 17402 10072 17408 10124
rect 17460 10072 17466 10124
rect 17512 10112 17540 10152
rect 18414 10140 18420 10192
rect 18472 10180 18478 10192
rect 18874 10180 18880 10192
rect 18472 10152 18880 10180
rect 18472 10140 18478 10152
rect 18874 10140 18880 10152
rect 18932 10140 18938 10192
rect 18601 10115 18659 10121
rect 17512 10084 18552 10112
rect 17678 10044 17684 10056
rect 15620 10016 16252 10044
rect 16316 10016 17684 10044
rect 15620 10004 15626 10016
rect 15746 9976 15752 9988
rect 11532 9948 15752 9976
rect 11532 9917 11560 9948
rect 15746 9936 15752 9948
rect 15804 9936 15810 9988
rect 10873 9911 10931 9917
rect 10873 9908 10885 9911
rect 10468 9880 10885 9908
rect 10468 9868 10474 9880
rect 10873 9877 10885 9880
rect 10919 9877 10931 9911
rect 10873 9871 10931 9877
rect 11517 9911 11575 9917
rect 11517 9877 11529 9911
rect 11563 9877 11575 9911
rect 11517 9871 11575 9877
rect 11882 9868 11888 9920
rect 11940 9868 11946 9920
rect 13081 9911 13139 9917
rect 13081 9877 13093 9911
rect 13127 9908 13139 9911
rect 13814 9908 13820 9920
rect 13127 9880 13820 9908
rect 13127 9877 13139 9880
rect 13081 9871 13139 9877
rect 13814 9868 13820 9880
rect 13872 9868 13878 9920
rect 13909 9911 13967 9917
rect 13909 9877 13921 9911
rect 13955 9908 13967 9911
rect 14090 9908 14096 9920
rect 13955 9880 14096 9908
rect 13955 9877 13967 9880
rect 13909 9871 13967 9877
rect 14090 9868 14096 9880
rect 14148 9908 14154 9920
rect 14921 9911 14979 9917
rect 14921 9908 14933 9911
rect 14148 9880 14933 9908
rect 14148 9868 14154 9880
rect 14921 9877 14933 9880
rect 14967 9877 14979 9911
rect 14921 9871 14979 9877
rect 16025 9911 16083 9917
rect 16025 9877 16037 9911
rect 16071 9908 16083 9911
rect 16316 9908 16344 10016
rect 17678 10004 17684 10016
rect 17736 10004 17742 10056
rect 18524 10053 18552 10084
rect 18601 10081 18613 10115
rect 18647 10112 18659 10115
rect 18690 10112 18696 10124
rect 18647 10084 18696 10112
rect 18647 10081 18659 10084
rect 18601 10075 18659 10081
rect 18690 10072 18696 10084
rect 18748 10072 18754 10124
rect 18785 10115 18843 10121
rect 18785 10081 18797 10115
rect 18831 10112 18843 10115
rect 19904 10112 19932 10220
rect 20070 10208 20076 10260
rect 20128 10208 20134 10260
rect 20162 10208 20168 10260
rect 20220 10248 20226 10260
rect 24394 10248 24400 10260
rect 20220 10220 24400 10248
rect 20220 10208 20226 10220
rect 24394 10208 24400 10220
rect 24452 10208 24458 10260
rect 25130 10208 25136 10260
rect 25188 10208 25194 10260
rect 19978 10140 19984 10192
rect 20036 10180 20042 10192
rect 20349 10183 20407 10189
rect 20349 10180 20361 10183
rect 20036 10152 20361 10180
rect 20036 10140 20042 10152
rect 20349 10149 20361 10152
rect 20395 10149 20407 10183
rect 20349 10143 20407 10149
rect 20806 10140 20812 10192
rect 20864 10140 20870 10192
rect 21910 10140 21916 10192
rect 21968 10140 21974 10192
rect 24118 10140 24124 10192
rect 24176 10180 24182 10192
rect 25148 10180 25176 10208
rect 24176 10152 25176 10180
rect 24176 10140 24182 10152
rect 21269 10115 21327 10121
rect 21269 10112 21281 10115
rect 18831 10084 19840 10112
rect 19904 10084 21281 10112
rect 18831 10081 18843 10084
rect 18785 10075 18843 10081
rect 18509 10047 18567 10053
rect 18509 10013 18521 10047
rect 18555 10013 18567 10047
rect 18509 10007 18567 10013
rect 18874 10004 18880 10056
rect 18932 10044 18938 10056
rect 19429 10047 19487 10053
rect 19429 10044 19441 10047
rect 18932 10016 19441 10044
rect 18932 10004 18938 10016
rect 19429 10013 19441 10016
rect 19475 10013 19487 10047
rect 19812 10044 19840 10084
rect 21269 10081 21281 10084
rect 21315 10081 21327 10115
rect 21269 10075 21327 10081
rect 21450 10072 21456 10124
rect 21508 10072 21514 10124
rect 22278 10072 22284 10124
rect 22336 10072 22342 10124
rect 22557 10115 22615 10121
rect 22557 10081 22569 10115
rect 22603 10112 22615 10115
rect 25222 10112 25228 10124
rect 22603 10084 25228 10112
rect 22603 10081 22615 10084
rect 22557 10075 22615 10081
rect 25222 10072 25228 10084
rect 25280 10072 25286 10124
rect 21082 10044 21088 10056
rect 19812 10016 21088 10044
rect 19429 10007 19487 10013
rect 21082 10004 21088 10016
rect 21140 10004 21146 10056
rect 21174 10004 21180 10056
rect 21232 10044 21238 10056
rect 21818 10044 21824 10056
rect 21232 10016 21824 10044
rect 21232 10004 21238 10016
rect 21818 10004 21824 10016
rect 21876 10004 21882 10056
rect 17221 9979 17279 9985
rect 17221 9945 17233 9979
rect 17267 9976 17279 9979
rect 20898 9976 20904 9988
rect 17267 9948 20904 9976
rect 17267 9945 17279 9948
rect 17221 9939 17279 9945
rect 20898 9936 20904 9948
rect 20956 9936 20962 9988
rect 21450 9976 21456 9988
rect 21376 9948 21456 9976
rect 16071 9880 16344 9908
rect 16071 9877 16083 9880
rect 16025 9871 16083 9877
rect 16574 9868 16580 9920
rect 16632 9908 16638 9920
rect 17310 9908 17316 9920
rect 16632 9880 17316 9908
rect 16632 9868 16638 9880
rect 17310 9868 17316 9880
rect 17368 9868 17374 9920
rect 18141 9911 18199 9917
rect 18141 9877 18153 9911
rect 18187 9908 18199 9911
rect 18414 9908 18420 9920
rect 18187 9880 18420 9908
rect 18187 9877 18199 9880
rect 18141 9871 18199 9877
rect 18414 9868 18420 9880
rect 18472 9868 18478 9920
rect 19242 9868 19248 9920
rect 19300 9908 19306 9920
rect 20622 9908 20628 9920
rect 19300 9880 20628 9908
rect 19300 9868 19306 9880
rect 20622 9868 20628 9880
rect 20680 9868 20686 9920
rect 21177 9911 21235 9917
rect 21177 9877 21189 9911
rect 21223 9908 21235 9911
rect 21376 9908 21404 9948
rect 21450 9936 21456 9948
rect 21508 9936 21514 9988
rect 21910 9936 21916 9988
rect 21968 9976 21974 9988
rect 21968 9948 23046 9976
rect 21968 9936 21974 9948
rect 21223 9880 21404 9908
rect 21223 9877 21235 9880
rect 21177 9871 21235 9877
rect 24026 9868 24032 9920
rect 24084 9868 24090 9920
rect 24578 9868 24584 9920
rect 24636 9868 24642 9920
rect 1104 9818 25852 9840
rect 1104 9766 7950 9818
rect 8002 9766 8014 9818
rect 8066 9766 8078 9818
rect 8130 9766 8142 9818
rect 8194 9766 8206 9818
rect 8258 9766 17950 9818
rect 18002 9766 18014 9818
rect 18066 9766 18078 9818
rect 18130 9766 18142 9818
rect 18194 9766 18206 9818
rect 18258 9766 25852 9818
rect 1104 9744 25852 9766
rect 3970 9664 3976 9716
rect 4028 9704 4034 9716
rect 9306 9704 9312 9716
rect 4028 9676 9312 9704
rect 4028 9664 4034 9676
rect 9306 9664 9312 9676
rect 9364 9664 9370 9716
rect 10502 9704 10508 9716
rect 9784 9676 10508 9704
rect 3326 9596 3332 9648
rect 3384 9636 3390 9648
rect 6270 9636 6276 9648
rect 3384 9608 6276 9636
rect 3384 9596 3390 9608
rect 6270 9596 6276 9608
rect 6328 9596 6334 9648
rect 9784 9636 9812 9676
rect 10502 9664 10508 9676
rect 10560 9664 10566 9716
rect 13538 9704 13544 9716
rect 12360 9676 13544 9704
rect 11514 9636 11520 9648
rect 9706 9608 9812 9636
rect 9876 9608 11520 9636
rect 7098 9460 7104 9512
rect 7156 9500 7162 9512
rect 8202 9500 8208 9512
rect 7156 9472 8208 9500
rect 7156 9460 7162 9472
rect 8202 9460 8208 9472
rect 8260 9460 8266 9512
rect 8481 9503 8539 9509
rect 8481 9500 8493 9503
rect 8312 9472 8493 9500
rect 7098 9324 7104 9376
rect 7156 9364 7162 9376
rect 7837 9367 7895 9373
rect 7837 9364 7849 9367
rect 7156 9336 7849 9364
rect 7156 9324 7162 9336
rect 7837 9333 7849 9336
rect 7883 9364 7895 9367
rect 8312 9364 8340 9472
rect 8481 9469 8493 9472
rect 8527 9500 8539 9503
rect 9876 9500 9904 9608
rect 11514 9596 11520 9608
rect 11572 9636 11578 9648
rect 12360 9636 12388 9676
rect 13538 9664 13544 9676
rect 13596 9664 13602 9716
rect 13814 9664 13820 9716
rect 13872 9704 13878 9716
rect 17218 9704 17224 9716
rect 13872 9676 17224 9704
rect 13872 9664 13878 9676
rect 17218 9664 17224 9676
rect 17276 9664 17282 9716
rect 17494 9664 17500 9716
rect 17552 9704 17558 9716
rect 21450 9704 21456 9716
rect 17552 9676 21456 9704
rect 17552 9664 17558 9676
rect 21450 9664 21456 9676
rect 21508 9664 21514 9716
rect 11572 9608 12388 9636
rect 11572 9596 11578 9608
rect 13262 9596 13268 9648
rect 13320 9636 13326 9648
rect 15105 9639 15163 9645
rect 15105 9636 15117 9639
rect 13320 9608 15117 9636
rect 13320 9596 13326 9608
rect 15105 9605 15117 9608
rect 15151 9636 15163 9639
rect 15151 9608 16252 9636
rect 15151 9605 15163 9608
rect 15105 9599 15163 9605
rect 11698 9528 11704 9580
rect 11756 9528 11762 9580
rect 13814 9568 13820 9580
rect 13110 9540 13820 9568
rect 13814 9528 13820 9540
rect 13872 9528 13878 9580
rect 15013 9571 15071 9577
rect 15013 9537 15025 9571
rect 15059 9568 15071 9571
rect 15194 9568 15200 9580
rect 15059 9540 15200 9568
rect 15059 9537 15071 9540
rect 15013 9531 15071 9537
rect 15194 9528 15200 9540
rect 15252 9528 15258 9580
rect 15470 9528 15476 9580
rect 15528 9568 15534 9580
rect 15746 9568 15752 9580
rect 15528 9540 15752 9568
rect 15528 9528 15534 9540
rect 15746 9528 15752 9540
rect 15804 9528 15810 9580
rect 16114 9528 16120 9580
rect 16172 9528 16178 9580
rect 16224 9568 16252 9608
rect 16942 9596 16948 9648
rect 17000 9596 17006 9648
rect 17862 9636 17868 9648
rect 17052 9608 17868 9636
rect 17052 9568 17080 9608
rect 17862 9596 17868 9608
rect 17920 9596 17926 9648
rect 19242 9636 19248 9648
rect 19182 9608 19248 9636
rect 19242 9596 19248 9608
rect 19300 9596 19306 9648
rect 19610 9596 19616 9648
rect 19668 9636 19674 9648
rect 20257 9639 20315 9645
rect 20257 9636 20269 9639
rect 19668 9608 20269 9636
rect 19668 9596 19674 9608
rect 20257 9605 20269 9608
rect 20303 9605 20315 9639
rect 20257 9599 20315 9605
rect 21177 9639 21235 9645
rect 21177 9605 21189 9639
rect 21223 9636 21235 9639
rect 21266 9636 21272 9648
rect 21223 9608 21272 9636
rect 21223 9605 21235 9608
rect 21177 9599 21235 9605
rect 21266 9596 21272 9608
rect 21324 9596 21330 9648
rect 23290 9596 23296 9648
rect 23348 9596 23354 9648
rect 16224 9540 17080 9568
rect 22094 9528 22100 9580
rect 22152 9528 22158 9580
rect 23014 9528 23020 9580
rect 23072 9568 23078 9580
rect 23937 9571 23995 9577
rect 23937 9568 23949 9571
rect 23072 9540 23949 9568
rect 23072 9528 23078 9540
rect 23937 9537 23949 9540
rect 23983 9537 23995 9571
rect 23937 9531 23995 9537
rect 8527 9472 9904 9500
rect 8527 9469 8539 9472
rect 8481 9463 8539 9469
rect 9950 9460 9956 9512
rect 10008 9460 10014 9512
rect 10594 9460 10600 9512
rect 10652 9460 10658 9512
rect 11977 9503 12035 9509
rect 11977 9469 11989 9503
rect 12023 9500 12035 9503
rect 12023 9472 13308 9500
rect 12023 9469 12035 9472
rect 11977 9463 12035 9469
rect 9766 9392 9772 9444
rect 9824 9432 9830 9444
rect 13280 9432 13308 9472
rect 13354 9460 13360 9512
rect 13412 9500 13418 9512
rect 13909 9503 13967 9509
rect 13909 9500 13921 9503
rect 13412 9472 13921 9500
rect 13412 9460 13418 9472
rect 13909 9469 13921 9472
rect 13955 9469 13967 9503
rect 13909 9463 13967 9469
rect 15289 9503 15347 9509
rect 15289 9469 15301 9503
rect 15335 9500 15347 9503
rect 16390 9500 16396 9512
rect 15335 9472 16396 9500
rect 15335 9469 15347 9472
rect 15289 9463 15347 9469
rect 16390 9460 16396 9472
rect 16448 9460 16454 9512
rect 17681 9503 17739 9509
rect 17681 9469 17693 9503
rect 17727 9500 17739 9503
rect 17727 9472 17816 9500
rect 17727 9469 17739 9472
rect 17681 9463 17739 9469
rect 13538 9432 13544 9444
rect 9824 9404 11376 9432
rect 13280 9404 13544 9432
rect 9824 9392 9830 9404
rect 7883 9336 8340 9364
rect 7883 9333 7895 9336
rect 7837 9327 7895 9333
rect 11054 9324 11060 9376
rect 11112 9364 11118 9376
rect 11241 9367 11299 9373
rect 11241 9364 11253 9367
rect 11112 9336 11253 9364
rect 11112 9324 11118 9336
rect 11241 9333 11253 9336
rect 11287 9333 11299 9367
rect 11348 9364 11376 9404
rect 13538 9392 13544 9404
rect 13596 9392 13602 9444
rect 14274 9392 14280 9444
rect 14332 9432 14338 9444
rect 14645 9435 14703 9441
rect 14645 9432 14657 9435
rect 14332 9404 14657 9432
rect 14332 9392 14338 9404
rect 14645 9401 14657 9404
rect 14691 9401 14703 9435
rect 14645 9395 14703 9401
rect 15562 9392 15568 9444
rect 15620 9432 15626 9444
rect 15657 9435 15715 9441
rect 15657 9432 15669 9435
rect 15620 9404 15669 9432
rect 15620 9392 15626 9404
rect 15657 9401 15669 9404
rect 15703 9401 15715 9435
rect 15657 9395 15715 9401
rect 16298 9392 16304 9444
rect 16356 9392 16362 9444
rect 13262 9364 13268 9376
rect 11348 9336 13268 9364
rect 11241 9327 11299 9333
rect 13262 9324 13268 9336
rect 13320 9324 13326 9376
rect 13449 9367 13507 9373
rect 13449 9333 13461 9367
rect 13495 9364 13507 9367
rect 15102 9364 15108 9376
rect 13495 9336 15108 9364
rect 13495 9333 13507 9336
rect 13449 9327 13507 9333
rect 15102 9324 15108 9336
rect 15160 9324 15166 9376
rect 17034 9324 17040 9376
rect 17092 9324 17098 9376
rect 17788 9364 17816 9472
rect 17954 9460 17960 9512
rect 18012 9460 18018 9512
rect 18046 9460 18052 9512
rect 18104 9500 18110 9512
rect 18966 9500 18972 9512
rect 18104 9472 18972 9500
rect 18104 9460 18110 9472
rect 18966 9460 18972 9472
rect 19024 9460 19030 9512
rect 20162 9460 20168 9512
rect 20220 9500 20226 9512
rect 20349 9503 20407 9509
rect 20349 9500 20361 9503
rect 20220 9472 20361 9500
rect 20220 9460 20226 9472
rect 20349 9469 20361 9472
rect 20395 9469 20407 9503
rect 20349 9463 20407 9469
rect 20533 9503 20591 9509
rect 20533 9469 20545 9503
rect 20579 9500 20591 9503
rect 24026 9500 24032 9512
rect 20579 9472 24032 9500
rect 20579 9469 20591 9472
rect 20533 9463 20591 9469
rect 24026 9460 24032 9472
rect 24084 9460 24090 9512
rect 24670 9460 24676 9512
rect 24728 9460 24734 9512
rect 20254 9432 20260 9444
rect 18984 9404 20260 9432
rect 18984 9364 19012 9404
rect 20254 9392 20260 9404
rect 20312 9432 20318 9444
rect 22278 9432 22284 9444
rect 20312 9404 22284 9432
rect 20312 9392 20318 9404
rect 22278 9392 22284 9404
rect 22336 9392 22342 9444
rect 17788 9336 19012 9364
rect 19058 9324 19064 9376
rect 19116 9364 19122 9376
rect 19429 9367 19487 9373
rect 19429 9364 19441 9367
rect 19116 9336 19441 9364
rect 19116 9324 19122 9336
rect 19429 9333 19441 9336
rect 19475 9333 19487 9367
rect 19429 9327 19487 9333
rect 19886 9324 19892 9376
rect 19944 9324 19950 9376
rect 20806 9324 20812 9376
rect 20864 9364 20870 9376
rect 21269 9367 21327 9373
rect 21269 9364 21281 9367
rect 20864 9336 21281 9364
rect 20864 9324 20870 9336
rect 21269 9333 21281 9336
rect 21315 9333 21327 9367
rect 21269 9327 21327 9333
rect 1104 9274 25852 9296
rect 1104 9222 2950 9274
rect 3002 9222 3014 9274
rect 3066 9222 3078 9274
rect 3130 9222 3142 9274
rect 3194 9222 3206 9274
rect 3258 9222 12950 9274
rect 13002 9222 13014 9274
rect 13066 9222 13078 9274
rect 13130 9222 13142 9274
rect 13194 9222 13206 9274
rect 13258 9222 22950 9274
rect 23002 9222 23014 9274
rect 23066 9222 23078 9274
rect 23130 9222 23142 9274
rect 23194 9222 23206 9274
rect 23258 9222 25852 9274
rect 1104 9200 25852 9222
rect 9674 9120 9680 9172
rect 9732 9160 9738 9172
rect 12345 9163 12403 9169
rect 12345 9160 12357 9163
rect 9732 9132 12357 9160
rect 9732 9120 9738 9132
rect 12345 9129 12357 9132
rect 12391 9129 12403 9163
rect 12345 9123 12403 9129
rect 12434 9120 12440 9172
rect 12492 9160 12498 9172
rect 12492 9132 13768 9160
rect 12492 9120 12498 9132
rect 11974 9052 11980 9104
rect 12032 9092 12038 9104
rect 12989 9095 13047 9101
rect 12989 9092 13001 9095
rect 12032 9064 13001 9092
rect 12032 9052 12038 9064
rect 12989 9061 13001 9064
rect 13035 9061 13047 9095
rect 13630 9092 13636 9104
rect 12989 9055 13047 9061
rect 13096 9064 13636 9092
rect 10321 9027 10379 9033
rect 10321 8993 10333 9027
rect 10367 9024 10379 9027
rect 13096 9024 13124 9064
rect 13630 9052 13636 9064
rect 13688 9052 13694 9104
rect 10367 8996 13124 9024
rect 10367 8993 10379 8996
rect 10321 8987 10379 8993
rect 13446 8984 13452 9036
rect 13504 9024 13510 9036
rect 13541 9027 13599 9033
rect 13541 9024 13553 9027
rect 13504 8996 13553 9024
rect 13504 8984 13510 8996
rect 13541 8993 13553 8996
rect 13587 8993 13599 9027
rect 13740 9024 13768 9132
rect 14090 9120 14096 9172
rect 14148 9160 14154 9172
rect 16850 9160 16856 9172
rect 14148 9132 16856 9160
rect 14148 9120 14154 9132
rect 16850 9120 16856 9132
rect 16908 9160 16914 9172
rect 17862 9160 17868 9172
rect 16908 9132 17868 9160
rect 16908 9120 16914 9132
rect 17862 9120 17868 9132
rect 17920 9120 17926 9172
rect 17954 9120 17960 9172
rect 18012 9160 18018 9172
rect 18877 9163 18935 9169
rect 18877 9160 18889 9163
rect 18012 9132 18889 9160
rect 18012 9120 18018 9132
rect 18877 9129 18889 9132
rect 18923 9129 18935 9163
rect 18877 9123 18935 9129
rect 19886 9120 19892 9172
rect 19944 9160 19950 9172
rect 25038 9160 25044 9172
rect 19944 9132 25044 9160
rect 19944 9120 19950 9132
rect 25038 9120 25044 9132
rect 25096 9120 25102 9172
rect 15194 9052 15200 9104
rect 15252 9092 15258 9104
rect 18690 9092 18696 9104
rect 15252 9064 18696 9092
rect 15252 9052 15258 9064
rect 18690 9052 18696 9064
rect 18748 9052 18754 9104
rect 15289 9027 15347 9033
rect 15289 9024 15301 9027
rect 13740 8996 15301 9024
rect 13541 8987 13599 8993
rect 15289 8993 15301 8996
rect 15335 9024 15347 9027
rect 16209 9027 16267 9033
rect 15335 8996 16068 9024
rect 15335 8993 15347 8996
rect 15289 8987 15347 8993
rect 9125 8959 9183 8965
rect 9125 8925 9137 8959
rect 9171 8956 9183 8959
rect 10410 8956 10416 8968
rect 9171 8928 10416 8956
rect 9171 8925 9183 8928
rect 9125 8919 9183 8925
rect 10410 8916 10416 8928
rect 10468 8916 10474 8968
rect 10597 8959 10655 8965
rect 10597 8925 10609 8959
rect 10643 8956 10655 8959
rect 11238 8956 11244 8968
rect 10643 8928 11244 8956
rect 10643 8925 10655 8928
rect 10597 8919 10655 8925
rect 11238 8916 11244 8928
rect 11296 8916 11302 8968
rect 11701 8959 11759 8965
rect 11701 8925 11713 8959
rect 11747 8956 11759 8959
rect 11882 8956 11888 8968
rect 11747 8928 11888 8956
rect 11747 8925 11759 8928
rect 11701 8919 11759 8925
rect 11882 8916 11888 8928
rect 11940 8916 11946 8968
rect 16040 8965 16068 8996
rect 16209 8993 16221 9027
rect 16255 9024 16267 9027
rect 16390 9024 16396 9036
rect 16255 8996 16396 9024
rect 16255 8993 16267 8996
rect 16209 8987 16267 8993
rect 16390 8984 16396 8996
rect 16448 8984 16454 9036
rect 18046 9024 18052 9036
rect 16500 8996 18052 9024
rect 12529 8959 12587 8965
rect 12529 8925 12541 8959
rect 12575 8925 12587 8959
rect 12529 8919 12587 8925
rect 13357 8959 13415 8965
rect 13357 8925 13369 8959
rect 13403 8956 13415 8959
rect 16025 8959 16083 8965
rect 13403 8928 15608 8956
rect 13403 8925 13415 8928
rect 13357 8919 13415 8925
rect 11422 8848 11428 8900
rect 11480 8888 11486 8900
rect 12342 8888 12348 8900
rect 11480 8860 12348 8888
rect 11480 8848 11486 8860
rect 12342 8848 12348 8860
rect 12400 8848 12406 8900
rect 12544 8888 12572 8919
rect 12544 8860 13768 8888
rect 13740 8832 13768 8860
rect 13906 8848 13912 8900
rect 13964 8888 13970 8900
rect 14369 8891 14427 8897
rect 14369 8888 14381 8891
rect 13964 8860 14381 8888
rect 13964 8848 13970 8860
rect 14369 8857 14381 8860
rect 14415 8857 14427 8891
rect 14369 8851 14427 8857
rect 8846 8780 8852 8832
rect 8904 8820 8910 8832
rect 9769 8823 9827 8829
rect 9769 8820 9781 8823
rect 8904 8792 9781 8820
rect 8904 8780 8910 8792
rect 9769 8789 9781 8792
rect 9815 8789 9827 8823
rect 9769 8783 9827 8789
rect 12250 8780 12256 8832
rect 12308 8820 12314 8832
rect 12434 8820 12440 8832
rect 12308 8792 12440 8820
rect 12308 8780 12314 8792
rect 12434 8780 12440 8792
rect 12492 8780 12498 8832
rect 13446 8780 13452 8832
rect 13504 8780 13510 8832
rect 13722 8780 13728 8832
rect 13780 8780 13786 8832
rect 14384 8820 14412 8851
rect 14550 8848 14556 8900
rect 14608 8848 14614 8900
rect 15580 8829 15608 8928
rect 16025 8925 16037 8959
rect 16071 8956 16083 8959
rect 16500 8956 16528 8996
rect 18046 8984 18052 8996
rect 18104 8984 18110 9036
rect 18414 8984 18420 9036
rect 18472 9024 18478 9036
rect 20073 9027 20131 9033
rect 20073 9024 20085 9027
rect 18472 8996 20085 9024
rect 18472 8984 18478 8996
rect 20073 8993 20085 8996
rect 20119 8993 20131 9027
rect 20073 8987 20131 8993
rect 20257 9027 20315 9033
rect 20257 8993 20269 9027
rect 20303 9024 20315 9027
rect 21450 9024 21456 9036
rect 20303 8996 21456 9024
rect 20303 8993 20315 8996
rect 20257 8987 20315 8993
rect 16071 8928 16528 8956
rect 16669 8959 16727 8965
rect 16071 8925 16083 8928
rect 16025 8919 16083 8925
rect 16669 8925 16681 8959
rect 16715 8956 16727 8959
rect 16850 8956 16856 8968
rect 16715 8928 16856 8956
rect 16715 8925 16727 8928
rect 16669 8919 16727 8925
rect 16850 8916 16856 8928
rect 16908 8916 16914 8968
rect 17129 8959 17187 8965
rect 17129 8925 17141 8959
rect 17175 8956 17187 8959
rect 17678 8956 17684 8968
rect 17175 8928 17684 8956
rect 17175 8925 17187 8928
rect 17129 8919 17187 8925
rect 17678 8916 17684 8928
rect 17736 8916 17742 8968
rect 18233 8959 18291 8965
rect 18233 8925 18245 8959
rect 18279 8956 18291 8959
rect 20272 8956 20300 8987
rect 21450 8984 21456 8996
rect 21508 8984 21514 9036
rect 18279 8928 20300 8956
rect 20993 8959 21051 8965
rect 18279 8925 18291 8928
rect 18233 8919 18291 8925
rect 20993 8925 21005 8959
rect 21039 8956 21051 8959
rect 21039 8928 22094 8956
rect 21039 8925 21051 8928
rect 20993 8919 21051 8925
rect 17218 8848 17224 8900
rect 17276 8888 17282 8900
rect 19981 8891 20039 8897
rect 19981 8888 19993 8891
rect 17276 8860 19993 8888
rect 17276 8848 17282 8860
rect 19981 8857 19993 8860
rect 20027 8857 20039 8891
rect 19981 8851 20039 8857
rect 21818 8848 21824 8900
rect 21876 8848 21882 8900
rect 22066 8888 22094 8928
rect 22370 8916 22376 8968
rect 22428 8956 22434 8968
rect 22649 8959 22707 8965
rect 22649 8956 22661 8959
rect 22428 8928 22661 8956
rect 22428 8916 22434 8928
rect 22649 8925 22661 8928
rect 22695 8925 22707 8959
rect 22649 8919 22707 8925
rect 24026 8916 24032 8968
rect 24084 8956 24090 8968
rect 24581 8959 24639 8965
rect 24581 8956 24593 8959
rect 24084 8928 24593 8956
rect 24084 8916 24090 8928
rect 24581 8925 24593 8928
rect 24627 8925 24639 8959
rect 24581 8919 24639 8925
rect 23474 8888 23480 8900
rect 22066 8860 23480 8888
rect 23474 8848 23480 8860
rect 23532 8848 23538 8900
rect 23845 8891 23903 8897
rect 23845 8857 23857 8891
rect 23891 8888 23903 8891
rect 24946 8888 24952 8900
rect 23891 8860 24952 8888
rect 23891 8857 23903 8860
rect 23845 8851 23903 8857
rect 24946 8848 24952 8860
rect 25004 8848 25010 8900
rect 14829 8823 14887 8829
rect 14829 8820 14841 8823
rect 14384 8792 14841 8820
rect 14829 8789 14841 8792
rect 14875 8789 14887 8823
rect 14829 8783 14887 8789
rect 15565 8823 15623 8829
rect 15565 8789 15577 8823
rect 15611 8789 15623 8823
rect 15565 8783 15623 8789
rect 15933 8823 15991 8829
rect 15933 8789 15945 8823
rect 15979 8820 15991 8823
rect 16482 8820 16488 8832
rect 15979 8792 16488 8820
rect 15979 8789 15991 8792
rect 15933 8783 15991 8789
rect 16482 8780 16488 8792
rect 16540 8780 16546 8832
rect 16853 8823 16911 8829
rect 16853 8789 16865 8823
rect 16899 8820 16911 8823
rect 17310 8820 17316 8832
rect 16899 8792 17316 8820
rect 16899 8789 16911 8792
rect 16853 8783 16911 8789
rect 17310 8780 17316 8792
rect 17368 8780 17374 8832
rect 17402 8780 17408 8832
rect 17460 8820 17466 8832
rect 17773 8823 17831 8829
rect 17773 8820 17785 8823
rect 17460 8792 17785 8820
rect 17460 8780 17466 8792
rect 17773 8789 17785 8792
rect 17819 8789 17831 8823
rect 17773 8783 17831 8789
rect 17862 8780 17868 8832
rect 17920 8820 17926 8832
rect 19058 8820 19064 8832
rect 17920 8792 19064 8820
rect 17920 8780 17926 8792
rect 19058 8780 19064 8792
rect 19116 8780 19122 8832
rect 19242 8780 19248 8832
rect 19300 8820 19306 8832
rect 19337 8823 19395 8829
rect 19337 8820 19349 8823
rect 19300 8792 19349 8820
rect 19300 8780 19306 8792
rect 19337 8789 19349 8792
rect 19383 8789 19395 8823
rect 19337 8783 19395 8789
rect 19610 8780 19616 8832
rect 19668 8780 19674 8832
rect 22646 8780 22652 8832
rect 22704 8820 22710 8832
rect 25225 8823 25283 8829
rect 25225 8820 25237 8823
rect 22704 8792 25237 8820
rect 22704 8780 22710 8792
rect 25225 8789 25237 8792
rect 25271 8789 25283 8823
rect 25225 8783 25283 8789
rect 1104 8730 25852 8752
rect 1104 8678 7950 8730
rect 8002 8678 8014 8730
rect 8066 8678 8078 8730
rect 8130 8678 8142 8730
rect 8194 8678 8206 8730
rect 8258 8678 17950 8730
rect 18002 8678 18014 8730
rect 18066 8678 18078 8730
rect 18130 8678 18142 8730
rect 18194 8678 18206 8730
rect 18258 8678 25852 8730
rect 1104 8656 25852 8678
rect 10594 8576 10600 8628
rect 10652 8616 10658 8628
rect 12069 8619 12127 8625
rect 12069 8616 12081 8619
rect 10652 8588 12081 8616
rect 10652 8576 10658 8588
rect 12069 8585 12081 8588
rect 12115 8585 12127 8619
rect 12069 8579 12127 8585
rect 12176 8588 13400 8616
rect 8846 8508 8852 8560
rect 8904 8508 8910 8560
rect 10410 8508 10416 8560
rect 10468 8548 10474 8560
rect 12176 8548 12204 8588
rect 13372 8548 13400 8588
rect 13446 8576 13452 8628
rect 13504 8616 13510 8628
rect 15565 8619 15623 8625
rect 15565 8616 15577 8619
rect 13504 8588 15577 8616
rect 13504 8576 13510 8588
rect 15565 8585 15577 8588
rect 15611 8585 15623 8619
rect 15565 8579 15623 8585
rect 15838 8576 15844 8628
rect 15896 8616 15902 8628
rect 15933 8619 15991 8625
rect 15933 8616 15945 8619
rect 15896 8588 15945 8616
rect 15896 8576 15902 8588
rect 15933 8585 15945 8588
rect 15979 8616 15991 8619
rect 17310 8616 17316 8628
rect 15979 8588 17316 8616
rect 15979 8585 15991 8588
rect 15933 8579 15991 8585
rect 17310 8576 17316 8588
rect 17368 8576 17374 8628
rect 17770 8576 17776 8628
rect 17828 8616 17834 8628
rect 17865 8619 17923 8625
rect 17865 8616 17877 8619
rect 17828 8588 17877 8616
rect 17828 8576 17834 8588
rect 17865 8585 17877 8588
rect 17911 8585 17923 8619
rect 17865 8579 17923 8585
rect 18414 8576 18420 8628
rect 18472 8616 18478 8628
rect 19242 8616 19248 8628
rect 18472 8588 19248 8616
rect 18472 8576 18478 8588
rect 19242 8576 19248 8588
rect 19300 8576 19306 8628
rect 19886 8616 19892 8628
rect 19628 8588 19892 8616
rect 16025 8551 16083 8557
rect 16025 8548 16037 8551
rect 10468 8520 12204 8548
rect 12360 8520 13308 8548
rect 13372 8520 16037 8548
rect 10468 8508 10474 8520
rect 8110 8440 8116 8492
rect 8168 8440 8174 8492
rect 9982 8452 10732 8480
rect 8294 8372 8300 8424
rect 8352 8412 8358 8424
rect 8573 8415 8631 8421
rect 8573 8412 8585 8415
rect 8352 8384 8585 8412
rect 8352 8372 8358 8384
rect 8573 8381 8585 8384
rect 8619 8381 8631 8415
rect 8573 8375 8631 8381
rect 7929 8347 7987 8353
rect 7929 8313 7941 8347
rect 7975 8344 7987 8347
rect 8478 8344 8484 8356
rect 7975 8316 8484 8344
rect 7975 8313 7987 8316
rect 7929 8307 7987 8313
rect 8478 8304 8484 8316
rect 8536 8304 8542 8356
rect 8588 8276 8616 8375
rect 10704 8353 10732 8452
rect 10965 8415 11023 8421
rect 10965 8381 10977 8415
rect 11011 8412 11023 8415
rect 11974 8412 11980 8424
rect 11011 8384 11980 8412
rect 11011 8381 11023 8384
rect 10965 8375 11023 8381
rect 11974 8372 11980 8384
rect 12032 8372 12038 8424
rect 12158 8372 12164 8424
rect 12216 8372 12222 8424
rect 12360 8421 12388 8520
rect 12802 8440 12808 8492
rect 12860 8480 12866 8492
rect 12897 8483 12955 8489
rect 12897 8480 12909 8483
rect 12860 8452 12909 8480
rect 12860 8440 12866 8452
rect 12897 8449 12909 8452
rect 12943 8449 12955 8483
rect 13280 8480 13308 8520
rect 16025 8517 16037 8520
rect 16071 8548 16083 8551
rect 18693 8551 18751 8557
rect 18693 8548 18705 8551
rect 16071 8520 18705 8548
rect 16071 8517 16083 8520
rect 16025 8511 16083 8517
rect 18693 8517 18705 8520
rect 18739 8517 18751 8551
rect 18693 8511 18751 8517
rect 18782 8508 18788 8560
rect 18840 8548 18846 8560
rect 19429 8551 19487 8557
rect 19429 8548 19441 8551
rect 18840 8520 19441 8548
rect 18840 8508 18846 8520
rect 19429 8517 19441 8520
rect 19475 8517 19487 8551
rect 19429 8511 19487 8517
rect 14090 8480 14096 8492
rect 13280 8452 14096 8480
rect 12897 8443 12955 8449
rect 14090 8440 14096 8452
rect 14148 8440 14154 8492
rect 17221 8483 17279 8489
rect 17221 8480 17233 8483
rect 14200 8452 17233 8480
rect 12345 8415 12403 8421
rect 12345 8381 12357 8415
rect 12391 8381 12403 8415
rect 12345 8375 12403 8381
rect 12618 8372 12624 8424
rect 12676 8412 12682 8424
rect 14200 8412 14228 8452
rect 17221 8449 17233 8452
rect 17267 8449 17279 8483
rect 17221 8443 17279 8449
rect 17313 8483 17371 8489
rect 17313 8449 17325 8483
rect 17359 8480 17371 8483
rect 17770 8480 17776 8492
rect 17359 8452 17776 8480
rect 17359 8449 17371 8452
rect 17313 8443 17371 8449
rect 17770 8440 17776 8452
rect 17828 8440 17834 8492
rect 19628 8480 19656 8588
rect 19886 8576 19892 8588
rect 19944 8576 19950 8628
rect 20162 8576 20168 8628
rect 20220 8616 20226 8628
rect 21821 8619 21879 8625
rect 21821 8616 21833 8619
rect 20220 8588 21833 8616
rect 20220 8576 20226 8588
rect 21821 8585 21833 8588
rect 21867 8585 21879 8619
rect 21821 8579 21879 8585
rect 22097 8619 22155 8625
rect 22097 8585 22109 8619
rect 22143 8616 22155 8619
rect 22143 8588 23980 8616
rect 22143 8585 22155 8588
rect 22097 8579 22155 8585
rect 20254 8548 20260 8560
rect 19720 8520 20260 8548
rect 19720 8492 19748 8520
rect 20254 8508 20260 8520
rect 20312 8508 20318 8560
rect 22002 8548 22008 8560
rect 21206 8520 22008 8548
rect 22002 8508 22008 8520
rect 22060 8548 22066 8560
rect 22112 8548 22140 8579
rect 22060 8520 22140 8548
rect 22060 8508 22066 8520
rect 22646 8508 22652 8560
rect 22704 8508 22710 8560
rect 23952 8548 23980 8588
rect 24026 8548 24032 8560
rect 23874 8520 24032 8548
rect 24026 8508 24032 8520
rect 24084 8508 24090 8560
rect 18248 8452 19656 8480
rect 12676 8384 14228 8412
rect 12676 8372 12682 8384
rect 14274 8372 14280 8424
rect 14332 8372 14338 8424
rect 14553 8415 14611 8421
rect 14553 8381 14565 8415
rect 14599 8412 14611 8415
rect 15102 8412 15108 8424
rect 14599 8384 15108 8412
rect 14599 8381 14611 8384
rect 14553 8375 14611 8381
rect 15102 8372 15108 8384
rect 15160 8372 15166 8424
rect 16209 8415 16267 8421
rect 16209 8381 16221 8415
rect 16255 8412 16267 8415
rect 16390 8412 16396 8424
rect 16255 8384 16396 8412
rect 16255 8381 16267 8384
rect 16209 8375 16267 8381
rect 16390 8372 16396 8384
rect 16448 8372 16454 8424
rect 16482 8372 16488 8424
rect 16540 8412 16546 8424
rect 17497 8415 17555 8421
rect 16540 8384 17264 8412
rect 16540 8372 16546 8384
rect 10689 8347 10747 8353
rect 10689 8313 10701 8347
rect 10735 8344 10747 8347
rect 11054 8344 11060 8356
rect 10735 8316 11060 8344
rect 10735 8313 10747 8316
rect 10689 8307 10747 8313
rect 11054 8304 11060 8316
rect 11112 8304 11118 8356
rect 11701 8347 11759 8353
rect 11701 8313 11713 8347
rect 11747 8344 11759 8347
rect 16758 8344 16764 8356
rect 11747 8316 16764 8344
rect 11747 8313 11759 8316
rect 11701 8307 11759 8313
rect 16758 8304 16764 8316
rect 16816 8304 16822 8356
rect 17236 8344 17264 8384
rect 17497 8381 17509 8415
rect 17543 8412 17555 8415
rect 17586 8412 17592 8424
rect 17543 8384 17592 8412
rect 17543 8381 17555 8384
rect 17497 8375 17555 8381
rect 17586 8372 17592 8384
rect 17644 8372 17650 8424
rect 18248 8344 18276 8452
rect 19702 8440 19708 8492
rect 19760 8440 19766 8492
rect 24581 8483 24639 8489
rect 24581 8480 24593 8483
rect 24136 8452 24593 8480
rect 18782 8372 18788 8424
rect 18840 8372 18846 8424
rect 18969 8415 19027 8421
rect 18969 8381 18981 8415
rect 19015 8412 19027 8415
rect 19981 8415 20039 8421
rect 19015 8384 19840 8412
rect 19015 8381 19027 8384
rect 18969 8375 19027 8381
rect 17236 8316 18276 8344
rect 18325 8347 18383 8353
rect 18325 8313 18337 8347
rect 18371 8344 18383 8347
rect 19242 8344 19248 8356
rect 18371 8316 19248 8344
rect 18371 8313 18383 8316
rect 18325 8307 18383 8313
rect 19242 8304 19248 8316
rect 19300 8304 19306 8356
rect 9030 8276 9036 8288
rect 8588 8248 9036 8276
rect 9030 8236 9036 8248
rect 9088 8236 9094 8288
rect 10318 8236 10324 8288
rect 10376 8236 10382 8288
rect 13538 8236 13544 8288
rect 13596 8236 13602 8288
rect 13814 8236 13820 8288
rect 13872 8236 13878 8288
rect 16853 8279 16911 8285
rect 16853 8245 16865 8279
rect 16899 8276 16911 8279
rect 17494 8276 17500 8288
rect 16899 8248 17500 8276
rect 16899 8245 16911 8248
rect 16853 8239 16911 8245
rect 17494 8236 17500 8248
rect 17552 8236 17558 8288
rect 19812 8276 19840 8384
rect 19981 8381 19993 8415
rect 20027 8412 20039 8415
rect 22186 8412 22192 8424
rect 20027 8384 22192 8412
rect 20027 8381 20039 8384
rect 19981 8375 20039 8381
rect 22186 8372 22192 8384
rect 22244 8372 22250 8424
rect 22278 8372 22284 8424
rect 22336 8412 22342 8424
rect 22373 8415 22431 8421
rect 22373 8412 22385 8415
rect 22336 8384 22385 8412
rect 22336 8372 22342 8384
rect 22373 8381 22385 8384
rect 22419 8381 22431 8415
rect 22738 8412 22744 8424
rect 22373 8375 22431 8381
rect 22480 8384 22744 8412
rect 22480 8344 22508 8384
rect 22738 8372 22744 8384
rect 22796 8372 22802 8424
rect 24136 8421 24164 8452
rect 24581 8449 24593 8452
rect 24627 8480 24639 8483
rect 24854 8480 24860 8492
rect 24627 8452 24860 8480
rect 24627 8449 24639 8452
rect 24581 8443 24639 8449
rect 24854 8440 24860 8452
rect 24912 8440 24918 8492
rect 24121 8415 24179 8421
rect 24121 8381 24133 8415
rect 24167 8381 24179 8415
rect 24121 8375 24179 8381
rect 21008 8316 22508 8344
rect 21008 8276 21036 8316
rect 19812 8248 21036 8276
rect 21450 8236 21456 8288
rect 21508 8236 21514 8288
rect 22186 8236 22192 8288
rect 22244 8276 22250 8288
rect 23382 8276 23388 8288
rect 22244 8248 23388 8276
rect 22244 8236 22250 8248
rect 23382 8236 23388 8248
rect 23440 8236 23446 8288
rect 25222 8236 25228 8288
rect 25280 8236 25286 8288
rect 1104 8186 25852 8208
rect 1104 8134 2950 8186
rect 3002 8134 3014 8186
rect 3066 8134 3078 8186
rect 3130 8134 3142 8186
rect 3194 8134 3206 8186
rect 3258 8134 12950 8186
rect 13002 8134 13014 8186
rect 13066 8134 13078 8186
rect 13130 8134 13142 8186
rect 13194 8134 13206 8186
rect 13258 8134 22950 8186
rect 23002 8134 23014 8186
rect 23066 8134 23078 8186
rect 23130 8134 23142 8186
rect 23194 8134 23206 8186
rect 23258 8134 25852 8186
rect 1104 8112 25852 8134
rect 10318 8032 10324 8084
rect 10376 8072 10382 8084
rect 10376 8044 10824 8072
rect 10376 8032 10382 8044
rect 10413 8007 10471 8013
rect 10413 7973 10425 8007
rect 10459 7973 10471 8007
rect 10413 7967 10471 7973
rect 9309 7871 9367 7877
rect 9309 7837 9321 7871
rect 9355 7868 9367 7871
rect 10318 7868 10324 7880
rect 9355 7840 10324 7868
rect 9355 7837 9367 7840
rect 9309 7831 9367 7837
rect 10318 7828 10324 7840
rect 10376 7828 10382 7880
rect 8386 7760 8392 7812
rect 8444 7800 8450 7812
rect 10428 7800 10456 7967
rect 10796 7868 10824 8044
rect 10870 8032 10876 8084
rect 10928 8072 10934 8084
rect 10928 8044 11652 8072
rect 10928 8032 10934 8044
rect 10888 7976 11560 8004
rect 10888 7945 10916 7976
rect 11532 7948 11560 7976
rect 10873 7939 10931 7945
rect 10873 7905 10885 7939
rect 10919 7905 10931 7939
rect 10873 7899 10931 7905
rect 10965 7939 11023 7945
rect 10965 7905 10977 7939
rect 11011 7905 11023 7939
rect 10965 7899 11023 7905
rect 10980 7868 11008 7899
rect 11514 7896 11520 7948
rect 11572 7896 11578 7948
rect 11624 7936 11652 8044
rect 11790 8032 11796 8084
rect 11848 8032 11854 8084
rect 14540 8075 14598 8081
rect 14540 8041 14552 8075
rect 14586 8072 14598 8075
rect 16666 8072 16672 8084
rect 14586 8044 16672 8072
rect 14586 8041 14598 8044
rect 14540 8035 14598 8041
rect 16666 8032 16672 8044
rect 16724 8032 16730 8084
rect 17236 8044 18460 8072
rect 15562 7964 15568 8016
rect 15620 8004 15626 8016
rect 17236 8004 17264 8044
rect 15620 7976 17264 8004
rect 18432 8004 18460 8044
rect 18874 8032 18880 8084
rect 18932 8032 18938 8084
rect 20162 8032 20168 8084
rect 20220 8072 20226 8084
rect 20530 8072 20536 8084
rect 20220 8044 20536 8072
rect 20220 8032 20226 8044
rect 20530 8032 20536 8044
rect 20588 8032 20594 8084
rect 21082 8032 21088 8084
rect 21140 8072 21146 8084
rect 21542 8072 21548 8084
rect 21140 8044 21548 8072
rect 21140 8032 21146 8044
rect 21542 8032 21548 8044
rect 21600 8072 21606 8084
rect 21600 8044 23336 8072
rect 21600 8032 21606 8044
rect 21726 8004 21732 8016
rect 18432 7976 21732 8004
rect 15620 7964 15626 7976
rect 21726 7964 21732 7976
rect 21784 7964 21790 8016
rect 23198 8004 23204 8016
rect 21836 7976 23204 8004
rect 12345 7939 12403 7945
rect 12345 7936 12357 7939
rect 11624 7908 12357 7936
rect 12345 7905 12357 7908
rect 12391 7905 12403 7939
rect 12345 7899 12403 7905
rect 12802 7896 12808 7948
rect 12860 7936 12866 7948
rect 13541 7939 13599 7945
rect 13541 7936 13553 7939
rect 12860 7908 13553 7936
rect 12860 7896 12866 7908
rect 13541 7905 13553 7908
rect 13587 7905 13599 7939
rect 13541 7899 13599 7905
rect 14277 7939 14335 7945
rect 14277 7905 14289 7939
rect 14323 7936 14335 7939
rect 15010 7936 15016 7948
rect 14323 7908 15016 7936
rect 14323 7905 14335 7908
rect 14277 7899 14335 7905
rect 15010 7896 15016 7908
rect 15068 7936 15074 7948
rect 16850 7936 16856 7948
rect 15068 7908 16856 7936
rect 15068 7896 15074 7908
rect 16850 7896 16856 7908
rect 16908 7936 16914 7948
rect 17129 7939 17187 7945
rect 17129 7936 17141 7939
rect 16908 7908 17141 7936
rect 16908 7896 16914 7908
rect 17129 7905 17141 7908
rect 17175 7905 17187 7939
rect 17129 7899 17187 7905
rect 17402 7896 17408 7948
rect 17460 7896 17466 7948
rect 18414 7896 18420 7948
rect 18472 7936 18478 7948
rect 19981 7939 20039 7945
rect 19981 7936 19993 7939
rect 18472 7908 19993 7936
rect 18472 7896 18478 7908
rect 19981 7905 19993 7908
rect 20027 7905 20039 7939
rect 19981 7899 20039 7905
rect 10796 7840 11008 7868
rect 11974 7828 11980 7880
rect 12032 7868 12038 7880
rect 12161 7871 12219 7877
rect 12161 7868 12173 7871
rect 12032 7840 12173 7868
rect 12032 7828 12038 7840
rect 12161 7837 12173 7840
rect 12207 7837 12219 7871
rect 12161 7831 12219 7837
rect 13354 7828 13360 7880
rect 13412 7828 13418 7880
rect 16666 7828 16672 7880
rect 16724 7828 16730 7880
rect 18690 7828 18696 7880
rect 18748 7868 18754 7880
rect 19521 7871 19579 7877
rect 19521 7868 19533 7871
rect 18748 7840 19533 7868
rect 18748 7828 18754 7840
rect 19521 7837 19533 7840
rect 19567 7837 19579 7871
rect 19521 7831 19579 7837
rect 20533 7871 20591 7877
rect 20533 7837 20545 7871
rect 20579 7868 20591 7871
rect 21836 7868 21864 7976
rect 23198 7964 23204 7976
rect 23256 7964 23262 8016
rect 22554 7896 22560 7948
rect 22612 7936 22618 7948
rect 22649 7939 22707 7945
rect 22649 7936 22661 7939
rect 22612 7908 22661 7936
rect 22612 7896 22618 7908
rect 22649 7905 22661 7908
rect 22695 7905 22707 7939
rect 22649 7899 22707 7905
rect 20579 7840 21864 7868
rect 20579 7837 20591 7840
rect 20533 7831 20591 7837
rect 22186 7828 22192 7880
rect 22244 7828 22250 7880
rect 23308 7868 23336 8044
rect 24581 7871 24639 7877
rect 24581 7868 24593 7871
rect 23308 7840 24593 7868
rect 24581 7837 24593 7840
rect 24627 7837 24639 7871
rect 24581 7831 24639 7837
rect 12253 7803 12311 7809
rect 12253 7800 12265 7803
rect 8444 7772 10088 7800
rect 10428 7772 12265 7800
rect 8444 7760 8450 7772
rect 9306 7692 9312 7744
rect 9364 7732 9370 7744
rect 9953 7735 10011 7741
rect 9953 7732 9965 7735
rect 9364 7704 9965 7732
rect 9364 7692 9370 7704
rect 9953 7701 9965 7704
rect 9999 7701 10011 7735
rect 10060 7732 10088 7772
rect 12253 7769 12265 7772
rect 12299 7769 12311 7803
rect 12253 7763 12311 7769
rect 12342 7760 12348 7812
rect 12400 7800 12406 7812
rect 13449 7803 13507 7809
rect 13449 7800 13461 7803
rect 12400 7772 13461 7800
rect 12400 7760 12406 7772
rect 13449 7769 13461 7772
rect 13495 7769 13507 7803
rect 13449 7763 13507 7769
rect 13814 7760 13820 7812
rect 13872 7800 13878 7812
rect 15010 7800 15016 7812
rect 13872 7772 15016 7800
rect 13872 7760 13878 7772
rect 15010 7760 15016 7772
rect 15068 7760 15074 7812
rect 18414 7760 18420 7812
rect 18472 7760 18478 7812
rect 19705 7803 19763 7809
rect 19705 7769 19717 7803
rect 19751 7800 19763 7803
rect 21545 7803 21603 7809
rect 19751 7772 20852 7800
rect 19751 7769 19763 7772
rect 19705 7763 19763 7769
rect 10781 7735 10839 7741
rect 10781 7732 10793 7735
rect 10060 7704 10793 7732
rect 9953 7695 10011 7701
rect 10781 7701 10793 7704
rect 10827 7701 10839 7735
rect 10781 7695 10839 7701
rect 12989 7735 13047 7741
rect 12989 7701 13001 7735
rect 13035 7732 13047 7735
rect 15562 7732 15568 7744
rect 13035 7704 15568 7732
rect 13035 7701 13047 7704
rect 12989 7695 13047 7701
rect 15562 7692 15568 7704
rect 15620 7692 15626 7744
rect 16022 7692 16028 7744
rect 16080 7692 16086 7744
rect 16485 7735 16543 7741
rect 16485 7701 16497 7735
rect 16531 7732 16543 7735
rect 18782 7732 18788 7744
rect 16531 7704 18788 7732
rect 16531 7701 16543 7704
rect 16485 7695 16543 7701
rect 18782 7692 18788 7704
rect 18840 7692 18846 7744
rect 20824 7732 20852 7772
rect 21545 7769 21557 7803
rect 21591 7800 21603 7803
rect 21591 7772 22968 7800
rect 21591 7769 21603 7772
rect 21545 7763 21603 7769
rect 22830 7732 22836 7744
rect 20824 7704 22836 7732
rect 22830 7692 22836 7704
rect 22888 7692 22894 7744
rect 22940 7732 22968 7772
rect 23382 7760 23388 7812
rect 23440 7800 23446 7812
rect 25225 7803 25283 7809
rect 25225 7800 25237 7803
rect 23440 7772 25237 7800
rect 23440 7760 23446 7772
rect 25225 7769 25237 7772
rect 25271 7769 25283 7803
rect 25225 7763 25283 7769
rect 23566 7732 23572 7744
rect 22940 7704 23572 7732
rect 23566 7692 23572 7704
rect 23624 7692 23630 7744
rect 24026 7692 24032 7744
rect 24084 7732 24090 7744
rect 24121 7735 24179 7741
rect 24121 7732 24133 7735
rect 24084 7704 24133 7732
rect 24084 7692 24090 7704
rect 24121 7701 24133 7704
rect 24167 7701 24179 7735
rect 24121 7695 24179 7701
rect 1104 7642 25852 7664
rect 1104 7590 7950 7642
rect 8002 7590 8014 7642
rect 8066 7590 8078 7642
rect 8130 7590 8142 7642
rect 8194 7590 8206 7642
rect 8258 7590 17950 7642
rect 18002 7590 18014 7642
rect 18066 7590 18078 7642
rect 18130 7590 18142 7642
rect 18194 7590 18206 7642
rect 18258 7590 25852 7642
rect 1104 7568 25852 7590
rect 10781 7531 10839 7537
rect 10781 7497 10793 7531
rect 10827 7528 10839 7531
rect 10870 7528 10876 7540
rect 10827 7500 10876 7528
rect 10827 7497 10839 7500
rect 10781 7491 10839 7497
rect 10870 7488 10876 7500
rect 10928 7488 10934 7540
rect 11701 7531 11759 7537
rect 11701 7497 11713 7531
rect 11747 7528 11759 7531
rect 12342 7528 12348 7540
rect 11747 7500 12348 7528
rect 11747 7497 11759 7500
rect 11701 7491 11759 7497
rect 12342 7488 12348 7500
rect 12400 7488 12406 7540
rect 12710 7488 12716 7540
rect 12768 7528 12774 7540
rect 15381 7531 15439 7537
rect 15381 7528 15393 7531
rect 12768 7500 15393 7528
rect 12768 7488 12774 7500
rect 15381 7497 15393 7500
rect 15427 7497 15439 7531
rect 15381 7491 15439 7497
rect 15470 7488 15476 7540
rect 15528 7528 15534 7540
rect 16301 7531 16359 7537
rect 16301 7528 16313 7531
rect 15528 7500 16313 7528
rect 15528 7488 15534 7500
rect 16301 7497 16313 7500
rect 16347 7528 16359 7531
rect 16390 7528 16396 7540
rect 16347 7500 16396 7528
rect 16347 7497 16359 7500
rect 16301 7491 16359 7497
rect 16390 7488 16396 7500
rect 16448 7488 16454 7540
rect 17494 7488 17500 7540
rect 17552 7488 17558 7540
rect 17770 7488 17776 7540
rect 17828 7528 17834 7540
rect 21910 7528 21916 7540
rect 17828 7500 21916 7528
rect 17828 7488 17834 7500
rect 21910 7488 21916 7500
rect 21968 7488 21974 7540
rect 23198 7488 23204 7540
rect 23256 7528 23262 7540
rect 24946 7528 24952 7540
rect 23256 7500 24952 7528
rect 23256 7488 23262 7500
rect 24946 7488 24952 7500
rect 25004 7488 25010 7540
rect 9306 7420 9312 7472
rect 9364 7420 9370 7472
rect 15102 7420 15108 7472
rect 15160 7460 15166 7472
rect 15160 7432 22140 7460
rect 15160 7420 15166 7432
rect 11054 7392 11060 7404
rect 10442 7364 11060 7392
rect 11054 7352 11060 7364
rect 11112 7392 11118 7404
rect 11112 7364 11192 7392
rect 11112 7352 11118 7364
rect 9030 7284 9036 7336
rect 9088 7284 9094 7336
rect 11164 7197 11192 7364
rect 12066 7352 12072 7404
rect 12124 7352 12130 7404
rect 13449 7395 13507 7401
rect 13449 7361 13461 7395
rect 13495 7392 13507 7395
rect 14277 7395 14335 7401
rect 14277 7392 14289 7395
rect 13495 7364 14289 7392
rect 13495 7361 13507 7364
rect 13449 7355 13507 7361
rect 14277 7361 14289 7364
rect 14323 7361 14335 7395
rect 14277 7355 14335 7361
rect 17405 7395 17463 7401
rect 17405 7361 17417 7395
rect 17451 7392 17463 7395
rect 18138 7392 18144 7404
rect 17451 7364 18144 7392
rect 17451 7361 17463 7364
rect 17405 7355 17463 7361
rect 18138 7352 18144 7364
rect 18196 7352 18202 7404
rect 18233 7395 18291 7401
rect 18233 7361 18245 7395
rect 18279 7361 18291 7395
rect 18233 7355 18291 7361
rect 12161 7327 12219 7333
rect 12161 7293 12173 7327
rect 12207 7293 12219 7327
rect 12161 7287 12219 7293
rect 12176 7256 12204 7287
rect 12250 7284 12256 7336
rect 12308 7284 12314 7336
rect 12342 7284 12348 7336
rect 12400 7324 12406 7336
rect 13541 7327 13599 7333
rect 13541 7324 13553 7327
rect 12400 7296 13553 7324
rect 12400 7284 12406 7296
rect 13541 7293 13553 7296
rect 13587 7293 13599 7327
rect 13541 7287 13599 7293
rect 13630 7284 13636 7336
rect 13688 7284 13694 7336
rect 15562 7284 15568 7336
rect 15620 7284 15626 7336
rect 16942 7284 16948 7336
rect 17000 7324 17006 7336
rect 17310 7324 17316 7336
rect 17000 7296 17316 7324
rect 17000 7284 17006 7296
rect 17310 7284 17316 7296
rect 17368 7284 17374 7336
rect 17678 7284 17684 7336
rect 17736 7284 17742 7336
rect 12805 7259 12863 7265
rect 12805 7256 12817 7259
rect 12176 7228 12817 7256
rect 12805 7225 12817 7228
rect 12851 7256 12863 7259
rect 13354 7256 13360 7268
rect 12851 7228 13360 7256
rect 12851 7225 12863 7228
rect 12805 7219 12863 7225
rect 13354 7216 13360 7228
rect 13412 7216 13418 7268
rect 13446 7216 13452 7268
rect 13504 7256 13510 7268
rect 18248 7256 18276 7355
rect 18782 7352 18788 7404
rect 18840 7392 18846 7404
rect 22112 7401 22140 7432
rect 25130 7420 25136 7472
rect 25188 7420 25194 7472
rect 20073 7395 20131 7401
rect 20073 7392 20085 7395
rect 18840 7364 20085 7392
rect 18840 7352 18846 7364
rect 20073 7361 20085 7364
rect 20119 7361 20131 7395
rect 20073 7355 20131 7361
rect 22097 7395 22155 7401
rect 22097 7361 22109 7395
rect 22143 7361 22155 7395
rect 22097 7355 22155 7361
rect 22462 7352 22468 7404
rect 22520 7392 22526 7404
rect 23937 7395 23995 7401
rect 23937 7392 23949 7395
rect 22520 7364 23949 7392
rect 22520 7352 22526 7364
rect 23937 7361 23949 7364
rect 23983 7361 23995 7395
rect 23937 7355 23995 7361
rect 19429 7327 19487 7333
rect 19429 7293 19441 7327
rect 19475 7293 19487 7327
rect 19429 7287 19487 7293
rect 21269 7327 21327 7333
rect 21269 7293 21281 7327
rect 21315 7324 21327 7327
rect 21910 7324 21916 7336
rect 21315 7296 21916 7324
rect 21315 7293 21327 7296
rect 21269 7287 21327 7293
rect 13504 7228 18276 7256
rect 19444 7256 19472 7287
rect 21910 7284 21916 7296
rect 21968 7284 21974 7336
rect 23290 7284 23296 7336
rect 23348 7284 23354 7336
rect 22002 7256 22008 7268
rect 19444 7228 22008 7256
rect 13504 7216 13510 7228
rect 22002 7216 22008 7228
rect 22060 7216 22066 7268
rect 11149 7191 11207 7197
rect 11149 7157 11161 7191
rect 11195 7188 11207 7191
rect 11974 7188 11980 7200
rect 11195 7160 11980 7188
rect 11195 7157 11207 7160
rect 11149 7151 11207 7157
rect 11974 7148 11980 7160
rect 12032 7148 12038 7200
rect 13081 7191 13139 7197
rect 13081 7157 13093 7191
rect 13127 7188 13139 7191
rect 13998 7188 14004 7200
rect 13127 7160 14004 7188
rect 13127 7157 13139 7160
rect 13081 7151 13139 7157
rect 13998 7148 14004 7160
rect 14056 7148 14062 7200
rect 15010 7148 15016 7200
rect 15068 7148 15074 7200
rect 15194 7148 15200 7200
rect 15252 7188 15258 7200
rect 16114 7188 16120 7200
rect 15252 7160 16120 7188
rect 15252 7148 15258 7160
rect 16114 7148 16120 7160
rect 16172 7148 16178 7200
rect 16390 7148 16396 7200
rect 16448 7188 16454 7200
rect 17037 7191 17095 7197
rect 17037 7188 17049 7191
rect 16448 7160 17049 7188
rect 16448 7148 16454 7160
rect 17037 7157 17049 7160
rect 17083 7157 17095 7191
rect 17037 7151 17095 7157
rect 18138 7148 18144 7200
rect 18196 7188 18202 7200
rect 21266 7188 21272 7200
rect 18196 7160 21272 7188
rect 18196 7148 18202 7160
rect 21266 7148 21272 7160
rect 21324 7148 21330 7200
rect 22094 7148 22100 7200
rect 22152 7188 22158 7200
rect 23750 7188 23756 7200
rect 22152 7160 23756 7188
rect 22152 7148 22158 7160
rect 23750 7148 23756 7160
rect 23808 7148 23814 7200
rect 1104 7098 25852 7120
rect 1104 7046 2950 7098
rect 3002 7046 3014 7098
rect 3066 7046 3078 7098
rect 3130 7046 3142 7098
rect 3194 7046 3206 7098
rect 3258 7046 12950 7098
rect 13002 7046 13014 7098
rect 13066 7046 13078 7098
rect 13130 7046 13142 7098
rect 13194 7046 13206 7098
rect 13258 7046 22950 7098
rect 23002 7046 23014 7098
rect 23066 7046 23078 7098
rect 23130 7046 23142 7098
rect 23194 7046 23206 7098
rect 23258 7046 25852 7098
rect 1104 7024 25852 7046
rect 9306 6944 9312 6996
rect 9364 6984 9370 6996
rect 12345 6987 12403 6993
rect 9364 6956 11928 6984
rect 9364 6944 9370 6956
rect 11900 6916 11928 6956
rect 12345 6953 12357 6987
rect 12391 6984 12403 6987
rect 12802 6984 12808 6996
rect 12391 6956 12808 6984
rect 12391 6953 12403 6956
rect 12345 6947 12403 6953
rect 12802 6944 12808 6956
rect 12860 6944 12866 6996
rect 15194 6944 15200 6996
rect 15252 6944 15258 6996
rect 17862 6984 17868 6996
rect 15304 6956 17868 6984
rect 12710 6916 12716 6928
rect 11900 6888 12716 6916
rect 12710 6876 12716 6888
rect 12768 6876 12774 6928
rect 13354 6876 13360 6928
rect 13412 6916 13418 6928
rect 15304 6916 15332 6956
rect 17862 6944 17868 6956
rect 17920 6944 17926 6996
rect 20060 6987 20118 6993
rect 20060 6953 20072 6987
rect 20106 6984 20118 6987
rect 22094 6984 22100 6996
rect 20106 6956 22100 6984
rect 20106 6953 20118 6956
rect 20060 6947 20118 6953
rect 22094 6944 22100 6956
rect 22152 6944 22158 6996
rect 22268 6987 22326 6993
rect 22268 6953 22280 6987
rect 22314 6984 22326 6987
rect 25222 6984 25228 6996
rect 22314 6956 25228 6984
rect 22314 6953 22326 6956
rect 22268 6947 22326 6953
rect 25222 6944 25228 6956
rect 25280 6944 25286 6996
rect 13412 6888 15332 6916
rect 13412 6876 13418 6888
rect 15838 6876 15844 6928
rect 15896 6916 15902 6928
rect 17770 6916 17776 6928
rect 15896 6888 17776 6916
rect 15896 6876 15902 6888
rect 17770 6876 17776 6888
rect 17828 6876 17834 6928
rect 21542 6876 21548 6928
rect 21600 6876 21606 6928
rect 23382 6876 23388 6928
rect 23440 6876 23446 6928
rect 24854 6876 24860 6928
rect 24912 6916 24918 6928
rect 24912 6888 25176 6916
rect 24912 6876 24918 6888
rect 5258 6808 5264 6860
rect 5316 6848 5322 6860
rect 10042 6848 10048 6860
rect 5316 6820 10048 6848
rect 5316 6808 5322 6820
rect 10042 6808 10048 6820
rect 10100 6808 10106 6860
rect 10597 6851 10655 6857
rect 10597 6817 10609 6851
rect 10643 6848 10655 6851
rect 11606 6848 11612 6860
rect 10643 6820 11612 6848
rect 10643 6817 10655 6820
rect 10597 6811 10655 6817
rect 11606 6808 11612 6820
rect 11664 6808 11670 6860
rect 12434 6808 12440 6860
rect 12492 6848 12498 6860
rect 12621 6851 12679 6857
rect 12621 6848 12633 6851
rect 12492 6820 12633 6848
rect 12492 6808 12498 6820
rect 12621 6817 12633 6820
rect 12667 6848 12679 6851
rect 13449 6851 13507 6857
rect 13449 6848 13461 6851
rect 12667 6820 13461 6848
rect 12667 6817 12679 6820
rect 12621 6811 12679 6817
rect 13449 6817 13461 6820
rect 13495 6817 13507 6851
rect 13449 6811 13507 6817
rect 13633 6851 13691 6857
rect 13633 6817 13645 6851
rect 13679 6848 13691 6851
rect 16022 6848 16028 6860
rect 13679 6820 16028 6848
rect 13679 6817 13691 6820
rect 13633 6811 13691 6817
rect 11974 6740 11980 6792
rect 12032 6740 12038 6792
rect 14292 6789 14320 6820
rect 16022 6808 16028 6820
rect 16080 6808 16086 6860
rect 16942 6808 16948 6860
rect 17000 6808 17006 6860
rect 19702 6808 19708 6860
rect 19760 6848 19766 6860
rect 19797 6851 19855 6857
rect 19797 6848 19809 6851
rect 19760 6820 19809 6848
rect 19760 6808 19766 6820
rect 19797 6817 19809 6820
rect 19843 6848 19855 6851
rect 22005 6851 22063 6857
rect 22005 6848 22017 6851
rect 19843 6820 22017 6848
rect 19843 6817 19855 6820
rect 19797 6811 19855 6817
rect 22005 6817 22017 6820
rect 22051 6848 22063 6851
rect 22278 6848 22284 6860
rect 22051 6820 22284 6848
rect 22051 6817 22063 6820
rect 22005 6811 22063 6817
rect 22278 6808 22284 6820
rect 22336 6808 22342 6860
rect 22738 6808 22744 6860
rect 22796 6848 22802 6860
rect 23400 6848 23428 6876
rect 23753 6851 23811 6857
rect 23753 6848 23765 6851
rect 22796 6820 23765 6848
rect 22796 6808 22802 6820
rect 23753 6817 23765 6820
rect 23799 6817 23811 6851
rect 23753 6811 23811 6817
rect 25038 6808 25044 6860
rect 25096 6808 25102 6860
rect 25148 6857 25176 6888
rect 25133 6851 25191 6857
rect 25133 6817 25145 6851
rect 25179 6817 25191 6851
rect 25133 6811 25191 6817
rect 14277 6783 14335 6789
rect 14277 6749 14289 6783
rect 14323 6749 14335 6783
rect 14277 6743 14335 6749
rect 15010 6740 15016 6792
rect 15068 6780 15074 6792
rect 16669 6783 16727 6789
rect 15068 6752 16160 6780
rect 15068 6740 15074 6752
rect 10873 6715 10931 6721
rect 10873 6681 10885 6715
rect 10919 6712 10931 6715
rect 11146 6712 11152 6724
rect 10919 6684 11152 6712
rect 10919 6681 10931 6684
rect 10873 6675 10931 6681
rect 11146 6672 11152 6684
rect 11204 6672 11210 6724
rect 15654 6672 15660 6724
rect 15712 6672 15718 6724
rect 15841 6715 15899 6721
rect 15841 6681 15853 6715
rect 15887 6712 15899 6715
rect 16022 6712 16028 6724
rect 15887 6684 16028 6712
rect 15887 6681 15899 6684
rect 15841 6675 15899 6681
rect 16022 6672 16028 6684
rect 16080 6672 16086 6724
rect 16132 6712 16160 6752
rect 16669 6749 16681 6783
rect 16715 6780 16727 6783
rect 16758 6780 16764 6792
rect 16715 6752 16764 6780
rect 16715 6749 16727 6752
rect 16669 6743 16727 6749
rect 16758 6740 16764 6752
rect 16816 6740 16822 6792
rect 17126 6740 17132 6792
rect 17184 6780 17190 6792
rect 17497 6783 17555 6789
rect 17497 6780 17509 6783
rect 17184 6752 17509 6780
rect 17184 6740 17190 6752
rect 17497 6749 17509 6752
rect 17543 6749 17555 6783
rect 17497 6743 17555 6749
rect 18693 6715 18751 6721
rect 16132 6684 16804 6712
rect 2038 6604 2044 6656
rect 2096 6644 2102 6656
rect 8754 6644 8760 6656
rect 2096 6616 8760 6644
rect 2096 6604 2102 6616
rect 8754 6604 8760 6616
rect 8812 6604 8818 6656
rect 12986 6604 12992 6656
rect 13044 6604 13050 6656
rect 13354 6604 13360 6656
rect 13412 6604 13418 6656
rect 13538 6604 13544 6656
rect 13596 6644 13602 6656
rect 14921 6647 14979 6653
rect 14921 6644 14933 6647
rect 13596 6616 14933 6644
rect 13596 6604 13602 6616
rect 14921 6613 14933 6616
rect 14967 6613 14979 6647
rect 14921 6607 14979 6613
rect 15286 6604 15292 6656
rect 15344 6644 15350 6656
rect 16776 6653 16804 6684
rect 18693 6681 18705 6715
rect 18739 6712 18751 6715
rect 18966 6712 18972 6724
rect 18739 6684 18972 6712
rect 18739 6681 18751 6684
rect 18693 6675 18751 6681
rect 18966 6672 18972 6684
rect 19024 6672 19030 6724
rect 19978 6672 19984 6724
rect 20036 6712 20042 6724
rect 20036 6684 20562 6712
rect 23506 6684 24072 6712
rect 20036 6672 20042 6684
rect 24044 6656 24072 6684
rect 16301 6647 16359 6653
rect 16301 6644 16313 6647
rect 15344 6616 16313 6644
rect 15344 6604 15350 6616
rect 16301 6613 16313 6616
rect 16347 6613 16359 6647
rect 16301 6607 16359 6613
rect 16761 6647 16819 6653
rect 16761 6613 16773 6647
rect 16807 6613 16819 6647
rect 16761 6607 16819 6613
rect 24026 6604 24032 6656
rect 24084 6604 24090 6656
rect 24578 6604 24584 6656
rect 24636 6604 24642 6656
rect 24946 6604 24952 6656
rect 25004 6604 25010 6656
rect 1104 6554 25852 6576
rect 1104 6502 7950 6554
rect 8002 6502 8014 6554
rect 8066 6502 8078 6554
rect 8130 6502 8142 6554
rect 8194 6502 8206 6554
rect 8258 6502 17950 6554
rect 18002 6502 18014 6554
rect 18066 6502 18078 6554
rect 18130 6502 18142 6554
rect 18194 6502 18206 6554
rect 18258 6502 25852 6554
rect 1104 6480 25852 6502
rect 11146 6400 11152 6452
rect 11204 6440 11210 6452
rect 12345 6443 12403 6449
rect 12345 6440 12357 6443
rect 11204 6412 12357 6440
rect 11204 6400 11210 6412
rect 12345 6409 12357 6412
rect 12391 6409 12403 6443
rect 12345 6403 12403 6409
rect 12986 6400 12992 6452
rect 13044 6440 13050 6452
rect 15565 6443 15623 6449
rect 13044 6412 14596 6440
rect 13044 6400 13050 6412
rect 13265 6375 13323 6381
rect 13265 6341 13277 6375
rect 13311 6372 13323 6375
rect 13538 6372 13544 6384
rect 13311 6344 13544 6372
rect 13311 6341 13323 6344
rect 13265 6335 13323 6341
rect 13538 6332 13544 6344
rect 13596 6332 13602 6384
rect 13814 6332 13820 6384
rect 13872 6332 13878 6384
rect 14568 6372 14596 6412
rect 15565 6409 15577 6443
rect 15611 6440 15623 6443
rect 19061 6443 19119 6449
rect 19061 6440 19073 6443
rect 15611 6412 19073 6440
rect 15611 6409 15623 6412
rect 15565 6403 15623 6409
rect 19061 6409 19073 6412
rect 19107 6409 19119 6443
rect 19061 6403 19119 6409
rect 22094 6400 22100 6452
rect 22152 6440 22158 6452
rect 22278 6440 22284 6452
rect 22152 6412 22284 6440
rect 22152 6400 22158 6412
rect 22278 6400 22284 6412
rect 22336 6400 22342 6452
rect 15657 6375 15715 6381
rect 15657 6372 15669 6375
rect 14568 6344 15669 6372
rect 15657 6341 15669 6344
rect 15703 6341 15715 6375
rect 17126 6372 17132 6384
rect 15657 6335 15715 6341
rect 15764 6344 17132 6372
rect 10505 6307 10563 6313
rect 10505 6273 10517 6307
rect 10551 6304 10563 6307
rect 10870 6304 10876 6316
rect 10551 6276 10876 6304
rect 10551 6273 10563 6276
rect 10505 6267 10563 6273
rect 10870 6264 10876 6276
rect 10928 6264 10934 6316
rect 11698 6264 11704 6316
rect 11756 6304 11762 6316
rect 12250 6304 12256 6316
rect 11756 6276 12256 6304
rect 11756 6264 11762 6276
rect 12250 6264 12256 6276
rect 12308 6264 12314 6316
rect 15010 6264 15016 6316
rect 15068 6304 15074 6316
rect 15764 6304 15792 6344
rect 17126 6332 17132 6344
rect 17184 6332 17190 6384
rect 18138 6332 18144 6384
rect 18196 6332 18202 6384
rect 24854 6372 24860 6384
rect 22204 6344 24860 6372
rect 15068 6276 15792 6304
rect 15068 6264 15074 6276
rect 16114 6264 16120 6316
rect 16172 6304 16178 6316
rect 16393 6307 16451 6313
rect 16393 6304 16405 6307
rect 16172 6276 16405 6304
rect 16172 6264 16178 6276
rect 16393 6273 16405 6276
rect 16439 6273 16451 6307
rect 16393 6267 16451 6273
rect 11606 6196 11612 6248
rect 11664 6236 11670 6248
rect 12989 6239 13047 6245
rect 12989 6236 13001 6239
rect 11664 6208 13001 6236
rect 11664 6196 11670 6208
rect 12989 6205 13001 6208
rect 13035 6205 13047 6239
rect 12989 6199 13047 6205
rect 2222 6128 2228 6180
rect 2280 6168 2286 6180
rect 12158 6168 12164 6180
rect 2280 6140 12164 6168
rect 2280 6128 2286 6140
rect 12158 6128 12164 6140
rect 12216 6128 12222 6180
rect 10226 6060 10232 6112
rect 10284 6100 10290 6112
rect 11149 6103 11207 6109
rect 11149 6100 11161 6103
rect 10284 6072 11161 6100
rect 10284 6060 10290 6072
rect 11149 6069 11161 6072
rect 11195 6069 11207 6103
rect 11149 6063 11207 6069
rect 11974 6060 11980 6112
rect 12032 6100 12038 6112
rect 12621 6103 12679 6109
rect 12621 6100 12633 6103
rect 12032 6072 12633 6100
rect 12032 6060 12038 6072
rect 12621 6069 12633 6072
rect 12667 6069 12679 6103
rect 13004 6100 13032 6199
rect 13722 6196 13728 6248
rect 13780 6236 13786 6248
rect 13780 6208 14320 6236
rect 13780 6196 13786 6208
rect 13722 6100 13728 6112
rect 13004 6072 13728 6100
rect 12621 6063 12679 6069
rect 13722 6060 13728 6072
rect 13780 6060 13786 6112
rect 14292 6100 14320 6208
rect 15194 6196 15200 6248
rect 15252 6236 15258 6248
rect 15562 6236 15568 6248
rect 15252 6208 15568 6236
rect 15252 6196 15258 6208
rect 15562 6196 15568 6208
rect 15620 6196 15626 6248
rect 15749 6239 15807 6245
rect 15749 6205 15761 6239
rect 15795 6205 15807 6239
rect 15749 6199 15807 6205
rect 14366 6128 14372 6180
rect 14424 6168 14430 6180
rect 14737 6171 14795 6177
rect 14737 6168 14749 6171
rect 14424 6140 14749 6168
rect 14424 6128 14430 6140
rect 14737 6137 14749 6140
rect 14783 6168 14795 6171
rect 15764 6168 15792 6199
rect 14783 6140 15792 6168
rect 14783 6137 14795 6140
rect 14737 6131 14795 6137
rect 15197 6103 15255 6109
rect 15197 6100 15209 6103
rect 14292 6072 15209 6100
rect 15197 6069 15209 6072
rect 15243 6069 15255 6103
rect 16408 6100 16436 6267
rect 16850 6264 16856 6316
rect 16908 6264 16914 6316
rect 19334 6264 19340 6316
rect 19392 6304 19398 6316
rect 22204 6313 22232 6344
rect 24854 6332 24860 6344
rect 24912 6332 24918 6384
rect 20073 6307 20131 6313
rect 20073 6304 20085 6307
rect 19392 6276 20085 6304
rect 19392 6264 19398 6276
rect 20073 6273 20085 6276
rect 20119 6273 20131 6307
rect 20073 6267 20131 6273
rect 22189 6307 22247 6313
rect 22189 6273 22201 6307
rect 22235 6273 22247 6307
rect 22189 6267 22247 6273
rect 23934 6264 23940 6316
rect 23992 6264 23998 6316
rect 17126 6196 17132 6248
rect 17184 6196 17190 6248
rect 17678 6196 17684 6248
rect 17736 6236 17742 6248
rect 18601 6239 18659 6245
rect 18601 6236 18613 6239
rect 17736 6208 18613 6236
rect 17736 6196 17742 6208
rect 18601 6205 18613 6208
rect 18647 6205 18659 6239
rect 18601 6199 18659 6205
rect 21269 6239 21327 6245
rect 21269 6205 21281 6239
rect 21315 6236 21327 6239
rect 21315 6208 22140 6236
rect 21315 6205 21327 6208
rect 21269 6199 21327 6205
rect 22112 6180 22140 6208
rect 22462 6196 22468 6248
rect 22520 6196 22526 6248
rect 24670 6196 24676 6248
rect 24728 6196 24734 6248
rect 19610 6128 19616 6180
rect 19668 6168 19674 6180
rect 20346 6168 20352 6180
rect 19668 6140 20352 6168
rect 19668 6128 19674 6140
rect 20346 6128 20352 6140
rect 20404 6128 20410 6180
rect 22094 6128 22100 6180
rect 22152 6128 22158 6180
rect 18138 6100 18144 6112
rect 16408 6072 18144 6100
rect 15197 6063 15255 6069
rect 18138 6060 18144 6072
rect 18196 6100 18202 6112
rect 18414 6100 18420 6112
rect 18196 6072 18420 6100
rect 18196 6060 18202 6072
rect 18414 6060 18420 6072
rect 18472 6100 18478 6112
rect 19521 6103 19579 6109
rect 19521 6100 19533 6103
rect 18472 6072 19533 6100
rect 18472 6060 18478 6072
rect 19521 6069 19533 6072
rect 19567 6100 19579 6103
rect 19978 6100 19984 6112
rect 19567 6072 19984 6100
rect 19567 6069 19579 6072
rect 19521 6063 19579 6069
rect 19978 6060 19984 6072
rect 20036 6060 20042 6112
rect 1104 6010 25852 6032
rect 1104 5958 2950 6010
rect 3002 5958 3014 6010
rect 3066 5958 3078 6010
rect 3130 5958 3142 6010
rect 3194 5958 3206 6010
rect 3258 5958 12950 6010
rect 13002 5958 13014 6010
rect 13066 5958 13078 6010
rect 13130 5958 13142 6010
rect 13194 5958 13206 6010
rect 13258 5958 22950 6010
rect 23002 5958 23014 6010
rect 23066 5958 23078 6010
rect 23130 5958 23142 6010
rect 23194 5958 23206 6010
rect 23258 5958 25852 6010
rect 1104 5936 25852 5958
rect 11698 5856 11704 5908
rect 11756 5856 11762 5908
rect 13725 5899 13783 5905
rect 13725 5865 13737 5899
rect 13771 5896 13783 5899
rect 17126 5896 17132 5908
rect 13771 5868 17132 5896
rect 13771 5865 13783 5868
rect 13725 5859 13783 5865
rect 17126 5856 17132 5868
rect 17184 5856 17190 5908
rect 23934 5896 23940 5908
rect 17236 5868 23940 5896
rect 10226 5720 10232 5772
rect 10284 5720 10290 5772
rect 11238 5720 11244 5772
rect 11296 5760 11302 5772
rect 17236 5760 17264 5868
rect 23934 5856 23940 5868
rect 23992 5856 23998 5908
rect 24213 5899 24271 5905
rect 24213 5865 24225 5899
rect 24259 5896 24271 5899
rect 24946 5896 24952 5908
rect 24259 5868 24952 5896
rect 24259 5865 24271 5868
rect 24213 5859 24271 5865
rect 17402 5788 17408 5840
rect 17460 5828 17466 5840
rect 24228 5828 24256 5859
rect 24946 5856 24952 5868
rect 25004 5856 25010 5908
rect 17460 5800 24256 5828
rect 17460 5788 17466 5800
rect 11296 5732 17264 5760
rect 11296 5720 11302 5732
rect 19978 5720 19984 5772
rect 20036 5720 20042 5772
rect 20254 5720 20260 5772
rect 20312 5760 20318 5772
rect 20809 5763 20867 5769
rect 20809 5760 20821 5763
rect 20312 5732 20821 5760
rect 20312 5720 20318 5732
rect 20809 5729 20821 5732
rect 20855 5729 20867 5763
rect 20809 5723 20867 5729
rect 22646 5720 22652 5772
rect 22704 5720 22710 5772
rect 8294 5652 8300 5704
rect 8352 5692 8358 5704
rect 9030 5692 9036 5704
rect 8352 5664 9036 5692
rect 8352 5652 8358 5664
rect 9030 5652 9036 5664
rect 9088 5692 9094 5704
rect 9953 5695 10011 5701
rect 9953 5692 9965 5695
rect 9088 5664 9965 5692
rect 9088 5652 9094 5664
rect 9953 5661 9965 5664
rect 9999 5661 10011 5695
rect 9953 5655 10011 5661
rect 12529 5695 12587 5701
rect 12529 5661 12541 5695
rect 12575 5692 12587 5695
rect 12710 5692 12716 5704
rect 12575 5664 12716 5692
rect 12575 5661 12587 5664
rect 12529 5655 12587 5661
rect 12710 5652 12716 5664
rect 12768 5652 12774 5704
rect 13081 5695 13139 5701
rect 13081 5661 13093 5695
rect 13127 5661 13139 5695
rect 13081 5655 13139 5661
rect 9582 5584 9588 5636
rect 9640 5624 9646 5636
rect 13096 5624 13124 5655
rect 14366 5652 14372 5704
rect 14424 5652 14430 5704
rect 15194 5652 15200 5704
rect 15252 5692 15258 5704
rect 15657 5695 15715 5701
rect 15657 5692 15669 5695
rect 15252 5664 15669 5692
rect 15252 5652 15258 5664
rect 15657 5661 15669 5664
rect 15703 5661 15715 5695
rect 17586 5692 17592 5704
rect 15657 5655 15715 5661
rect 16776 5664 17592 5692
rect 16776 5624 16804 5664
rect 17586 5652 17592 5664
rect 17644 5652 17650 5704
rect 17681 5695 17739 5701
rect 17681 5661 17693 5695
rect 17727 5692 17739 5695
rect 20346 5692 20352 5704
rect 17727 5664 20352 5692
rect 17727 5661 17739 5664
rect 17681 5655 17739 5661
rect 20346 5652 20352 5664
rect 20404 5652 20410 5704
rect 20533 5695 20591 5701
rect 20533 5661 20545 5695
rect 20579 5661 20591 5695
rect 20533 5655 20591 5661
rect 9640 5596 10718 5624
rect 13096 5596 16804 5624
rect 16853 5627 16911 5633
rect 9640 5584 9646 5596
rect 10612 5556 10640 5596
rect 16853 5593 16865 5627
rect 16899 5624 16911 5627
rect 17218 5624 17224 5636
rect 16899 5596 17224 5624
rect 16899 5593 16911 5596
rect 16853 5587 16911 5593
rect 17218 5584 17224 5596
rect 17276 5584 17282 5636
rect 17604 5624 17632 5652
rect 17862 5624 17868 5636
rect 17604 5596 17868 5624
rect 17862 5584 17868 5596
rect 17920 5584 17926 5636
rect 18690 5584 18696 5636
rect 18748 5584 18754 5636
rect 19521 5627 19579 5633
rect 19521 5593 19533 5627
rect 19567 5593 19579 5627
rect 19521 5587 19579 5593
rect 19705 5627 19763 5633
rect 19705 5593 19717 5627
rect 19751 5624 19763 5627
rect 20438 5624 20444 5636
rect 19751 5596 20444 5624
rect 19751 5593 19763 5596
rect 19705 5587 19763 5593
rect 11974 5556 11980 5568
rect 10612 5528 11980 5556
rect 11974 5516 11980 5528
rect 12032 5516 12038 5568
rect 12342 5516 12348 5568
rect 12400 5516 12406 5568
rect 13998 5516 14004 5568
rect 14056 5556 14062 5568
rect 15013 5559 15071 5565
rect 15013 5556 15025 5559
rect 14056 5528 15025 5556
rect 14056 5516 14062 5528
rect 15013 5525 15025 5528
rect 15059 5525 15071 5559
rect 15013 5519 15071 5525
rect 15102 5516 15108 5568
rect 15160 5556 15166 5568
rect 15289 5559 15347 5565
rect 15289 5556 15301 5559
rect 15160 5528 15301 5556
rect 15160 5516 15166 5528
rect 15289 5525 15301 5528
rect 15335 5525 15347 5559
rect 15289 5519 15347 5525
rect 16298 5516 16304 5568
rect 16356 5556 16362 5568
rect 18506 5556 18512 5568
rect 16356 5528 18512 5556
rect 16356 5516 16362 5528
rect 18506 5516 18512 5528
rect 18564 5516 18570 5568
rect 19536 5556 19564 5587
rect 20438 5584 20444 5596
rect 20496 5584 20502 5636
rect 20548 5624 20576 5655
rect 22278 5652 22284 5704
rect 22336 5652 22342 5704
rect 23382 5652 23388 5704
rect 23440 5692 23446 5704
rect 24581 5695 24639 5701
rect 24581 5692 24593 5695
rect 23440 5664 24593 5692
rect 23440 5652 23446 5664
rect 24581 5661 24593 5664
rect 24627 5661 24639 5695
rect 24581 5655 24639 5661
rect 20898 5624 20904 5636
rect 20548 5596 20904 5624
rect 20898 5584 20904 5596
rect 20956 5584 20962 5636
rect 19794 5556 19800 5568
rect 19536 5528 19800 5556
rect 19794 5516 19800 5528
rect 19852 5516 19858 5568
rect 20070 5516 20076 5568
rect 20128 5556 20134 5568
rect 21542 5556 21548 5568
rect 20128 5528 21548 5556
rect 20128 5516 20134 5528
rect 21542 5516 21548 5528
rect 21600 5516 21606 5568
rect 23937 5559 23995 5565
rect 23937 5525 23949 5559
rect 23983 5556 23995 5559
rect 24026 5556 24032 5568
rect 23983 5528 24032 5556
rect 23983 5525 23995 5528
rect 23937 5519 23995 5525
rect 24026 5516 24032 5528
rect 24084 5516 24090 5568
rect 24210 5516 24216 5568
rect 24268 5556 24274 5568
rect 25225 5559 25283 5565
rect 25225 5556 25237 5559
rect 24268 5528 25237 5556
rect 24268 5516 24274 5528
rect 25225 5525 25237 5528
rect 25271 5525 25283 5559
rect 25225 5519 25283 5525
rect 1104 5466 25852 5488
rect 1104 5414 7950 5466
rect 8002 5414 8014 5466
rect 8066 5414 8078 5466
rect 8130 5414 8142 5466
rect 8194 5414 8206 5466
rect 8258 5414 17950 5466
rect 18002 5414 18014 5466
rect 18066 5414 18078 5466
rect 18130 5414 18142 5466
rect 18194 5414 18206 5466
rect 18258 5414 25852 5466
rect 1104 5392 25852 5414
rect 10321 5355 10379 5361
rect 10321 5321 10333 5355
rect 10367 5352 10379 5355
rect 13538 5352 13544 5364
rect 10367 5324 13544 5352
rect 10367 5321 10379 5324
rect 10321 5315 10379 5321
rect 13538 5312 13544 5324
rect 13596 5312 13602 5364
rect 19061 5355 19119 5361
rect 19061 5352 19073 5355
rect 13648 5324 19073 5352
rect 10502 5244 10508 5296
rect 10560 5284 10566 5296
rect 10560 5256 12434 5284
rect 10560 5244 10566 5256
rect 10873 5219 10931 5225
rect 10873 5185 10885 5219
rect 10919 5216 10931 5219
rect 11146 5216 11152 5228
rect 10919 5188 11152 5216
rect 10919 5185 10931 5188
rect 10873 5179 10931 5185
rect 11146 5176 11152 5188
rect 11204 5176 11210 5228
rect 12406 5216 12434 5256
rect 13262 5244 13268 5296
rect 13320 5284 13326 5296
rect 13648 5284 13676 5324
rect 19061 5321 19073 5324
rect 19107 5321 19119 5355
rect 24210 5352 24216 5364
rect 19061 5315 19119 5321
rect 19996 5324 24216 5352
rect 13320 5256 13676 5284
rect 13320 5244 13326 5256
rect 13998 5244 14004 5296
rect 14056 5244 14062 5296
rect 15378 5244 15384 5296
rect 15436 5284 15442 5296
rect 16117 5287 16175 5293
rect 16117 5284 16129 5287
rect 15436 5256 16129 5284
rect 15436 5244 15442 5256
rect 16117 5253 16129 5256
rect 16163 5253 16175 5287
rect 16117 5247 16175 5253
rect 16408 5256 17618 5284
rect 13173 5219 13231 5225
rect 13173 5216 13185 5219
rect 12406 5188 13185 5216
rect 13173 5185 13185 5188
rect 13219 5185 13231 5219
rect 13173 5179 13231 5185
rect 13722 5176 13728 5228
rect 13780 5176 13786 5228
rect 15102 5176 15108 5228
rect 15160 5216 15166 5228
rect 16408 5216 16436 5256
rect 18598 5244 18604 5296
rect 18656 5284 18662 5296
rect 19996 5293 20024 5324
rect 24210 5312 24216 5324
rect 24268 5312 24274 5364
rect 19981 5287 20039 5293
rect 18656 5256 19288 5284
rect 18656 5244 18662 5256
rect 15160 5188 16436 5216
rect 15160 5176 15166 5188
rect 16850 5176 16856 5228
rect 16908 5176 16914 5228
rect 19260 5225 19288 5256
rect 19981 5253 19993 5287
rect 20027 5253 20039 5287
rect 19981 5247 20039 5253
rect 20070 5244 20076 5296
rect 20128 5284 20134 5296
rect 20128 5256 20470 5284
rect 20128 5244 20134 5256
rect 19245 5219 19303 5225
rect 19245 5185 19257 5219
rect 19291 5185 19303 5219
rect 19245 5179 19303 5185
rect 19702 5176 19708 5228
rect 19760 5176 19766 5228
rect 22005 5219 22063 5225
rect 22005 5185 22017 5219
rect 22051 5185 22063 5219
rect 22005 5179 22063 5185
rect 10962 5108 10968 5160
rect 11020 5148 11026 5160
rect 11701 5151 11759 5157
rect 11701 5148 11713 5151
rect 11020 5120 11713 5148
rect 11020 5108 11026 5120
rect 11701 5117 11713 5120
rect 11747 5117 11759 5151
rect 11701 5111 11759 5117
rect 11977 5151 12035 5157
rect 11977 5117 11989 5151
rect 12023 5148 12035 5151
rect 15838 5148 15844 5160
rect 12023 5120 15844 5148
rect 12023 5117 12035 5120
rect 11977 5111 12035 5117
rect 15838 5108 15844 5120
rect 15896 5108 15902 5160
rect 17129 5151 17187 5157
rect 17129 5117 17141 5151
rect 17175 5148 17187 5151
rect 18598 5148 18604 5160
rect 17175 5120 18604 5148
rect 17175 5117 17187 5120
rect 17129 5111 17187 5117
rect 18598 5108 18604 5120
rect 18656 5108 18662 5160
rect 20438 5108 20444 5160
rect 20496 5148 20502 5160
rect 22020 5148 22048 5179
rect 23658 5176 23664 5228
rect 23716 5216 23722 5228
rect 23937 5219 23995 5225
rect 23937 5216 23949 5219
rect 23716 5188 23949 5216
rect 23716 5176 23722 5188
rect 23937 5185 23949 5188
rect 23983 5185 23995 5219
rect 23937 5179 23995 5185
rect 20496 5120 22048 5148
rect 22465 5151 22523 5157
rect 20496 5108 20502 5120
rect 22465 5117 22477 5151
rect 22511 5117 22523 5151
rect 22465 5111 22523 5117
rect 9490 5040 9496 5092
rect 9548 5080 9554 5092
rect 13262 5080 13268 5092
rect 9548 5052 13268 5080
rect 9548 5040 9554 5052
rect 13262 5040 13268 5052
rect 13320 5040 13326 5092
rect 19334 5080 19340 5092
rect 18156 5052 19340 5080
rect 10965 5015 11023 5021
rect 10965 4981 10977 5015
rect 11011 5012 11023 5015
rect 12802 5012 12808 5024
rect 11011 4984 12808 5012
rect 11011 4981 11023 4984
rect 10965 4975 11023 4981
rect 12802 4972 12808 4984
rect 12860 4972 12866 5024
rect 12989 5015 13047 5021
rect 12989 4981 13001 5015
rect 13035 5012 13047 5015
rect 15194 5012 15200 5024
rect 13035 4984 15200 5012
rect 13035 4981 13047 4984
rect 12989 4975 13047 4981
rect 15194 4972 15200 4984
rect 15252 4972 15258 5024
rect 15470 4972 15476 5024
rect 15528 4972 15534 5024
rect 16209 5015 16267 5021
rect 16209 4981 16221 5015
rect 16255 5012 16267 5015
rect 18156 5012 18184 5052
rect 19334 5040 19340 5052
rect 19392 5040 19398 5092
rect 22480 5080 22508 5111
rect 24762 5108 24768 5160
rect 24820 5108 24826 5160
rect 21008 5052 22508 5080
rect 16255 4984 18184 5012
rect 16255 4981 16267 4984
rect 16209 4975 16267 4981
rect 18230 4972 18236 5024
rect 18288 5012 18294 5024
rect 18601 5015 18659 5021
rect 18601 5012 18613 5015
rect 18288 4984 18613 5012
rect 18288 4972 18294 4984
rect 18601 4981 18613 4984
rect 18647 4981 18659 5015
rect 18601 4975 18659 4981
rect 20714 4972 20720 5024
rect 20772 5012 20778 5024
rect 21008 5012 21036 5052
rect 20772 4984 21036 5012
rect 20772 4972 20778 4984
rect 21450 4972 21456 5024
rect 21508 4972 21514 5024
rect 1104 4922 25852 4944
rect 1104 4870 2950 4922
rect 3002 4870 3014 4922
rect 3066 4870 3078 4922
rect 3130 4870 3142 4922
rect 3194 4870 3206 4922
rect 3258 4870 12950 4922
rect 13002 4870 13014 4922
rect 13066 4870 13078 4922
rect 13130 4870 13142 4922
rect 13194 4870 13206 4922
rect 13258 4870 22950 4922
rect 23002 4870 23014 4922
rect 23066 4870 23078 4922
rect 23130 4870 23142 4922
rect 23194 4870 23206 4922
rect 23258 4870 25852 4922
rect 1104 4848 25852 4870
rect 8846 4768 8852 4820
rect 8904 4808 8910 4820
rect 9033 4811 9091 4817
rect 9033 4808 9045 4811
rect 8904 4780 9045 4808
rect 8904 4768 8910 4780
rect 9033 4777 9045 4780
rect 9079 4808 9091 4811
rect 9079 4780 12756 4808
rect 9079 4777 9091 4780
rect 9033 4771 9091 4777
rect 9677 4743 9735 4749
rect 9677 4709 9689 4743
rect 9723 4740 9735 4743
rect 9766 4740 9772 4752
rect 9723 4712 9772 4740
rect 9723 4709 9735 4712
rect 9677 4703 9735 4709
rect 9766 4700 9772 4712
rect 9824 4700 9830 4752
rect 10321 4743 10379 4749
rect 10321 4709 10333 4743
rect 10367 4740 10379 4743
rect 12728 4740 12756 4780
rect 12802 4768 12808 4820
rect 12860 4808 12866 4820
rect 16666 4808 16672 4820
rect 12860 4780 16672 4808
rect 12860 4768 12866 4780
rect 16666 4768 16672 4780
rect 16724 4768 16730 4820
rect 16853 4811 16911 4817
rect 16853 4777 16865 4811
rect 16899 4808 16911 4811
rect 16942 4808 16948 4820
rect 16899 4780 16948 4808
rect 16899 4777 16911 4780
rect 16853 4771 16911 4777
rect 16942 4768 16948 4780
rect 17000 4768 17006 4820
rect 23750 4768 23756 4820
rect 23808 4768 23814 4820
rect 14185 4743 14243 4749
rect 10367 4712 12434 4740
rect 12728 4712 13584 4740
rect 10367 4709 10379 4712
rect 10321 4703 10379 4709
rect 5077 4675 5135 4681
rect 5077 4641 5089 4675
rect 5123 4672 5135 4675
rect 8202 4672 8208 4684
rect 5123 4644 8208 4672
rect 5123 4641 5135 4644
rect 5077 4635 5135 4641
rect 8202 4632 8208 4644
rect 8260 4632 8266 4684
rect 8478 4632 8484 4684
rect 8536 4672 8542 4684
rect 11609 4675 11667 4681
rect 11609 4672 11621 4675
rect 8536 4644 11621 4672
rect 8536 4632 8542 4644
rect 11609 4641 11621 4644
rect 11655 4641 11667 4675
rect 11609 4635 11667 4641
rect 11882 4632 11888 4684
rect 11940 4632 11946 4684
rect 12406 4672 12434 4712
rect 12897 4675 12955 4681
rect 12897 4672 12909 4675
rect 12406 4644 12909 4672
rect 12897 4641 12909 4644
rect 12943 4641 12955 4675
rect 12897 4635 12955 4641
rect 13173 4675 13231 4681
rect 13173 4641 13185 4675
rect 13219 4672 13231 4675
rect 13446 4672 13452 4684
rect 13219 4644 13452 4672
rect 13219 4641 13231 4644
rect 13173 4635 13231 4641
rect 13446 4632 13452 4644
rect 13504 4632 13510 4684
rect 13556 4672 13584 4712
rect 14185 4709 14197 4743
rect 14231 4740 14243 4743
rect 14642 4740 14648 4752
rect 14231 4712 14648 4740
rect 14231 4709 14243 4712
rect 14185 4703 14243 4709
rect 14642 4700 14648 4712
rect 14700 4700 14706 4752
rect 16482 4700 16488 4752
rect 16540 4740 16546 4752
rect 21082 4740 21088 4752
rect 16540 4712 21088 4740
rect 16540 4700 16546 4712
rect 21082 4700 21088 4712
rect 21140 4700 21146 4752
rect 24857 4743 24915 4749
rect 24857 4709 24869 4743
rect 24903 4740 24915 4743
rect 25038 4740 25044 4752
rect 24903 4712 25044 4740
rect 24903 4709 24915 4712
rect 24857 4703 24915 4709
rect 25038 4700 25044 4712
rect 25096 4700 25102 4752
rect 14366 4672 14372 4684
rect 13556 4644 14372 4672
rect 14366 4632 14372 4644
rect 14424 4632 14430 4684
rect 7098 4564 7104 4616
rect 7156 4564 7162 4616
rect 9861 4607 9919 4613
rect 9861 4573 9873 4607
rect 9907 4604 9919 4607
rect 9950 4604 9956 4616
rect 9907 4576 9956 4604
rect 9907 4573 9919 4576
rect 9861 4567 9919 4573
rect 9950 4564 9956 4576
rect 10008 4564 10014 4616
rect 10229 4607 10287 4613
rect 10229 4573 10241 4607
rect 10275 4604 10287 4607
rect 10410 4604 10416 4616
rect 10275 4576 10416 4604
rect 10275 4573 10287 4576
rect 10229 4567 10287 4573
rect 10410 4564 10416 4576
rect 10468 4604 10474 4616
rect 14660 4613 14688 4700
rect 15105 4675 15163 4681
rect 15105 4641 15117 4675
rect 15151 4672 15163 4675
rect 16850 4672 16856 4684
rect 15151 4644 16856 4672
rect 15151 4641 15163 4644
rect 15105 4635 15163 4641
rect 16850 4632 16856 4644
rect 16908 4632 16914 4684
rect 18322 4672 18328 4684
rect 16960 4644 18328 4672
rect 10505 4607 10563 4613
rect 10505 4604 10517 4607
rect 10468 4576 10517 4604
rect 10468 4564 10474 4576
rect 10505 4573 10517 4576
rect 10551 4573 10563 4607
rect 10505 4567 10563 4573
rect 11149 4607 11207 4613
rect 11149 4573 11161 4607
rect 11195 4573 11207 4607
rect 11149 4567 11207 4573
rect 14645 4607 14703 4613
rect 14645 4573 14657 4607
rect 14691 4573 14703 4607
rect 14645 4567 14703 4573
rect 5350 4496 5356 4548
rect 5408 4496 5414 4548
rect 7377 4539 7435 4545
rect 7377 4536 7389 4539
rect 6578 4508 7389 4536
rect 7377 4505 7389 4508
rect 7423 4536 7435 4539
rect 9582 4536 9588 4548
rect 7423 4508 9588 4536
rect 7423 4505 7435 4508
rect 7377 4499 7435 4505
rect 9582 4496 9588 4508
rect 9640 4496 9646 4548
rect 11164 4536 11192 4567
rect 16666 4564 16672 4616
rect 16724 4604 16730 4616
rect 16960 4604 16988 4644
rect 18322 4632 18328 4644
rect 18380 4632 18386 4684
rect 18782 4632 18788 4684
rect 18840 4672 18846 4684
rect 19889 4675 19947 4681
rect 19889 4672 19901 4675
rect 18840 4644 19901 4672
rect 18840 4632 18846 4644
rect 19889 4641 19901 4644
rect 19935 4641 19947 4675
rect 19889 4635 19947 4641
rect 21726 4632 21732 4684
rect 21784 4632 21790 4684
rect 16724 4576 16988 4604
rect 17589 4607 17647 4613
rect 16724 4564 16730 4576
rect 17589 4573 17601 4607
rect 17635 4604 17647 4607
rect 19150 4604 19156 4616
rect 17635 4576 19156 4604
rect 17635 4573 17647 4576
rect 17589 4567 17647 4573
rect 19150 4564 19156 4576
rect 19208 4564 19214 4616
rect 19613 4607 19671 4613
rect 19613 4573 19625 4607
rect 19659 4604 19671 4607
rect 20530 4604 20536 4616
rect 19659 4576 20536 4604
rect 19659 4573 19671 4576
rect 19613 4567 19671 4573
rect 20530 4564 20536 4576
rect 20588 4564 20594 4616
rect 21358 4564 21364 4616
rect 21416 4564 21422 4616
rect 21450 4564 21456 4616
rect 21508 4604 21514 4616
rect 23109 4607 23167 4613
rect 23109 4604 23121 4607
rect 21508 4576 23121 4604
rect 21508 4564 21514 4576
rect 23109 4573 23121 4576
rect 23155 4573 23167 4607
rect 23109 4567 23167 4573
rect 15286 4536 15292 4548
rect 11164 4508 15292 4536
rect 15286 4496 15292 4508
rect 15344 4496 15350 4548
rect 15378 4496 15384 4548
rect 15436 4496 15442 4548
rect 15764 4508 15870 4536
rect 1486 4428 1492 4480
rect 1544 4428 1550 4480
rect 10962 4428 10968 4480
rect 11020 4428 11026 4480
rect 14458 4428 14464 4480
rect 14516 4428 14522 4480
rect 15102 4428 15108 4480
rect 15160 4468 15166 4480
rect 15764 4468 15792 4508
rect 18322 4496 18328 4548
rect 18380 4496 18386 4548
rect 19058 4496 19064 4548
rect 19116 4536 19122 4548
rect 24673 4539 24731 4545
rect 24673 4536 24685 4539
rect 19116 4508 24685 4536
rect 19116 4496 19122 4508
rect 24673 4505 24685 4508
rect 24719 4536 24731 4539
rect 25133 4539 25191 4545
rect 25133 4536 25145 4539
rect 24719 4508 25145 4536
rect 24719 4505 24731 4508
rect 24673 4499 24731 4505
rect 25133 4505 25145 4508
rect 25179 4505 25191 4539
rect 25133 4499 25191 4505
rect 15160 4440 15792 4468
rect 15160 4428 15166 4440
rect 1104 4378 25852 4400
rect 1104 4326 7950 4378
rect 8002 4326 8014 4378
rect 8066 4326 8078 4378
rect 8130 4326 8142 4378
rect 8194 4326 8206 4378
rect 8258 4326 17950 4378
rect 18002 4326 18014 4378
rect 18066 4326 18078 4378
rect 18130 4326 18142 4378
rect 18194 4326 18206 4378
rect 18258 4326 25852 4378
rect 1104 4304 25852 4326
rect 11146 4224 11152 4276
rect 11204 4264 11210 4276
rect 11204 4236 13492 4264
rect 11204 4224 11210 4236
rect 7282 4156 7288 4208
rect 7340 4156 7346 4208
rect 13464 4196 13492 4236
rect 13538 4224 13544 4276
rect 13596 4264 13602 4276
rect 21174 4264 21180 4276
rect 13596 4236 21180 4264
rect 13596 4224 13602 4236
rect 21174 4224 21180 4236
rect 21232 4224 21238 4276
rect 21358 4224 21364 4276
rect 21416 4264 21422 4276
rect 22278 4264 22284 4276
rect 21416 4236 22284 4264
rect 21416 4224 21422 4236
rect 22278 4224 22284 4236
rect 22336 4224 22342 4276
rect 15562 4196 15568 4208
rect 12912 4168 13124 4196
rect 13464 4168 15568 4196
rect 1486 4088 1492 4140
rect 1544 4128 1550 4140
rect 1765 4131 1823 4137
rect 1765 4128 1777 4131
rect 1544 4100 1777 4128
rect 1544 4088 1550 4100
rect 1765 4097 1777 4100
rect 1811 4097 1823 4131
rect 1765 4091 1823 4097
rect 1854 4088 1860 4140
rect 1912 4128 1918 4140
rect 2409 4131 2467 4137
rect 2409 4128 2421 4131
rect 1912 4100 2421 4128
rect 1912 4088 1918 4100
rect 2409 4097 2421 4100
rect 2455 4128 2467 4131
rect 2685 4131 2743 4137
rect 2685 4128 2697 4131
rect 2455 4100 2697 4128
rect 2455 4097 2467 4100
rect 2409 4091 2467 4097
rect 2685 4097 2697 4100
rect 2731 4097 2743 4131
rect 2685 4091 2743 4097
rect 4062 4088 4068 4140
rect 4120 4128 4126 4140
rect 4341 4131 4399 4137
rect 4341 4128 4353 4131
rect 4120 4100 4353 4128
rect 4120 4088 4126 4100
rect 4341 4097 4353 4100
rect 4387 4128 4399 4131
rect 4617 4131 4675 4137
rect 4617 4128 4629 4131
rect 4387 4100 4629 4128
rect 4387 4097 4399 4100
rect 4341 4091 4399 4097
rect 4617 4097 4629 4100
rect 4663 4097 4675 4131
rect 4617 4091 4675 4097
rect 6638 4088 6644 4140
rect 6696 4128 6702 4140
rect 6733 4131 6791 4137
rect 6733 4128 6745 4131
rect 6696 4100 6745 4128
rect 6696 4088 6702 4100
rect 6733 4097 6745 4100
rect 6779 4128 6791 4131
rect 7101 4131 7159 4137
rect 7101 4128 7113 4131
rect 6779 4100 7113 4128
rect 6779 4097 6791 4100
rect 6733 4091 6791 4097
rect 7101 4097 7113 4100
rect 7147 4097 7159 4131
rect 7101 4091 7159 4097
rect 7208 4100 8524 4128
rect 1581 3995 1639 4001
rect 1581 3961 1593 3995
rect 1627 3992 1639 3995
rect 5350 3992 5356 4004
rect 1627 3964 5356 3992
rect 1627 3961 1639 3964
rect 1581 3955 1639 3961
rect 5350 3952 5356 3964
rect 5408 3952 5414 4004
rect 6178 3992 6184 4004
rect 5460 3964 6184 3992
rect 2222 3884 2228 3936
rect 2280 3884 2286 3936
rect 2866 3884 2872 3936
rect 2924 3884 2930 3936
rect 4157 3927 4215 3933
rect 4157 3893 4169 3927
rect 4203 3924 4215 3927
rect 5460 3924 5488 3964
rect 6178 3952 6184 3964
rect 6236 3952 6242 4004
rect 6549 3995 6607 4001
rect 6549 3961 6561 3995
rect 6595 3992 6607 3995
rect 7208 3992 7236 4100
rect 8386 4060 8392 4072
rect 6595 3964 7236 3992
rect 7300 4032 8392 4060
rect 6595 3961 6607 3964
rect 6549 3955 6607 3961
rect 4203 3896 5488 3924
rect 4203 3893 4215 3896
rect 4157 3887 4215 3893
rect 6086 3884 6092 3936
rect 6144 3884 6150 3936
rect 6362 3884 6368 3936
rect 6420 3924 6426 3936
rect 7300 3924 7328 4032
rect 8386 4020 8392 4032
rect 8444 4020 8450 4072
rect 8496 3992 8524 4100
rect 8846 4088 8852 4140
rect 8904 4088 8910 4140
rect 9214 4088 9220 4140
rect 9272 4128 9278 4140
rect 9493 4131 9551 4137
rect 9493 4128 9505 4131
rect 9272 4100 9505 4128
rect 9272 4088 9278 4100
rect 9493 4097 9505 4100
rect 9539 4128 9551 4131
rect 9769 4131 9827 4137
rect 9769 4128 9781 4131
rect 9539 4100 9781 4128
rect 9539 4097 9551 4100
rect 9493 4091 9551 4097
rect 9769 4097 9781 4100
rect 9815 4097 9827 4131
rect 9769 4091 9827 4097
rect 9876 4100 10548 4128
rect 8570 4020 8576 4072
rect 8628 4060 8634 4072
rect 9876 4060 9904 4100
rect 8628 4032 9904 4060
rect 10321 4063 10379 4069
rect 8628 4020 8634 4032
rect 10321 4029 10333 4063
rect 10367 4060 10379 4063
rect 10410 4060 10416 4072
rect 10367 4032 10416 4060
rect 10367 4029 10379 4032
rect 10321 4023 10379 4029
rect 10410 4020 10416 4032
rect 10468 4020 10474 4072
rect 10520 4060 10548 4100
rect 10594 4088 10600 4140
rect 10652 4088 10658 4140
rect 11885 4131 11943 4137
rect 11885 4097 11897 4131
rect 11931 4128 11943 4131
rect 12912 4128 12940 4168
rect 11931 4100 12940 4128
rect 11931 4097 11943 4100
rect 11885 4091 11943 4097
rect 12986 4088 12992 4140
rect 13044 4088 13050 4140
rect 13096 4128 13124 4168
rect 15562 4156 15568 4168
rect 15620 4156 15626 4208
rect 18414 4156 18420 4208
rect 18472 4156 18478 4208
rect 19058 4156 19064 4208
rect 19116 4196 19122 4208
rect 20901 4199 20959 4205
rect 20901 4196 20913 4199
rect 19116 4168 20913 4196
rect 19116 4156 19122 4168
rect 20901 4165 20913 4168
rect 20947 4165 20959 4199
rect 20901 4159 20959 4165
rect 21082 4156 21088 4208
rect 21140 4196 21146 4208
rect 21140 4168 22311 4196
rect 21140 4156 21146 4168
rect 15105 4131 15163 4137
rect 13096 4100 15056 4128
rect 12250 4060 12256 4072
rect 10520 4032 12256 4060
rect 12250 4020 12256 4032
rect 12308 4020 12314 4072
rect 12802 4020 12808 4072
rect 12860 4060 12866 4072
rect 13449 4063 13507 4069
rect 13449 4060 13461 4063
rect 12860 4032 13461 4060
rect 12860 4020 12866 4032
rect 13449 4029 13461 4032
rect 13495 4029 13507 4063
rect 13449 4023 13507 4029
rect 13906 4020 13912 4072
rect 13964 4060 13970 4072
rect 14366 4060 14372 4072
rect 13964 4032 14372 4060
rect 13964 4020 13970 4032
rect 14366 4020 14372 4032
rect 14424 4020 14430 4072
rect 15028 4060 15056 4100
rect 15105 4097 15117 4131
rect 15151 4128 15163 4131
rect 17037 4131 17095 4137
rect 15151 4100 15976 4128
rect 15151 4097 15163 4100
rect 15105 4091 15163 4097
rect 15470 4060 15476 4072
rect 15028 4032 15476 4060
rect 15470 4020 15476 4032
rect 15528 4020 15534 4072
rect 12066 3992 12072 4004
rect 8496 3964 12072 3992
rect 12066 3952 12072 3964
rect 12124 3952 12130 4004
rect 12529 3995 12587 4001
rect 12529 3961 12541 3995
rect 12575 3992 12587 3995
rect 15378 3992 15384 4004
rect 12575 3964 15384 3992
rect 12575 3961 12587 3964
rect 12529 3955 12587 3961
rect 15378 3952 15384 3964
rect 15436 3952 15442 4004
rect 15948 3992 15976 4100
rect 17037 4097 17049 4131
rect 17083 4128 17095 4131
rect 18432 4128 18460 4156
rect 17083 4100 18460 4128
rect 17083 4097 17095 4100
rect 17037 4091 17095 4097
rect 18506 4088 18512 4140
rect 18564 4128 18570 4140
rect 18693 4131 18751 4137
rect 18693 4128 18705 4131
rect 18564 4100 18705 4128
rect 18564 4088 18570 4100
rect 18693 4097 18705 4100
rect 18739 4097 18751 4131
rect 18693 4091 18751 4097
rect 21542 4088 21548 4140
rect 21600 4088 21606 4140
rect 22094 4088 22100 4140
rect 22152 4088 22158 4140
rect 16114 4020 16120 4072
rect 16172 4020 16178 4072
rect 16206 4020 16212 4072
rect 16264 4060 16270 4072
rect 17313 4063 17371 4069
rect 17313 4060 17325 4063
rect 16264 4032 17325 4060
rect 16264 4020 16270 4032
rect 17313 4029 17325 4032
rect 17359 4029 17371 4063
rect 17313 4023 17371 4029
rect 18414 4020 18420 4072
rect 18472 4060 18478 4072
rect 19153 4063 19211 4069
rect 19153 4060 19165 4063
rect 18472 4032 19165 4060
rect 18472 4020 18478 4032
rect 19153 4029 19165 4032
rect 19199 4029 19211 4063
rect 19153 4023 19211 4029
rect 19242 4020 19248 4072
rect 19300 4060 19306 4072
rect 20993 4063 21051 4069
rect 20993 4060 21005 4063
rect 19300 4032 21005 4060
rect 19300 4020 19306 4032
rect 20993 4029 21005 4032
rect 21039 4029 21051 4063
rect 20993 4023 21051 4029
rect 21177 4063 21235 4069
rect 21177 4029 21189 4063
rect 21223 4060 21235 4063
rect 21450 4060 21456 4072
rect 21223 4032 21456 4060
rect 21223 4029 21235 4032
rect 21177 4023 21235 4029
rect 21450 4020 21456 4032
rect 21508 4020 21514 4072
rect 22283 4060 22311 4168
rect 22922 4156 22928 4208
rect 22980 4156 22986 4208
rect 22830 4088 22836 4140
rect 22888 4128 22894 4140
rect 23845 4131 23903 4137
rect 23845 4128 23857 4131
rect 22888 4100 23857 4128
rect 22888 4088 22894 4100
rect 23845 4097 23857 4100
rect 23891 4097 23903 4131
rect 23845 4091 23903 4097
rect 24305 4063 24363 4069
rect 24305 4060 24317 4063
rect 22283 4032 24317 4060
rect 24305 4029 24317 4032
rect 24351 4029 24363 4063
rect 24305 4023 24363 4029
rect 16850 3992 16856 4004
rect 15948 3964 16856 3992
rect 16850 3952 16856 3964
rect 16908 3952 16914 4004
rect 19978 3952 19984 4004
rect 20036 3992 20042 4004
rect 22922 3992 22928 4004
rect 20036 3964 22928 3992
rect 20036 3952 20042 3964
rect 22922 3952 22928 3964
rect 22980 3952 22986 4004
rect 6420 3896 7328 3924
rect 6420 3884 6426 3896
rect 7374 3884 7380 3936
rect 7432 3924 7438 3936
rect 7469 3927 7527 3933
rect 7469 3924 7481 3927
rect 7432 3896 7481 3924
rect 7432 3884 7438 3896
rect 7469 3893 7481 3896
rect 7515 3893 7527 3927
rect 7469 3887 7527 3893
rect 8662 3884 8668 3936
rect 8720 3884 8726 3936
rect 9306 3884 9312 3936
rect 9364 3884 9370 3936
rect 9950 3884 9956 3936
rect 10008 3884 10014 3936
rect 11606 3884 11612 3936
rect 11664 3884 11670 3936
rect 12710 3884 12716 3936
rect 12768 3924 12774 3936
rect 20533 3927 20591 3933
rect 20533 3924 20545 3927
rect 12768 3896 20545 3924
rect 12768 3884 12774 3896
rect 20533 3893 20545 3896
rect 20579 3893 20591 3927
rect 20533 3887 20591 3893
rect 21542 3884 21548 3936
rect 21600 3924 21606 3936
rect 24026 3924 24032 3936
rect 21600 3896 24032 3924
rect 21600 3884 21606 3896
rect 24026 3884 24032 3896
rect 24084 3884 24090 3936
rect 1104 3834 25852 3856
rect 1104 3782 2950 3834
rect 3002 3782 3014 3834
rect 3066 3782 3078 3834
rect 3130 3782 3142 3834
rect 3194 3782 3206 3834
rect 3258 3782 12950 3834
rect 13002 3782 13014 3834
rect 13066 3782 13078 3834
rect 13130 3782 13142 3834
rect 13194 3782 13206 3834
rect 13258 3782 22950 3834
rect 23002 3782 23014 3834
rect 23066 3782 23078 3834
rect 23130 3782 23142 3834
rect 23194 3782 23206 3834
rect 23258 3782 25852 3834
rect 1104 3760 25852 3782
rect 2869 3723 2927 3729
rect 2869 3689 2881 3723
rect 2915 3720 2927 3723
rect 3786 3720 3792 3732
rect 2915 3692 3792 3720
rect 2915 3689 2927 3692
rect 2869 3683 2927 3689
rect 3786 3680 3792 3692
rect 3844 3680 3850 3732
rect 4249 3723 4307 3729
rect 4249 3689 4261 3723
rect 4295 3720 4307 3723
rect 6914 3720 6920 3732
rect 4295 3692 6920 3720
rect 4295 3689 4307 3692
rect 4249 3683 4307 3689
rect 6914 3680 6920 3692
rect 6972 3680 6978 3732
rect 8662 3680 8668 3732
rect 8720 3720 8726 3732
rect 14274 3720 14280 3732
rect 8720 3692 14280 3720
rect 8720 3680 8726 3692
rect 14274 3680 14280 3692
rect 14332 3680 14338 3732
rect 18598 3680 18604 3732
rect 18656 3680 18662 3732
rect 19518 3680 19524 3732
rect 19576 3720 19582 3732
rect 21726 3720 21732 3732
rect 19576 3692 21732 3720
rect 19576 3680 19582 3692
rect 21726 3680 21732 3692
rect 21784 3680 21790 3732
rect 22738 3680 22744 3732
rect 22796 3720 22802 3732
rect 23293 3723 23351 3729
rect 23293 3720 23305 3723
rect 22796 3692 23305 3720
rect 22796 3680 22802 3692
rect 23293 3689 23305 3692
rect 23339 3689 23351 3723
rect 23293 3683 23351 3689
rect 6362 3612 6368 3664
rect 6420 3612 6426 3664
rect 6454 3612 6460 3664
rect 6512 3652 6518 3664
rect 10134 3652 10140 3664
rect 6512 3624 10140 3652
rect 6512 3612 6518 3624
rect 10134 3612 10140 3624
rect 10192 3612 10198 3664
rect 10413 3655 10471 3661
rect 10413 3621 10425 3655
rect 10459 3652 10471 3655
rect 10502 3652 10508 3664
rect 10459 3624 10508 3652
rect 10459 3621 10471 3624
rect 10413 3615 10471 3621
rect 10502 3612 10508 3624
rect 10560 3612 10566 3664
rect 15010 3652 15016 3664
rect 12406 3624 15016 3652
rect 1857 3587 1915 3593
rect 1857 3553 1869 3587
rect 1903 3584 1915 3587
rect 2038 3584 2044 3596
rect 1903 3556 2044 3584
rect 1903 3553 1915 3556
rect 1857 3547 1915 3553
rect 2038 3544 2044 3556
rect 2096 3544 2102 3596
rect 2866 3584 2872 3596
rect 2148 3556 2872 3584
rect 1581 3519 1639 3525
rect 1581 3485 1593 3519
rect 1627 3516 1639 3519
rect 2148 3516 2176 3556
rect 2866 3544 2872 3556
rect 2924 3584 2930 3596
rect 3694 3584 3700 3596
rect 2924 3556 3700 3584
rect 2924 3544 2930 3556
rect 3694 3544 3700 3556
rect 3752 3544 3758 3596
rect 5166 3544 5172 3596
rect 5224 3544 5230 3596
rect 8113 3587 8171 3593
rect 8113 3553 8125 3587
rect 8159 3584 8171 3587
rect 8159 3556 9352 3584
rect 8159 3553 8171 3556
rect 8113 3547 8171 3553
rect 1627 3488 2176 3516
rect 1627 3485 1639 3488
rect 1581 3479 1639 3485
rect 2222 3476 2228 3528
rect 2280 3516 2286 3528
rect 3053 3519 3111 3525
rect 3053 3516 3065 3519
rect 2280 3488 3065 3516
rect 2280 3476 2286 3488
rect 3053 3485 3065 3488
rect 3099 3516 3111 3519
rect 3513 3519 3571 3525
rect 3513 3516 3525 3519
rect 3099 3488 3525 3516
rect 3099 3485 3111 3488
rect 3053 3479 3111 3485
rect 3513 3485 3525 3488
rect 3559 3485 3571 3519
rect 3513 3479 3571 3485
rect 4430 3476 4436 3528
rect 4488 3476 4494 3528
rect 4890 3476 4896 3528
rect 4948 3476 4954 3528
rect 6089 3519 6147 3525
rect 6089 3485 6101 3519
rect 6135 3516 6147 3519
rect 6270 3516 6276 3528
rect 6135 3488 6276 3516
rect 6135 3485 6147 3488
rect 6089 3479 6147 3485
rect 6270 3476 6276 3488
rect 6328 3516 6334 3528
rect 6549 3519 6607 3525
rect 6549 3516 6561 3519
rect 6328 3488 6561 3516
rect 6328 3476 6334 3488
rect 6549 3485 6561 3488
rect 6595 3485 6607 3519
rect 6549 3479 6607 3485
rect 7006 3476 7012 3528
rect 7064 3516 7070 3528
rect 7282 3516 7288 3528
rect 7064 3488 7288 3516
rect 7064 3476 7070 3488
rect 7282 3476 7288 3488
rect 7340 3476 7346 3528
rect 7929 3519 7987 3525
rect 7929 3485 7941 3519
rect 7975 3516 7987 3519
rect 8478 3516 8484 3528
rect 7975 3488 8484 3516
rect 7975 3485 7987 3488
rect 7929 3479 7987 3485
rect 8478 3476 8484 3488
rect 8536 3516 8542 3528
rect 9324 3525 9352 3556
rect 9766 3544 9772 3596
rect 9824 3544 9830 3596
rect 11333 3587 11391 3593
rect 11333 3553 11345 3587
rect 11379 3584 11391 3587
rect 12406 3584 12434 3624
rect 15010 3612 15016 3624
rect 15068 3612 15074 3664
rect 17402 3612 17408 3664
rect 17460 3652 17466 3664
rect 18322 3652 18328 3664
rect 17460 3624 18328 3652
rect 17460 3612 17466 3624
rect 18322 3612 18328 3624
rect 18380 3612 18386 3664
rect 18690 3612 18696 3664
rect 18748 3652 18754 3664
rect 18748 3624 21864 3652
rect 18748 3612 18754 3624
rect 11379 3556 12434 3584
rect 11379 3553 11391 3556
rect 11333 3547 11391 3553
rect 13998 3544 14004 3596
rect 14056 3584 14062 3596
rect 14737 3587 14795 3593
rect 14737 3584 14749 3587
rect 14056 3556 14749 3584
rect 14056 3544 14062 3556
rect 14737 3553 14749 3556
rect 14783 3553 14795 3587
rect 14737 3547 14795 3553
rect 15470 3544 15476 3596
rect 15528 3584 15534 3596
rect 16577 3587 16635 3593
rect 16577 3584 16589 3587
rect 15528 3556 16589 3584
rect 15528 3544 15534 3556
rect 16577 3553 16589 3556
rect 16623 3553 16635 3587
rect 16577 3547 16635 3553
rect 17678 3544 17684 3596
rect 17736 3584 17742 3596
rect 19889 3587 19947 3593
rect 19889 3584 19901 3587
rect 17736 3556 19901 3584
rect 17736 3544 17742 3556
rect 19889 3553 19901 3556
rect 19935 3553 19947 3587
rect 19889 3547 19947 3553
rect 21729 3587 21787 3593
rect 21729 3553 21741 3587
rect 21775 3553 21787 3587
rect 21836 3584 21864 3624
rect 22830 3584 22836 3596
rect 21836 3556 22836 3584
rect 21729 3547 21787 3553
rect 8573 3519 8631 3525
rect 8573 3516 8585 3519
rect 8536 3488 8585 3516
rect 8536 3476 8542 3488
rect 8573 3485 8585 3488
rect 8619 3485 8631 3519
rect 8573 3479 8631 3485
rect 9309 3519 9367 3525
rect 9309 3485 9321 3519
rect 9355 3516 9367 3519
rect 9582 3516 9588 3528
rect 9355 3488 9588 3516
rect 9355 3485 9367 3488
rect 9309 3479 9367 3485
rect 9582 3476 9588 3488
rect 9640 3476 9646 3528
rect 10321 3519 10379 3525
rect 10321 3485 10333 3519
rect 10367 3516 10379 3519
rect 10594 3516 10600 3528
rect 10367 3488 10600 3516
rect 10367 3485 10379 3488
rect 10321 3479 10379 3485
rect 10594 3476 10600 3488
rect 10652 3476 10658 3528
rect 11057 3519 11115 3525
rect 11057 3485 11069 3519
rect 11103 3516 11115 3519
rect 12342 3516 12348 3528
rect 11103 3488 12348 3516
rect 11103 3485 11115 3488
rect 11057 3479 11115 3485
rect 12342 3476 12348 3488
rect 12400 3476 12406 3528
rect 12529 3519 12587 3525
rect 12529 3485 12541 3519
rect 12575 3516 12587 3519
rect 13906 3516 13912 3528
rect 12575 3488 13912 3516
rect 12575 3485 12587 3488
rect 12529 3479 12587 3485
rect 13906 3476 13912 3488
rect 13964 3476 13970 3528
rect 14461 3519 14519 3525
rect 14461 3485 14473 3519
rect 14507 3516 14519 3519
rect 14642 3516 14648 3528
rect 14507 3488 14648 3516
rect 14507 3485 14519 3488
rect 14461 3479 14519 3485
rect 14642 3476 14648 3488
rect 14700 3476 14706 3528
rect 16301 3519 16359 3525
rect 16301 3485 16313 3519
rect 16347 3516 16359 3519
rect 16666 3516 16672 3528
rect 16347 3488 16672 3516
rect 16347 3485 16359 3488
rect 16301 3479 16359 3485
rect 16666 3476 16672 3488
rect 16724 3476 16730 3528
rect 16942 3476 16948 3528
rect 17000 3516 17006 3528
rect 17957 3519 18015 3525
rect 17957 3516 17969 3519
rect 17000 3488 17969 3516
rect 17000 3476 17006 3488
rect 17957 3485 17969 3488
rect 18003 3485 18015 3519
rect 17957 3479 18015 3485
rect 19613 3519 19671 3525
rect 19613 3485 19625 3519
rect 19659 3516 19671 3519
rect 20806 3516 20812 3528
rect 19659 3488 20812 3516
rect 19659 3485 19671 3488
rect 19613 3479 19671 3485
rect 20806 3476 20812 3488
rect 20864 3476 20870 3528
rect 20990 3476 20996 3528
rect 21048 3516 21054 3528
rect 21269 3519 21327 3525
rect 21269 3516 21281 3519
rect 21048 3488 21281 3516
rect 21048 3476 21054 3488
rect 21269 3485 21281 3488
rect 21315 3485 21327 3519
rect 21269 3479 21327 3485
rect 12618 3448 12624 3460
rect 9140 3420 12624 3448
rect 3326 3340 3332 3392
rect 3384 3340 3390 3392
rect 7101 3383 7159 3389
rect 7101 3349 7113 3383
rect 7147 3380 7159 3383
rect 7190 3380 7196 3392
rect 7147 3352 7196 3380
rect 7147 3349 7159 3352
rect 7101 3343 7159 3349
rect 7190 3340 7196 3352
rect 7248 3340 7254 3392
rect 7742 3340 7748 3392
rect 7800 3340 7806 3392
rect 8389 3383 8447 3389
rect 8389 3349 8401 3383
rect 8435 3380 8447 3383
rect 8570 3380 8576 3392
rect 8435 3352 8576 3380
rect 8435 3349 8447 3352
rect 8389 3343 8447 3349
rect 8570 3340 8576 3352
rect 8628 3340 8634 3392
rect 9140 3389 9168 3420
rect 12618 3408 12624 3420
rect 12676 3408 12682 3460
rect 13541 3451 13599 3457
rect 13541 3417 13553 3451
rect 13587 3448 13599 3451
rect 17586 3448 17592 3460
rect 13587 3420 17592 3448
rect 13587 3417 13599 3420
rect 13541 3411 13599 3417
rect 17586 3408 17592 3420
rect 17644 3408 17650 3460
rect 19150 3408 19156 3460
rect 19208 3448 19214 3460
rect 21744 3448 21772 3547
rect 22830 3544 22836 3556
rect 22888 3544 22894 3596
rect 23308 3516 23336 3683
rect 23474 3680 23480 3732
rect 23532 3720 23538 3732
rect 23661 3723 23719 3729
rect 23661 3720 23673 3723
rect 23532 3692 23673 3720
rect 23532 3680 23538 3692
rect 23661 3689 23673 3692
rect 23707 3689 23719 3723
rect 23661 3683 23719 3689
rect 24854 3612 24860 3664
rect 24912 3612 24918 3664
rect 23569 3519 23627 3525
rect 23569 3516 23581 3519
rect 23308 3488 23581 3516
rect 23569 3485 23581 3488
rect 23615 3485 23627 3519
rect 23569 3479 23627 3485
rect 24394 3476 24400 3528
rect 24452 3516 24458 3528
rect 24673 3519 24731 3525
rect 24673 3516 24685 3519
rect 24452 3488 24685 3516
rect 24452 3476 24458 3488
rect 24673 3485 24685 3488
rect 24719 3516 24731 3519
rect 25133 3519 25191 3525
rect 25133 3516 25145 3519
rect 24719 3488 25145 3516
rect 24719 3485 24731 3488
rect 24673 3479 24731 3485
rect 25133 3485 25145 3488
rect 25179 3485 25191 3519
rect 25133 3479 25191 3485
rect 19208 3420 21772 3448
rect 19208 3408 19214 3420
rect 9125 3383 9183 3389
rect 9125 3349 9137 3383
rect 9171 3349 9183 3383
rect 9125 3343 9183 3349
rect 9306 3340 9312 3392
rect 9364 3380 9370 3392
rect 13354 3380 13360 3392
rect 9364 3352 13360 3380
rect 9364 3340 9370 3352
rect 13354 3340 13360 3352
rect 13412 3340 13418 3392
rect 17310 3340 17316 3392
rect 17368 3380 17374 3392
rect 18874 3380 18880 3392
rect 17368 3352 18880 3380
rect 17368 3340 17374 3352
rect 18874 3340 18880 3352
rect 18932 3340 18938 3392
rect 18966 3340 18972 3392
rect 19024 3380 19030 3392
rect 23198 3380 23204 3392
rect 19024 3352 23204 3380
rect 19024 3340 19030 3352
rect 23198 3340 23204 3352
rect 23256 3340 23262 3392
rect 1104 3290 25852 3312
rect 1104 3238 7950 3290
rect 8002 3238 8014 3290
rect 8066 3238 8078 3290
rect 8130 3238 8142 3290
rect 8194 3238 8206 3290
rect 8258 3238 17950 3290
rect 18002 3238 18014 3290
rect 18066 3238 18078 3290
rect 18130 3238 18142 3290
rect 18194 3238 18206 3290
rect 18258 3238 25852 3290
rect 1104 3216 25852 3238
rect 4430 3136 4436 3188
rect 4488 3176 4494 3188
rect 4525 3179 4583 3185
rect 4525 3176 4537 3179
rect 4488 3148 4537 3176
rect 4488 3136 4494 3148
rect 4525 3145 4537 3148
rect 4571 3145 4583 3179
rect 4525 3139 4583 3145
rect 4801 3179 4859 3185
rect 4801 3145 4813 3179
rect 4847 3176 4859 3179
rect 4890 3176 4896 3188
rect 4847 3148 4896 3176
rect 4847 3145 4859 3148
rect 4801 3139 4859 3145
rect 4890 3136 4896 3148
rect 4948 3136 4954 3188
rect 6549 3179 6607 3185
rect 6549 3145 6561 3179
rect 6595 3145 6607 3179
rect 6549 3139 6607 3145
rect 7193 3179 7251 3185
rect 7193 3145 7205 3179
rect 7239 3176 7251 3179
rect 8938 3176 8944 3188
rect 7239 3148 8944 3176
rect 7239 3145 7251 3148
rect 7193 3139 7251 3145
rect 6564 3108 6592 3139
rect 8938 3136 8944 3148
rect 8996 3136 9002 3188
rect 9217 3179 9275 3185
rect 9217 3145 9229 3179
rect 9263 3176 9275 3179
rect 10965 3179 11023 3185
rect 9263 3148 9996 3176
rect 9263 3145 9275 3148
rect 9217 3139 9275 3145
rect 9306 3108 9312 3120
rect 6564 3080 9312 3108
rect 9306 3068 9312 3080
rect 9364 3068 9370 3120
rect 9401 3111 9459 3117
rect 9401 3077 9413 3111
rect 9447 3108 9459 3111
rect 9766 3108 9772 3120
rect 9447 3080 9772 3108
rect 9447 3077 9459 3080
rect 9401 3071 9459 3077
rect 9766 3068 9772 3080
rect 9824 3068 9830 3120
rect 2133 3043 2191 3049
rect 2133 3009 2145 3043
rect 2179 3040 2191 3043
rect 2590 3040 2596 3052
rect 2179 3012 2596 3040
rect 2179 3009 2191 3012
rect 2133 3003 2191 3009
rect 2590 3000 2596 3012
rect 2648 3000 2654 3052
rect 3326 3000 3332 3052
rect 3384 3040 3390 3052
rect 3421 3043 3479 3049
rect 3421 3040 3433 3043
rect 3384 3012 3433 3040
rect 3384 3000 3390 3012
rect 3421 3009 3433 3012
rect 3467 3009 3479 3043
rect 3421 3003 3479 3009
rect 3697 3043 3755 3049
rect 3697 3009 3709 3043
rect 3743 3040 3755 3043
rect 5074 3040 5080 3052
rect 3743 3012 5080 3040
rect 3743 3009 3755 3012
rect 3697 3003 3755 3009
rect 5074 3000 5080 3012
rect 5132 3000 5138 3052
rect 5442 3000 5448 3052
rect 5500 3000 5506 3052
rect 6733 3043 6791 3049
rect 6733 3009 6745 3043
rect 6779 3009 6791 3043
rect 6733 3003 6791 3009
rect 2409 2975 2467 2981
rect 2409 2941 2421 2975
rect 2455 2941 2467 2975
rect 2409 2935 2467 2941
rect 2424 2904 2452 2935
rect 5166 2932 5172 2984
rect 5224 2932 5230 2984
rect 6748 2916 6776 3003
rect 7374 3000 7380 3052
rect 7432 3000 7438 3052
rect 7742 3000 7748 3052
rect 7800 3040 7806 3052
rect 7837 3043 7895 3049
rect 7837 3040 7849 3043
rect 7800 3012 7849 3040
rect 7800 3000 7806 3012
rect 7837 3009 7849 3012
rect 7883 3009 7895 3043
rect 7837 3003 7895 3009
rect 9033 3043 9091 3049
rect 9033 3009 9045 3043
rect 9079 3040 9091 3043
rect 9861 3043 9919 3049
rect 9861 3040 9873 3043
rect 9079 3012 9873 3040
rect 9079 3009 9091 3012
rect 9033 3003 9091 3009
rect 9861 3009 9873 3012
rect 9907 3009 9919 3043
rect 9968 3040 9996 3148
rect 10965 3145 10977 3179
rect 11011 3176 11023 3179
rect 13630 3176 13636 3188
rect 11011 3148 13636 3176
rect 11011 3145 11023 3148
rect 10965 3139 11023 3145
rect 13630 3136 13636 3148
rect 13688 3136 13694 3188
rect 16114 3136 16120 3188
rect 16172 3176 16178 3188
rect 16172 3148 19380 3176
rect 16172 3136 16178 3148
rect 16574 3068 16580 3120
rect 16632 3108 16638 3120
rect 16632 3080 17540 3108
rect 16632 3068 16638 3080
rect 11149 3052 11207 3053
rect 10505 3043 10563 3049
rect 10505 3040 10517 3043
rect 9968 3012 10517 3040
rect 9861 3003 9919 3009
rect 10505 3009 10517 3012
rect 10551 3040 10563 3043
rect 10551 3012 10824 3040
rect 10551 3009 10563 3012
rect 10505 3003 10563 3009
rect 7650 2932 7656 2984
rect 7708 2972 7714 2984
rect 8113 2975 8171 2981
rect 8113 2972 8125 2975
rect 7708 2944 8125 2972
rect 7708 2932 7714 2944
rect 8113 2941 8125 2944
rect 8159 2941 8171 2975
rect 9876 2972 9904 3003
rect 10686 2972 10692 2984
rect 9876 2944 10692 2972
rect 8113 2935 8171 2941
rect 10686 2932 10692 2944
rect 10744 2932 10750 2984
rect 10796 2972 10824 3012
rect 11146 3000 11152 3052
rect 11204 3044 11210 3052
rect 11204 3016 11245 3044
rect 11204 3000 11210 3016
rect 11606 3000 11612 3052
rect 11664 3040 11670 3052
rect 11701 3043 11759 3049
rect 11701 3040 11713 3043
rect 11664 3012 11713 3040
rect 11664 3000 11670 3012
rect 11701 3009 11713 3012
rect 11747 3009 11759 3043
rect 11701 3003 11759 3009
rect 11977 3043 12035 3049
rect 11977 3009 11989 3043
rect 12023 3040 12035 3043
rect 12526 3040 12532 3052
rect 12023 3012 12532 3040
rect 12023 3009 12035 3012
rect 11977 3003 12035 3009
rect 12526 3000 12532 3012
rect 12584 3000 12590 3052
rect 13170 3000 13176 3052
rect 13228 3000 13234 3052
rect 14550 3000 14556 3052
rect 14608 3040 14614 3052
rect 14829 3043 14887 3049
rect 14829 3040 14841 3043
rect 14608 3012 14841 3040
rect 14608 3000 14614 3012
rect 14829 3009 14841 3012
rect 14875 3009 14887 3043
rect 14829 3003 14887 3009
rect 17037 3043 17095 3049
rect 17037 3009 17049 3043
rect 17083 3040 17095 3043
rect 17126 3040 17132 3052
rect 17083 3012 17132 3040
rect 17083 3009 17095 3012
rect 17037 3003 17095 3009
rect 17126 3000 17132 3012
rect 17184 3000 17190 3052
rect 12158 2972 12164 2984
rect 10796 2944 12164 2972
rect 12158 2932 12164 2944
rect 12216 2932 12222 2984
rect 13630 2932 13636 2984
rect 13688 2932 13694 2984
rect 14734 2932 14740 2984
rect 14792 2972 14798 2984
rect 15289 2975 15347 2981
rect 15289 2972 15301 2975
rect 14792 2944 15301 2972
rect 14792 2932 14798 2944
rect 15289 2941 15301 2944
rect 15335 2941 15347 2975
rect 15289 2935 15347 2941
rect 15838 2932 15844 2984
rect 15896 2972 15902 2984
rect 17405 2975 17463 2981
rect 17405 2972 17417 2975
rect 15896 2944 17417 2972
rect 15896 2932 15902 2944
rect 17405 2941 17417 2944
rect 17451 2941 17463 2975
rect 17512 2972 17540 3080
rect 18877 3043 18935 3049
rect 18877 3009 18889 3043
rect 18923 3040 18935 3043
rect 19242 3040 19248 3052
rect 18923 3012 19248 3040
rect 18923 3009 18935 3012
rect 18877 3003 18935 3009
rect 19242 3000 19248 3012
rect 19300 3000 19306 3052
rect 19153 2975 19211 2981
rect 19153 2972 19165 2975
rect 17512 2944 19165 2972
rect 17405 2935 17463 2941
rect 19153 2941 19165 2944
rect 19199 2941 19211 2975
rect 19153 2935 19211 2941
rect 6454 2904 6460 2916
rect 2424 2876 6460 2904
rect 6454 2864 6460 2876
rect 6512 2864 6518 2916
rect 6730 2864 6736 2916
rect 6788 2904 6794 2916
rect 8846 2904 8852 2916
rect 6788 2876 8852 2904
rect 6788 2864 6794 2876
rect 8846 2864 8852 2876
rect 8904 2864 8910 2916
rect 9677 2907 9735 2913
rect 9677 2873 9689 2907
rect 9723 2904 9735 2907
rect 9723 2876 12434 2904
rect 9723 2873 9735 2876
rect 9677 2867 9735 2873
rect 10318 2796 10324 2848
rect 10376 2796 10382 2848
rect 11146 2796 11152 2848
rect 11204 2836 11210 2848
rect 11790 2836 11796 2848
rect 11204 2808 11796 2836
rect 11204 2796 11210 2808
rect 11790 2796 11796 2808
rect 11848 2796 11854 2848
rect 12406 2836 12434 2876
rect 15102 2864 15108 2916
rect 15160 2904 15166 2916
rect 17310 2904 17316 2916
rect 15160 2876 17316 2904
rect 15160 2864 15166 2876
rect 17310 2864 17316 2876
rect 17368 2864 17374 2916
rect 19352 2904 19380 3148
rect 19886 3136 19892 3188
rect 19944 3176 19950 3188
rect 19944 3148 20760 3176
rect 19944 3136 19950 3148
rect 20162 3068 20168 3120
rect 20220 3108 20226 3120
rect 20625 3111 20683 3117
rect 20625 3108 20637 3111
rect 20220 3080 20637 3108
rect 20220 3068 20226 3080
rect 20625 3077 20637 3080
rect 20671 3077 20683 3111
rect 20732 3108 20760 3148
rect 21266 3136 21272 3188
rect 21324 3136 21330 3188
rect 22186 3136 22192 3188
rect 22244 3136 22250 3188
rect 22922 3136 22928 3188
rect 22980 3136 22986 3188
rect 24026 3136 24032 3188
rect 24084 3176 24090 3188
rect 24857 3179 24915 3185
rect 24857 3176 24869 3179
rect 24084 3148 24869 3176
rect 24084 3136 24090 3148
rect 24857 3145 24869 3148
rect 24903 3145 24915 3179
rect 24857 3139 24915 3145
rect 22097 3111 22155 3117
rect 22097 3108 22109 3111
rect 20732 3080 22109 3108
rect 20625 3071 20683 3077
rect 22097 3077 22109 3080
rect 22143 3077 22155 3111
rect 22097 3071 22155 3077
rect 22833 3111 22891 3117
rect 22833 3077 22845 3111
rect 22879 3108 22891 3111
rect 23382 3108 23388 3120
rect 22879 3080 23388 3108
rect 22879 3077 22891 3080
rect 22833 3071 22891 3077
rect 23382 3068 23388 3080
rect 23440 3068 23446 3120
rect 20809 3043 20867 3049
rect 20809 3009 20821 3043
rect 20855 3040 20867 3043
rect 21358 3040 21364 3052
rect 20855 3012 21364 3040
rect 20855 3009 20867 3012
rect 20809 3003 20867 3009
rect 21358 3000 21364 3012
rect 21416 3000 21422 3052
rect 23569 3043 23627 3049
rect 23569 3009 23581 3043
rect 23615 3040 23627 3043
rect 24302 3040 24308 3052
rect 23615 3012 24308 3040
rect 23615 3009 23627 3012
rect 23569 3003 23627 3009
rect 24302 3000 24308 3012
rect 24360 3040 24366 3052
rect 24762 3040 24768 3052
rect 24360 3012 24768 3040
rect 24360 3000 24366 3012
rect 24762 3000 24768 3012
rect 24820 3000 24826 3052
rect 21726 2932 21732 2984
rect 21784 2972 21790 2984
rect 22462 2972 22468 2984
rect 21784 2944 22468 2972
rect 21784 2932 21790 2944
rect 22462 2932 22468 2944
rect 22520 2932 22526 2984
rect 23290 2904 23296 2916
rect 19352 2876 23296 2904
rect 23290 2864 23296 2876
rect 23348 2864 23354 2916
rect 15746 2836 15752 2848
rect 12406 2808 15752 2836
rect 15746 2796 15752 2808
rect 15804 2796 15810 2848
rect 16942 2796 16948 2848
rect 17000 2836 17006 2848
rect 19886 2836 19892 2848
rect 17000 2808 19892 2836
rect 17000 2796 17006 2808
rect 19886 2796 19892 2808
rect 19944 2796 19950 2848
rect 21358 2796 21364 2848
rect 21416 2836 21422 2848
rect 22646 2836 22652 2848
rect 21416 2808 22652 2836
rect 21416 2796 21422 2808
rect 22646 2796 22652 2808
rect 22704 2796 22710 2848
rect 1104 2746 25852 2768
rect 1104 2694 2950 2746
rect 3002 2694 3014 2746
rect 3066 2694 3078 2746
rect 3130 2694 3142 2746
rect 3194 2694 3206 2746
rect 3258 2694 12950 2746
rect 13002 2694 13014 2746
rect 13066 2694 13078 2746
rect 13130 2694 13142 2746
rect 13194 2694 13206 2746
rect 13258 2694 22950 2746
rect 23002 2694 23014 2746
rect 23066 2694 23078 2746
rect 23130 2694 23142 2746
rect 23194 2694 23206 2746
rect 23258 2694 25852 2746
rect 1104 2672 25852 2694
rect 6641 2635 6699 2641
rect 6641 2601 6653 2635
rect 6687 2632 6699 2635
rect 6730 2632 6736 2644
rect 6687 2604 6736 2632
rect 6687 2601 6699 2604
rect 6641 2595 6699 2601
rect 6730 2592 6736 2604
rect 6788 2592 6794 2644
rect 10042 2632 10048 2644
rect 7300 2604 10048 2632
rect 4525 2567 4583 2573
rect 4525 2533 4537 2567
rect 4571 2564 4583 2567
rect 7300 2564 7328 2604
rect 10042 2592 10048 2604
rect 10100 2592 10106 2644
rect 10551 2635 10609 2641
rect 10551 2601 10563 2635
rect 10597 2632 10609 2635
rect 13814 2632 13820 2644
rect 10597 2604 13820 2632
rect 10597 2601 10609 2604
rect 10551 2595 10609 2601
rect 13814 2592 13820 2604
rect 13872 2592 13878 2644
rect 13906 2592 13912 2644
rect 13964 2632 13970 2644
rect 14093 2635 14151 2641
rect 14093 2632 14105 2635
rect 13964 2604 14105 2632
rect 13964 2592 13970 2604
rect 14093 2601 14105 2604
rect 14139 2601 14151 2635
rect 14093 2595 14151 2601
rect 18693 2635 18751 2641
rect 18693 2601 18705 2635
rect 18739 2632 18751 2635
rect 20898 2632 20904 2644
rect 18739 2604 20904 2632
rect 18739 2601 18751 2604
rect 18693 2595 18751 2601
rect 20898 2592 20904 2604
rect 20956 2592 20962 2644
rect 21266 2592 21272 2644
rect 21324 2592 21330 2644
rect 23842 2592 23848 2644
rect 23900 2592 23906 2644
rect 24762 2592 24768 2644
rect 24820 2632 24826 2644
rect 25409 2635 25467 2641
rect 25409 2632 25421 2635
rect 24820 2604 25421 2632
rect 24820 2592 24826 2604
rect 25409 2601 25421 2604
rect 25455 2601 25467 2635
rect 25409 2595 25467 2601
rect 4571 2536 7328 2564
rect 7745 2567 7803 2573
rect 4571 2533 4583 2536
rect 4525 2527 4583 2533
rect 7745 2533 7757 2567
rect 7791 2564 7803 2567
rect 8202 2564 8208 2576
rect 7791 2536 8208 2564
rect 7791 2533 7803 2536
rect 7745 2527 7803 2533
rect 8202 2524 8208 2536
rect 8260 2524 8266 2576
rect 9692 2536 16344 2564
rect 5258 2456 5264 2508
rect 5316 2496 5322 2508
rect 9692 2505 9720 2536
rect 5445 2499 5503 2505
rect 5445 2496 5457 2499
rect 5316 2468 5457 2496
rect 5316 2456 5322 2468
rect 5445 2465 5457 2468
rect 5491 2465 5503 2499
rect 5445 2459 5503 2465
rect 9677 2499 9735 2505
rect 9677 2465 9689 2499
rect 9723 2465 9735 2499
rect 9677 2459 9735 2465
rect 11701 2499 11759 2505
rect 11701 2465 11713 2499
rect 11747 2496 11759 2499
rect 11747 2468 16252 2496
rect 11747 2465 11759 2468
rect 11701 2459 11759 2465
rect 2593 2431 2651 2437
rect 2593 2397 2605 2431
rect 2639 2428 2651 2431
rect 2639 2400 2774 2428
rect 2639 2397 2651 2400
rect 2593 2391 2651 2397
rect 2746 2360 2774 2400
rect 2866 2388 2872 2440
rect 2924 2388 2930 2440
rect 4709 2431 4767 2437
rect 4709 2397 4721 2431
rect 4755 2397 4767 2431
rect 4709 2391 4767 2397
rect 5169 2431 5227 2437
rect 5169 2397 5181 2431
rect 5215 2428 5227 2431
rect 6086 2428 6092 2440
rect 5215 2400 6092 2428
rect 5215 2397 5227 2400
rect 5169 2391 5227 2397
rect 2958 2360 2964 2372
rect 2746 2332 2964 2360
rect 2958 2320 2964 2332
rect 3016 2360 3022 2372
rect 3973 2363 4031 2369
rect 3973 2360 3985 2363
rect 3016 2332 3985 2360
rect 3016 2320 3022 2332
rect 3973 2329 3985 2332
rect 4019 2329 4031 2363
rect 3973 2323 4031 2329
rect 4249 2363 4307 2369
rect 4249 2329 4261 2363
rect 4295 2360 4307 2363
rect 4724 2360 4752 2391
rect 6086 2388 6092 2400
rect 6144 2388 6150 2440
rect 6825 2431 6883 2437
rect 6825 2397 6837 2431
rect 6871 2428 6883 2431
rect 7285 2431 7343 2437
rect 7285 2428 7297 2431
rect 6871 2400 7297 2428
rect 6871 2397 6883 2400
rect 6825 2391 6883 2397
rect 7285 2397 7297 2400
rect 7331 2428 7343 2431
rect 7834 2428 7840 2440
rect 7331 2400 7840 2428
rect 7331 2397 7343 2400
rect 7285 2391 7343 2397
rect 7834 2388 7840 2400
rect 7892 2388 7898 2440
rect 7929 2431 7987 2437
rect 7929 2397 7941 2431
rect 7975 2428 7987 2431
rect 8573 2431 8631 2437
rect 7975 2400 8524 2428
rect 7975 2397 7987 2400
rect 7929 2391 7987 2397
rect 5902 2360 5908 2372
rect 4295 2332 5908 2360
rect 4295 2329 4307 2332
rect 4249 2323 4307 2329
rect 5902 2320 5908 2332
rect 5960 2320 5966 2372
rect 2590 2252 2596 2304
rect 2648 2292 2654 2304
rect 3789 2295 3847 2301
rect 3789 2292 3801 2295
rect 2648 2264 3801 2292
rect 2648 2252 2654 2264
rect 3789 2261 3801 2264
rect 3835 2261 3847 2295
rect 3789 2255 3847 2261
rect 5166 2252 5172 2304
rect 5224 2292 5230 2304
rect 6365 2295 6423 2301
rect 6365 2292 6377 2295
rect 5224 2264 6377 2292
rect 5224 2252 5230 2264
rect 6365 2261 6377 2264
rect 6411 2261 6423 2295
rect 6365 2255 6423 2261
rect 7098 2252 7104 2304
rect 7156 2252 7162 2304
rect 8386 2252 8392 2304
rect 8444 2252 8450 2304
rect 8496 2292 8524 2400
rect 8573 2397 8585 2431
rect 8619 2428 8631 2431
rect 9401 2431 9459 2437
rect 8619 2400 9076 2428
rect 8619 2397 8631 2400
rect 8573 2391 8631 2397
rect 9048 2369 9076 2400
rect 9401 2397 9413 2431
rect 9447 2428 9459 2431
rect 10321 2431 10379 2437
rect 10321 2428 10333 2431
rect 9447 2400 10333 2428
rect 9447 2397 9459 2400
rect 9401 2391 9459 2397
rect 10321 2397 10333 2400
rect 10367 2428 10379 2431
rect 12342 2428 12348 2440
rect 10367 2400 12348 2428
rect 10367 2397 10379 2400
rect 10321 2391 10379 2397
rect 12342 2388 12348 2400
rect 12400 2388 12406 2440
rect 12529 2431 12587 2437
rect 12529 2397 12541 2431
rect 12575 2428 12587 2431
rect 12575 2400 14320 2428
rect 12575 2397 12587 2400
rect 12529 2391 12587 2397
rect 9033 2363 9091 2369
rect 9033 2329 9045 2363
rect 9079 2360 9091 2363
rect 10962 2360 10968 2372
rect 9079 2332 10968 2360
rect 9079 2329 9091 2332
rect 9033 2323 9091 2329
rect 10962 2320 10968 2332
rect 11020 2320 11026 2372
rect 13262 2320 13268 2372
rect 13320 2320 13326 2372
rect 13814 2320 13820 2372
rect 13872 2360 13878 2372
rect 14182 2360 14188 2372
rect 13872 2332 14188 2360
rect 13872 2320 13878 2332
rect 14182 2320 14188 2332
rect 14240 2320 14246 2372
rect 9217 2295 9275 2301
rect 9217 2292 9229 2295
rect 8496 2264 9229 2292
rect 9217 2261 9229 2264
rect 9263 2292 9275 2295
rect 10318 2292 10324 2304
rect 9263 2264 10324 2292
rect 9263 2261 9275 2264
rect 9217 2255 9275 2261
rect 10318 2252 10324 2264
rect 10376 2252 10382 2304
rect 14292 2292 14320 2400
rect 14458 2388 14464 2440
rect 14516 2388 14522 2440
rect 14366 2320 14372 2372
rect 14424 2360 14430 2372
rect 15381 2363 15439 2369
rect 15381 2360 15393 2363
rect 14424 2332 15393 2360
rect 14424 2320 14430 2332
rect 15381 2329 15393 2332
rect 15427 2329 15439 2363
rect 15381 2323 15439 2329
rect 16114 2292 16120 2304
rect 14292 2264 16120 2292
rect 16114 2252 16120 2264
rect 16172 2252 16178 2304
rect 16224 2292 16252 2468
rect 16316 2428 16344 2536
rect 16390 2524 16396 2576
rect 16448 2564 16454 2576
rect 16448 2536 21496 2564
rect 16448 2524 16454 2536
rect 17310 2456 17316 2508
rect 17368 2456 17374 2508
rect 17420 2468 19564 2496
rect 16758 2428 16764 2440
rect 16316 2400 16764 2428
rect 16758 2388 16764 2400
rect 16816 2388 16822 2440
rect 17034 2388 17040 2440
rect 17092 2388 17098 2440
rect 17218 2388 17224 2440
rect 17276 2428 17282 2440
rect 17420 2428 17448 2468
rect 17276 2400 17448 2428
rect 17276 2388 17282 2400
rect 18874 2388 18880 2440
rect 18932 2388 18938 2440
rect 17494 2320 17500 2372
rect 17552 2360 17558 2372
rect 19536 2360 19564 2468
rect 19886 2456 19892 2508
rect 19944 2456 19950 2508
rect 19610 2388 19616 2440
rect 19668 2388 19674 2440
rect 21468 2437 21496 2536
rect 21634 2524 21640 2576
rect 21692 2564 21698 2576
rect 21692 2536 24072 2564
rect 21692 2524 21698 2536
rect 21542 2456 21548 2508
rect 21600 2496 21606 2508
rect 22465 2499 22523 2505
rect 22465 2496 22477 2499
rect 21600 2468 22477 2496
rect 21600 2456 21606 2468
rect 22465 2465 22477 2468
rect 22511 2465 22523 2499
rect 22465 2459 22523 2465
rect 21453 2431 21511 2437
rect 21453 2397 21465 2431
rect 21499 2397 21511 2431
rect 21453 2391 21511 2397
rect 22002 2388 22008 2440
rect 22060 2388 22066 2440
rect 24044 2437 24072 2536
rect 24029 2431 24087 2437
rect 24029 2397 24041 2431
rect 24075 2397 24087 2431
rect 24029 2391 24087 2397
rect 22094 2360 22100 2372
rect 17552 2332 19472 2360
rect 19536 2332 22100 2360
rect 17552 2320 17558 2332
rect 19058 2292 19064 2304
rect 16224 2264 19064 2292
rect 19058 2252 19064 2264
rect 19116 2252 19122 2304
rect 19444 2292 19472 2332
rect 22094 2320 22100 2332
rect 22152 2320 22158 2372
rect 24673 2363 24731 2369
rect 24673 2329 24685 2363
rect 24719 2360 24731 2363
rect 25133 2363 25191 2369
rect 25133 2360 25145 2363
rect 24719 2332 25145 2360
rect 24719 2329 24731 2332
rect 24673 2323 24731 2329
rect 25133 2329 25145 2332
rect 25179 2329 25191 2363
rect 25133 2323 25191 2329
rect 24688 2292 24716 2323
rect 19444 2264 24716 2292
rect 24762 2252 24768 2304
rect 24820 2252 24826 2304
rect 1104 2202 25852 2224
rect 1104 2150 7950 2202
rect 8002 2150 8014 2202
rect 8066 2150 8078 2202
rect 8130 2150 8142 2202
rect 8194 2150 8206 2202
rect 8258 2150 17950 2202
rect 18002 2150 18014 2202
rect 18066 2150 18078 2202
rect 18130 2150 18142 2202
rect 18194 2150 18206 2202
rect 18258 2150 25852 2202
rect 1104 2128 25852 2150
rect 8386 2048 8392 2100
rect 8444 2088 8450 2100
rect 11330 2088 11336 2100
rect 8444 2060 11336 2088
rect 8444 2048 8450 2060
rect 11330 2048 11336 2060
rect 11388 2048 11394 2100
rect 16850 2048 16856 2100
rect 16908 2088 16914 2100
rect 24762 2088 24768 2100
rect 16908 2060 24768 2088
rect 16908 2048 16914 2060
rect 24762 2048 24768 2060
rect 24820 2048 24826 2100
rect 2866 1980 2872 2032
rect 2924 2020 2930 2032
rect 10870 2020 10876 2032
rect 2924 1992 10876 2020
rect 2924 1980 2930 1992
rect 10870 1980 10876 1992
rect 10928 1980 10934 2032
rect 16022 1912 16028 1964
rect 16080 1952 16086 1964
rect 22002 1952 22008 1964
rect 16080 1924 22008 1952
rect 16080 1912 16086 1924
rect 22002 1912 22008 1924
rect 22060 1912 22066 1964
rect 10410 1844 10416 1896
rect 10468 1884 10474 1896
rect 21266 1884 21272 1896
rect 10468 1856 21272 1884
rect 10468 1844 10474 1856
rect 21266 1844 21272 1856
rect 21324 1844 21330 1896
rect 18506 1776 18512 1828
rect 18564 1816 18570 1828
rect 21542 1816 21548 1828
rect 18564 1788 21548 1816
rect 18564 1776 18570 1788
rect 21542 1776 21548 1788
rect 21600 1776 21606 1828
rect 5534 1708 5540 1760
rect 5592 1748 5598 1760
rect 6086 1748 6092 1760
rect 5592 1720 6092 1748
rect 5592 1708 5598 1720
rect 6086 1708 6092 1720
rect 6144 1708 6150 1760
rect 22278 892 22284 944
rect 22336 932 22342 944
rect 22462 932 22468 944
rect 22336 904 22468 932
rect 22336 892 22342 904
rect 22462 892 22468 904
rect 22520 892 22526 944
<< via1 >>
rect 7950 54374 8002 54426
rect 8014 54374 8066 54426
rect 8078 54374 8130 54426
rect 8142 54374 8194 54426
rect 8206 54374 8258 54426
rect 17950 54374 18002 54426
rect 18014 54374 18066 54426
rect 18078 54374 18130 54426
rect 18142 54374 18194 54426
rect 18206 54374 18258 54426
rect 18972 54315 19024 54324
rect 18972 54281 18981 54315
rect 18981 54281 19015 54315
rect 19015 54281 19024 54315
rect 18972 54272 19024 54281
rect 24492 54315 24544 54324
rect 24492 54281 24501 54315
rect 24501 54281 24535 54315
rect 24535 54281 24544 54315
rect 24492 54272 24544 54281
rect 3884 54136 3936 54188
rect 6552 54136 6604 54188
rect 6736 54179 6788 54188
rect 6736 54145 6745 54179
rect 6745 54145 6779 54179
rect 6779 54145 6788 54179
rect 6736 54136 6788 54145
rect 13452 54136 13504 54188
rect 14832 54136 14884 54188
rect 16580 54136 16632 54188
rect 17592 54136 17644 54188
rect 2412 54068 2464 54120
rect 4068 54068 4120 54120
rect 6920 54068 6972 54120
rect 8484 54068 8536 54120
rect 23480 54136 23532 54188
rect 24768 54179 24820 54188
rect 24768 54145 24777 54179
rect 24777 54145 24811 54179
rect 24811 54145 24820 54179
rect 24768 54136 24820 54145
rect 18972 54068 19024 54120
rect 18788 54000 18840 54052
rect 12624 53932 12676 53984
rect 14924 53975 14976 53984
rect 14924 53941 14933 53975
rect 14933 53941 14967 53975
rect 14967 53941 14976 53975
rect 14924 53932 14976 53941
rect 15476 53932 15528 53984
rect 17132 53932 17184 53984
rect 20720 53932 20772 53984
rect 26792 53932 26844 53984
rect 2950 53830 3002 53882
rect 3014 53830 3066 53882
rect 3078 53830 3130 53882
rect 3142 53830 3194 53882
rect 3206 53830 3258 53882
rect 12950 53830 13002 53882
rect 13014 53830 13066 53882
rect 13078 53830 13130 53882
rect 13142 53830 13194 53882
rect 13206 53830 13258 53882
rect 22950 53830 23002 53882
rect 23014 53830 23066 53882
rect 23078 53830 23130 53882
rect 23142 53830 23194 53882
rect 23206 53830 23258 53882
rect 23480 53771 23532 53780
rect 23480 53737 23489 53771
rect 23489 53737 23523 53771
rect 23523 53737 23532 53771
rect 23480 53728 23532 53737
rect 25872 53728 25924 53780
rect 1032 53592 1084 53644
rect 5172 53592 5224 53644
rect 7656 53524 7708 53576
rect 23388 53524 23440 53576
rect 24676 53567 24728 53576
rect 24676 53533 24685 53567
rect 24685 53533 24719 53567
rect 24719 53533 24728 53567
rect 24676 53524 24728 53533
rect 7564 53456 7616 53508
rect 23940 53431 23992 53440
rect 23940 53397 23949 53431
rect 23949 53397 23983 53431
rect 23983 53397 23992 53431
rect 23940 53388 23992 53397
rect 24860 53388 24912 53440
rect 7950 53286 8002 53338
rect 8014 53286 8066 53338
rect 8078 53286 8130 53338
rect 8142 53286 8194 53338
rect 8206 53286 8258 53338
rect 17950 53286 18002 53338
rect 18014 53286 18066 53338
rect 18078 53286 18130 53338
rect 18142 53286 18194 53338
rect 18206 53286 18258 53338
rect 3884 53184 3936 53236
rect 6552 53227 6604 53236
rect 6552 53193 6561 53227
rect 6561 53193 6595 53227
rect 6595 53193 6604 53227
rect 6552 53184 6604 53193
rect 9588 53048 9640 53100
rect 25044 53091 25096 53100
rect 25044 53057 25053 53091
rect 25053 53057 25087 53091
rect 25087 53057 25096 53091
rect 25044 53048 25096 53057
rect 7748 52980 7800 53032
rect 26056 52844 26108 52896
rect 2950 52742 3002 52794
rect 3014 52742 3066 52794
rect 3078 52742 3130 52794
rect 3142 52742 3194 52794
rect 3206 52742 3258 52794
rect 12950 52742 13002 52794
rect 13014 52742 13066 52794
rect 13078 52742 13130 52794
rect 13142 52742 13194 52794
rect 13206 52742 13258 52794
rect 22950 52742 23002 52794
rect 23014 52742 23066 52794
rect 23078 52742 23130 52794
rect 23142 52742 23194 52794
rect 23206 52742 23258 52794
rect 7656 52683 7708 52692
rect 7656 52649 7665 52683
rect 7665 52649 7699 52683
rect 7699 52649 7708 52683
rect 7656 52640 7708 52649
rect 7840 52572 7892 52624
rect 8392 52572 8444 52624
rect 9496 52436 9548 52488
rect 16948 52436 17000 52488
rect 20352 52436 20404 52488
rect 26516 52436 26568 52488
rect 24952 52411 25004 52420
rect 24952 52377 24961 52411
rect 24961 52377 24995 52411
rect 24995 52377 25004 52411
rect 24952 52368 25004 52377
rect 7950 52198 8002 52250
rect 8014 52198 8066 52250
rect 8078 52198 8130 52250
rect 8142 52198 8194 52250
rect 8206 52198 8258 52250
rect 17950 52198 18002 52250
rect 18014 52198 18066 52250
rect 18078 52198 18130 52250
rect 18142 52198 18194 52250
rect 18206 52198 18258 52250
rect 6736 52096 6788 52148
rect 10324 51960 10376 52012
rect 25504 51799 25556 51808
rect 25504 51765 25513 51799
rect 25513 51765 25547 51799
rect 25547 51765 25556 51799
rect 25504 51756 25556 51765
rect 2950 51654 3002 51706
rect 3014 51654 3066 51706
rect 3078 51654 3130 51706
rect 3142 51654 3194 51706
rect 3206 51654 3258 51706
rect 12950 51654 13002 51706
rect 13014 51654 13066 51706
rect 13078 51654 13130 51706
rect 13142 51654 13194 51706
rect 13206 51654 13258 51706
rect 22950 51654 23002 51706
rect 23014 51654 23066 51706
rect 23078 51654 23130 51706
rect 23142 51654 23194 51706
rect 23206 51654 23258 51706
rect 7656 51595 7708 51604
rect 7656 51561 7665 51595
rect 7665 51561 7699 51595
rect 7699 51561 7708 51595
rect 7656 51552 7708 51561
rect 7748 51552 7800 51604
rect 8484 51595 8536 51604
rect 8484 51561 8493 51595
rect 8493 51561 8527 51595
rect 8527 51561 8536 51595
rect 8484 51552 8536 51561
rect 8484 51348 8536 51400
rect 25504 51348 25556 51400
rect 21364 51212 21416 51264
rect 7950 51110 8002 51162
rect 8014 51110 8066 51162
rect 8078 51110 8130 51162
rect 8142 51110 8194 51162
rect 8206 51110 8258 51162
rect 17950 51110 18002 51162
rect 18014 51110 18066 51162
rect 18078 51110 18130 51162
rect 18142 51110 18194 51162
rect 18206 51110 18258 51162
rect 24952 50915 25004 50924
rect 24952 50881 24961 50915
rect 24961 50881 24995 50915
rect 24995 50881 25004 50915
rect 24952 50872 25004 50881
rect 25044 50711 25096 50720
rect 25044 50677 25053 50711
rect 25053 50677 25087 50711
rect 25087 50677 25096 50711
rect 25044 50668 25096 50677
rect 2950 50566 3002 50618
rect 3014 50566 3066 50618
rect 3078 50566 3130 50618
rect 3142 50566 3194 50618
rect 3206 50566 3258 50618
rect 12950 50566 13002 50618
rect 13014 50566 13066 50618
rect 13078 50566 13130 50618
rect 13142 50566 13194 50618
rect 13206 50566 13258 50618
rect 22950 50566 23002 50618
rect 23014 50566 23066 50618
rect 23078 50566 23130 50618
rect 23142 50566 23194 50618
rect 23206 50566 23258 50618
rect 16028 50464 16080 50516
rect 25044 50464 25096 50516
rect 17224 50396 17276 50448
rect 24400 50396 24452 50448
rect 25504 50167 25556 50176
rect 25504 50133 25513 50167
rect 25513 50133 25547 50167
rect 25547 50133 25556 50167
rect 25504 50124 25556 50133
rect 7950 50022 8002 50074
rect 8014 50022 8066 50074
rect 8078 50022 8130 50074
rect 8142 50022 8194 50074
rect 8206 50022 8258 50074
rect 17950 50022 18002 50074
rect 18014 50022 18066 50074
rect 18078 50022 18130 50074
rect 18142 50022 18194 50074
rect 18206 50022 18258 50074
rect 25504 49784 25556 49836
rect 20904 49716 20956 49768
rect 2950 49478 3002 49530
rect 3014 49478 3066 49530
rect 3078 49478 3130 49530
rect 3142 49478 3194 49530
rect 3206 49478 3258 49530
rect 12950 49478 13002 49530
rect 13014 49478 13066 49530
rect 13078 49478 13130 49530
rect 13142 49478 13194 49530
rect 13206 49478 13258 49530
rect 22950 49478 23002 49530
rect 23014 49478 23066 49530
rect 23078 49478 23130 49530
rect 23142 49478 23194 49530
rect 23206 49478 23258 49530
rect 7656 49376 7708 49428
rect 9128 49376 9180 49428
rect 9588 49376 9640 49428
rect 8484 49308 8536 49360
rect 8760 49240 8812 49292
rect 10968 49308 11020 49360
rect 9680 49104 9732 49156
rect 25136 49147 25188 49156
rect 25136 49113 25145 49147
rect 25145 49113 25179 49147
rect 25179 49113 25188 49147
rect 25136 49104 25188 49113
rect 8300 49036 8352 49088
rect 8760 49079 8812 49088
rect 8760 49045 8769 49079
rect 8769 49045 8803 49079
rect 8803 49045 8812 49079
rect 8760 49036 8812 49045
rect 25228 49079 25280 49088
rect 25228 49045 25237 49079
rect 25237 49045 25271 49079
rect 25271 49045 25280 49079
rect 25228 49036 25280 49045
rect 7950 48934 8002 48986
rect 8014 48934 8066 48986
rect 8078 48934 8130 48986
rect 8142 48934 8194 48986
rect 8206 48934 8258 48986
rect 17950 48934 18002 48986
rect 18014 48934 18066 48986
rect 18078 48934 18130 48986
rect 18142 48934 18194 48986
rect 18206 48934 18258 48986
rect 7748 48764 7800 48816
rect 7748 48671 7800 48680
rect 7748 48637 7757 48671
rect 7757 48637 7791 48671
rect 7791 48637 7800 48671
rect 7748 48628 7800 48637
rect 8392 48671 8444 48680
rect 8392 48637 8401 48671
rect 8401 48637 8435 48671
rect 8435 48637 8444 48671
rect 8392 48628 8444 48637
rect 12348 48492 12400 48544
rect 25136 48492 25188 48544
rect 2950 48390 3002 48442
rect 3014 48390 3066 48442
rect 3078 48390 3130 48442
rect 3142 48390 3194 48442
rect 3206 48390 3258 48442
rect 12950 48390 13002 48442
rect 13014 48390 13066 48442
rect 13078 48390 13130 48442
rect 13142 48390 13194 48442
rect 13206 48390 13258 48442
rect 22950 48390 23002 48442
rect 23014 48390 23066 48442
rect 23078 48390 23130 48442
rect 23142 48390 23194 48442
rect 23206 48390 23258 48442
rect 9588 48288 9640 48340
rect 8300 48220 8352 48272
rect 9128 48127 9180 48136
rect 9128 48093 9137 48127
rect 9137 48093 9171 48127
rect 9171 48093 9180 48127
rect 9128 48084 9180 48093
rect 25136 48127 25188 48136
rect 25136 48093 25145 48127
rect 25145 48093 25179 48127
rect 25179 48093 25188 48127
rect 25136 48084 25188 48093
rect 14464 47948 14516 48000
rect 17592 47948 17644 48000
rect 7950 47846 8002 47898
rect 8014 47846 8066 47898
rect 8078 47846 8130 47898
rect 8142 47846 8194 47898
rect 8206 47846 8258 47898
rect 17950 47846 18002 47898
rect 18014 47846 18066 47898
rect 18078 47846 18130 47898
rect 18142 47846 18194 47898
rect 18206 47846 18258 47898
rect 9588 47676 9640 47728
rect 12348 47676 12400 47728
rect 12624 47651 12676 47660
rect 12624 47617 12633 47651
rect 12633 47617 12667 47651
rect 12667 47617 12676 47651
rect 12624 47608 12676 47617
rect 25320 47651 25372 47660
rect 25320 47617 25329 47651
rect 25329 47617 25363 47651
rect 25363 47617 25372 47651
rect 25320 47608 25372 47617
rect 9312 47583 9364 47592
rect 9312 47549 9321 47583
rect 9321 47549 9355 47583
rect 9355 47549 9364 47583
rect 9312 47540 9364 47549
rect 14832 47540 14884 47592
rect 9036 47472 9088 47524
rect 25964 47404 26016 47456
rect 2950 47302 3002 47354
rect 3014 47302 3066 47354
rect 3078 47302 3130 47354
rect 3142 47302 3194 47354
rect 3206 47302 3258 47354
rect 12950 47302 13002 47354
rect 13014 47302 13066 47354
rect 13078 47302 13130 47354
rect 13142 47302 13194 47354
rect 13206 47302 13258 47354
rect 22950 47302 23002 47354
rect 23014 47302 23066 47354
rect 23078 47302 23130 47354
rect 23142 47302 23194 47354
rect 23206 47302 23258 47354
rect 10692 47200 10744 47252
rect 10968 47200 11020 47252
rect 18972 47200 19024 47252
rect 25228 47200 25280 47252
rect 9496 47132 9548 47184
rect 11520 47064 11572 47116
rect 14924 47064 14976 47116
rect 14188 46996 14240 47048
rect 10968 46928 11020 46980
rect 14280 46928 14332 46980
rect 14464 46971 14516 46980
rect 14464 46937 14473 46971
rect 14473 46937 14507 46971
rect 14507 46937 14516 46971
rect 14464 46928 14516 46937
rect 16120 46971 16172 46980
rect 16120 46937 16129 46971
rect 16129 46937 16163 46971
rect 16163 46937 16172 46971
rect 16120 46928 16172 46937
rect 25320 46860 25372 46912
rect 7950 46758 8002 46810
rect 8014 46758 8066 46810
rect 8078 46758 8130 46810
rect 8142 46758 8194 46810
rect 8206 46758 8258 46810
rect 17950 46758 18002 46810
rect 18014 46758 18066 46810
rect 18078 46758 18130 46810
rect 18142 46758 18194 46810
rect 18206 46758 18258 46810
rect 9128 46656 9180 46708
rect 9680 46588 9732 46640
rect 14280 46588 14332 46640
rect 25320 46563 25372 46572
rect 25320 46529 25329 46563
rect 25329 46529 25363 46563
rect 25363 46529 25372 46563
rect 25320 46520 25372 46529
rect 8760 46452 8812 46504
rect 10600 46452 10652 46504
rect 15476 46452 15528 46504
rect 16304 46495 16356 46504
rect 16304 46461 16313 46495
rect 16313 46461 16347 46495
rect 16347 46461 16356 46495
rect 16304 46452 16356 46461
rect 9220 46316 9272 46368
rect 9680 46316 9732 46368
rect 11152 46384 11204 46436
rect 10968 46359 11020 46368
rect 10968 46325 10977 46359
rect 10977 46325 11011 46359
rect 11011 46325 11020 46359
rect 10968 46316 11020 46325
rect 23296 46316 23348 46368
rect 2950 46214 3002 46266
rect 3014 46214 3066 46266
rect 3078 46214 3130 46266
rect 3142 46214 3194 46266
rect 3206 46214 3258 46266
rect 12950 46214 13002 46266
rect 13014 46214 13066 46266
rect 13078 46214 13130 46266
rect 13142 46214 13194 46266
rect 13206 46214 13258 46266
rect 22950 46214 23002 46266
rect 23014 46214 23066 46266
rect 23078 46214 23130 46266
rect 23142 46214 23194 46266
rect 23206 46214 23258 46266
rect 24216 46044 24268 46096
rect 10324 45976 10376 46028
rect 11520 45976 11572 46028
rect 12072 46019 12124 46028
rect 12072 45985 12081 46019
rect 12081 45985 12115 46019
rect 12115 45985 12124 46019
rect 12072 45976 12124 45985
rect 14188 45976 14240 46028
rect 10416 45951 10468 45960
rect 10416 45917 10425 45951
rect 10425 45917 10459 45951
rect 10459 45917 10468 45951
rect 10416 45908 10468 45917
rect 25320 45951 25372 45960
rect 25320 45917 25329 45951
rect 25329 45917 25363 45951
rect 25363 45917 25372 45951
rect 25320 45908 25372 45917
rect 17132 45840 17184 45892
rect 17500 45883 17552 45892
rect 17500 45849 17509 45883
rect 17509 45849 17543 45883
rect 17543 45849 17552 45883
rect 17500 45840 17552 45849
rect 7950 45670 8002 45722
rect 8014 45670 8066 45722
rect 8078 45670 8130 45722
rect 8142 45670 8194 45722
rect 8206 45670 8258 45722
rect 17950 45670 18002 45722
rect 18014 45670 18066 45722
rect 18078 45670 18130 45722
rect 18142 45670 18194 45722
rect 18206 45670 18258 45722
rect 9496 45543 9548 45552
rect 9496 45509 9505 45543
rect 9505 45509 9539 45543
rect 9539 45509 9548 45543
rect 9496 45500 9548 45509
rect 8944 45364 8996 45416
rect 10876 45407 10928 45416
rect 10876 45373 10885 45407
rect 10885 45373 10919 45407
rect 10919 45373 10928 45407
rect 10876 45364 10928 45373
rect 25320 45228 25372 45280
rect 2950 45126 3002 45178
rect 3014 45126 3066 45178
rect 3078 45126 3130 45178
rect 3142 45126 3194 45178
rect 3206 45126 3258 45178
rect 12950 45126 13002 45178
rect 13014 45126 13066 45178
rect 13078 45126 13130 45178
rect 13142 45126 13194 45178
rect 13206 45126 13258 45178
rect 22950 45126 23002 45178
rect 23014 45126 23066 45178
rect 23078 45126 23130 45178
rect 23142 45126 23194 45178
rect 23206 45126 23258 45178
rect 10600 45067 10652 45076
rect 10600 45033 10609 45067
rect 10609 45033 10643 45067
rect 10643 45033 10652 45067
rect 10600 45024 10652 45033
rect 11336 45067 11388 45076
rect 11336 45033 11345 45067
rect 11345 45033 11379 45067
rect 11379 45033 11388 45067
rect 11336 45024 11388 45033
rect 11520 45067 11572 45076
rect 11520 45033 11529 45067
rect 11529 45033 11563 45067
rect 11563 45033 11572 45067
rect 11520 45024 11572 45033
rect 15752 45024 15804 45076
rect 21364 45024 21416 45076
rect 20720 44931 20772 44940
rect 20720 44897 20729 44931
rect 20729 44897 20763 44931
rect 20763 44897 20772 44931
rect 20720 44888 20772 44897
rect 21272 44888 21324 44940
rect 9956 44863 10008 44872
rect 9956 44829 9965 44863
rect 9965 44829 9999 44863
rect 9999 44829 10008 44863
rect 9956 44820 10008 44829
rect 10692 44820 10744 44872
rect 11060 44863 11112 44872
rect 11060 44829 11069 44863
rect 11069 44829 11103 44863
rect 11103 44829 11112 44863
rect 11060 44820 11112 44829
rect 19432 44820 19484 44872
rect 25320 44863 25372 44872
rect 25320 44829 25329 44863
rect 25329 44829 25363 44863
rect 25363 44829 25372 44863
rect 25320 44820 25372 44829
rect 21272 44752 21324 44804
rect 22192 44727 22244 44736
rect 22192 44693 22201 44727
rect 22201 44693 22235 44727
rect 22235 44693 22244 44727
rect 22192 44684 22244 44693
rect 23480 44684 23532 44736
rect 7950 44582 8002 44634
rect 8014 44582 8066 44634
rect 8078 44582 8130 44634
rect 8142 44582 8194 44634
rect 8206 44582 8258 44634
rect 17950 44582 18002 44634
rect 18014 44582 18066 44634
rect 18078 44582 18130 44634
rect 18142 44582 18194 44634
rect 18206 44582 18258 44634
rect 24768 44387 24820 44396
rect 24768 44353 24777 44387
rect 24777 44353 24811 44387
rect 24811 44353 24820 44387
rect 24768 44344 24820 44353
rect 25780 44208 25832 44260
rect 2950 44038 3002 44090
rect 3014 44038 3066 44090
rect 3078 44038 3130 44090
rect 3142 44038 3194 44090
rect 3206 44038 3258 44090
rect 12950 44038 13002 44090
rect 13014 44038 13066 44090
rect 13078 44038 13130 44090
rect 13142 44038 13194 44090
rect 13206 44038 13258 44090
rect 22950 44038 23002 44090
rect 23014 44038 23066 44090
rect 23078 44038 23130 44090
rect 23142 44038 23194 44090
rect 23206 44038 23258 44090
rect 25504 43639 25556 43648
rect 25504 43605 25513 43639
rect 25513 43605 25547 43639
rect 25547 43605 25556 43639
rect 25504 43596 25556 43605
rect 7950 43494 8002 43546
rect 8014 43494 8066 43546
rect 8078 43494 8130 43546
rect 8142 43494 8194 43546
rect 8206 43494 8258 43546
rect 17950 43494 18002 43546
rect 18014 43494 18066 43546
rect 18078 43494 18130 43546
rect 18142 43494 18194 43546
rect 18206 43494 18258 43546
rect 9956 43392 10008 43444
rect 25504 43324 25556 43376
rect 11152 43256 11204 43308
rect 11704 43299 11756 43308
rect 11704 43265 11713 43299
rect 11713 43265 11747 43299
rect 11747 43265 11756 43299
rect 11704 43256 11756 43265
rect 9220 43188 9272 43240
rect 12348 43188 12400 43240
rect 11060 43120 11112 43172
rect 25596 43120 25648 43172
rect 11612 43095 11664 43104
rect 11612 43061 11621 43095
rect 11621 43061 11655 43095
rect 11655 43061 11664 43095
rect 11612 43052 11664 43061
rect 2950 42950 3002 43002
rect 3014 42950 3066 43002
rect 3078 42950 3130 43002
rect 3142 42950 3194 43002
rect 3206 42950 3258 43002
rect 12950 42950 13002 43002
rect 13014 42950 13066 43002
rect 13078 42950 13130 43002
rect 13142 42950 13194 43002
rect 13206 42950 13258 43002
rect 22950 42950 23002 43002
rect 23014 42950 23066 43002
rect 23078 42950 23130 43002
rect 23142 42950 23194 43002
rect 23206 42950 23258 43002
rect 25136 42619 25188 42628
rect 25136 42585 25145 42619
rect 25145 42585 25179 42619
rect 25179 42585 25188 42619
rect 25136 42576 25188 42585
rect 26148 42576 26200 42628
rect 7950 42406 8002 42458
rect 8014 42406 8066 42458
rect 8078 42406 8130 42458
rect 8142 42406 8194 42458
rect 8206 42406 8258 42458
rect 17950 42406 18002 42458
rect 18014 42406 18066 42458
rect 18078 42406 18130 42458
rect 18142 42406 18194 42458
rect 18206 42406 18258 42458
rect 25136 41964 25188 42016
rect 2950 41862 3002 41914
rect 3014 41862 3066 41914
rect 3078 41862 3130 41914
rect 3142 41862 3194 41914
rect 3206 41862 3258 41914
rect 12950 41862 13002 41914
rect 13014 41862 13066 41914
rect 13078 41862 13130 41914
rect 13142 41862 13194 41914
rect 13206 41862 13258 41914
rect 22950 41862 23002 41914
rect 23014 41862 23066 41914
rect 23078 41862 23130 41914
rect 23142 41862 23194 41914
rect 23206 41862 23258 41914
rect 25136 41599 25188 41608
rect 25136 41565 25145 41599
rect 25145 41565 25179 41599
rect 25179 41565 25188 41599
rect 25136 41556 25188 41565
rect 25872 41488 25924 41540
rect 16856 41420 16908 41472
rect 23940 41420 23992 41472
rect 7950 41318 8002 41370
rect 8014 41318 8066 41370
rect 8078 41318 8130 41370
rect 8142 41318 8194 41370
rect 8206 41318 8258 41370
rect 17950 41318 18002 41370
rect 18014 41318 18066 41370
rect 18078 41318 18130 41370
rect 18142 41318 18194 41370
rect 18206 41318 18258 41370
rect 25320 41123 25372 41132
rect 25320 41089 25329 41123
rect 25329 41089 25363 41123
rect 25363 41089 25372 41123
rect 25320 41080 25372 41089
rect 25228 40876 25280 40928
rect 2950 40774 3002 40826
rect 3014 40774 3066 40826
rect 3078 40774 3130 40826
rect 3142 40774 3194 40826
rect 3206 40774 3258 40826
rect 12950 40774 13002 40826
rect 13014 40774 13066 40826
rect 13078 40774 13130 40826
rect 13142 40774 13194 40826
rect 13206 40774 13258 40826
rect 22950 40774 23002 40826
rect 23014 40774 23066 40826
rect 23078 40774 23130 40826
rect 23142 40774 23194 40826
rect 23206 40774 23258 40826
rect 25412 40375 25464 40384
rect 25412 40341 25421 40375
rect 25421 40341 25455 40375
rect 25455 40341 25464 40375
rect 25412 40332 25464 40341
rect 7950 40230 8002 40282
rect 8014 40230 8066 40282
rect 8078 40230 8130 40282
rect 8142 40230 8194 40282
rect 8206 40230 8258 40282
rect 17950 40230 18002 40282
rect 18014 40230 18066 40282
rect 18078 40230 18130 40282
rect 18142 40230 18194 40282
rect 18206 40230 18258 40282
rect 12348 40171 12400 40180
rect 12348 40137 12357 40171
rect 12357 40137 12391 40171
rect 12391 40137 12400 40171
rect 12348 40128 12400 40137
rect 25044 40128 25096 40180
rect 11336 39992 11388 40044
rect 21180 39992 21232 40044
rect 23296 39992 23348 40044
rect 25412 40060 25464 40112
rect 2950 39686 3002 39738
rect 3014 39686 3066 39738
rect 3078 39686 3130 39738
rect 3142 39686 3194 39738
rect 3206 39686 3258 39738
rect 12950 39686 13002 39738
rect 13014 39686 13066 39738
rect 13078 39686 13130 39738
rect 13142 39686 13194 39738
rect 13206 39686 13258 39738
rect 22950 39686 23002 39738
rect 23014 39686 23066 39738
rect 23078 39686 23130 39738
rect 23142 39686 23194 39738
rect 23206 39686 23258 39738
rect 7748 39584 7800 39636
rect 9772 39380 9824 39432
rect 25320 39423 25372 39432
rect 25320 39389 25329 39423
rect 25329 39389 25363 39423
rect 25363 39389 25372 39423
rect 25320 39380 25372 39389
rect 22008 39244 22060 39296
rect 7950 39142 8002 39194
rect 8014 39142 8066 39194
rect 8078 39142 8130 39194
rect 8142 39142 8194 39194
rect 8206 39142 8258 39194
rect 17950 39142 18002 39194
rect 18014 39142 18066 39194
rect 18078 39142 18130 39194
rect 18142 39142 18194 39194
rect 18206 39142 18258 39194
rect 25320 38700 25372 38752
rect 2950 38598 3002 38650
rect 3014 38598 3066 38650
rect 3078 38598 3130 38650
rect 3142 38598 3194 38650
rect 3206 38598 3258 38650
rect 12950 38598 13002 38650
rect 13014 38598 13066 38650
rect 13078 38598 13130 38650
rect 13142 38598 13194 38650
rect 13206 38598 13258 38650
rect 22950 38598 23002 38650
rect 23014 38598 23066 38650
rect 23078 38598 23130 38650
rect 23142 38598 23194 38650
rect 23206 38598 23258 38650
rect 22468 38496 22520 38548
rect 24216 38496 24268 38548
rect 16672 38292 16724 38344
rect 22192 38292 22244 38344
rect 25320 38335 25372 38344
rect 25320 38301 25329 38335
rect 25329 38301 25363 38335
rect 25363 38301 25372 38335
rect 25320 38292 25372 38301
rect 16764 38156 16816 38208
rect 20536 38156 20588 38208
rect 7950 38054 8002 38106
rect 8014 38054 8066 38106
rect 8078 38054 8130 38106
rect 8142 38054 8194 38106
rect 8206 38054 8258 38106
rect 17950 38054 18002 38106
rect 18014 38054 18066 38106
rect 18078 38054 18130 38106
rect 18142 38054 18194 38106
rect 18206 38054 18258 38106
rect 25136 37859 25188 37868
rect 25136 37825 25145 37859
rect 25145 37825 25179 37859
rect 25179 37825 25188 37859
rect 25136 37816 25188 37825
rect 26608 37680 26660 37732
rect 2950 37510 3002 37562
rect 3014 37510 3066 37562
rect 3078 37510 3130 37562
rect 3142 37510 3194 37562
rect 3206 37510 3258 37562
rect 12950 37510 13002 37562
rect 13014 37510 13066 37562
rect 13078 37510 13130 37562
rect 13142 37510 13194 37562
rect 13206 37510 13258 37562
rect 22950 37510 23002 37562
rect 23014 37510 23066 37562
rect 23078 37510 23130 37562
rect 23142 37510 23194 37562
rect 23206 37510 23258 37562
rect 25320 37247 25372 37256
rect 25320 37213 25329 37247
rect 25329 37213 25363 37247
rect 25363 37213 25372 37247
rect 25320 37204 25372 37213
rect 25688 37068 25740 37120
rect 7950 36966 8002 37018
rect 8014 36966 8066 37018
rect 8078 36966 8130 37018
rect 8142 36966 8194 37018
rect 8206 36966 8258 37018
rect 17950 36966 18002 37018
rect 18014 36966 18066 37018
rect 18078 36966 18130 37018
rect 18142 36966 18194 37018
rect 18206 36966 18258 37018
rect 11336 36864 11388 36916
rect 11704 36907 11756 36916
rect 11704 36873 11713 36907
rect 11713 36873 11747 36907
rect 11747 36873 11756 36907
rect 11704 36864 11756 36873
rect 11244 36796 11296 36848
rect 25136 36771 25188 36780
rect 25136 36737 25145 36771
rect 25145 36737 25179 36771
rect 25179 36737 25188 36771
rect 25136 36728 25188 36737
rect 9680 36703 9732 36712
rect 9680 36669 9689 36703
rect 9689 36669 9723 36703
rect 9723 36669 9732 36703
rect 9680 36660 9732 36669
rect 26700 36592 26752 36644
rect 11612 36567 11664 36576
rect 11612 36533 11621 36567
rect 11621 36533 11655 36567
rect 11655 36533 11664 36567
rect 11612 36524 11664 36533
rect 2950 36422 3002 36474
rect 3014 36422 3066 36474
rect 3078 36422 3130 36474
rect 3142 36422 3194 36474
rect 3206 36422 3258 36474
rect 12950 36422 13002 36474
rect 13014 36422 13066 36474
rect 13078 36422 13130 36474
rect 13142 36422 13194 36474
rect 13206 36422 13258 36474
rect 22950 36422 23002 36474
rect 23014 36422 23066 36474
rect 23078 36422 23130 36474
rect 23142 36422 23194 36474
rect 23206 36422 23258 36474
rect 9036 36320 9088 36372
rect 9220 36116 9272 36168
rect 24768 35980 24820 36032
rect 25504 35980 25556 36032
rect 7950 35878 8002 35930
rect 8014 35878 8066 35930
rect 8078 35878 8130 35930
rect 8142 35878 8194 35930
rect 8206 35878 8258 35930
rect 17950 35878 18002 35930
rect 18014 35878 18066 35930
rect 18078 35878 18130 35930
rect 18142 35878 18194 35930
rect 18206 35878 18258 35930
rect 16120 35776 16172 35828
rect 21180 35819 21232 35828
rect 21180 35785 21189 35819
rect 21189 35785 21223 35819
rect 21223 35785 21232 35819
rect 21180 35776 21232 35785
rect 22468 35819 22520 35828
rect 22468 35785 22477 35819
rect 22477 35785 22511 35819
rect 22511 35785 22520 35819
rect 22468 35776 22520 35785
rect 22836 35776 22888 35828
rect 24952 35708 25004 35760
rect 16304 35640 16356 35692
rect 21824 35640 21876 35692
rect 21272 35615 21324 35624
rect 21272 35581 21281 35615
rect 21281 35581 21315 35615
rect 21315 35581 21324 35615
rect 21272 35572 21324 35581
rect 22100 35572 22152 35624
rect 19892 35504 19944 35556
rect 20628 35436 20680 35488
rect 24768 35436 24820 35488
rect 2950 35334 3002 35386
rect 3014 35334 3066 35386
rect 3078 35334 3130 35386
rect 3142 35334 3194 35386
rect 3206 35334 3258 35386
rect 12950 35334 13002 35386
rect 13014 35334 13066 35386
rect 13078 35334 13130 35386
rect 13142 35334 13194 35386
rect 13206 35334 13258 35386
rect 22950 35334 23002 35386
rect 23014 35334 23066 35386
rect 23078 35334 23130 35386
rect 23142 35334 23194 35386
rect 23206 35334 23258 35386
rect 17500 35232 17552 35284
rect 21364 35207 21416 35216
rect 21364 35173 21373 35207
rect 21373 35173 21407 35207
rect 21407 35173 21416 35207
rect 21364 35164 21416 35173
rect 21824 35207 21876 35216
rect 21824 35173 21833 35207
rect 21833 35173 21867 35207
rect 21867 35173 21876 35207
rect 21824 35164 21876 35173
rect 19616 35071 19668 35080
rect 19616 35037 19625 35071
rect 19625 35037 19659 35071
rect 19659 35037 19668 35071
rect 19616 35028 19668 35037
rect 22192 35028 22244 35080
rect 24952 35232 25004 35284
rect 25320 35232 25372 35284
rect 24124 35164 24176 35216
rect 23296 35139 23348 35148
rect 23296 35105 23305 35139
rect 23305 35105 23339 35139
rect 23339 35105 23348 35139
rect 23296 35096 23348 35105
rect 23388 35028 23440 35080
rect 24584 35028 24636 35080
rect 24676 34960 24728 35012
rect 19708 34892 19760 34944
rect 22468 34892 22520 34944
rect 24584 34935 24636 34944
rect 24584 34901 24593 34935
rect 24593 34901 24627 34935
rect 24627 34901 24636 34935
rect 24584 34892 24636 34901
rect 7950 34790 8002 34842
rect 8014 34790 8066 34842
rect 8078 34790 8130 34842
rect 8142 34790 8194 34842
rect 8206 34790 8258 34842
rect 17950 34790 18002 34842
rect 18014 34790 18066 34842
rect 18078 34790 18130 34842
rect 18142 34790 18194 34842
rect 18206 34790 18258 34842
rect 23664 34688 23716 34740
rect 11612 34620 11664 34672
rect 19340 34552 19392 34604
rect 21272 34552 21324 34604
rect 22100 34552 22152 34604
rect 23296 34552 23348 34604
rect 24676 34595 24728 34604
rect 24676 34561 24685 34595
rect 24685 34561 24719 34595
rect 24719 34561 24728 34595
rect 24676 34552 24728 34561
rect 20076 34527 20128 34536
rect 20076 34493 20085 34527
rect 20085 34493 20119 34527
rect 20119 34493 20128 34527
rect 20076 34484 20128 34493
rect 20260 34484 20312 34536
rect 21548 34484 21600 34536
rect 24492 34484 24544 34536
rect 16580 34416 16632 34468
rect 23756 34391 23808 34400
rect 23756 34357 23765 34391
rect 23765 34357 23799 34391
rect 23799 34357 23808 34391
rect 23756 34348 23808 34357
rect 25136 34391 25188 34400
rect 25136 34357 25145 34391
rect 25145 34357 25179 34391
rect 25179 34357 25188 34391
rect 25136 34348 25188 34357
rect 2950 34246 3002 34298
rect 3014 34246 3066 34298
rect 3078 34246 3130 34298
rect 3142 34246 3194 34298
rect 3206 34246 3258 34298
rect 12950 34246 13002 34298
rect 13014 34246 13066 34298
rect 13078 34246 13130 34298
rect 13142 34246 13194 34298
rect 13206 34246 13258 34298
rect 22950 34246 23002 34298
rect 23014 34246 23066 34298
rect 23078 34246 23130 34298
rect 23142 34246 23194 34298
rect 23206 34246 23258 34298
rect 21272 34144 21324 34196
rect 22100 34144 22152 34196
rect 19432 34076 19484 34128
rect 22284 34008 22336 34060
rect 17408 33940 17460 33992
rect 23480 33940 23532 33992
rect 16580 33804 16632 33856
rect 19708 33915 19760 33924
rect 19708 33881 19717 33915
rect 19717 33881 19751 33915
rect 19751 33881 19760 33915
rect 19708 33872 19760 33881
rect 21364 33872 21416 33924
rect 22376 33872 22428 33924
rect 23572 33804 23624 33856
rect 24400 33804 24452 33856
rect 7950 33702 8002 33754
rect 8014 33702 8066 33754
rect 8078 33702 8130 33754
rect 8142 33702 8194 33754
rect 8206 33702 8258 33754
rect 17950 33702 18002 33754
rect 18014 33702 18066 33754
rect 18078 33702 18130 33754
rect 18142 33702 18194 33754
rect 18206 33702 18258 33754
rect 9680 33600 9732 33652
rect 19616 33600 19668 33652
rect 20444 33600 20496 33652
rect 21364 33600 21416 33652
rect 22376 33600 22428 33652
rect 10232 33464 10284 33516
rect 19432 33507 19484 33516
rect 19432 33473 19441 33507
rect 19441 33473 19475 33507
rect 19475 33473 19484 33507
rect 19432 33464 19484 33473
rect 22284 33532 22336 33584
rect 23572 33600 23624 33652
rect 24400 33600 24452 33652
rect 25228 33600 25280 33652
rect 21548 33396 21600 33448
rect 23756 33396 23808 33448
rect 24768 33439 24820 33448
rect 24768 33405 24777 33439
rect 24777 33405 24811 33439
rect 24811 33405 24820 33439
rect 24768 33396 24820 33405
rect 23480 33260 23532 33312
rect 24952 33260 25004 33312
rect 2950 33158 3002 33210
rect 3014 33158 3066 33210
rect 3078 33158 3130 33210
rect 3142 33158 3194 33210
rect 3206 33158 3258 33210
rect 12950 33158 13002 33210
rect 13014 33158 13066 33210
rect 13078 33158 13130 33210
rect 13142 33158 13194 33210
rect 13206 33158 13258 33210
rect 22950 33158 23002 33210
rect 23014 33158 23066 33210
rect 23078 33158 23130 33210
rect 23142 33158 23194 33210
rect 23206 33158 23258 33210
rect 10416 33056 10468 33108
rect 21364 33056 21416 33108
rect 23296 33056 23348 33108
rect 20260 32920 20312 32972
rect 22284 32963 22336 32972
rect 22284 32929 22293 32963
rect 22293 32929 22327 32963
rect 22327 32929 22336 32963
rect 22284 32920 22336 32929
rect 25044 32963 25096 32972
rect 25044 32929 25053 32963
rect 25053 32929 25087 32963
rect 25087 32929 25096 32963
rect 25044 32920 25096 32929
rect 9312 32895 9364 32904
rect 9312 32861 9321 32895
rect 9321 32861 9355 32895
rect 9355 32861 9364 32895
rect 9312 32852 9364 32861
rect 18604 32852 18656 32904
rect 19432 32895 19484 32904
rect 19432 32861 19441 32895
rect 19441 32861 19475 32895
rect 19475 32861 19484 32895
rect 19432 32852 19484 32861
rect 23940 32852 23992 32904
rect 26056 32920 26108 32972
rect 26240 32920 26292 32972
rect 21364 32784 21416 32836
rect 22560 32827 22612 32836
rect 22560 32793 22569 32827
rect 22569 32793 22603 32827
rect 22603 32793 22612 32827
rect 22560 32784 22612 32793
rect 23572 32784 23624 32836
rect 25320 32784 25372 32836
rect 26056 32784 26108 32836
rect 17684 32716 17736 32768
rect 19524 32716 19576 32768
rect 24032 32716 24084 32768
rect 7950 32614 8002 32666
rect 8014 32614 8066 32666
rect 8078 32614 8130 32666
rect 8142 32614 8194 32666
rect 8206 32614 8258 32666
rect 17950 32614 18002 32666
rect 18014 32614 18066 32666
rect 18078 32614 18130 32666
rect 18142 32614 18194 32666
rect 18206 32614 18258 32666
rect 8944 32555 8996 32564
rect 8944 32521 8953 32555
rect 8953 32521 8987 32555
rect 8987 32521 8996 32555
rect 8944 32512 8996 32521
rect 17040 32512 17092 32564
rect 17132 32555 17184 32564
rect 17132 32521 17141 32555
rect 17141 32521 17175 32555
rect 17175 32521 17184 32555
rect 17132 32512 17184 32521
rect 18420 32512 18472 32564
rect 17684 32487 17736 32496
rect 17684 32453 17693 32487
rect 17693 32453 17727 32487
rect 17727 32453 17736 32487
rect 17684 32444 17736 32453
rect 8668 32376 8720 32428
rect 16856 32376 16908 32428
rect 17408 32419 17460 32428
rect 17408 32385 17417 32419
rect 17417 32385 17451 32419
rect 17451 32385 17460 32419
rect 17408 32376 17460 32385
rect 18972 32512 19024 32564
rect 19432 32444 19484 32496
rect 21088 32512 21140 32564
rect 26516 32512 26568 32564
rect 16672 32308 16724 32360
rect 17316 32308 17368 32360
rect 18972 32308 19024 32360
rect 21364 32308 21416 32360
rect 13452 32172 13504 32224
rect 17868 32172 17920 32224
rect 21088 32240 21140 32292
rect 19340 32172 19392 32224
rect 22100 32419 22152 32428
rect 22100 32385 22109 32419
rect 22109 32385 22143 32419
rect 22143 32385 22152 32419
rect 22100 32376 22152 32385
rect 22100 32172 22152 32224
rect 22284 32444 22336 32496
rect 23756 32444 23808 32496
rect 25320 32308 25372 32360
rect 24860 32172 24912 32224
rect 25228 32215 25280 32224
rect 25228 32181 25237 32215
rect 25237 32181 25271 32215
rect 25271 32181 25280 32215
rect 25228 32172 25280 32181
rect 2950 32070 3002 32122
rect 3014 32070 3066 32122
rect 3078 32070 3130 32122
rect 3142 32070 3194 32122
rect 3206 32070 3258 32122
rect 12950 32070 13002 32122
rect 13014 32070 13066 32122
rect 13078 32070 13130 32122
rect 13142 32070 13194 32122
rect 13206 32070 13258 32122
rect 22950 32070 23002 32122
rect 23014 32070 23066 32122
rect 23078 32070 23130 32122
rect 23142 32070 23194 32122
rect 23206 32070 23258 32122
rect 13360 31900 13412 31952
rect 17868 31968 17920 32020
rect 18604 32011 18656 32020
rect 18604 31977 18613 32011
rect 18613 31977 18647 32011
rect 18647 31977 18656 32011
rect 18604 31968 18656 31977
rect 19340 31968 19392 32020
rect 21180 31900 21232 31952
rect 22560 31968 22612 32020
rect 16672 31832 16724 31884
rect 16856 31875 16908 31884
rect 16856 31841 16865 31875
rect 16865 31841 16899 31875
rect 16899 31841 16908 31875
rect 16856 31832 16908 31841
rect 19432 31875 19484 31884
rect 19432 31841 19441 31875
rect 19441 31841 19475 31875
rect 19475 31841 19484 31875
rect 19432 31832 19484 31841
rect 20076 31832 20128 31884
rect 11520 31764 11572 31816
rect 22008 31832 22060 31884
rect 23296 31764 23348 31816
rect 25228 31764 25280 31816
rect 14280 31739 14332 31748
rect 14280 31705 14289 31739
rect 14289 31705 14323 31739
rect 14323 31705 14332 31739
rect 14280 31696 14332 31705
rect 17132 31739 17184 31748
rect 17132 31705 17141 31739
rect 17141 31705 17175 31739
rect 17175 31705 17184 31739
rect 17132 31696 17184 31705
rect 18420 31696 18472 31748
rect 18880 31696 18932 31748
rect 16672 31628 16724 31680
rect 17316 31628 17368 31680
rect 20076 31628 20128 31680
rect 21180 31671 21232 31680
rect 21180 31637 21189 31671
rect 21189 31637 21223 31671
rect 21223 31637 21232 31671
rect 21180 31628 21232 31637
rect 21272 31628 21324 31680
rect 22008 31671 22060 31680
rect 22008 31637 22017 31671
rect 22017 31637 22051 31671
rect 22051 31637 22060 31671
rect 22008 31628 22060 31637
rect 23848 31628 23900 31680
rect 7950 31526 8002 31578
rect 8014 31526 8066 31578
rect 8078 31526 8130 31578
rect 8142 31526 8194 31578
rect 8206 31526 8258 31578
rect 17950 31526 18002 31578
rect 18014 31526 18066 31578
rect 18078 31526 18130 31578
rect 18142 31526 18194 31578
rect 18206 31526 18258 31578
rect 16856 31424 16908 31476
rect 17132 31424 17184 31476
rect 20536 31424 20588 31476
rect 22008 31424 22060 31476
rect 22284 31424 22336 31476
rect 15476 31356 15528 31408
rect 21364 31399 21416 31408
rect 21364 31365 21373 31399
rect 21373 31365 21407 31399
rect 21407 31365 21416 31399
rect 21364 31356 21416 31365
rect 21732 31356 21784 31408
rect 16764 31220 16816 31272
rect 19524 31288 19576 31340
rect 19984 31288 20036 31340
rect 20352 31288 20404 31340
rect 22192 31288 22244 31340
rect 22376 31288 22428 31340
rect 23756 31288 23808 31340
rect 25320 31467 25372 31476
rect 25320 31433 25329 31467
rect 25329 31433 25363 31467
rect 25363 31433 25372 31467
rect 25320 31424 25372 31433
rect 24768 31288 24820 31340
rect 18696 31220 18748 31272
rect 19432 31152 19484 31204
rect 20536 31152 20588 31204
rect 22744 31263 22796 31272
rect 22744 31229 22753 31263
rect 22753 31229 22787 31263
rect 22787 31229 22796 31263
rect 22744 31220 22796 31229
rect 13912 31084 13964 31136
rect 15476 31127 15528 31136
rect 15476 31093 15485 31127
rect 15485 31093 15519 31127
rect 15519 31093 15528 31127
rect 15476 31084 15528 31093
rect 16580 31084 16632 31136
rect 17684 31084 17736 31136
rect 20076 31084 20128 31136
rect 23940 31084 23992 31136
rect 2950 30982 3002 31034
rect 3014 30982 3066 31034
rect 3078 30982 3130 31034
rect 3142 30982 3194 31034
rect 3206 30982 3258 31034
rect 12950 30982 13002 31034
rect 13014 30982 13066 31034
rect 13078 30982 13130 31034
rect 13142 30982 13194 31034
rect 13206 30982 13258 31034
rect 22950 30982 23002 31034
rect 23014 30982 23066 31034
rect 23078 30982 23130 31034
rect 23142 30982 23194 31034
rect 23206 30982 23258 31034
rect 18696 30880 18748 30932
rect 18880 30923 18932 30932
rect 18880 30889 18889 30923
rect 18889 30889 18923 30923
rect 18923 30889 18932 30923
rect 18880 30880 18932 30889
rect 20352 30923 20404 30932
rect 20352 30889 20361 30923
rect 20361 30889 20395 30923
rect 20395 30889 20404 30923
rect 20352 30880 20404 30889
rect 22744 30880 22796 30932
rect 19340 30744 19392 30796
rect 20536 30744 20588 30796
rect 23296 30744 23348 30796
rect 15476 30676 15528 30728
rect 18880 30676 18932 30728
rect 14280 30608 14332 30660
rect 15108 30608 15160 30660
rect 16580 30540 16632 30592
rect 17316 30540 17368 30592
rect 18420 30608 18472 30660
rect 21732 30608 21784 30660
rect 23848 30676 23900 30728
rect 23940 30676 23992 30728
rect 23572 30608 23624 30660
rect 23756 30540 23808 30592
rect 24584 30540 24636 30592
rect 7950 30438 8002 30490
rect 8014 30438 8066 30490
rect 8078 30438 8130 30490
rect 8142 30438 8194 30490
rect 8206 30438 8258 30490
rect 17950 30438 18002 30490
rect 18014 30438 18066 30490
rect 18078 30438 18130 30490
rect 18142 30438 18194 30490
rect 18206 30438 18258 30490
rect 20260 30336 20312 30388
rect 21272 30336 21324 30388
rect 22376 30336 22428 30388
rect 24492 30336 24544 30388
rect 24584 30336 24636 30388
rect 11244 30268 11296 30320
rect 10324 30200 10376 30252
rect 14372 30200 14424 30252
rect 15844 30200 15896 30252
rect 10232 30175 10284 30184
rect 10232 30141 10241 30175
rect 10241 30141 10275 30175
rect 10275 30141 10284 30175
rect 10232 30132 10284 30141
rect 9772 30064 9824 30116
rect 10048 30064 10100 30116
rect 20628 30268 20680 30320
rect 22468 30311 22520 30320
rect 22468 30277 22477 30311
rect 22477 30277 22511 30311
rect 22511 30277 22520 30311
rect 22468 30268 22520 30277
rect 18788 30200 18840 30252
rect 16028 30175 16080 30184
rect 16028 30141 16037 30175
rect 16037 30141 16071 30175
rect 16071 30141 16080 30175
rect 16028 30132 16080 30141
rect 16120 30175 16172 30184
rect 16120 30141 16129 30175
rect 16129 30141 16163 30175
rect 16163 30141 16172 30175
rect 16120 30132 16172 30141
rect 20444 30175 20496 30184
rect 20444 30141 20453 30175
rect 20453 30141 20487 30175
rect 20487 30141 20496 30175
rect 20444 30132 20496 30141
rect 23480 30268 23532 30320
rect 23572 30311 23624 30320
rect 23572 30277 23581 30311
rect 23581 30277 23615 30311
rect 23615 30277 23624 30311
rect 23572 30268 23624 30277
rect 23296 30175 23348 30184
rect 23296 30141 23305 30175
rect 23305 30141 23339 30175
rect 23339 30141 23348 30175
rect 23296 30132 23348 30141
rect 24768 30132 24820 30184
rect 16948 30064 17000 30116
rect 12532 29996 12584 30048
rect 13728 29996 13780 30048
rect 14556 29996 14608 30048
rect 16028 29996 16080 30048
rect 16212 29996 16264 30048
rect 17408 29996 17460 30048
rect 19616 29996 19668 30048
rect 21456 29996 21508 30048
rect 26792 29996 26844 30048
rect 2950 29894 3002 29946
rect 3014 29894 3066 29946
rect 3078 29894 3130 29946
rect 3142 29894 3194 29946
rect 3206 29894 3258 29946
rect 12950 29894 13002 29946
rect 13014 29894 13066 29946
rect 13078 29894 13130 29946
rect 13142 29894 13194 29946
rect 13206 29894 13258 29946
rect 22950 29894 23002 29946
rect 23014 29894 23066 29946
rect 23078 29894 23130 29946
rect 23142 29894 23194 29946
rect 23206 29894 23258 29946
rect 11244 29835 11296 29844
rect 11244 29801 11253 29835
rect 11253 29801 11287 29835
rect 11287 29801 11296 29835
rect 11244 29792 11296 29801
rect 14372 29792 14424 29844
rect 16304 29792 16356 29844
rect 11520 29699 11572 29708
rect 11520 29665 11529 29699
rect 11529 29665 11563 29699
rect 11563 29665 11572 29699
rect 11520 29656 11572 29665
rect 12532 29656 12584 29708
rect 15108 29656 15160 29708
rect 17408 29699 17460 29708
rect 17408 29665 17417 29699
rect 17417 29665 17451 29699
rect 17451 29665 17460 29699
rect 17408 29656 17460 29665
rect 22652 29792 22704 29844
rect 9128 29631 9180 29640
rect 9128 29597 9137 29631
rect 9137 29597 9171 29631
rect 9171 29597 9180 29631
rect 9128 29588 9180 29597
rect 11244 29520 11296 29572
rect 11796 29563 11848 29572
rect 11796 29529 11805 29563
rect 11805 29529 11839 29563
rect 11839 29529 11848 29563
rect 11796 29520 11848 29529
rect 9588 29452 9640 29504
rect 10232 29452 10284 29504
rect 14832 29520 14884 29572
rect 13544 29495 13596 29504
rect 13544 29461 13553 29495
rect 13553 29461 13587 29495
rect 13587 29461 13596 29495
rect 13544 29452 13596 29461
rect 15200 29452 15252 29504
rect 15476 29452 15528 29504
rect 18420 29520 18472 29572
rect 16028 29495 16080 29504
rect 16028 29461 16037 29495
rect 16037 29461 16071 29495
rect 16071 29461 16080 29495
rect 16028 29452 16080 29461
rect 16580 29495 16632 29504
rect 16580 29461 16589 29495
rect 16589 29461 16623 29495
rect 16623 29461 16632 29495
rect 16580 29452 16632 29461
rect 16856 29452 16908 29504
rect 19892 29699 19944 29708
rect 19892 29665 19901 29699
rect 19901 29665 19935 29699
rect 19935 29665 19944 29699
rect 19892 29656 19944 29665
rect 19984 29699 20036 29708
rect 19984 29665 19993 29699
rect 19993 29665 20027 29699
rect 20027 29665 20036 29699
rect 19984 29656 20036 29665
rect 22836 29724 22888 29776
rect 18788 29588 18840 29640
rect 22100 29699 22152 29708
rect 22100 29665 22109 29699
rect 22109 29665 22143 29699
rect 22143 29665 22152 29699
rect 22100 29656 22152 29665
rect 22468 29588 22520 29640
rect 25320 29631 25372 29640
rect 20444 29520 20496 29572
rect 25320 29597 25329 29631
rect 25329 29597 25363 29631
rect 25363 29597 25372 29631
rect 25320 29588 25372 29597
rect 24860 29520 24912 29572
rect 18880 29495 18932 29504
rect 18880 29461 18889 29495
rect 18889 29461 18923 29495
rect 18923 29461 18932 29495
rect 18880 29452 18932 29461
rect 19800 29495 19852 29504
rect 19800 29461 19809 29495
rect 19809 29461 19843 29495
rect 19843 29461 19852 29495
rect 19800 29452 19852 29461
rect 19984 29452 20036 29504
rect 22560 29495 22612 29504
rect 22560 29461 22569 29495
rect 22569 29461 22603 29495
rect 22603 29461 22612 29495
rect 22560 29452 22612 29461
rect 23664 29452 23716 29504
rect 23756 29452 23808 29504
rect 24584 29495 24636 29504
rect 24584 29461 24593 29495
rect 24593 29461 24627 29495
rect 24627 29461 24636 29495
rect 24584 29452 24636 29461
rect 25044 29452 25096 29504
rect 7950 29350 8002 29402
rect 8014 29350 8066 29402
rect 8078 29350 8130 29402
rect 8142 29350 8194 29402
rect 8206 29350 8258 29402
rect 17950 29350 18002 29402
rect 18014 29350 18066 29402
rect 18078 29350 18130 29402
rect 18142 29350 18194 29402
rect 18206 29350 18258 29402
rect 13360 29291 13412 29300
rect 13360 29257 13369 29291
rect 13369 29257 13403 29291
rect 13403 29257 13412 29291
rect 13360 29248 13412 29257
rect 13452 29291 13504 29300
rect 13452 29257 13461 29291
rect 13461 29257 13495 29291
rect 13495 29257 13504 29291
rect 13452 29248 13504 29257
rect 14556 29291 14608 29300
rect 14556 29257 14565 29291
rect 14565 29257 14599 29291
rect 14599 29257 14608 29291
rect 14556 29248 14608 29257
rect 16488 29248 16540 29300
rect 16580 29248 16632 29300
rect 17040 29248 17092 29300
rect 18420 29248 18472 29300
rect 19800 29248 19852 29300
rect 23112 29291 23164 29300
rect 23112 29257 23121 29291
rect 23121 29257 23155 29291
rect 23155 29257 23164 29291
rect 23112 29248 23164 29257
rect 25964 29248 26016 29300
rect 14924 29180 14976 29232
rect 20444 29223 20496 29232
rect 20444 29189 20453 29223
rect 20453 29189 20487 29223
rect 20487 29189 20496 29223
rect 20444 29180 20496 29189
rect 24400 29180 24452 29232
rect 10784 29112 10836 29164
rect 12624 29112 12676 29164
rect 13728 29112 13780 29164
rect 13912 29044 13964 29096
rect 15384 29112 15436 29164
rect 15752 29155 15804 29164
rect 15752 29121 15761 29155
rect 15761 29121 15795 29155
rect 15795 29121 15804 29155
rect 15752 29112 15804 29121
rect 17224 29155 17276 29164
rect 17224 29121 17233 29155
rect 17233 29121 17267 29155
rect 17267 29121 17276 29155
rect 17224 29112 17276 29121
rect 22652 29112 22704 29164
rect 25412 29112 25464 29164
rect 16120 29044 16172 29096
rect 17040 29044 17092 29096
rect 17408 29044 17460 29096
rect 19800 29044 19852 29096
rect 9496 28976 9548 29028
rect 12164 28976 12216 29028
rect 13636 28976 13688 29028
rect 21180 28976 21232 29028
rect 12440 28908 12492 28960
rect 22560 28908 22612 28960
rect 24860 29044 24912 29096
rect 25320 28976 25372 29028
rect 2950 28806 3002 28858
rect 3014 28806 3066 28858
rect 3078 28806 3130 28858
rect 3142 28806 3194 28858
rect 3206 28806 3258 28858
rect 12950 28806 13002 28858
rect 13014 28806 13066 28858
rect 13078 28806 13130 28858
rect 13142 28806 13194 28858
rect 13206 28806 13258 28858
rect 22950 28806 23002 28858
rect 23014 28806 23066 28858
rect 23078 28806 23130 28858
rect 23142 28806 23194 28858
rect 23206 28806 23258 28858
rect 10232 28704 10284 28756
rect 13912 28747 13964 28756
rect 13912 28713 13921 28747
rect 13921 28713 13955 28747
rect 13955 28713 13964 28747
rect 13912 28704 13964 28713
rect 18788 28704 18840 28756
rect 9128 28568 9180 28620
rect 9404 28568 9456 28620
rect 11520 28568 11572 28620
rect 12440 28568 12492 28620
rect 13544 28636 13596 28688
rect 15108 28636 15160 28688
rect 20168 28636 20220 28688
rect 22836 28636 22888 28688
rect 13084 28500 13136 28552
rect 9772 28475 9824 28484
rect 9772 28441 9781 28475
rect 9781 28441 9815 28475
rect 9815 28441 9824 28475
rect 9772 28432 9824 28441
rect 10140 28364 10192 28416
rect 11980 28364 12032 28416
rect 20076 28568 20128 28620
rect 24952 28568 25004 28620
rect 25228 28611 25280 28620
rect 25228 28577 25237 28611
rect 25237 28577 25271 28611
rect 25271 28577 25280 28611
rect 25228 28568 25280 28577
rect 15936 28500 15988 28552
rect 16396 28500 16448 28552
rect 19800 28543 19852 28552
rect 19800 28509 19809 28543
rect 19809 28509 19843 28543
rect 19843 28509 19852 28543
rect 19800 28500 19852 28509
rect 19892 28500 19944 28552
rect 17408 28475 17460 28484
rect 17408 28441 17417 28475
rect 17417 28441 17451 28475
rect 17451 28441 17460 28475
rect 17408 28432 17460 28441
rect 18420 28432 18472 28484
rect 22192 28432 22244 28484
rect 23296 28432 23348 28484
rect 13452 28407 13504 28416
rect 13452 28373 13461 28407
rect 13461 28373 13495 28407
rect 13495 28373 13504 28407
rect 13452 28364 13504 28373
rect 14740 28407 14792 28416
rect 14740 28373 14749 28407
rect 14749 28373 14783 28407
rect 14783 28373 14792 28407
rect 14740 28364 14792 28373
rect 15200 28407 15252 28416
rect 15200 28373 15209 28407
rect 15209 28373 15243 28407
rect 15243 28373 15252 28407
rect 15200 28364 15252 28373
rect 15936 28407 15988 28416
rect 15936 28373 15945 28407
rect 15945 28373 15979 28407
rect 15979 28373 15988 28407
rect 15936 28364 15988 28373
rect 16212 28364 16264 28416
rect 16488 28364 16540 28416
rect 19156 28364 19208 28416
rect 20260 28364 20312 28416
rect 22560 28364 22612 28416
rect 24860 28432 24912 28484
rect 24308 28364 24360 28416
rect 7950 28262 8002 28314
rect 8014 28262 8066 28314
rect 8078 28262 8130 28314
rect 8142 28262 8194 28314
rect 8206 28262 8258 28314
rect 17950 28262 18002 28314
rect 18014 28262 18066 28314
rect 18078 28262 18130 28314
rect 18142 28262 18194 28314
rect 18206 28262 18258 28314
rect 9772 28160 9824 28212
rect 11796 28160 11848 28212
rect 12716 28203 12768 28212
rect 12716 28169 12725 28203
rect 12725 28169 12759 28203
rect 12759 28169 12768 28203
rect 12716 28160 12768 28169
rect 13084 28160 13136 28212
rect 14740 28160 14792 28212
rect 14832 28160 14884 28212
rect 17408 28160 17460 28212
rect 20168 28160 20220 28212
rect 23204 28160 23256 28212
rect 25136 28160 25188 28212
rect 25412 28160 25464 28212
rect 11980 28092 12032 28144
rect 15936 28092 15988 28144
rect 19432 28092 19484 28144
rect 11152 28024 11204 28076
rect 13452 28024 13504 28076
rect 16028 28024 16080 28076
rect 16672 28024 16724 28076
rect 17684 28024 17736 28076
rect 18420 28067 18472 28076
rect 18420 28033 18429 28067
rect 18429 28033 18463 28067
rect 18463 28033 18472 28067
rect 18420 28024 18472 28033
rect 19248 28067 19300 28076
rect 19248 28033 19257 28067
rect 19257 28033 19291 28067
rect 19291 28033 19300 28067
rect 19248 28024 19300 28033
rect 22192 28092 22244 28144
rect 24308 28092 24360 28144
rect 10232 27888 10284 27940
rect 17408 27956 17460 28008
rect 17500 27999 17552 28008
rect 17500 27965 17509 27999
rect 17509 27965 17543 27999
rect 17543 27965 17552 27999
rect 17500 27956 17552 27965
rect 18604 27999 18656 28008
rect 18604 27965 18613 27999
rect 18613 27965 18647 27999
rect 18647 27965 18656 27999
rect 18604 27956 18656 27965
rect 14832 27888 14884 27940
rect 24584 28067 24636 28076
rect 24584 28033 24593 28067
rect 24593 28033 24627 28067
rect 24627 28033 24636 28067
rect 24584 28024 24636 28033
rect 19892 27956 19944 28008
rect 21916 27956 21968 28008
rect 12808 27820 12860 27872
rect 14004 27820 14056 27872
rect 16396 27863 16448 27872
rect 16396 27829 16405 27863
rect 16405 27829 16439 27863
rect 16439 27829 16448 27863
rect 16396 27820 16448 27829
rect 17316 27820 17368 27872
rect 17960 27820 18012 27872
rect 19064 27820 19116 27872
rect 20444 27820 20496 27872
rect 23480 27888 23532 27940
rect 24768 27999 24820 28008
rect 24768 27965 24777 27999
rect 24777 27965 24811 27999
rect 24811 27965 24820 27999
rect 24768 27956 24820 27965
rect 25228 27888 25280 27940
rect 23296 27820 23348 27872
rect 23388 27820 23440 27872
rect 25136 27820 25188 27872
rect 2950 27718 3002 27770
rect 3014 27718 3066 27770
rect 3078 27718 3130 27770
rect 3142 27718 3194 27770
rect 3206 27718 3258 27770
rect 12950 27718 13002 27770
rect 13014 27718 13066 27770
rect 13078 27718 13130 27770
rect 13142 27718 13194 27770
rect 13206 27718 13258 27770
rect 22950 27718 23002 27770
rect 23014 27718 23066 27770
rect 23078 27718 23130 27770
rect 23142 27718 23194 27770
rect 23206 27718 23258 27770
rect 14648 27659 14700 27668
rect 14648 27625 14657 27659
rect 14657 27625 14691 27659
rect 14691 27625 14700 27659
rect 14648 27616 14700 27625
rect 15108 27616 15160 27668
rect 21180 27616 21232 27668
rect 11980 27591 12032 27600
rect 11980 27557 11989 27591
rect 11989 27557 12023 27591
rect 12023 27557 12032 27591
rect 11980 27548 12032 27557
rect 18696 27548 18748 27600
rect 15108 27480 15160 27532
rect 9128 27412 9180 27464
rect 12072 27412 12124 27464
rect 16212 27412 16264 27464
rect 17132 27480 17184 27532
rect 18420 27480 18472 27532
rect 16488 27412 16540 27464
rect 17500 27412 17552 27464
rect 17960 27412 18012 27464
rect 20168 27480 20220 27532
rect 20260 27480 20312 27532
rect 22652 27523 22704 27532
rect 22652 27489 22661 27523
rect 22661 27489 22695 27523
rect 22695 27489 22704 27523
rect 22652 27480 22704 27489
rect 23388 27480 23440 27532
rect 23940 27523 23992 27532
rect 23940 27489 23949 27523
rect 23949 27489 23983 27523
rect 23983 27489 23992 27523
rect 23940 27480 23992 27489
rect 25228 27591 25280 27600
rect 25228 27557 25237 27591
rect 25237 27557 25271 27591
rect 25271 27557 25280 27591
rect 25228 27548 25280 27557
rect 26240 27480 26292 27532
rect 19432 27412 19484 27464
rect 19892 27455 19944 27464
rect 19892 27421 19901 27455
rect 19901 27421 19935 27455
rect 19935 27421 19944 27455
rect 19892 27412 19944 27421
rect 22284 27412 22336 27464
rect 23664 27455 23716 27464
rect 23664 27421 23673 27455
rect 23673 27421 23707 27455
rect 23707 27421 23716 27455
rect 23664 27412 23716 27421
rect 24032 27412 24084 27464
rect 24492 27412 24544 27464
rect 12716 27344 12768 27396
rect 18604 27344 18656 27396
rect 20260 27344 20312 27396
rect 21548 27344 21600 27396
rect 24124 27344 24176 27396
rect 11336 27276 11388 27328
rect 15476 27319 15528 27328
rect 15476 27285 15485 27319
rect 15485 27285 15519 27319
rect 15519 27285 15528 27319
rect 15476 27276 15528 27285
rect 16488 27319 16540 27328
rect 16488 27285 16497 27319
rect 16497 27285 16531 27319
rect 16531 27285 16540 27319
rect 16488 27276 16540 27285
rect 17132 27276 17184 27328
rect 17408 27276 17460 27328
rect 17684 27319 17736 27328
rect 17684 27285 17693 27319
rect 17693 27285 17727 27319
rect 17727 27285 17736 27319
rect 17684 27276 17736 27285
rect 20996 27276 21048 27328
rect 21180 27276 21232 27328
rect 22284 27276 22336 27328
rect 22744 27276 22796 27328
rect 7950 27174 8002 27226
rect 8014 27174 8066 27226
rect 8078 27174 8130 27226
rect 8142 27174 8194 27226
rect 8206 27174 8258 27226
rect 17950 27174 18002 27226
rect 18014 27174 18066 27226
rect 18078 27174 18130 27226
rect 18142 27174 18194 27226
rect 18206 27174 18258 27226
rect 12256 27072 12308 27124
rect 10140 27004 10192 27056
rect 9404 26979 9456 26988
rect 9404 26945 9413 26979
rect 9413 26945 9447 26979
rect 9447 26945 9456 26979
rect 9404 26936 9456 26945
rect 11520 26936 11572 26988
rect 15016 27072 15068 27124
rect 18604 27072 18656 27124
rect 14648 27004 14700 27056
rect 15200 27004 15252 27056
rect 15936 27004 15988 27056
rect 18512 27004 18564 27056
rect 23572 27072 23624 27124
rect 24308 27072 24360 27124
rect 21640 27004 21692 27056
rect 25136 27072 25188 27124
rect 25412 27072 25464 27124
rect 26056 27072 26108 27124
rect 14740 26936 14792 26988
rect 16396 26936 16448 26988
rect 10232 26868 10284 26920
rect 11336 26868 11388 26920
rect 12348 26868 12400 26920
rect 14004 26868 14056 26920
rect 9680 26732 9732 26784
rect 11152 26775 11204 26784
rect 11152 26741 11161 26775
rect 11161 26741 11195 26775
rect 11195 26741 11204 26775
rect 11152 26732 11204 26741
rect 12256 26732 12308 26784
rect 12716 26732 12768 26784
rect 14096 26800 14148 26852
rect 15108 26800 15160 26852
rect 14280 26732 14332 26784
rect 14372 26732 14424 26784
rect 15936 26732 15988 26784
rect 16488 26732 16540 26784
rect 20076 26868 20128 26920
rect 19248 26800 19300 26852
rect 21180 26936 21232 26988
rect 21272 26911 21324 26920
rect 21272 26877 21281 26911
rect 21281 26877 21315 26911
rect 21315 26877 21324 26911
rect 21272 26868 21324 26877
rect 23204 26911 23256 26920
rect 23204 26877 23213 26911
rect 23213 26877 23247 26911
rect 23247 26877 23256 26911
rect 23204 26868 23256 26877
rect 25228 26868 25280 26920
rect 19432 26732 19484 26784
rect 20904 26732 20956 26784
rect 21640 26732 21692 26784
rect 22652 26775 22704 26784
rect 22652 26741 22661 26775
rect 22661 26741 22695 26775
rect 22695 26741 22704 26775
rect 22652 26732 22704 26741
rect 23572 26732 23624 26784
rect 23664 26732 23716 26784
rect 24492 26732 24544 26784
rect 2950 26630 3002 26682
rect 3014 26630 3066 26682
rect 3078 26630 3130 26682
rect 3142 26630 3194 26682
rect 3206 26630 3258 26682
rect 12950 26630 13002 26682
rect 13014 26630 13066 26682
rect 13078 26630 13130 26682
rect 13142 26630 13194 26682
rect 13206 26630 13258 26682
rect 22950 26630 23002 26682
rect 23014 26630 23066 26682
rect 23078 26630 23130 26682
rect 23142 26630 23194 26682
rect 23206 26630 23258 26682
rect 12072 26528 12124 26580
rect 14004 26528 14056 26580
rect 22652 26528 22704 26580
rect 23572 26528 23624 26580
rect 25412 26528 25464 26580
rect 12900 26460 12952 26512
rect 15108 26460 15160 26512
rect 9128 26435 9180 26444
rect 9128 26401 9137 26435
rect 9137 26401 9171 26435
rect 9171 26401 9180 26435
rect 9128 26392 9180 26401
rect 9496 26392 9548 26444
rect 10140 26392 10192 26444
rect 11152 26392 11204 26444
rect 13452 26392 13504 26444
rect 14648 26392 14700 26444
rect 15016 26435 15068 26444
rect 15016 26401 15025 26435
rect 15025 26401 15059 26435
rect 15059 26401 15068 26435
rect 15016 26392 15068 26401
rect 11244 26367 11296 26376
rect 11244 26333 11253 26367
rect 11253 26333 11287 26367
rect 11287 26333 11296 26367
rect 11244 26324 11296 26333
rect 12808 26324 12860 26376
rect 14280 26324 14332 26376
rect 24676 26460 24728 26512
rect 18880 26392 18932 26444
rect 20444 26392 20496 26444
rect 20720 26392 20772 26444
rect 21272 26392 21324 26444
rect 21548 26392 21600 26444
rect 25044 26435 25096 26444
rect 25044 26401 25053 26435
rect 25053 26401 25087 26435
rect 25087 26401 25096 26435
rect 25044 26392 25096 26401
rect 25136 26435 25188 26444
rect 25136 26401 25145 26435
rect 25145 26401 25179 26435
rect 25179 26401 25188 26435
rect 25136 26392 25188 26401
rect 17960 26324 18012 26376
rect 18328 26324 18380 26376
rect 20996 26324 21048 26376
rect 10140 26256 10192 26308
rect 10692 26256 10744 26308
rect 12532 26256 12584 26308
rect 13636 26256 13688 26308
rect 14832 26299 14884 26308
rect 14832 26265 14841 26299
rect 14841 26265 14875 26299
rect 14875 26265 14884 26299
rect 14832 26256 14884 26265
rect 16580 26256 16632 26308
rect 14464 26231 14516 26240
rect 14464 26197 14473 26231
rect 14473 26197 14507 26231
rect 14507 26197 14516 26231
rect 14464 26188 14516 26197
rect 16028 26231 16080 26240
rect 16028 26197 16037 26231
rect 16037 26197 16071 26231
rect 16071 26197 16080 26231
rect 16028 26188 16080 26197
rect 16672 26188 16724 26240
rect 19984 26256 20036 26308
rect 21916 26299 21968 26308
rect 21916 26265 21925 26299
rect 21925 26265 21959 26299
rect 21959 26265 21968 26299
rect 21916 26256 21968 26265
rect 22376 26256 22428 26308
rect 25320 26324 25372 26376
rect 21640 26188 21692 26240
rect 22192 26188 22244 26240
rect 22560 26188 22612 26240
rect 23020 26231 23072 26240
rect 23020 26197 23029 26231
rect 23029 26197 23063 26231
rect 23063 26197 23072 26231
rect 23020 26188 23072 26197
rect 23848 26299 23900 26308
rect 23848 26265 23857 26299
rect 23857 26265 23891 26299
rect 23891 26265 23900 26299
rect 23848 26256 23900 26265
rect 25044 26256 25096 26308
rect 25412 26256 25464 26308
rect 7950 26086 8002 26138
rect 8014 26086 8066 26138
rect 8078 26086 8130 26138
rect 8142 26086 8194 26138
rect 8206 26086 8258 26138
rect 17950 26086 18002 26138
rect 18014 26086 18066 26138
rect 18078 26086 18130 26138
rect 18142 26086 18194 26138
rect 18206 26086 18258 26138
rect 12900 25984 12952 26036
rect 12716 25916 12768 25968
rect 11520 25848 11572 25900
rect 12348 25891 12400 25900
rect 12348 25857 12357 25891
rect 12357 25857 12391 25891
rect 12391 25857 12400 25891
rect 12348 25848 12400 25857
rect 16028 25984 16080 26036
rect 16120 25984 16172 26036
rect 18328 25984 18380 26036
rect 20076 25984 20128 26036
rect 23756 25984 23808 26036
rect 24768 25984 24820 26036
rect 15108 25916 15160 25968
rect 24124 25916 24176 25968
rect 24308 25916 24360 25968
rect 12624 25823 12676 25832
rect 12624 25789 12633 25823
rect 12633 25789 12667 25823
rect 12667 25789 12676 25823
rect 12624 25780 12676 25789
rect 12716 25780 12768 25832
rect 14004 25780 14056 25832
rect 11152 25687 11204 25696
rect 11152 25653 11161 25687
rect 11161 25653 11195 25687
rect 11195 25653 11204 25687
rect 11152 25644 11204 25653
rect 11704 25644 11756 25696
rect 20720 25848 20772 25900
rect 20812 25891 20864 25900
rect 20812 25857 20821 25891
rect 20821 25857 20855 25891
rect 20855 25857 20864 25891
rect 20812 25848 20864 25857
rect 22192 25848 22244 25900
rect 15016 25823 15068 25832
rect 15016 25789 15025 25823
rect 15025 25789 15059 25823
rect 15059 25789 15068 25823
rect 15016 25780 15068 25789
rect 15108 25823 15160 25832
rect 15108 25789 15117 25823
rect 15117 25789 15151 25823
rect 15151 25789 15160 25823
rect 15108 25780 15160 25789
rect 18880 25823 18932 25832
rect 18880 25789 18889 25823
rect 18889 25789 18923 25823
rect 18923 25789 18932 25823
rect 18880 25780 18932 25789
rect 22468 25780 22520 25832
rect 23020 25823 23072 25832
rect 23020 25789 23029 25823
rect 23029 25789 23063 25823
rect 23063 25789 23072 25823
rect 23020 25780 23072 25789
rect 15844 25712 15896 25764
rect 21916 25712 21968 25764
rect 14096 25687 14148 25696
rect 14096 25653 14105 25687
rect 14105 25653 14139 25687
rect 14139 25653 14148 25687
rect 14096 25644 14148 25653
rect 15016 25644 15068 25696
rect 16120 25644 16172 25696
rect 16488 25687 16540 25696
rect 16488 25653 16497 25687
rect 16497 25653 16531 25687
rect 16531 25653 16540 25687
rect 16488 25644 16540 25653
rect 18972 25644 19024 25696
rect 21640 25644 21692 25696
rect 22008 25687 22060 25696
rect 22008 25653 22017 25687
rect 22017 25653 22051 25687
rect 22051 25653 22060 25687
rect 22008 25644 22060 25653
rect 23296 25780 23348 25832
rect 23572 25823 23624 25832
rect 23572 25789 23581 25823
rect 23581 25789 23615 25823
rect 23615 25789 23624 25823
rect 23572 25780 23624 25789
rect 24584 25780 24636 25832
rect 23940 25644 23992 25696
rect 2950 25542 3002 25594
rect 3014 25542 3066 25594
rect 3078 25542 3130 25594
rect 3142 25542 3194 25594
rect 3206 25542 3258 25594
rect 12950 25542 13002 25594
rect 13014 25542 13066 25594
rect 13078 25542 13130 25594
rect 13142 25542 13194 25594
rect 13206 25542 13258 25594
rect 22950 25542 23002 25594
rect 23014 25542 23066 25594
rect 23078 25542 23130 25594
rect 23142 25542 23194 25594
rect 23206 25542 23258 25594
rect 10324 25483 10376 25492
rect 10324 25449 10333 25483
rect 10333 25449 10367 25483
rect 10367 25449 10376 25483
rect 10324 25440 10376 25449
rect 12624 25440 12676 25492
rect 25228 25483 25280 25492
rect 25228 25449 25237 25483
rect 25237 25449 25271 25483
rect 25271 25449 25280 25483
rect 25228 25440 25280 25449
rect 9588 25304 9640 25356
rect 12072 25347 12124 25356
rect 12072 25313 12081 25347
rect 12081 25313 12115 25347
rect 12115 25313 12124 25347
rect 12072 25304 12124 25313
rect 12716 25304 12768 25356
rect 12256 25236 12308 25288
rect 15108 25304 15160 25356
rect 13452 25236 13504 25288
rect 17316 25279 17368 25288
rect 17316 25245 17325 25279
rect 17325 25245 17359 25279
rect 17359 25245 17368 25279
rect 17316 25236 17368 25245
rect 12164 25168 12216 25220
rect 10324 25100 10376 25152
rect 11060 25100 11112 25152
rect 12072 25100 12124 25152
rect 15292 25100 15344 25152
rect 15384 25143 15436 25152
rect 15384 25109 15393 25143
rect 15393 25109 15427 25143
rect 15427 25109 15436 25143
rect 15384 25100 15436 25109
rect 19708 25279 19760 25288
rect 19708 25245 19717 25279
rect 19717 25245 19751 25279
rect 19751 25245 19760 25279
rect 19708 25236 19760 25245
rect 21088 25236 21140 25288
rect 21456 25236 21508 25288
rect 21548 25279 21600 25288
rect 21548 25245 21557 25279
rect 21557 25245 21591 25279
rect 21591 25245 21600 25279
rect 21548 25236 21600 25245
rect 24768 25236 24820 25288
rect 24952 25168 25004 25220
rect 19340 25143 19392 25152
rect 19340 25109 19349 25143
rect 19349 25109 19383 25143
rect 19383 25109 19392 25143
rect 19340 25100 19392 25109
rect 19984 25100 20036 25152
rect 20996 25143 21048 25152
rect 20996 25109 21005 25143
rect 21005 25109 21039 25143
rect 21039 25109 21048 25143
rect 20996 25100 21048 25109
rect 22192 25143 22244 25152
rect 22192 25109 22201 25143
rect 22201 25109 22235 25143
rect 22235 25109 22244 25143
rect 22192 25100 22244 25109
rect 7950 24998 8002 25050
rect 8014 24998 8066 25050
rect 8078 24998 8130 25050
rect 8142 24998 8194 25050
rect 8206 24998 8258 25050
rect 17950 24998 18002 25050
rect 18014 24998 18066 25050
rect 18078 24998 18130 25050
rect 18142 24998 18194 25050
rect 18206 24998 18258 25050
rect 10876 24896 10928 24948
rect 12256 24896 12308 24948
rect 15476 24896 15528 24948
rect 16396 24896 16448 24948
rect 17408 24896 17460 24948
rect 20168 24896 20220 24948
rect 20812 24896 20864 24948
rect 25412 24896 25464 24948
rect 9772 24828 9824 24880
rect 11152 24828 11204 24880
rect 12716 24828 12768 24880
rect 17132 24828 17184 24880
rect 11244 24803 11296 24812
rect 11244 24769 11253 24803
rect 11253 24769 11287 24803
rect 11287 24769 11296 24803
rect 11244 24760 11296 24769
rect 14372 24803 14424 24812
rect 14372 24769 14381 24803
rect 14381 24769 14415 24803
rect 14415 24769 14424 24803
rect 14372 24760 14424 24769
rect 15292 24803 15344 24812
rect 15292 24769 15301 24803
rect 15301 24769 15335 24803
rect 15335 24769 15344 24803
rect 19984 24871 20036 24880
rect 19984 24837 19993 24871
rect 19993 24837 20027 24871
rect 20027 24837 20036 24871
rect 19984 24828 20036 24837
rect 21272 24828 21324 24880
rect 24124 24828 24176 24880
rect 15292 24760 15344 24769
rect 18788 24760 18840 24812
rect 21640 24760 21692 24812
rect 23480 24760 23532 24812
rect 8576 24735 8628 24744
rect 8576 24701 8585 24735
rect 8585 24701 8619 24735
rect 8619 24701 8628 24735
rect 8576 24692 8628 24701
rect 8392 24624 8444 24676
rect 9128 24556 9180 24608
rect 10968 24692 11020 24744
rect 11152 24692 11204 24744
rect 12348 24692 12400 24744
rect 16028 24735 16080 24744
rect 16028 24701 16037 24735
rect 16037 24701 16071 24735
rect 16071 24701 16080 24735
rect 16028 24692 16080 24701
rect 16856 24692 16908 24744
rect 10876 24556 10928 24608
rect 13452 24599 13504 24608
rect 13452 24565 13461 24599
rect 13461 24565 13495 24599
rect 13495 24565 13504 24599
rect 13452 24556 13504 24565
rect 13544 24556 13596 24608
rect 14004 24556 14056 24608
rect 15384 24556 15436 24608
rect 15844 24556 15896 24608
rect 17408 24735 17460 24744
rect 17408 24701 17417 24735
rect 17417 24701 17451 24735
rect 17451 24701 17460 24735
rect 17408 24692 17460 24701
rect 18512 24735 18564 24744
rect 18512 24701 18521 24735
rect 18521 24701 18555 24735
rect 18555 24701 18564 24735
rect 18512 24692 18564 24701
rect 18604 24735 18656 24744
rect 18604 24701 18613 24735
rect 18613 24701 18647 24735
rect 18647 24701 18656 24735
rect 18604 24692 18656 24701
rect 19432 24692 19484 24744
rect 21548 24692 21600 24744
rect 17040 24624 17092 24676
rect 17776 24556 17828 24608
rect 17868 24556 17920 24608
rect 18788 24556 18840 24608
rect 21640 24624 21692 24676
rect 23296 24692 23348 24744
rect 23572 24735 23624 24744
rect 23572 24701 23581 24735
rect 23581 24701 23615 24735
rect 23615 24701 23624 24735
rect 23572 24692 23624 24701
rect 25320 24692 25372 24744
rect 21824 24556 21876 24608
rect 22100 24599 22152 24608
rect 22100 24565 22109 24599
rect 22109 24565 22143 24599
rect 22143 24565 22152 24599
rect 22100 24556 22152 24565
rect 23480 24556 23532 24608
rect 23664 24556 23716 24608
rect 2950 24454 3002 24506
rect 3014 24454 3066 24506
rect 3078 24454 3130 24506
rect 3142 24454 3194 24506
rect 3206 24454 3258 24506
rect 12950 24454 13002 24506
rect 13014 24454 13066 24506
rect 13078 24454 13130 24506
rect 13142 24454 13194 24506
rect 13206 24454 13258 24506
rect 22950 24454 23002 24506
rect 23014 24454 23066 24506
rect 23078 24454 23130 24506
rect 23142 24454 23194 24506
rect 23206 24454 23258 24506
rect 9404 24352 9456 24404
rect 12348 24395 12400 24404
rect 7748 24216 7800 24268
rect 9220 24148 9272 24200
rect 12348 24361 12357 24395
rect 12357 24361 12391 24395
rect 12391 24361 12400 24395
rect 12348 24352 12400 24361
rect 12716 24352 12768 24404
rect 15016 24352 15068 24404
rect 16396 24395 16448 24404
rect 16396 24361 16405 24395
rect 16405 24361 16439 24395
rect 16439 24361 16448 24395
rect 16396 24352 16448 24361
rect 19340 24352 19392 24404
rect 19708 24352 19760 24404
rect 20076 24352 20128 24404
rect 21456 24395 21508 24404
rect 21456 24361 21465 24395
rect 21465 24361 21499 24395
rect 21499 24361 21508 24395
rect 21456 24352 21508 24361
rect 16028 24284 16080 24336
rect 18512 24284 18564 24336
rect 8944 24123 8996 24132
rect 8944 24089 8953 24123
rect 8953 24089 8987 24123
rect 8987 24089 8996 24123
rect 8944 24080 8996 24089
rect 10508 24080 10560 24132
rect 9680 24012 9732 24064
rect 10140 24055 10192 24064
rect 10140 24021 10149 24055
rect 10149 24021 10183 24055
rect 10183 24021 10192 24055
rect 10140 24012 10192 24021
rect 11336 24080 11388 24132
rect 19248 24216 19300 24268
rect 23296 24284 23348 24336
rect 23940 24327 23992 24336
rect 23940 24293 23949 24327
rect 23949 24293 23983 24327
rect 23983 24293 23992 24327
rect 23940 24284 23992 24293
rect 24952 24284 25004 24336
rect 20904 24216 20956 24268
rect 23480 24216 23532 24268
rect 24124 24216 24176 24268
rect 14096 24148 14148 24200
rect 17040 24191 17092 24200
rect 17040 24157 17049 24191
rect 17049 24157 17083 24191
rect 17083 24157 17092 24191
rect 17040 24148 17092 24157
rect 18236 24148 18288 24200
rect 18880 24148 18932 24200
rect 19432 24191 19484 24200
rect 19432 24157 19441 24191
rect 19441 24157 19475 24191
rect 19475 24157 19484 24191
rect 19432 24148 19484 24157
rect 11152 24012 11204 24064
rect 17684 24012 17736 24064
rect 18236 24012 18288 24064
rect 19064 24012 19116 24064
rect 19708 24123 19760 24132
rect 19708 24089 19717 24123
rect 19717 24089 19751 24123
rect 19751 24089 19760 24123
rect 19708 24080 19760 24089
rect 21640 24080 21692 24132
rect 22192 24123 22244 24132
rect 22192 24089 22201 24123
rect 22201 24089 22235 24123
rect 22235 24089 22244 24123
rect 22192 24080 22244 24089
rect 21088 24012 21140 24064
rect 22836 24012 22888 24064
rect 24124 24055 24176 24064
rect 24124 24021 24133 24055
rect 24133 24021 24167 24055
rect 24167 24021 24176 24055
rect 24124 24012 24176 24021
rect 25228 24055 25280 24064
rect 25228 24021 25237 24055
rect 25237 24021 25271 24055
rect 25271 24021 25280 24055
rect 25228 24012 25280 24021
rect 7950 23910 8002 23962
rect 8014 23910 8066 23962
rect 8078 23910 8130 23962
rect 8142 23910 8194 23962
rect 8206 23910 8258 23962
rect 17950 23910 18002 23962
rect 18014 23910 18066 23962
rect 18078 23910 18130 23962
rect 18142 23910 18194 23962
rect 18206 23910 18258 23962
rect 10140 23808 10192 23860
rect 12716 23808 12768 23860
rect 8944 23740 8996 23792
rect 14464 23808 14516 23860
rect 17592 23808 17644 23860
rect 17776 23808 17828 23860
rect 18236 23808 18288 23860
rect 19708 23808 19760 23860
rect 7748 23672 7800 23724
rect 12624 23672 12676 23724
rect 16120 23672 16172 23724
rect 10600 23604 10652 23656
rect 13452 23604 13504 23656
rect 11888 23536 11940 23588
rect 16948 23604 17000 23656
rect 17132 23604 17184 23656
rect 16212 23536 16264 23588
rect 18512 23672 18564 23724
rect 17776 23604 17828 23656
rect 19800 23740 19852 23792
rect 22284 23740 22336 23792
rect 20352 23672 20404 23724
rect 20812 23715 20864 23724
rect 20812 23681 20821 23715
rect 20821 23681 20855 23715
rect 20855 23681 20864 23715
rect 20812 23672 20864 23681
rect 22468 23672 22520 23724
rect 23388 23740 23440 23792
rect 25228 23808 25280 23860
rect 20996 23647 21048 23656
rect 20996 23613 21005 23647
rect 21005 23613 21039 23647
rect 21039 23613 21048 23647
rect 20996 23604 21048 23613
rect 21088 23604 21140 23656
rect 22192 23604 22244 23656
rect 22284 23604 22336 23656
rect 22652 23604 22704 23656
rect 23204 23647 23256 23656
rect 23204 23613 23213 23647
rect 23213 23613 23247 23647
rect 23247 23613 23256 23647
rect 23204 23604 23256 23613
rect 23848 23604 23900 23656
rect 10232 23468 10284 23520
rect 11336 23468 11388 23520
rect 12716 23468 12768 23520
rect 14648 23511 14700 23520
rect 14648 23477 14657 23511
rect 14657 23477 14691 23511
rect 14691 23477 14700 23511
rect 14648 23468 14700 23477
rect 15108 23468 15160 23520
rect 16120 23468 16172 23520
rect 16948 23468 17000 23520
rect 18328 23468 18380 23520
rect 19892 23468 19944 23520
rect 20536 23468 20588 23520
rect 20996 23468 21048 23520
rect 21364 23468 21416 23520
rect 21640 23468 21692 23520
rect 22468 23468 22520 23520
rect 22928 23468 22980 23520
rect 24124 23468 24176 23520
rect 25136 23604 25188 23656
rect 2950 23366 3002 23418
rect 3014 23366 3066 23418
rect 3078 23366 3130 23418
rect 3142 23366 3194 23418
rect 3206 23366 3258 23418
rect 12950 23366 13002 23418
rect 13014 23366 13066 23418
rect 13078 23366 13130 23418
rect 13142 23366 13194 23418
rect 13206 23366 13258 23418
rect 22950 23366 23002 23418
rect 23014 23366 23066 23418
rect 23078 23366 23130 23418
rect 23142 23366 23194 23418
rect 23206 23366 23258 23418
rect 10968 23264 11020 23316
rect 10876 23128 10928 23180
rect 10600 23103 10652 23112
rect 10600 23069 10609 23103
rect 10609 23069 10643 23103
rect 10643 23069 10652 23103
rect 10600 23060 10652 23069
rect 9128 22992 9180 23044
rect 17132 23264 17184 23316
rect 19064 23264 19116 23316
rect 15108 23196 15160 23248
rect 18512 23196 18564 23248
rect 22652 23196 22704 23248
rect 15016 23128 15068 23180
rect 18236 23128 18288 23180
rect 18880 23128 18932 23180
rect 20076 23171 20128 23180
rect 20076 23137 20085 23171
rect 20085 23137 20119 23171
rect 20119 23137 20128 23171
rect 20076 23128 20128 23137
rect 23756 23171 23808 23180
rect 23756 23137 23765 23171
rect 23765 23137 23799 23171
rect 23799 23137 23808 23171
rect 23756 23128 23808 23137
rect 25044 23171 25096 23180
rect 25044 23137 25053 23171
rect 25053 23137 25087 23171
rect 25087 23137 25096 23171
rect 25044 23128 25096 23137
rect 25228 23171 25280 23180
rect 25228 23137 25237 23171
rect 25237 23137 25271 23171
rect 25271 23137 25280 23171
rect 25228 23128 25280 23137
rect 18788 22992 18840 23044
rect 19892 23103 19944 23112
rect 19892 23069 19901 23103
rect 19901 23069 19935 23103
rect 19935 23069 19944 23103
rect 19892 23060 19944 23069
rect 19984 23060 20036 23112
rect 22284 23060 22336 23112
rect 23848 23060 23900 23112
rect 26056 23060 26108 23112
rect 21364 22992 21416 23044
rect 25044 22992 25096 23044
rect 8484 22924 8536 22976
rect 12348 22924 12400 22976
rect 17040 22924 17092 22976
rect 18604 22924 18656 22976
rect 19524 22967 19576 22976
rect 19524 22933 19533 22967
rect 19533 22933 19567 22967
rect 19567 22933 19576 22967
rect 19524 22924 19576 22933
rect 22008 22924 22060 22976
rect 23572 22924 23624 22976
rect 24492 22924 24544 22976
rect 7950 22822 8002 22874
rect 8014 22822 8066 22874
rect 8078 22822 8130 22874
rect 8142 22822 8194 22874
rect 8206 22822 8258 22874
rect 17950 22822 18002 22874
rect 18014 22822 18066 22874
rect 18078 22822 18130 22874
rect 18142 22822 18194 22874
rect 18206 22822 18258 22874
rect 8484 22695 8536 22704
rect 8484 22661 8493 22695
rect 8493 22661 8527 22695
rect 8527 22661 8536 22695
rect 8484 22652 8536 22661
rect 9864 22720 9916 22772
rect 10232 22763 10284 22772
rect 10232 22729 10241 22763
rect 10241 22729 10275 22763
rect 10275 22729 10284 22763
rect 10232 22720 10284 22729
rect 8944 22652 8996 22704
rect 10600 22652 10652 22704
rect 7748 22584 7800 22636
rect 11796 22584 11848 22636
rect 15016 22652 15068 22704
rect 16304 22652 16356 22704
rect 17132 22720 17184 22772
rect 19708 22720 19760 22772
rect 21088 22763 21140 22772
rect 21088 22729 21097 22763
rect 21097 22729 21131 22763
rect 21131 22729 21140 22763
rect 21088 22720 21140 22729
rect 18420 22695 18472 22704
rect 18420 22661 18429 22695
rect 18429 22661 18463 22695
rect 18463 22661 18472 22695
rect 18420 22652 18472 22661
rect 19340 22652 19392 22704
rect 24860 22652 24912 22704
rect 13360 22448 13412 22500
rect 7288 22380 7340 22432
rect 9956 22423 10008 22432
rect 9956 22389 9965 22423
rect 9965 22389 9999 22423
rect 9999 22389 10008 22423
rect 9956 22380 10008 22389
rect 12808 22423 12860 22432
rect 12808 22389 12817 22423
rect 12817 22389 12851 22423
rect 12851 22389 12860 22423
rect 12808 22380 12860 22389
rect 13728 22559 13780 22568
rect 13728 22525 13737 22559
rect 13737 22525 13771 22559
rect 13771 22525 13780 22559
rect 13728 22516 13780 22525
rect 14464 22516 14516 22568
rect 19248 22584 19300 22636
rect 20076 22584 20128 22636
rect 22376 22584 22428 22636
rect 17592 22516 17644 22568
rect 18788 22516 18840 22568
rect 20628 22516 20680 22568
rect 16120 22448 16172 22500
rect 19984 22448 20036 22500
rect 20904 22448 20956 22500
rect 24768 22559 24820 22568
rect 24768 22525 24777 22559
rect 24777 22525 24811 22559
rect 24811 22525 24820 22559
rect 24768 22516 24820 22525
rect 15200 22423 15252 22432
rect 15200 22389 15209 22423
rect 15209 22389 15243 22423
rect 15243 22389 15252 22423
rect 15200 22380 15252 22389
rect 17408 22380 17460 22432
rect 17776 22380 17828 22432
rect 18236 22423 18288 22432
rect 18236 22389 18245 22423
rect 18245 22389 18279 22423
rect 18279 22389 18288 22423
rect 18236 22380 18288 22389
rect 18420 22380 18472 22432
rect 19064 22380 19116 22432
rect 20352 22380 20404 22432
rect 20720 22423 20772 22432
rect 20720 22389 20729 22423
rect 20729 22389 20763 22423
rect 20763 22389 20772 22423
rect 20720 22380 20772 22389
rect 2950 22278 3002 22330
rect 3014 22278 3066 22330
rect 3078 22278 3130 22330
rect 3142 22278 3194 22330
rect 3206 22278 3258 22330
rect 12950 22278 13002 22330
rect 13014 22278 13066 22330
rect 13078 22278 13130 22330
rect 13142 22278 13194 22330
rect 13206 22278 13258 22330
rect 22950 22278 23002 22330
rect 23014 22278 23066 22330
rect 23078 22278 23130 22330
rect 23142 22278 23194 22330
rect 23206 22278 23258 22330
rect 9404 22176 9456 22228
rect 9956 22176 10008 22228
rect 9496 22108 9548 22160
rect 12440 22176 12492 22228
rect 12716 22176 12768 22228
rect 13728 22176 13780 22228
rect 15660 22176 15712 22228
rect 18236 22176 18288 22228
rect 7564 22040 7616 22092
rect 9864 22040 9916 22092
rect 12440 22040 12492 22092
rect 12808 22040 12860 22092
rect 15200 22108 15252 22160
rect 18420 22151 18472 22160
rect 18420 22117 18429 22151
rect 18429 22117 18463 22151
rect 18463 22117 18472 22151
rect 18420 22108 18472 22117
rect 18788 22176 18840 22228
rect 21180 22176 21232 22228
rect 23388 22176 23440 22228
rect 23848 22219 23900 22228
rect 23848 22185 23857 22219
rect 23857 22185 23891 22219
rect 23891 22185 23900 22219
rect 23848 22176 23900 22185
rect 15384 22083 15436 22092
rect 15384 22049 15393 22083
rect 15393 22049 15427 22083
rect 15427 22049 15436 22083
rect 15384 22040 15436 22049
rect 15476 22083 15528 22092
rect 15476 22049 15485 22083
rect 15485 22049 15519 22083
rect 15519 22049 15528 22083
rect 15476 22040 15528 22049
rect 16028 22040 16080 22092
rect 17040 22040 17092 22092
rect 17592 22054 17644 22106
rect 20444 22108 20496 22160
rect 8208 21972 8260 22024
rect 6276 21836 6328 21888
rect 11704 22015 11756 22024
rect 11704 21981 11713 22015
rect 11713 21981 11747 22015
rect 11747 21981 11756 22015
rect 11704 21972 11756 21981
rect 11980 21972 12032 22024
rect 20812 22040 20864 22092
rect 23296 22040 23348 22092
rect 24676 22040 24728 22092
rect 25412 22108 25464 22160
rect 8484 21836 8536 21888
rect 9496 21879 9548 21888
rect 9496 21845 9505 21879
rect 9505 21845 9539 21879
rect 9539 21845 9548 21879
rect 9496 21836 9548 21845
rect 10048 21836 10100 21888
rect 10600 21879 10652 21888
rect 10600 21845 10609 21879
rect 10609 21845 10643 21879
rect 10643 21845 10652 21879
rect 10600 21836 10652 21845
rect 11244 21836 11296 21888
rect 13360 21904 13412 21956
rect 11612 21836 11664 21888
rect 12532 21879 12584 21888
rect 12532 21845 12541 21879
rect 12541 21845 12575 21879
rect 12575 21845 12584 21879
rect 12532 21836 12584 21845
rect 14924 21879 14976 21888
rect 14924 21845 14933 21879
rect 14933 21845 14967 21879
rect 14967 21845 14976 21879
rect 14924 21836 14976 21845
rect 15292 21879 15344 21888
rect 15292 21845 15301 21879
rect 15301 21845 15335 21879
rect 15335 21845 15344 21879
rect 15292 21836 15344 21845
rect 18420 21904 18472 21956
rect 17776 21836 17828 21888
rect 21272 21972 21324 22024
rect 23112 21972 23164 22024
rect 18604 21836 18656 21888
rect 19340 21879 19392 21888
rect 19340 21845 19349 21879
rect 19349 21845 19383 21879
rect 19383 21845 19392 21879
rect 19340 21836 19392 21845
rect 20352 21904 20404 21956
rect 21824 21947 21876 21956
rect 21824 21913 21833 21947
rect 21833 21913 21867 21947
rect 21867 21913 21876 21947
rect 21824 21904 21876 21913
rect 23204 21904 23256 21956
rect 20168 21836 20220 21888
rect 20628 21836 20680 21888
rect 24584 21879 24636 21888
rect 24584 21845 24593 21879
rect 24593 21845 24627 21879
rect 24627 21845 24636 21879
rect 24584 21836 24636 21845
rect 7950 21734 8002 21786
rect 8014 21734 8066 21786
rect 8078 21734 8130 21786
rect 8142 21734 8194 21786
rect 8206 21734 8258 21786
rect 17950 21734 18002 21786
rect 18014 21734 18066 21786
rect 18078 21734 18130 21786
rect 18142 21734 18194 21786
rect 18206 21734 18258 21786
rect 9772 21632 9824 21684
rect 14648 21632 14700 21684
rect 15660 21675 15712 21684
rect 15660 21641 15669 21675
rect 15669 21641 15703 21675
rect 15703 21641 15712 21675
rect 15660 21632 15712 21641
rect 19248 21675 19300 21684
rect 19248 21641 19257 21675
rect 19257 21641 19291 21675
rect 19291 21641 19300 21675
rect 19248 21632 19300 21641
rect 20168 21632 20220 21684
rect 20536 21632 20588 21684
rect 22560 21632 22612 21684
rect 22744 21632 22796 21684
rect 8300 21564 8352 21616
rect 9864 21607 9916 21616
rect 9864 21573 9873 21607
rect 9873 21573 9907 21607
rect 9907 21573 9916 21607
rect 9864 21564 9916 21573
rect 13636 21564 13688 21616
rect 14924 21564 14976 21616
rect 12716 21496 12768 21548
rect 7564 21471 7616 21480
rect 7564 21437 7573 21471
rect 7573 21437 7607 21471
rect 7607 21437 7616 21471
rect 7564 21428 7616 21437
rect 8576 21428 8628 21480
rect 9588 21471 9640 21480
rect 9588 21437 9597 21471
rect 9597 21437 9631 21471
rect 9631 21437 9640 21471
rect 9588 21428 9640 21437
rect 10416 21428 10468 21480
rect 9404 21360 9456 21412
rect 11152 21428 11204 21480
rect 12624 21428 12676 21480
rect 13820 21428 13872 21480
rect 14096 21428 14148 21480
rect 15476 21496 15528 21548
rect 16580 21496 16632 21548
rect 19064 21564 19116 21616
rect 18972 21496 19024 21548
rect 23112 21564 23164 21616
rect 23204 21564 23256 21616
rect 24032 21564 24084 21616
rect 24124 21564 24176 21616
rect 22008 21496 22060 21548
rect 22560 21496 22612 21548
rect 23296 21539 23348 21548
rect 23296 21505 23305 21539
rect 23305 21505 23339 21539
rect 23339 21505 23348 21539
rect 23296 21496 23348 21505
rect 15108 21428 15160 21480
rect 19340 21428 19392 21480
rect 20904 21428 20956 21480
rect 11796 21360 11848 21412
rect 12716 21292 12768 21344
rect 15384 21360 15436 21412
rect 14740 21292 14792 21344
rect 15476 21292 15528 21344
rect 18604 21360 18656 21412
rect 21088 21360 21140 21412
rect 22928 21428 22980 21480
rect 25412 21428 25464 21480
rect 20444 21292 20496 21344
rect 21732 21292 21784 21344
rect 23388 21292 23440 21344
rect 24124 21292 24176 21344
rect 2950 21190 3002 21242
rect 3014 21190 3066 21242
rect 3078 21190 3130 21242
rect 3142 21190 3194 21242
rect 3206 21190 3258 21242
rect 12950 21190 13002 21242
rect 13014 21190 13066 21242
rect 13078 21190 13130 21242
rect 13142 21190 13194 21242
rect 13206 21190 13258 21242
rect 22950 21190 23002 21242
rect 23014 21190 23066 21242
rect 23078 21190 23130 21242
rect 23142 21190 23194 21242
rect 23206 21190 23258 21242
rect 8576 21131 8628 21140
rect 8576 21097 8585 21131
rect 8585 21097 8619 21131
rect 8619 21097 8628 21131
rect 8576 21088 8628 21097
rect 10692 21088 10744 21140
rect 5264 21020 5316 21072
rect 12808 21088 12860 21140
rect 13544 21088 13596 21140
rect 15200 21088 15252 21140
rect 16120 21088 16172 21140
rect 16488 21088 16540 21140
rect 17040 21088 17092 21140
rect 19984 21088 20036 21140
rect 20260 21088 20312 21140
rect 22008 21131 22060 21140
rect 22008 21097 22017 21131
rect 22017 21097 22051 21131
rect 22051 21097 22060 21131
rect 22008 21088 22060 21097
rect 15108 21020 15160 21072
rect 10232 20995 10284 21004
rect 10232 20961 10241 20995
rect 10241 20961 10275 20995
rect 10275 20961 10284 20995
rect 10232 20952 10284 20961
rect 11152 20995 11204 21004
rect 11152 20961 11161 20995
rect 11161 20961 11195 20995
rect 11195 20961 11204 20995
rect 11152 20952 11204 20961
rect 13360 20995 13412 21004
rect 13360 20961 13369 20995
rect 13369 20961 13403 20995
rect 13403 20961 13412 20995
rect 13360 20952 13412 20961
rect 15476 20995 15528 21004
rect 15476 20961 15485 20995
rect 15485 20961 15519 20995
rect 15519 20961 15528 20995
rect 15476 20952 15528 20961
rect 16028 20952 16080 21004
rect 18328 20952 18380 21004
rect 19984 20995 20036 21004
rect 19984 20961 19993 20995
rect 19993 20961 20027 20995
rect 20027 20961 20036 20995
rect 19984 20952 20036 20961
rect 8484 20884 8536 20936
rect 9496 20884 9548 20936
rect 15200 20927 15252 20936
rect 15200 20893 15209 20927
rect 15209 20893 15243 20927
rect 15243 20893 15252 20927
rect 15200 20884 15252 20893
rect 18420 20884 18472 20936
rect 19892 20884 19944 20936
rect 21088 20884 21140 20936
rect 22192 21020 22244 21072
rect 11428 20859 11480 20868
rect 11428 20825 11437 20859
rect 11437 20825 11471 20859
rect 11471 20825 11480 20859
rect 11428 20816 11480 20825
rect 8300 20748 8352 20800
rect 8484 20748 8536 20800
rect 10232 20748 10284 20800
rect 10968 20748 11020 20800
rect 13360 20816 13412 20868
rect 13636 20816 13688 20868
rect 19708 20816 19760 20868
rect 14096 20748 14148 20800
rect 14740 20748 14792 20800
rect 19340 20748 19392 20800
rect 19800 20748 19852 20800
rect 22008 20816 22060 20868
rect 20904 20748 20956 20800
rect 21088 20791 21140 20800
rect 21088 20757 21097 20791
rect 21097 20757 21131 20791
rect 21131 20757 21140 20791
rect 21088 20748 21140 20757
rect 21364 20748 21416 20800
rect 24860 20952 24912 21004
rect 22652 20927 22704 20936
rect 22652 20893 22661 20927
rect 22661 20893 22695 20927
rect 22695 20893 22704 20927
rect 22652 20884 22704 20893
rect 23940 20884 23992 20936
rect 23756 20816 23808 20868
rect 25504 20816 25556 20868
rect 22652 20748 22704 20800
rect 24860 20748 24912 20800
rect 24952 20791 25004 20800
rect 24952 20757 24961 20791
rect 24961 20757 24995 20791
rect 24995 20757 25004 20791
rect 24952 20748 25004 20757
rect 25872 20748 25924 20800
rect 7950 20646 8002 20698
rect 8014 20646 8066 20698
rect 8078 20646 8130 20698
rect 8142 20646 8194 20698
rect 8206 20646 8258 20698
rect 17950 20646 18002 20698
rect 18014 20646 18066 20698
rect 18078 20646 18130 20698
rect 18142 20646 18194 20698
rect 18206 20646 18258 20698
rect 9312 20544 9364 20596
rect 11428 20544 11480 20596
rect 10140 20476 10192 20528
rect 12716 20476 12768 20528
rect 13360 20476 13412 20528
rect 15844 20544 15896 20596
rect 19248 20544 19300 20596
rect 19892 20544 19944 20596
rect 21824 20544 21876 20596
rect 25228 20544 25280 20596
rect 8300 20408 8352 20460
rect 9036 20408 9088 20460
rect 11704 20451 11756 20460
rect 11704 20417 11713 20451
rect 11713 20417 11747 20451
rect 11747 20417 11756 20451
rect 11704 20408 11756 20417
rect 7656 20272 7708 20324
rect 12624 20340 12676 20392
rect 13544 20340 13596 20392
rect 18604 20408 18656 20460
rect 19616 20476 19668 20528
rect 22008 20519 22060 20528
rect 22008 20485 22017 20519
rect 22017 20485 22051 20519
rect 22051 20485 22060 20519
rect 22008 20476 22060 20485
rect 24124 20476 24176 20528
rect 14648 20340 14700 20392
rect 7196 20204 7248 20256
rect 18788 20340 18840 20392
rect 19340 20408 19392 20460
rect 21180 20408 21232 20460
rect 22744 20408 22796 20460
rect 19616 20340 19668 20392
rect 23204 20340 23256 20392
rect 23296 20340 23348 20392
rect 19432 20272 19484 20324
rect 19892 20272 19944 20324
rect 18696 20204 18748 20256
rect 18972 20204 19024 20256
rect 19064 20247 19116 20256
rect 19064 20213 19073 20247
rect 19073 20213 19107 20247
rect 19107 20213 19116 20247
rect 19064 20204 19116 20213
rect 19616 20247 19668 20256
rect 19616 20213 19625 20247
rect 19625 20213 19659 20247
rect 19659 20213 19668 20247
rect 19616 20204 19668 20213
rect 25044 20204 25096 20256
rect 2950 20102 3002 20154
rect 3014 20102 3066 20154
rect 3078 20102 3130 20154
rect 3142 20102 3194 20154
rect 3206 20102 3258 20154
rect 12950 20102 13002 20154
rect 13014 20102 13066 20154
rect 13078 20102 13130 20154
rect 13142 20102 13194 20154
rect 13206 20102 13258 20154
rect 22950 20102 23002 20154
rect 23014 20102 23066 20154
rect 23078 20102 23130 20154
rect 23142 20102 23194 20154
rect 23206 20102 23258 20154
rect 8484 20043 8536 20052
rect 8484 20009 8493 20043
rect 8493 20009 8527 20043
rect 8527 20009 8536 20043
rect 8484 20000 8536 20009
rect 9864 20000 9916 20052
rect 10968 20000 11020 20052
rect 6736 19864 6788 19916
rect 8484 19728 8536 19780
rect 9128 19932 9180 19984
rect 11704 19864 11756 19916
rect 9128 19839 9180 19848
rect 9128 19805 9137 19839
rect 9137 19805 9171 19839
rect 9171 19805 9180 19839
rect 9128 19796 9180 19805
rect 12348 19839 12400 19848
rect 12348 19805 12357 19839
rect 12357 19805 12391 19839
rect 12391 19805 12400 19839
rect 12348 19796 12400 19805
rect 12624 19796 12676 19848
rect 15936 19932 15988 19984
rect 22192 20000 22244 20052
rect 24952 20000 25004 20052
rect 25320 20000 25372 20052
rect 17408 19932 17460 19984
rect 17776 19932 17828 19984
rect 16580 19864 16632 19916
rect 17868 19864 17920 19916
rect 19892 19907 19944 19916
rect 19892 19873 19901 19907
rect 19901 19873 19935 19907
rect 19935 19873 19944 19907
rect 19892 19864 19944 19873
rect 19156 19796 19208 19848
rect 9864 19728 9916 19780
rect 7012 19660 7064 19712
rect 7288 19660 7340 19712
rect 8300 19660 8352 19712
rect 8392 19660 8444 19712
rect 9496 19660 9548 19712
rect 9680 19660 9732 19712
rect 14556 19771 14608 19780
rect 14556 19737 14565 19771
rect 14565 19737 14599 19771
rect 14599 19737 14608 19771
rect 14556 19728 14608 19737
rect 10968 19660 11020 19712
rect 13084 19660 13136 19712
rect 13360 19660 13412 19712
rect 18420 19728 18472 19780
rect 20168 19771 20220 19780
rect 20168 19737 20177 19771
rect 20177 19737 20211 19771
rect 20211 19737 20220 19771
rect 20168 19728 20220 19737
rect 25136 19796 25188 19848
rect 16764 19660 16816 19712
rect 19616 19703 19668 19712
rect 19616 19669 19625 19703
rect 19625 19669 19659 19703
rect 19659 19669 19668 19703
rect 22284 19728 22336 19780
rect 22376 19771 22428 19780
rect 22376 19737 22385 19771
rect 22385 19737 22419 19771
rect 22419 19737 22428 19771
rect 22376 19728 22428 19737
rect 24124 19728 24176 19780
rect 19616 19660 19668 19669
rect 22008 19660 22060 19712
rect 23940 19660 23992 19712
rect 7950 19558 8002 19610
rect 8014 19558 8066 19610
rect 8078 19558 8130 19610
rect 8142 19558 8194 19610
rect 8206 19558 8258 19610
rect 17950 19558 18002 19610
rect 18014 19558 18066 19610
rect 18078 19558 18130 19610
rect 18142 19558 18194 19610
rect 18206 19558 18258 19610
rect 6828 19320 6880 19372
rect 7564 19456 7616 19508
rect 9128 19456 9180 19508
rect 9312 19456 9364 19508
rect 9496 19499 9548 19508
rect 9496 19465 9505 19499
rect 9505 19465 9539 19499
rect 9539 19465 9548 19499
rect 9496 19456 9548 19465
rect 10324 19456 10376 19508
rect 12716 19456 12768 19508
rect 12808 19456 12860 19508
rect 10324 19320 10376 19372
rect 12624 19388 12676 19440
rect 13084 19388 13136 19440
rect 13912 19388 13964 19440
rect 14648 19388 14700 19440
rect 16028 19456 16080 19508
rect 16396 19456 16448 19508
rect 16764 19456 16816 19508
rect 16948 19456 17000 19508
rect 18788 19499 18840 19508
rect 18788 19465 18797 19499
rect 18797 19465 18831 19499
rect 18831 19465 18840 19499
rect 18788 19456 18840 19465
rect 18972 19456 19024 19508
rect 20444 19499 20496 19508
rect 20444 19465 20453 19499
rect 20453 19465 20487 19499
rect 20487 19465 20496 19499
rect 20444 19456 20496 19465
rect 20720 19456 20772 19508
rect 21456 19456 21508 19508
rect 24492 19456 24544 19508
rect 9772 19252 9824 19304
rect 11152 19295 11204 19304
rect 3516 19116 3568 19168
rect 10508 19184 10560 19236
rect 11152 19261 11161 19295
rect 11161 19261 11195 19295
rect 11195 19261 11204 19295
rect 11152 19252 11204 19261
rect 20260 19388 20312 19440
rect 24124 19388 24176 19440
rect 10968 19184 11020 19236
rect 14096 19184 14148 19236
rect 17776 19320 17828 19372
rect 19248 19320 19300 19372
rect 22468 19320 22520 19372
rect 22560 19363 22612 19372
rect 22560 19329 22569 19363
rect 22569 19329 22603 19363
rect 22603 19329 22612 19363
rect 22560 19320 22612 19329
rect 16580 19252 16632 19304
rect 22008 19252 22060 19304
rect 22744 19295 22796 19304
rect 22744 19261 22753 19295
rect 22753 19261 22787 19295
rect 22787 19261 22796 19295
rect 22744 19252 22796 19261
rect 23296 19252 23348 19304
rect 25228 19252 25280 19304
rect 21088 19184 21140 19236
rect 11336 19116 11388 19168
rect 14372 19116 14424 19168
rect 18788 19116 18840 19168
rect 19248 19159 19300 19168
rect 19248 19125 19257 19159
rect 19257 19125 19291 19159
rect 19291 19125 19300 19159
rect 19248 19116 19300 19125
rect 19708 19159 19760 19168
rect 19708 19125 19717 19159
rect 19717 19125 19751 19159
rect 19751 19125 19760 19159
rect 19708 19116 19760 19125
rect 21272 19159 21324 19168
rect 21272 19125 21281 19159
rect 21281 19125 21315 19159
rect 21315 19125 21324 19159
rect 21272 19116 21324 19125
rect 22744 19116 22796 19168
rect 23756 19116 23808 19168
rect 24124 19116 24176 19168
rect 25136 19159 25188 19168
rect 25136 19125 25145 19159
rect 25145 19125 25179 19159
rect 25179 19125 25188 19159
rect 25136 19116 25188 19125
rect 2950 19014 3002 19066
rect 3014 19014 3066 19066
rect 3078 19014 3130 19066
rect 3142 19014 3194 19066
rect 3206 19014 3258 19066
rect 12950 19014 13002 19066
rect 13014 19014 13066 19066
rect 13078 19014 13130 19066
rect 13142 19014 13194 19066
rect 13206 19014 13258 19066
rect 22950 19014 23002 19066
rect 23014 19014 23066 19066
rect 23078 19014 23130 19066
rect 23142 19014 23194 19066
rect 23206 19014 23258 19066
rect 11336 18912 11388 18964
rect 22192 18912 22244 18964
rect 25412 18912 25464 18964
rect 6828 18819 6880 18828
rect 6828 18785 6837 18819
rect 6837 18785 6871 18819
rect 6871 18785 6880 18819
rect 6828 18776 6880 18785
rect 7196 18776 7248 18828
rect 8300 18776 8352 18828
rect 14096 18844 14148 18896
rect 8392 18708 8444 18760
rect 8760 18708 8812 18760
rect 10784 18708 10836 18760
rect 10968 18708 11020 18760
rect 11520 18819 11572 18828
rect 11520 18785 11529 18819
rect 11529 18785 11563 18819
rect 11563 18785 11572 18819
rect 11520 18776 11572 18785
rect 7380 18572 7432 18624
rect 11244 18640 11296 18692
rect 12532 18708 12584 18760
rect 19064 18844 19116 18896
rect 20168 18844 20220 18896
rect 14740 18776 14792 18828
rect 16304 18776 16356 18828
rect 17132 18776 17184 18828
rect 17224 18819 17276 18828
rect 17224 18785 17233 18819
rect 17233 18785 17267 18819
rect 17267 18785 17276 18819
rect 17224 18776 17276 18785
rect 17776 18776 17828 18828
rect 15292 18708 15344 18760
rect 17500 18708 17552 18760
rect 17592 18708 17644 18760
rect 18788 18776 18840 18828
rect 18604 18708 18656 18760
rect 18696 18708 18748 18760
rect 20720 18751 20772 18760
rect 20720 18717 20729 18751
rect 20729 18717 20763 18751
rect 20763 18717 20772 18751
rect 20720 18708 20772 18717
rect 21180 18708 21232 18760
rect 22560 18776 22612 18828
rect 23388 18776 23440 18828
rect 25320 18708 25372 18760
rect 8484 18572 8536 18624
rect 9496 18572 9548 18624
rect 11704 18572 11756 18624
rect 12624 18640 12676 18692
rect 15752 18640 15804 18692
rect 20812 18640 20864 18692
rect 21916 18640 21968 18692
rect 22744 18640 22796 18692
rect 13452 18615 13504 18624
rect 13452 18581 13461 18615
rect 13461 18581 13495 18615
rect 13495 18581 13504 18615
rect 13452 18572 13504 18581
rect 13636 18615 13688 18624
rect 13636 18581 13645 18615
rect 13645 18581 13679 18615
rect 13679 18581 13688 18615
rect 13636 18572 13688 18581
rect 14004 18572 14056 18624
rect 14648 18615 14700 18624
rect 14648 18581 14657 18615
rect 14657 18581 14691 18615
rect 14691 18581 14700 18615
rect 14648 18572 14700 18581
rect 16120 18572 16172 18624
rect 17040 18572 17092 18624
rect 17132 18615 17184 18624
rect 17132 18581 17141 18615
rect 17141 18581 17175 18615
rect 17175 18581 17184 18615
rect 17132 18572 17184 18581
rect 19708 18572 19760 18624
rect 20076 18615 20128 18624
rect 20076 18581 20085 18615
rect 20085 18581 20119 18615
rect 20119 18581 20128 18615
rect 20076 18572 20128 18581
rect 20444 18615 20496 18624
rect 20444 18581 20453 18615
rect 20453 18581 20487 18615
rect 20487 18581 20496 18615
rect 20444 18572 20496 18581
rect 22192 18572 22244 18624
rect 7950 18470 8002 18522
rect 8014 18470 8066 18522
rect 8078 18470 8130 18522
rect 8142 18470 8194 18522
rect 8206 18470 8258 18522
rect 17950 18470 18002 18522
rect 18014 18470 18066 18522
rect 18078 18470 18130 18522
rect 18142 18470 18194 18522
rect 18206 18470 18258 18522
rect 8668 18368 8720 18420
rect 9588 18368 9640 18420
rect 11520 18368 11572 18420
rect 11704 18411 11756 18420
rect 11704 18377 11713 18411
rect 11713 18377 11747 18411
rect 11747 18377 11756 18411
rect 11704 18368 11756 18377
rect 12716 18368 12768 18420
rect 13636 18411 13688 18420
rect 13636 18377 13645 18411
rect 13645 18377 13679 18411
rect 13679 18377 13688 18411
rect 13636 18368 13688 18377
rect 14556 18368 14608 18420
rect 15200 18368 15252 18420
rect 9864 18300 9916 18352
rect 11152 18343 11204 18352
rect 11152 18309 11161 18343
rect 11161 18309 11195 18343
rect 11195 18309 11204 18343
rect 11152 18300 11204 18309
rect 8300 18275 8352 18284
rect 8300 18241 8309 18275
rect 8309 18241 8343 18275
rect 8343 18241 8352 18275
rect 8300 18232 8352 18241
rect 8392 18207 8444 18216
rect 8392 18173 8401 18207
rect 8401 18173 8435 18207
rect 8435 18173 8444 18207
rect 8392 18164 8444 18173
rect 7748 18096 7800 18148
rect 9128 18207 9180 18216
rect 9128 18173 9137 18207
rect 9137 18173 9171 18207
rect 9171 18173 9180 18207
rect 9128 18164 9180 18173
rect 9404 18164 9456 18216
rect 5172 18028 5224 18080
rect 13636 18232 13688 18284
rect 13912 18232 13964 18284
rect 16212 18300 16264 18352
rect 20076 18368 20128 18420
rect 22376 18368 22428 18420
rect 17868 18300 17920 18352
rect 18604 18300 18656 18352
rect 13820 18096 13872 18148
rect 11520 18028 11572 18080
rect 12532 18028 12584 18080
rect 15752 18207 15804 18216
rect 15752 18173 15761 18207
rect 15761 18173 15795 18207
rect 15795 18173 15804 18207
rect 15752 18164 15804 18173
rect 16856 18275 16908 18284
rect 16856 18241 16865 18275
rect 16865 18241 16899 18275
rect 16899 18241 16908 18275
rect 16856 18232 16908 18241
rect 20996 18300 21048 18352
rect 21640 18300 21692 18352
rect 25688 18368 25740 18420
rect 23572 18343 23624 18352
rect 23572 18309 23581 18343
rect 23581 18309 23615 18343
rect 23615 18309 23624 18343
rect 23572 18300 23624 18309
rect 20260 18275 20312 18284
rect 20260 18241 20269 18275
rect 20269 18241 20303 18275
rect 20303 18241 20312 18275
rect 20260 18232 20312 18241
rect 22008 18275 22060 18284
rect 22008 18241 22017 18275
rect 22017 18241 22051 18275
rect 22051 18241 22060 18275
rect 22008 18232 22060 18241
rect 19248 18164 19300 18216
rect 20444 18164 20496 18216
rect 20996 18164 21048 18216
rect 22192 18164 22244 18216
rect 22284 18164 22336 18216
rect 23296 18207 23348 18216
rect 23296 18173 23305 18207
rect 23305 18173 23339 18207
rect 23339 18173 23348 18207
rect 23296 18164 23348 18173
rect 17224 18028 17276 18080
rect 21916 18096 21968 18148
rect 24124 18164 24176 18216
rect 18604 18071 18656 18080
rect 18604 18037 18613 18071
rect 18613 18037 18647 18071
rect 18647 18037 18656 18071
rect 18604 18028 18656 18037
rect 18880 18028 18932 18080
rect 19616 18028 19668 18080
rect 20076 18071 20128 18080
rect 20076 18037 20085 18071
rect 20085 18037 20119 18071
rect 20119 18037 20128 18071
rect 20076 18028 20128 18037
rect 20996 18028 21048 18080
rect 21364 18071 21416 18080
rect 21364 18037 21373 18071
rect 21373 18037 21407 18071
rect 21407 18037 21416 18071
rect 21364 18028 21416 18037
rect 23388 18028 23440 18080
rect 2950 17926 3002 17978
rect 3014 17926 3066 17978
rect 3078 17926 3130 17978
rect 3142 17926 3194 17978
rect 3206 17926 3258 17978
rect 12950 17926 13002 17978
rect 13014 17926 13066 17978
rect 13078 17926 13130 17978
rect 13142 17926 13194 17978
rect 13206 17926 13258 17978
rect 22950 17926 23002 17978
rect 23014 17926 23066 17978
rect 23078 17926 23130 17978
rect 23142 17926 23194 17978
rect 23206 17926 23258 17978
rect 8760 17867 8812 17876
rect 8760 17833 8769 17867
rect 8769 17833 8803 17867
rect 8803 17833 8812 17867
rect 8760 17824 8812 17833
rect 10692 17824 10744 17876
rect 10876 17824 10928 17876
rect 11060 17756 11112 17808
rect 11244 17824 11296 17876
rect 13452 17824 13504 17876
rect 17316 17824 17368 17876
rect 11336 17756 11388 17808
rect 12164 17756 12216 17808
rect 12440 17756 12492 17808
rect 9404 17688 9456 17740
rect 10876 17620 10928 17672
rect 11060 17620 11112 17672
rect 12808 17663 12860 17672
rect 12808 17629 12817 17663
rect 12817 17629 12851 17663
rect 12851 17629 12860 17663
rect 12808 17620 12860 17629
rect 3792 17484 3844 17536
rect 11244 17552 11296 17604
rect 12072 17552 12124 17604
rect 12164 17552 12216 17604
rect 13820 17756 13872 17808
rect 19432 17824 19484 17876
rect 21180 17867 21232 17876
rect 21180 17833 21189 17867
rect 21189 17833 21223 17867
rect 21223 17833 21232 17867
rect 21180 17824 21232 17833
rect 21640 17867 21692 17876
rect 21640 17833 21649 17867
rect 21649 17833 21683 17867
rect 21683 17833 21692 17867
rect 21640 17824 21692 17833
rect 21824 17824 21876 17876
rect 26148 17824 26200 17876
rect 14648 17688 14700 17740
rect 16672 17688 16724 17740
rect 17868 17756 17920 17808
rect 19156 17756 19208 17808
rect 18512 17688 18564 17740
rect 18604 17731 18656 17740
rect 18604 17697 18613 17731
rect 18613 17697 18647 17731
rect 18647 17697 18656 17731
rect 18604 17688 18656 17697
rect 18788 17688 18840 17740
rect 24860 17688 24912 17740
rect 24952 17688 25004 17740
rect 25136 17731 25188 17740
rect 25136 17697 25145 17731
rect 25145 17697 25179 17731
rect 25179 17697 25188 17731
rect 25136 17688 25188 17697
rect 16764 17620 16816 17672
rect 18328 17620 18380 17672
rect 21916 17620 21968 17672
rect 22652 17663 22704 17672
rect 22652 17629 22661 17663
rect 22661 17629 22695 17663
rect 22695 17629 22704 17663
rect 22652 17620 22704 17629
rect 14004 17552 14056 17604
rect 15200 17552 15252 17604
rect 15568 17552 15620 17604
rect 7840 17484 7892 17536
rect 9772 17484 9824 17536
rect 11520 17527 11572 17536
rect 11520 17493 11529 17527
rect 11529 17493 11563 17527
rect 11563 17493 11572 17527
rect 11520 17484 11572 17493
rect 13452 17527 13504 17536
rect 13452 17493 13461 17527
rect 13461 17493 13495 17527
rect 13495 17493 13504 17527
rect 13452 17484 13504 17493
rect 13912 17484 13964 17536
rect 15660 17527 15712 17536
rect 15660 17493 15669 17527
rect 15669 17493 15703 17527
rect 15703 17493 15712 17527
rect 15660 17484 15712 17493
rect 16764 17484 16816 17536
rect 19248 17552 19300 17604
rect 19340 17552 19392 17604
rect 20996 17552 21048 17604
rect 21364 17552 21416 17604
rect 18788 17484 18840 17536
rect 22100 17527 22152 17536
rect 22100 17493 22109 17527
rect 22109 17493 22143 17527
rect 22143 17493 22152 17527
rect 22100 17484 22152 17493
rect 24584 17527 24636 17536
rect 24584 17493 24593 17527
rect 24593 17493 24627 17527
rect 24627 17493 24636 17527
rect 24584 17484 24636 17493
rect 24952 17527 25004 17536
rect 24952 17493 24961 17527
rect 24961 17493 24995 17527
rect 24995 17493 25004 17527
rect 24952 17484 25004 17493
rect 7950 17382 8002 17434
rect 8014 17382 8066 17434
rect 8078 17382 8130 17434
rect 8142 17382 8194 17434
rect 8206 17382 8258 17434
rect 17950 17382 18002 17434
rect 18014 17382 18066 17434
rect 18078 17382 18130 17434
rect 18142 17382 18194 17434
rect 18206 17382 18258 17434
rect 7840 17280 7892 17332
rect 9496 17323 9548 17332
rect 9496 17289 9505 17323
rect 9505 17289 9539 17323
rect 9539 17289 9548 17323
rect 9496 17280 9548 17289
rect 8576 17212 8628 17264
rect 11612 17280 11664 17332
rect 12256 17212 12308 17264
rect 13912 17280 13964 17332
rect 13544 17212 13596 17264
rect 7656 17144 7708 17196
rect 9220 17144 9272 17196
rect 11704 17144 11756 17196
rect 12072 17187 12124 17196
rect 12072 17153 12081 17187
rect 12081 17153 12115 17187
rect 12115 17153 12124 17187
rect 12072 17144 12124 17153
rect 15108 17280 15160 17332
rect 19248 17280 19300 17332
rect 21180 17323 21232 17332
rect 21180 17289 21189 17323
rect 21189 17289 21223 17323
rect 21223 17289 21232 17323
rect 21180 17280 21232 17289
rect 15200 17212 15252 17264
rect 17316 17255 17368 17264
rect 17316 17221 17325 17255
rect 17325 17221 17359 17255
rect 17359 17221 17368 17255
rect 17316 17212 17368 17221
rect 19524 17212 19576 17264
rect 20812 17212 20864 17264
rect 16856 17144 16908 17196
rect 18328 17144 18380 17196
rect 18604 17144 18656 17196
rect 19248 17144 19300 17196
rect 9312 17008 9364 17060
rect 12164 17119 12216 17128
rect 12164 17085 12173 17119
rect 12173 17085 12207 17119
rect 12207 17085 12216 17119
rect 12164 17076 12216 17085
rect 11152 17008 11204 17060
rect 13360 17119 13412 17128
rect 13360 17085 13369 17119
rect 13369 17085 13403 17119
rect 13403 17085 13412 17119
rect 13360 17076 13412 17085
rect 13728 17076 13780 17128
rect 15476 17076 15528 17128
rect 16304 17076 16356 17128
rect 22192 17187 22244 17196
rect 22192 17153 22201 17187
rect 22201 17153 22235 17187
rect 22235 17153 22244 17187
rect 22192 17144 22244 17153
rect 24860 17212 24912 17264
rect 12348 17008 12400 17060
rect 16212 17051 16264 17060
rect 16212 17017 16221 17051
rect 16221 17017 16255 17051
rect 16255 17017 16264 17051
rect 16212 17008 16264 17017
rect 16580 17008 16632 17060
rect 23388 17076 23440 17128
rect 24768 17119 24820 17128
rect 24768 17085 24777 17119
rect 24777 17085 24811 17119
rect 24811 17085 24820 17119
rect 24768 17076 24820 17085
rect 24584 17008 24636 17060
rect 7840 16940 7892 16992
rect 8852 16983 8904 16992
rect 8852 16949 8861 16983
rect 8861 16949 8895 16983
rect 8895 16949 8904 16983
rect 8852 16940 8904 16949
rect 11980 16940 12032 16992
rect 15200 16940 15252 16992
rect 16672 16983 16724 16992
rect 16672 16949 16681 16983
rect 16681 16949 16715 16983
rect 16715 16949 16724 16983
rect 16672 16940 16724 16949
rect 16856 16940 16908 16992
rect 22376 16940 22428 16992
rect 2950 16838 3002 16890
rect 3014 16838 3066 16890
rect 3078 16838 3130 16890
rect 3142 16838 3194 16890
rect 3206 16838 3258 16890
rect 12950 16838 13002 16890
rect 13014 16838 13066 16890
rect 13078 16838 13130 16890
rect 13142 16838 13194 16890
rect 13206 16838 13258 16890
rect 22950 16838 23002 16890
rect 23014 16838 23066 16890
rect 23078 16838 23130 16890
rect 23142 16838 23194 16890
rect 23206 16838 23258 16890
rect 7656 16779 7708 16788
rect 7656 16745 7665 16779
rect 7665 16745 7699 16779
rect 7699 16745 7708 16779
rect 7656 16736 7708 16745
rect 8760 16736 8812 16788
rect 9588 16736 9640 16788
rect 11152 16736 11204 16788
rect 12440 16736 12492 16788
rect 14004 16736 14056 16788
rect 16672 16736 16724 16788
rect 17316 16736 17368 16788
rect 18328 16736 18380 16788
rect 6828 16600 6880 16652
rect 7472 16600 7524 16652
rect 9680 16600 9732 16652
rect 11244 16600 11296 16652
rect 12348 16643 12400 16652
rect 12348 16609 12357 16643
rect 12357 16609 12391 16643
rect 12391 16609 12400 16643
rect 12348 16600 12400 16609
rect 10600 16532 10652 16584
rect 11060 16532 11112 16584
rect 13360 16600 13412 16652
rect 13544 16643 13596 16652
rect 13544 16609 13553 16643
rect 13553 16609 13587 16643
rect 13587 16609 13596 16643
rect 13544 16600 13596 16609
rect 14096 16643 14148 16652
rect 14096 16609 14105 16643
rect 14105 16609 14139 16643
rect 14139 16609 14148 16643
rect 14096 16600 14148 16609
rect 15752 16643 15804 16652
rect 15752 16609 15761 16643
rect 15761 16609 15795 16643
rect 15795 16609 15804 16643
rect 15752 16600 15804 16609
rect 16488 16600 16540 16652
rect 15660 16575 15712 16584
rect 15660 16541 15669 16575
rect 15669 16541 15703 16575
rect 15703 16541 15712 16575
rect 15660 16532 15712 16541
rect 17684 16532 17736 16584
rect 6184 16507 6236 16516
rect 6184 16473 6193 16507
rect 6193 16473 6227 16507
rect 6227 16473 6236 16507
rect 6184 16464 6236 16473
rect 10416 16396 10468 16448
rect 10692 16396 10744 16448
rect 10968 16396 11020 16448
rect 13636 16464 13688 16516
rect 18420 16668 18472 16720
rect 18604 16575 18656 16584
rect 18604 16541 18613 16575
rect 18613 16541 18647 16575
rect 18647 16541 18656 16575
rect 18604 16532 18656 16541
rect 19432 16736 19484 16788
rect 25780 16736 25832 16788
rect 20720 16532 20772 16584
rect 20996 16532 21048 16584
rect 22560 16532 22612 16584
rect 22744 16575 22796 16584
rect 22744 16541 22753 16575
rect 22753 16541 22787 16575
rect 22787 16541 22796 16575
rect 22744 16532 22796 16541
rect 23940 16532 23992 16584
rect 25228 16575 25280 16584
rect 25228 16541 25237 16575
rect 25237 16541 25271 16575
rect 25271 16541 25280 16575
rect 25228 16532 25280 16541
rect 12440 16396 12492 16448
rect 14096 16396 14148 16448
rect 16396 16396 16448 16448
rect 17408 16396 17460 16448
rect 19708 16464 19760 16516
rect 20628 16464 20680 16516
rect 24952 16464 25004 16516
rect 18880 16396 18932 16448
rect 19248 16396 19300 16448
rect 19984 16396 20036 16448
rect 21548 16396 21600 16448
rect 24860 16396 24912 16448
rect 7950 16294 8002 16346
rect 8014 16294 8066 16346
rect 8078 16294 8130 16346
rect 8142 16294 8194 16346
rect 8206 16294 8258 16346
rect 17950 16294 18002 16346
rect 18014 16294 18066 16346
rect 18078 16294 18130 16346
rect 18142 16294 18194 16346
rect 18206 16294 18258 16346
rect 5448 16192 5500 16244
rect 11060 16192 11112 16244
rect 11612 16192 11664 16244
rect 12624 16192 12676 16244
rect 7840 16167 7892 16176
rect 7840 16133 7849 16167
rect 7849 16133 7883 16167
rect 7883 16133 7892 16167
rect 7840 16124 7892 16133
rect 9588 16124 9640 16176
rect 11520 16124 11572 16176
rect 12440 16124 12492 16176
rect 15476 16192 15528 16244
rect 18604 16192 18656 16244
rect 19340 16192 19392 16244
rect 17224 16167 17276 16176
rect 17224 16133 17233 16167
rect 17233 16133 17267 16167
rect 17267 16133 17276 16167
rect 17224 16124 17276 16133
rect 21548 16192 21600 16244
rect 21640 16192 21692 16244
rect 19984 16167 20036 16176
rect 19984 16133 19993 16167
rect 19993 16133 20027 16167
rect 20027 16133 20036 16167
rect 19984 16124 20036 16133
rect 21364 16124 21416 16176
rect 21916 16124 21968 16176
rect 25044 16192 25096 16244
rect 25872 16124 25924 16176
rect 6920 16056 6972 16108
rect 11612 16056 11664 16108
rect 15292 16056 15344 16108
rect 15844 16056 15896 16108
rect 18604 16099 18656 16108
rect 18604 16065 18613 16099
rect 18613 16065 18647 16099
rect 18647 16065 18656 16099
rect 18604 16056 18656 16065
rect 9588 16031 9640 16040
rect 9588 15997 9597 16031
rect 9597 15997 9631 16031
rect 9631 15997 9640 16031
rect 9588 15988 9640 15997
rect 13452 15988 13504 16040
rect 14556 16031 14608 16040
rect 14556 15997 14565 16031
rect 14565 15997 14599 16031
rect 14599 15997 14608 16031
rect 14556 15988 14608 15997
rect 12440 15852 12492 15904
rect 13912 15920 13964 15972
rect 19708 16031 19760 16040
rect 19708 15997 19717 16031
rect 19717 15997 19751 16031
rect 19751 15997 19760 16031
rect 19708 15988 19760 15997
rect 13452 15895 13504 15904
rect 13452 15861 13461 15895
rect 13461 15861 13495 15895
rect 13495 15861 13504 15895
rect 17500 15920 17552 15972
rect 20444 15988 20496 16040
rect 20628 15988 20680 16040
rect 22284 15988 22336 16040
rect 25136 16056 25188 16108
rect 13452 15852 13504 15861
rect 17316 15895 17368 15904
rect 17316 15861 17325 15895
rect 17325 15861 17359 15895
rect 17359 15861 17368 15895
rect 17316 15852 17368 15861
rect 19340 15852 19392 15904
rect 20168 15852 20220 15904
rect 20536 15852 20588 15904
rect 23572 15920 23624 15972
rect 23756 15895 23808 15904
rect 23756 15861 23765 15895
rect 23765 15861 23799 15895
rect 23799 15861 23808 15895
rect 23756 15852 23808 15861
rect 2950 15750 3002 15802
rect 3014 15750 3066 15802
rect 3078 15750 3130 15802
rect 3142 15750 3194 15802
rect 3206 15750 3258 15802
rect 12950 15750 13002 15802
rect 13014 15750 13066 15802
rect 13078 15750 13130 15802
rect 13142 15750 13194 15802
rect 13206 15750 13258 15802
rect 22950 15750 23002 15802
rect 23014 15750 23066 15802
rect 23078 15750 23130 15802
rect 23142 15750 23194 15802
rect 23206 15750 23258 15802
rect 7748 15648 7800 15700
rect 8760 15648 8812 15700
rect 9312 15648 9364 15700
rect 14556 15648 14608 15700
rect 17776 15648 17828 15700
rect 21640 15648 21692 15700
rect 9404 15512 9456 15564
rect 6368 15487 6420 15496
rect 6368 15453 6377 15487
rect 6377 15453 6411 15487
rect 6411 15453 6420 15487
rect 6368 15444 6420 15453
rect 8760 15376 8812 15428
rect 11244 15512 11296 15564
rect 11980 15555 12032 15564
rect 11980 15521 11989 15555
rect 11989 15521 12023 15555
rect 12023 15521 12032 15555
rect 11980 15512 12032 15521
rect 12440 15512 12492 15564
rect 12808 15512 12860 15564
rect 15292 15555 15344 15564
rect 15292 15521 15301 15555
rect 15301 15521 15335 15555
rect 15335 15521 15344 15555
rect 15292 15512 15344 15521
rect 19708 15512 19760 15564
rect 20444 15512 20496 15564
rect 9956 15487 10008 15496
rect 9956 15453 9965 15487
rect 9965 15453 9999 15487
rect 9999 15453 10008 15487
rect 9956 15444 10008 15453
rect 19340 15444 19392 15496
rect 22284 15555 22336 15564
rect 22284 15521 22293 15555
rect 22293 15521 22327 15555
rect 22327 15521 22336 15555
rect 22284 15512 22336 15521
rect 23848 15444 23900 15496
rect 10232 15419 10284 15428
rect 10232 15385 10241 15419
rect 10241 15385 10275 15419
rect 10275 15385 10284 15419
rect 10232 15376 10284 15385
rect 12716 15351 12768 15360
rect 12716 15317 12725 15351
rect 12725 15317 12759 15351
rect 12759 15317 12768 15351
rect 13360 15351 13412 15360
rect 12716 15308 12768 15317
rect 13360 15317 13369 15351
rect 13369 15317 13403 15351
rect 13403 15317 13412 15351
rect 13360 15308 13412 15317
rect 14280 15351 14332 15360
rect 14280 15317 14289 15351
rect 14289 15317 14323 15351
rect 14323 15317 14332 15351
rect 14280 15308 14332 15317
rect 16028 15308 16080 15360
rect 16580 15376 16632 15428
rect 16948 15376 17000 15428
rect 21916 15376 21968 15428
rect 23572 15376 23624 15428
rect 17224 15308 17276 15360
rect 18788 15308 18840 15360
rect 19524 15308 19576 15360
rect 19892 15308 19944 15360
rect 20996 15308 21048 15360
rect 21640 15351 21692 15360
rect 21640 15317 21649 15351
rect 21649 15317 21683 15351
rect 21683 15317 21692 15351
rect 21640 15308 21692 15317
rect 22468 15308 22520 15360
rect 7950 15206 8002 15258
rect 8014 15206 8066 15258
rect 8078 15206 8130 15258
rect 8142 15206 8194 15258
rect 8206 15206 8258 15258
rect 17950 15206 18002 15258
rect 18014 15206 18066 15258
rect 18078 15206 18130 15258
rect 18142 15206 18194 15258
rect 18206 15206 18258 15258
rect 6184 15104 6236 15156
rect 8760 15036 8812 15088
rect 10232 15036 10284 15088
rect 11336 15147 11388 15156
rect 11336 15113 11345 15147
rect 11345 15113 11379 15147
rect 11379 15113 11388 15147
rect 11336 15104 11388 15113
rect 11520 15036 11572 15088
rect 3424 14968 3476 15020
rect 5264 14968 5316 15020
rect 7564 14968 7616 15020
rect 9680 14968 9732 15020
rect 6368 14900 6420 14952
rect 8576 14900 8628 14952
rect 10968 14968 11020 15020
rect 12716 15104 12768 15156
rect 13728 15104 13780 15156
rect 14280 15104 14332 15156
rect 15292 15104 15344 15156
rect 19800 15104 19852 15156
rect 20352 15104 20404 15156
rect 21916 15147 21968 15156
rect 21916 15113 21925 15147
rect 21925 15113 21959 15147
rect 21959 15113 21968 15147
rect 21916 15104 21968 15113
rect 23572 15104 23624 15156
rect 12624 15079 12676 15088
rect 12624 15045 12633 15079
rect 12633 15045 12667 15079
rect 12667 15045 12676 15079
rect 12624 15036 12676 15045
rect 14188 15036 14240 15088
rect 14464 15036 14516 15088
rect 13452 14968 13504 15020
rect 14556 14968 14608 15020
rect 16212 15036 16264 15088
rect 16948 15036 17000 15088
rect 18972 15036 19024 15088
rect 20812 15036 20864 15088
rect 10140 14832 10192 14884
rect 16028 14943 16080 14952
rect 16028 14909 16037 14943
rect 16037 14909 16071 14943
rect 16071 14909 16080 14943
rect 16028 14900 16080 14909
rect 18696 14968 18748 15020
rect 18880 14968 18932 15020
rect 21088 15011 21140 15020
rect 21088 14977 21097 15011
rect 21097 14977 21131 15011
rect 21131 14977 21140 15011
rect 21088 14968 21140 14977
rect 21456 15036 21508 15088
rect 22468 15011 22520 15020
rect 22468 14977 22477 15011
rect 22477 14977 22511 15011
rect 22511 14977 22520 15011
rect 22468 14968 22520 14977
rect 11428 14832 11480 14884
rect 13452 14832 13504 14884
rect 15568 14875 15620 14884
rect 15568 14841 15577 14875
rect 15577 14841 15611 14875
rect 15611 14841 15620 14875
rect 15568 14832 15620 14841
rect 19800 14900 19852 14952
rect 20996 14900 21048 14952
rect 23756 14900 23808 14952
rect 24768 14943 24820 14952
rect 24768 14909 24777 14943
rect 24777 14909 24811 14943
rect 24811 14909 24820 14943
rect 24768 14900 24820 14909
rect 19432 14832 19484 14884
rect 19708 14832 19760 14884
rect 25596 14832 25648 14884
rect 9956 14764 10008 14816
rect 10324 14764 10376 14816
rect 13544 14764 13596 14816
rect 18696 14807 18748 14816
rect 18696 14773 18705 14807
rect 18705 14773 18739 14807
rect 18739 14773 18748 14807
rect 18696 14764 18748 14773
rect 19064 14764 19116 14816
rect 22560 14764 22612 14816
rect 23572 14764 23624 14816
rect 23848 14764 23900 14816
rect 2950 14662 3002 14714
rect 3014 14662 3066 14714
rect 3078 14662 3130 14714
rect 3142 14662 3194 14714
rect 3206 14662 3258 14714
rect 12950 14662 13002 14714
rect 13014 14662 13066 14714
rect 13078 14662 13130 14714
rect 13142 14662 13194 14714
rect 13206 14662 13258 14714
rect 22950 14662 23002 14714
rect 23014 14662 23066 14714
rect 23078 14662 23130 14714
rect 23142 14662 23194 14714
rect 23206 14662 23258 14714
rect 8576 14603 8628 14612
rect 8576 14569 8585 14603
rect 8585 14569 8619 14603
rect 8619 14569 8628 14603
rect 8576 14560 8628 14569
rect 9036 14560 9088 14612
rect 11704 14603 11756 14612
rect 11704 14569 11713 14603
rect 11713 14569 11747 14603
rect 11747 14569 11756 14603
rect 11704 14560 11756 14569
rect 14372 14603 14424 14612
rect 14372 14569 14381 14603
rect 14381 14569 14415 14603
rect 14415 14569 14424 14603
rect 14372 14560 14424 14569
rect 14740 14560 14792 14612
rect 16856 14560 16908 14612
rect 18328 14603 18380 14612
rect 18328 14569 18337 14603
rect 18337 14569 18371 14603
rect 18371 14569 18380 14603
rect 18328 14560 18380 14569
rect 19432 14560 19484 14612
rect 22652 14560 22704 14612
rect 12348 14492 12400 14544
rect 15108 14492 15160 14544
rect 19064 14492 19116 14544
rect 19340 14492 19392 14544
rect 20076 14492 20128 14544
rect 22284 14492 22336 14544
rect 7564 14424 7616 14476
rect 9680 14467 9732 14476
rect 9680 14433 9689 14467
rect 9689 14433 9723 14467
rect 9723 14433 9732 14467
rect 9680 14424 9732 14433
rect 9956 14424 10008 14476
rect 11980 14424 12032 14476
rect 13452 14467 13504 14476
rect 13452 14433 13461 14467
rect 13461 14433 13495 14467
rect 13495 14433 13504 14467
rect 13452 14424 13504 14433
rect 7748 14356 7800 14408
rect 8944 14356 8996 14408
rect 9588 14356 9640 14408
rect 11336 14356 11388 14408
rect 15384 14424 15436 14476
rect 15568 14467 15620 14476
rect 15568 14433 15577 14467
rect 15577 14433 15611 14467
rect 15611 14433 15620 14467
rect 15568 14424 15620 14433
rect 18328 14424 18380 14476
rect 19156 14424 19208 14476
rect 15200 14356 15252 14408
rect 12532 14288 12584 14340
rect 13544 14288 13596 14340
rect 19340 14356 19392 14408
rect 19800 14424 19852 14476
rect 22192 14424 22244 14476
rect 22560 14467 22612 14476
rect 22560 14433 22569 14467
rect 22569 14433 22603 14467
rect 22603 14433 22612 14467
rect 22560 14424 22612 14433
rect 9496 14263 9548 14272
rect 9496 14229 9505 14263
rect 9505 14229 9539 14263
rect 9539 14229 9548 14263
rect 9496 14220 9548 14229
rect 9588 14263 9640 14272
rect 9588 14229 9597 14263
rect 9597 14229 9631 14263
rect 9631 14229 9640 14263
rect 9588 14220 9640 14229
rect 10232 14220 10284 14272
rect 10968 14220 11020 14272
rect 12716 14220 12768 14272
rect 12808 14220 12860 14272
rect 19800 14288 19852 14340
rect 20720 14356 20772 14408
rect 21732 14356 21784 14408
rect 22284 14399 22336 14408
rect 22284 14365 22293 14399
rect 22293 14365 22327 14399
rect 22327 14365 22336 14399
rect 22284 14356 22336 14365
rect 24676 14356 24728 14408
rect 16028 14263 16080 14272
rect 16028 14229 16037 14263
rect 16037 14229 16071 14263
rect 16071 14229 16080 14263
rect 16028 14220 16080 14229
rect 16304 14263 16356 14272
rect 16304 14229 16313 14263
rect 16313 14229 16347 14263
rect 16347 14229 16356 14263
rect 16304 14220 16356 14229
rect 16580 14263 16632 14272
rect 16580 14229 16589 14263
rect 16589 14229 16623 14263
rect 16623 14229 16632 14263
rect 16580 14220 16632 14229
rect 19432 14220 19484 14272
rect 19892 14220 19944 14272
rect 20352 14220 20404 14272
rect 23848 14288 23900 14340
rect 21364 14220 21416 14272
rect 22100 14220 22152 14272
rect 24032 14263 24084 14272
rect 24032 14229 24041 14263
rect 24041 14229 24075 14263
rect 24075 14229 24084 14263
rect 24032 14220 24084 14229
rect 24492 14220 24544 14272
rect 25044 14263 25096 14272
rect 25044 14229 25053 14263
rect 25053 14229 25087 14263
rect 25087 14229 25096 14263
rect 25044 14220 25096 14229
rect 7950 14118 8002 14170
rect 8014 14118 8066 14170
rect 8078 14118 8130 14170
rect 8142 14118 8194 14170
rect 8206 14118 8258 14170
rect 17950 14118 18002 14170
rect 18014 14118 18066 14170
rect 18078 14118 18130 14170
rect 18142 14118 18194 14170
rect 18206 14118 18258 14170
rect 8300 14016 8352 14068
rect 9496 14016 9548 14068
rect 12256 14016 12308 14068
rect 14648 14016 14700 14068
rect 6368 13880 6420 13932
rect 7104 13948 7156 14000
rect 8760 13948 8812 14000
rect 10140 13948 10192 14000
rect 12624 13948 12676 14000
rect 9772 13880 9824 13932
rect 13452 13880 13504 13932
rect 14924 13880 14976 13932
rect 15568 13923 15620 13932
rect 7564 13812 7616 13864
rect 9404 13812 9456 13864
rect 9496 13676 9548 13728
rect 11980 13744 12032 13796
rect 13544 13855 13596 13864
rect 13544 13821 13553 13855
rect 13553 13821 13587 13855
rect 13587 13821 13596 13855
rect 13544 13812 13596 13821
rect 14372 13812 14424 13864
rect 15568 13889 15577 13923
rect 15577 13889 15611 13923
rect 15611 13889 15620 13923
rect 15568 13880 15620 13889
rect 15844 13812 15896 13864
rect 14924 13744 14976 13796
rect 16488 14016 16540 14068
rect 16948 14016 17000 14068
rect 17132 13948 17184 14000
rect 18604 14059 18656 14068
rect 18604 14025 18613 14059
rect 18613 14025 18647 14059
rect 18647 14025 18656 14059
rect 18604 14016 18656 14025
rect 19800 14016 19852 14068
rect 18420 13948 18472 14000
rect 19432 13948 19484 14000
rect 21364 13880 21416 13932
rect 24860 13948 24912 14000
rect 25136 13991 25188 14000
rect 25136 13957 25145 13991
rect 25145 13957 25179 13991
rect 25179 13957 25188 13991
rect 25136 13948 25188 13957
rect 17868 13812 17920 13864
rect 20260 13812 20312 13864
rect 22836 13812 22888 13864
rect 11888 13676 11940 13728
rect 15200 13676 15252 13728
rect 15936 13676 15988 13728
rect 16304 13676 16356 13728
rect 17224 13676 17276 13728
rect 17592 13676 17644 13728
rect 17684 13676 17736 13728
rect 21916 13744 21968 13796
rect 26608 13744 26660 13796
rect 19340 13676 19392 13728
rect 20536 13676 20588 13728
rect 20628 13719 20680 13728
rect 20628 13685 20637 13719
rect 20637 13685 20671 13719
rect 20671 13685 20680 13719
rect 20628 13676 20680 13685
rect 21272 13719 21324 13728
rect 21272 13685 21281 13719
rect 21281 13685 21315 13719
rect 21315 13685 21324 13719
rect 21272 13676 21324 13685
rect 2950 13574 3002 13626
rect 3014 13574 3066 13626
rect 3078 13574 3130 13626
rect 3142 13574 3194 13626
rect 3206 13574 3258 13626
rect 12950 13574 13002 13626
rect 13014 13574 13066 13626
rect 13078 13574 13130 13626
rect 13142 13574 13194 13626
rect 13206 13574 13258 13626
rect 22950 13574 23002 13626
rect 23014 13574 23066 13626
rect 23078 13574 23130 13626
rect 23142 13574 23194 13626
rect 23206 13574 23258 13626
rect 7380 13472 7432 13524
rect 13912 13472 13964 13524
rect 14188 13472 14240 13524
rect 15016 13472 15068 13524
rect 20536 13472 20588 13524
rect 7012 13336 7064 13388
rect 9220 13268 9272 13320
rect 11704 13336 11756 13388
rect 13544 13336 13596 13388
rect 14924 13336 14976 13388
rect 15384 13336 15436 13388
rect 11336 13268 11388 13320
rect 15292 13268 15344 13320
rect 15844 13336 15896 13388
rect 16396 13268 16448 13320
rect 16580 13268 16632 13320
rect 17592 13311 17644 13320
rect 17592 13277 17601 13311
rect 17601 13277 17635 13311
rect 17635 13277 17644 13311
rect 17592 13268 17644 13277
rect 17776 13268 17828 13320
rect 18328 13268 18380 13320
rect 19248 13336 19300 13388
rect 24768 13404 24820 13456
rect 6184 13200 6236 13252
rect 8760 13200 8812 13252
rect 7380 13175 7432 13184
rect 7380 13141 7389 13175
rect 7389 13141 7423 13175
rect 7423 13141 7432 13175
rect 7380 13132 7432 13141
rect 9128 13175 9180 13184
rect 9128 13141 9137 13175
rect 9137 13141 9171 13175
rect 9171 13141 9180 13175
rect 9128 13132 9180 13141
rect 10324 13200 10376 13252
rect 10508 13200 10560 13252
rect 17500 13200 17552 13252
rect 11060 13132 11112 13184
rect 13452 13132 13504 13184
rect 15384 13132 15436 13184
rect 15568 13175 15620 13184
rect 15568 13141 15577 13175
rect 15577 13141 15611 13175
rect 15611 13141 15620 13175
rect 15568 13132 15620 13141
rect 15660 13175 15712 13184
rect 15660 13141 15669 13175
rect 15669 13141 15703 13175
rect 15703 13141 15712 13175
rect 15660 13132 15712 13141
rect 15752 13132 15804 13184
rect 18328 13132 18380 13184
rect 19524 13243 19576 13252
rect 19524 13209 19533 13243
rect 19533 13209 19567 13243
rect 19567 13209 19576 13243
rect 19524 13200 19576 13209
rect 19340 13132 19392 13184
rect 20076 13132 20128 13184
rect 20168 13175 20220 13184
rect 20168 13141 20177 13175
rect 20177 13141 20211 13175
rect 20211 13141 20220 13175
rect 20168 13132 20220 13141
rect 20536 13175 20588 13184
rect 20536 13141 20545 13175
rect 20545 13141 20579 13175
rect 20579 13141 20588 13175
rect 20536 13132 20588 13141
rect 24032 13336 24084 13388
rect 20904 13268 20956 13320
rect 20720 13200 20772 13252
rect 23756 13268 23808 13320
rect 24952 13200 25004 13252
rect 20996 13132 21048 13184
rect 21732 13132 21784 13184
rect 23296 13132 23348 13184
rect 7950 13030 8002 13082
rect 8014 13030 8066 13082
rect 8078 13030 8130 13082
rect 8142 13030 8194 13082
rect 8206 13030 8258 13082
rect 17950 13030 18002 13082
rect 18014 13030 18066 13082
rect 18078 13030 18130 13082
rect 18142 13030 18194 13082
rect 18206 13030 18258 13082
rect 7380 12928 7432 12980
rect 8392 12928 8444 12980
rect 8760 12860 8812 12912
rect 14004 12928 14056 12980
rect 15752 12928 15804 12980
rect 20904 12971 20956 12980
rect 7104 12792 7156 12844
rect 12624 12860 12676 12912
rect 9404 12792 9456 12844
rect 11980 12792 12032 12844
rect 15108 12860 15160 12912
rect 12992 12835 13044 12844
rect 12992 12801 13001 12835
rect 13001 12801 13035 12835
rect 13035 12801 13044 12835
rect 12992 12792 13044 12801
rect 13360 12792 13412 12844
rect 14280 12792 14332 12844
rect 16212 12860 16264 12912
rect 20904 12937 20913 12971
rect 20913 12937 20947 12971
rect 20947 12937 20956 12971
rect 20904 12928 20956 12937
rect 20996 12928 21048 12980
rect 24768 12971 24820 12980
rect 24768 12937 24777 12971
rect 24777 12937 24811 12971
rect 24811 12937 24820 12971
rect 24768 12928 24820 12937
rect 8576 12656 8628 12708
rect 7656 12588 7708 12640
rect 11612 12724 11664 12776
rect 14372 12724 14424 12776
rect 15108 12724 15160 12776
rect 9404 12656 9456 12708
rect 9680 12656 9732 12708
rect 14004 12656 14056 12708
rect 15292 12656 15344 12708
rect 15752 12792 15804 12844
rect 15568 12724 15620 12776
rect 15936 12724 15988 12776
rect 16948 12792 17000 12844
rect 18420 12792 18472 12844
rect 19064 12835 19116 12844
rect 19064 12801 19073 12835
rect 19073 12801 19107 12835
rect 19107 12801 19116 12835
rect 19064 12792 19116 12801
rect 20076 12860 20128 12912
rect 20536 12860 20588 12912
rect 21456 12903 21508 12912
rect 21456 12869 21465 12903
rect 21465 12869 21499 12903
rect 21499 12869 21508 12903
rect 21456 12860 21508 12869
rect 20352 12792 20404 12844
rect 21548 12792 21600 12844
rect 22376 12860 22428 12912
rect 23296 12903 23348 12912
rect 23296 12869 23305 12903
rect 23305 12869 23339 12903
rect 23339 12869 23348 12903
rect 23296 12860 23348 12869
rect 25136 12860 25188 12912
rect 22284 12792 22336 12844
rect 22836 12792 22888 12844
rect 17868 12724 17920 12776
rect 18512 12724 18564 12776
rect 19248 12767 19300 12776
rect 19248 12733 19257 12767
rect 19257 12733 19291 12767
rect 19291 12733 19300 12767
rect 19248 12724 19300 12733
rect 11612 12631 11664 12640
rect 11612 12597 11621 12631
rect 11621 12597 11655 12631
rect 11655 12597 11664 12631
rect 11612 12588 11664 12597
rect 12348 12588 12400 12640
rect 12992 12588 13044 12640
rect 13728 12631 13780 12640
rect 13728 12597 13737 12631
rect 13737 12597 13771 12631
rect 13771 12597 13780 12631
rect 13728 12588 13780 12597
rect 15844 12588 15896 12640
rect 15936 12588 15988 12640
rect 17684 12588 17736 12640
rect 17776 12588 17828 12640
rect 21088 12656 21140 12708
rect 20076 12631 20128 12640
rect 20076 12597 20085 12631
rect 20085 12597 20119 12631
rect 20119 12597 20128 12631
rect 20076 12588 20128 12597
rect 22284 12588 22336 12640
rect 25136 12631 25188 12640
rect 25136 12597 25145 12631
rect 25145 12597 25179 12631
rect 25179 12597 25188 12631
rect 25136 12588 25188 12597
rect 2950 12486 3002 12538
rect 3014 12486 3066 12538
rect 3078 12486 3130 12538
rect 3142 12486 3194 12538
rect 3206 12486 3258 12538
rect 12950 12486 13002 12538
rect 13014 12486 13066 12538
rect 13078 12486 13130 12538
rect 13142 12486 13194 12538
rect 13206 12486 13258 12538
rect 22950 12486 23002 12538
rect 23014 12486 23066 12538
rect 23078 12486 23130 12538
rect 23142 12486 23194 12538
rect 23206 12486 23258 12538
rect 7472 12384 7524 12436
rect 9772 12427 9824 12436
rect 9772 12393 9781 12427
rect 9781 12393 9815 12427
rect 9815 12393 9824 12427
rect 9772 12384 9824 12393
rect 11428 12427 11480 12436
rect 11428 12393 11437 12427
rect 11437 12393 11471 12427
rect 11471 12393 11480 12427
rect 11428 12384 11480 12393
rect 12072 12384 12124 12436
rect 13636 12384 13688 12436
rect 18420 12384 18472 12436
rect 8484 12291 8536 12300
rect 8484 12257 8493 12291
rect 8493 12257 8527 12291
rect 8527 12257 8536 12291
rect 8484 12248 8536 12257
rect 10784 12248 10836 12300
rect 15660 12316 15712 12368
rect 12072 12291 12124 12300
rect 12072 12257 12081 12291
rect 12081 12257 12115 12291
rect 12115 12257 12124 12291
rect 12072 12248 12124 12257
rect 12440 12248 12492 12300
rect 14188 12248 14240 12300
rect 15016 12248 15068 12300
rect 15292 12248 15344 12300
rect 16764 12248 16816 12300
rect 9128 12180 9180 12232
rect 12808 12180 12860 12232
rect 5080 12112 5132 12164
rect 10876 12112 10928 12164
rect 12440 12112 12492 12164
rect 14280 12180 14332 12232
rect 14372 12180 14424 12232
rect 16304 12180 16356 12232
rect 17684 12316 17736 12368
rect 18788 12316 18840 12368
rect 18604 12248 18656 12300
rect 18972 12180 19024 12232
rect 20352 12384 20404 12436
rect 21732 12316 21784 12368
rect 21916 12316 21968 12368
rect 20260 12248 20312 12300
rect 22192 12180 22244 12232
rect 24768 12180 24820 12232
rect 6920 12044 6972 12096
rect 8760 12044 8812 12096
rect 9036 12044 9088 12096
rect 9128 12044 9180 12096
rect 13360 12044 13412 12096
rect 13636 12087 13688 12096
rect 13636 12053 13645 12087
rect 13645 12053 13679 12087
rect 13679 12053 13688 12087
rect 13636 12044 13688 12053
rect 14372 12044 14424 12096
rect 14740 12087 14792 12096
rect 14740 12053 14749 12087
rect 14749 12053 14783 12087
rect 14783 12053 14792 12087
rect 14740 12044 14792 12053
rect 14924 12044 14976 12096
rect 18328 12112 18380 12164
rect 18420 12112 18472 12164
rect 19156 12112 19208 12164
rect 20352 12112 20404 12164
rect 20628 12155 20680 12164
rect 20628 12121 20637 12155
rect 20637 12121 20671 12155
rect 20671 12121 20680 12155
rect 20628 12112 20680 12121
rect 21916 12112 21968 12164
rect 22284 12112 22336 12164
rect 24952 12112 25004 12164
rect 16120 12044 16172 12096
rect 16212 12087 16264 12096
rect 16212 12053 16221 12087
rect 16221 12053 16255 12087
rect 16255 12053 16264 12087
rect 16212 12044 16264 12053
rect 16764 12044 16816 12096
rect 18512 12044 18564 12096
rect 18972 12044 19024 12096
rect 19432 12044 19484 12096
rect 23388 12044 23440 12096
rect 7950 11942 8002 11994
rect 8014 11942 8066 11994
rect 8078 11942 8130 11994
rect 8142 11942 8194 11994
rect 8206 11942 8258 11994
rect 17950 11942 18002 11994
rect 18014 11942 18066 11994
rect 18078 11942 18130 11994
rect 18142 11942 18194 11994
rect 18206 11942 18258 11994
rect 9680 11840 9732 11892
rect 10140 11883 10192 11892
rect 10140 11849 10149 11883
rect 10149 11849 10183 11883
rect 10183 11849 10192 11883
rect 10140 11840 10192 11849
rect 9588 11772 9640 11824
rect 8760 11704 8812 11756
rect 11060 11840 11112 11892
rect 11520 11840 11572 11892
rect 12164 11840 12216 11892
rect 13268 11840 13320 11892
rect 13820 11840 13872 11892
rect 14464 11840 14516 11892
rect 14832 11840 14884 11892
rect 15200 11840 15252 11892
rect 17040 11840 17092 11892
rect 18880 11840 18932 11892
rect 19156 11840 19208 11892
rect 11428 11704 11480 11756
rect 12256 11704 12308 11756
rect 12440 11747 12492 11756
rect 12440 11713 12449 11747
rect 12449 11713 12483 11747
rect 12483 11713 12492 11747
rect 12440 11704 12492 11713
rect 9496 11636 9548 11688
rect 9956 11636 10008 11688
rect 9404 11568 9456 11620
rect 7196 11500 7248 11552
rect 9128 11500 9180 11552
rect 10784 11679 10836 11688
rect 10784 11645 10793 11679
rect 10793 11645 10827 11679
rect 10827 11645 10836 11679
rect 10784 11636 10836 11645
rect 11060 11636 11112 11688
rect 11888 11636 11940 11688
rect 12072 11636 12124 11688
rect 14004 11772 14056 11824
rect 14832 11747 14884 11756
rect 14832 11713 14841 11747
rect 14841 11713 14875 11747
rect 14875 11713 14884 11747
rect 14832 11704 14884 11713
rect 15108 11704 15160 11756
rect 16120 11772 16172 11824
rect 20628 11840 20680 11892
rect 20720 11772 20772 11824
rect 21732 11772 21784 11824
rect 23388 11815 23440 11824
rect 23388 11781 23397 11815
rect 23397 11781 23431 11815
rect 23431 11781 23440 11815
rect 23388 11772 23440 11781
rect 25136 11772 25188 11824
rect 11244 11543 11296 11552
rect 11244 11509 11253 11543
rect 11253 11509 11287 11543
rect 11287 11509 11296 11543
rect 11244 11500 11296 11509
rect 12808 11500 12860 11552
rect 13268 11500 13320 11552
rect 14188 11636 14240 11688
rect 17408 11679 17460 11688
rect 17408 11645 17417 11679
rect 17417 11645 17451 11679
rect 17451 11645 17460 11679
rect 17408 11636 17460 11645
rect 14096 11568 14148 11620
rect 19064 11704 19116 11756
rect 20444 11704 20496 11756
rect 21456 11704 21508 11756
rect 22284 11704 22336 11756
rect 22836 11704 22888 11756
rect 18512 11679 18564 11688
rect 18512 11645 18521 11679
rect 18521 11645 18555 11679
rect 18555 11645 18564 11679
rect 18512 11636 18564 11645
rect 19432 11636 19484 11688
rect 20812 11636 20864 11688
rect 19156 11568 19208 11620
rect 19708 11568 19760 11620
rect 14188 11500 14240 11552
rect 15292 11500 15344 11552
rect 18604 11500 18656 11552
rect 20720 11500 20772 11552
rect 24584 11500 24636 11552
rect 25136 11543 25188 11552
rect 25136 11509 25145 11543
rect 25145 11509 25179 11543
rect 25179 11509 25188 11543
rect 25136 11500 25188 11509
rect 2950 11398 3002 11450
rect 3014 11398 3066 11450
rect 3078 11398 3130 11450
rect 3142 11398 3194 11450
rect 3206 11398 3258 11450
rect 12950 11398 13002 11450
rect 13014 11398 13066 11450
rect 13078 11398 13130 11450
rect 13142 11398 13194 11450
rect 13206 11398 13258 11450
rect 22950 11398 23002 11450
rect 23014 11398 23066 11450
rect 23078 11398 23130 11450
rect 23142 11398 23194 11450
rect 23206 11398 23258 11450
rect 8576 11339 8628 11348
rect 8576 11305 8585 11339
rect 8585 11305 8619 11339
rect 8619 11305 8628 11339
rect 8576 11296 8628 11305
rect 10784 11296 10836 11348
rect 9496 11160 9548 11212
rect 10048 11160 10100 11212
rect 10876 11092 10928 11144
rect 11796 11203 11848 11212
rect 11796 11169 11805 11203
rect 11805 11169 11839 11203
rect 11839 11169 11848 11203
rect 11796 11160 11848 11169
rect 11888 11203 11940 11212
rect 11888 11169 11897 11203
rect 11897 11169 11931 11203
rect 11931 11169 11940 11203
rect 11888 11160 11940 11169
rect 12624 11339 12676 11348
rect 12624 11305 12633 11339
rect 12633 11305 12667 11339
rect 12667 11305 12676 11339
rect 12624 11296 12676 11305
rect 12992 11296 13044 11348
rect 15384 11296 15436 11348
rect 17224 11296 17276 11348
rect 17408 11296 17460 11348
rect 18328 11296 18380 11348
rect 18420 11296 18472 11348
rect 18696 11296 18748 11348
rect 19064 11339 19116 11348
rect 19064 11305 19073 11339
rect 19073 11305 19107 11339
rect 19107 11305 19116 11339
rect 19064 11296 19116 11305
rect 19432 11296 19484 11348
rect 21548 11339 21600 11348
rect 21548 11305 21557 11339
rect 21557 11305 21591 11339
rect 21591 11305 21600 11339
rect 21548 11296 21600 11305
rect 12900 11228 12952 11280
rect 13452 11160 13504 11212
rect 13820 11228 13872 11280
rect 14556 11228 14608 11280
rect 14372 11160 14424 11212
rect 15016 11160 15068 11212
rect 13636 11092 13688 11144
rect 14188 11135 14240 11144
rect 14188 11101 14197 11135
rect 14197 11101 14231 11135
rect 14231 11101 14240 11135
rect 14188 11092 14240 11101
rect 10784 11024 10836 11076
rect 11336 10999 11388 11008
rect 11336 10965 11345 10999
rect 11345 10965 11379 10999
rect 11379 10965 11388 10999
rect 11336 10956 11388 10965
rect 12624 11024 12676 11076
rect 12900 11024 12952 11076
rect 12992 11067 13044 11076
rect 12992 11033 13001 11067
rect 13001 11033 13035 11067
rect 13035 11033 13044 11067
rect 12992 11024 13044 11033
rect 14280 11024 14332 11076
rect 14464 11024 14516 11076
rect 14924 11067 14976 11076
rect 14924 11033 14933 11067
rect 14933 11033 14967 11067
rect 14967 11033 14976 11067
rect 14924 11024 14976 11033
rect 16488 11024 16540 11076
rect 14096 10956 14148 11008
rect 16672 10956 16724 11008
rect 16948 10956 17000 11008
rect 17408 11135 17460 11144
rect 17408 11101 17417 11135
rect 17417 11101 17451 11135
rect 17451 11101 17460 11135
rect 17408 11092 17460 11101
rect 18512 11228 18564 11280
rect 18972 11228 19024 11280
rect 18144 11160 18196 11212
rect 19156 11160 19208 11212
rect 19340 11160 19392 11212
rect 17868 11092 17920 11144
rect 19708 11228 19760 11280
rect 20812 11228 20864 11280
rect 19984 11160 20036 11212
rect 20168 11160 20220 11212
rect 18420 11024 18472 11076
rect 18696 11024 18748 11076
rect 20996 11092 21048 11144
rect 21364 11092 21416 11144
rect 21732 11135 21784 11144
rect 21732 11101 21741 11135
rect 21741 11101 21775 11135
rect 21775 11101 21784 11135
rect 21732 11092 21784 11101
rect 24584 11135 24636 11144
rect 24584 11101 24593 11135
rect 24593 11101 24627 11135
rect 24627 11101 24636 11135
rect 24584 11092 24636 11101
rect 17868 10956 17920 11008
rect 19340 10956 19392 11008
rect 19800 10956 19852 11008
rect 20444 10956 20496 11008
rect 20904 10999 20956 11008
rect 20904 10965 20913 10999
rect 20913 10965 20947 10999
rect 20947 10965 20956 10999
rect 20904 10956 20956 10965
rect 21364 10956 21416 11008
rect 23480 11024 23532 11076
rect 25228 10999 25280 11008
rect 25228 10965 25237 10999
rect 25237 10965 25271 10999
rect 25271 10965 25280 10999
rect 25228 10956 25280 10965
rect 7950 10854 8002 10906
rect 8014 10854 8066 10906
rect 8078 10854 8130 10906
rect 8142 10854 8194 10906
rect 8206 10854 8258 10906
rect 17950 10854 18002 10906
rect 18014 10854 18066 10906
rect 18078 10854 18130 10906
rect 18142 10854 18194 10906
rect 18206 10854 18258 10906
rect 10784 10752 10836 10804
rect 11428 10752 11480 10804
rect 11796 10752 11848 10804
rect 12256 10752 12308 10804
rect 12532 10795 12584 10804
rect 12532 10761 12541 10795
rect 12541 10761 12575 10795
rect 12575 10761 12584 10795
rect 12532 10752 12584 10761
rect 13728 10752 13780 10804
rect 14372 10795 14424 10804
rect 14372 10761 14381 10795
rect 14381 10761 14415 10795
rect 14415 10761 14424 10795
rect 14372 10752 14424 10761
rect 15568 10752 15620 10804
rect 15936 10795 15988 10804
rect 15936 10761 15945 10795
rect 15945 10761 15979 10795
rect 15979 10761 15988 10795
rect 15936 10752 15988 10761
rect 16120 10752 16172 10804
rect 20628 10752 20680 10804
rect 20904 10752 20956 10804
rect 8944 10684 8996 10736
rect 10508 10684 10560 10736
rect 9220 10659 9272 10668
rect 9220 10625 9229 10659
rect 9229 10625 9263 10659
rect 9263 10625 9272 10659
rect 9220 10616 9272 10625
rect 8944 10548 8996 10600
rect 13820 10684 13872 10736
rect 13728 10616 13780 10668
rect 13360 10548 13412 10600
rect 14740 10616 14792 10668
rect 15384 10480 15436 10532
rect 15568 10480 15620 10532
rect 16672 10684 16724 10736
rect 17224 10616 17276 10668
rect 17316 10616 17368 10668
rect 19616 10684 19668 10736
rect 21456 10795 21508 10804
rect 21456 10761 21465 10795
rect 21465 10761 21499 10795
rect 21499 10761 21508 10795
rect 21456 10752 21508 10761
rect 22744 10752 22796 10804
rect 23388 10684 23440 10736
rect 17408 10548 17460 10600
rect 18696 10616 18748 10668
rect 19064 10659 19116 10668
rect 19064 10625 19073 10659
rect 19073 10625 19107 10659
rect 19107 10625 19116 10659
rect 19064 10616 19116 10625
rect 19708 10659 19760 10668
rect 19708 10625 19717 10659
rect 19717 10625 19751 10659
rect 19751 10625 19760 10659
rect 19708 10616 19760 10625
rect 21916 10616 21968 10668
rect 23480 10659 23532 10668
rect 23480 10625 23489 10659
rect 23489 10625 23523 10659
rect 23523 10625 23532 10659
rect 23480 10616 23532 10625
rect 23940 10659 23992 10668
rect 23940 10625 23949 10659
rect 23949 10625 23983 10659
rect 23983 10625 23992 10659
rect 23940 10616 23992 10625
rect 20076 10548 20128 10600
rect 22008 10591 22060 10600
rect 22008 10557 22017 10591
rect 22017 10557 22051 10591
rect 22051 10557 22060 10591
rect 22008 10548 22060 10557
rect 23664 10548 23716 10600
rect 24768 10591 24820 10600
rect 24768 10557 24777 10591
rect 24777 10557 24811 10591
rect 24811 10557 24820 10591
rect 24768 10548 24820 10557
rect 13544 10455 13596 10464
rect 13544 10421 13553 10455
rect 13553 10421 13587 10455
rect 13587 10421 13596 10455
rect 13544 10412 13596 10421
rect 14188 10412 14240 10464
rect 14832 10412 14884 10464
rect 16488 10412 16540 10464
rect 16672 10412 16724 10464
rect 18328 10412 18380 10464
rect 18696 10455 18748 10464
rect 18696 10421 18705 10455
rect 18705 10421 18739 10455
rect 18739 10421 18748 10455
rect 18696 10412 18748 10421
rect 19156 10455 19208 10464
rect 19156 10421 19165 10455
rect 19165 10421 19199 10455
rect 19199 10421 19208 10455
rect 19156 10412 19208 10421
rect 19708 10480 19760 10532
rect 20168 10412 20220 10464
rect 2950 10310 3002 10362
rect 3014 10310 3066 10362
rect 3078 10310 3130 10362
rect 3142 10310 3194 10362
rect 3206 10310 3258 10362
rect 12950 10310 13002 10362
rect 13014 10310 13066 10362
rect 13078 10310 13130 10362
rect 13142 10310 13194 10362
rect 13206 10310 13258 10362
rect 22950 10310 23002 10362
rect 23014 10310 23066 10362
rect 23078 10310 23130 10362
rect 23142 10310 23194 10362
rect 23206 10310 23258 10362
rect 12716 10251 12768 10260
rect 12716 10217 12725 10251
rect 12725 10217 12759 10251
rect 12759 10217 12768 10251
rect 12716 10208 12768 10217
rect 13728 10208 13780 10260
rect 15568 10208 15620 10260
rect 15660 10251 15712 10260
rect 15660 10217 15669 10251
rect 15669 10217 15703 10251
rect 15703 10217 15712 10251
rect 15660 10208 15712 10217
rect 16580 10208 16632 10260
rect 17316 10208 17368 10260
rect 19616 10208 19668 10260
rect 19800 10208 19852 10260
rect 12440 10140 12492 10192
rect 9128 10115 9180 10124
rect 9128 10081 9137 10115
rect 9137 10081 9171 10115
rect 9171 10081 9180 10115
rect 9128 10072 9180 10081
rect 9404 10115 9456 10124
rect 9404 10081 9413 10115
rect 9413 10081 9447 10115
rect 9447 10081 9456 10115
rect 9404 10072 9456 10081
rect 11060 10072 11112 10124
rect 11336 10072 11388 10124
rect 10508 10004 10560 10056
rect 13360 10115 13412 10124
rect 13360 10081 13369 10115
rect 13369 10081 13403 10115
rect 13403 10081 13412 10115
rect 13360 10072 13412 10081
rect 9680 9936 9732 9988
rect 8392 9911 8444 9920
rect 8392 9877 8401 9911
rect 8401 9877 8435 9911
rect 8435 9877 8444 9911
rect 8392 9868 8444 9877
rect 10416 9868 10468 9920
rect 12624 10004 12676 10056
rect 13544 10004 13596 10056
rect 14924 10072 14976 10124
rect 16028 10140 16080 10192
rect 16488 10140 16540 10192
rect 15568 10004 15620 10056
rect 17408 10115 17460 10124
rect 17408 10081 17417 10115
rect 17417 10081 17451 10115
rect 17451 10081 17460 10115
rect 17408 10072 17460 10081
rect 18420 10140 18472 10192
rect 18880 10140 18932 10192
rect 15752 9936 15804 9988
rect 11888 9911 11940 9920
rect 11888 9877 11897 9911
rect 11897 9877 11931 9911
rect 11931 9877 11940 9911
rect 11888 9868 11940 9877
rect 13820 9868 13872 9920
rect 14096 9868 14148 9920
rect 17684 10004 17736 10056
rect 18696 10072 18748 10124
rect 20076 10251 20128 10260
rect 20076 10217 20085 10251
rect 20085 10217 20119 10251
rect 20119 10217 20128 10251
rect 20076 10208 20128 10217
rect 20168 10208 20220 10260
rect 24400 10208 24452 10260
rect 25136 10251 25188 10260
rect 25136 10217 25145 10251
rect 25145 10217 25179 10251
rect 25179 10217 25188 10251
rect 25136 10208 25188 10217
rect 19984 10140 20036 10192
rect 20812 10183 20864 10192
rect 20812 10149 20821 10183
rect 20821 10149 20855 10183
rect 20855 10149 20864 10183
rect 20812 10140 20864 10149
rect 21916 10183 21968 10192
rect 21916 10149 21925 10183
rect 21925 10149 21959 10183
rect 21959 10149 21968 10183
rect 21916 10140 21968 10149
rect 24124 10140 24176 10192
rect 18880 10004 18932 10056
rect 21456 10115 21508 10124
rect 21456 10081 21465 10115
rect 21465 10081 21499 10115
rect 21499 10081 21508 10115
rect 21456 10072 21508 10081
rect 22284 10115 22336 10124
rect 22284 10081 22293 10115
rect 22293 10081 22327 10115
rect 22327 10081 22336 10115
rect 22284 10072 22336 10081
rect 25228 10072 25280 10124
rect 21088 10004 21140 10056
rect 21180 10004 21232 10056
rect 21824 10004 21876 10056
rect 20904 9936 20956 9988
rect 16580 9868 16632 9920
rect 17316 9911 17368 9920
rect 17316 9877 17325 9911
rect 17325 9877 17359 9911
rect 17359 9877 17368 9911
rect 17316 9868 17368 9877
rect 18420 9868 18472 9920
rect 19248 9868 19300 9920
rect 20628 9868 20680 9920
rect 21456 9936 21508 9988
rect 21916 9936 21968 9988
rect 24032 9911 24084 9920
rect 24032 9877 24041 9911
rect 24041 9877 24075 9911
rect 24075 9877 24084 9911
rect 24032 9868 24084 9877
rect 24584 9911 24636 9920
rect 24584 9877 24593 9911
rect 24593 9877 24627 9911
rect 24627 9877 24636 9911
rect 24584 9868 24636 9877
rect 7950 9766 8002 9818
rect 8014 9766 8066 9818
rect 8078 9766 8130 9818
rect 8142 9766 8194 9818
rect 8206 9766 8258 9818
rect 17950 9766 18002 9818
rect 18014 9766 18066 9818
rect 18078 9766 18130 9818
rect 18142 9766 18194 9818
rect 18206 9766 18258 9818
rect 3976 9664 4028 9716
rect 9312 9664 9364 9716
rect 3332 9596 3384 9648
rect 6276 9596 6328 9648
rect 10508 9664 10560 9716
rect 7104 9460 7156 9512
rect 8208 9503 8260 9512
rect 8208 9469 8217 9503
rect 8217 9469 8251 9503
rect 8251 9469 8260 9503
rect 8208 9460 8260 9469
rect 7104 9324 7156 9376
rect 11520 9596 11572 9648
rect 13544 9664 13596 9716
rect 13820 9664 13872 9716
rect 17224 9664 17276 9716
rect 17500 9664 17552 9716
rect 21456 9664 21508 9716
rect 13268 9596 13320 9648
rect 11704 9571 11756 9580
rect 11704 9537 11713 9571
rect 11713 9537 11747 9571
rect 11747 9537 11756 9571
rect 11704 9528 11756 9537
rect 13820 9528 13872 9580
rect 15200 9528 15252 9580
rect 15476 9528 15528 9580
rect 15752 9528 15804 9580
rect 16120 9571 16172 9580
rect 16120 9537 16129 9571
rect 16129 9537 16163 9571
rect 16163 9537 16172 9571
rect 16120 9528 16172 9537
rect 16948 9639 17000 9648
rect 16948 9605 16957 9639
rect 16957 9605 16991 9639
rect 16991 9605 17000 9639
rect 16948 9596 17000 9605
rect 17868 9596 17920 9648
rect 19248 9596 19300 9648
rect 19616 9596 19668 9648
rect 21272 9596 21324 9648
rect 23296 9639 23348 9648
rect 23296 9605 23305 9639
rect 23305 9605 23339 9639
rect 23339 9605 23348 9639
rect 23296 9596 23348 9605
rect 22100 9571 22152 9580
rect 22100 9537 22109 9571
rect 22109 9537 22143 9571
rect 22143 9537 22152 9571
rect 22100 9528 22152 9537
rect 23020 9528 23072 9580
rect 9956 9503 10008 9512
rect 9956 9469 9965 9503
rect 9965 9469 9999 9503
rect 9999 9469 10008 9503
rect 9956 9460 10008 9469
rect 10600 9503 10652 9512
rect 10600 9469 10609 9503
rect 10609 9469 10643 9503
rect 10643 9469 10652 9503
rect 10600 9460 10652 9469
rect 9772 9392 9824 9444
rect 13360 9460 13412 9512
rect 16396 9460 16448 9512
rect 11060 9367 11112 9376
rect 11060 9333 11069 9367
rect 11069 9333 11103 9367
rect 11103 9333 11112 9367
rect 11060 9324 11112 9333
rect 13544 9392 13596 9444
rect 14280 9392 14332 9444
rect 15568 9392 15620 9444
rect 16304 9435 16356 9444
rect 16304 9401 16313 9435
rect 16313 9401 16347 9435
rect 16347 9401 16356 9435
rect 16304 9392 16356 9401
rect 13268 9324 13320 9376
rect 15108 9324 15160 9376
rect 17040 9367 17092 9376
rect 17040 9333 17049 9367
rect 17049 9333 17083 9367
rect 17083 9333 17092 9367
rect 17040 9324 17092 9333
rect 17960 9503 18012 9512
rect 17960 9469 17969 9503
rect 17969 9469 18003 9503
rect 18003 9469 18012 9503
rect 17960 9460 18012 9469
rect 18052 9460 18104 9512
rect 18972 9460 19024 9512
rect 20168 9460 20220 9512
rect 24032 9460 24084 9512
rect 24676 9503 24728 9512
rect 24676 9469 24685 9503
rect 24685 9469 24719 9503
rect 24719 9469 24728 9503
rect 24676 9460 24728 9469
rect 20260 9392 20312 9444
rect 22284 9392 22336 9444
rect 19064 9324 19116 9376
rect 19892 9367 19944 9376
rect 19892 9333 19901 9367
rect 19901 9333 19935 9367
rect 19935 9333 19944 9367
rect 19892 9324 19944 9333
rect 20812 9324 20864 9376
rect 2950 9222 3002 9274
rect 3014 9222 3066 9274
rect 3078 9222 3130 9274
rect 3142 9222 3194 9274
rect 3206 9222 3258 9274
rect 12950 9222 13002 9274
rect 13014 9222 13066 9274
rect 13078 9222 13130 9274
rect 13142 9222 13194 9274
rect 13206 9222 13258 9274
rect 22950 9222 23002 9274
rect 23014 9222 23066 9274
rect 23078 9222 23130 9274
rect 23142 9222 23194 9274
rect 23206 9222 23258 9274
rect 9680 9120 9732 9172
rect 12440 9120 12492 9172
rect 11980 9052 12032 9104
rect 13636 9052 13688 9104
rect 13452 8984 13504 9036
rect 14096 9120 14148 9172
rect 16856 9120 16908 9172
rect 17868 9120 17920 9172
rect 17960 9120 18012 9172
rect 19892 9120 19944 9172
rect 25044 9120 25096 9172
rect 15200 9052 15252 9104
rect 18696 9052 18748 9104
rect 10416 8916 10468 8968
rect 11244 8916 11296 8968
rect 11888 8916 11940 8968
rect 16396 8984 16448 9036
rect 11428 8848 11480 8900
rect 12348 8848 12400 8900
rect 13912 8848 13964 8900
rect 8852 8780 8904 8832
rect 12256 8780 12308 8832
rect 12440 8780 12492 8832
rect 13452 8823 13504 8832
rect 13452 8789 13461 8823
rect 13461 8789 13495 8823
rect 13495 8789 13504 8823
rect 13452 8780 13504 8789
rect 13728 8780 13780 8832
rect 14556 8891 14608 8900
rect 14556 8857 14565 8891
rect 14565 8857 14599 8891
rect 14599 8857 14608 8891
rect 14556 8848 14608 8857
rect 18052 8984 18104 9036
rect 18420 8984 18472 9036
rect 16856 8916 16908 8968
rect 17684 8916 17736 8968
rect 21456 8984 21508 9036
rect 17224 8848 17276 8900
rect 21824 8891 21876 8900
rect 21824 8857 21833 8891
rect 21833 8857 21867 8891
rect 21867 8857 21876 8891
rect 21824 8848 21876 8857
rect 22376 8916 22428 8968
rect 24032 8916 24084 8968
rect 23480 8848 23532 8900
rect 24952 8848 25004 8900
rect 16488 8780 16540 8832
rect 17316 8780 17368 8832
rect 17408 8780 17460 8832
rect 17868 8780 17920 8832
rect 19064 8780 19116 8832
rect 19248 8780 19300 8832
rect 19616 8823 19668 8832
rect 19616 8789 19625 8823
rect 19625 8789 19659 8823
rect 19659 8789 19668 8823
rect 19616 8780 19668 8789
rect 22652 8780 22704 8832
rect 7950 8678 8002 8730
rect 8014 8678 8066 8730
rect 8078 8678 8130 8730
rect 8142 8678 8194 8730
rect 8206 8678 8258 8730
rect 17950 8678 18002 8730
rect 18014 8678 18066 8730
rect 18078 8678 18130 8730
rect 18142 8678 18194 8730
rect 18206 8678 18258 8730
rect 10600 8576 10652 8628
rect 8852 8551 8904 8560
rect 8852 8517 8861 8551
rect 8861 8517 8895 8551
rect 8895 8517 8904 8551
rect 8852 8508 8904 8517
rect 10416 8508 10468 8560
rect 13452 8576 13504 8628
rect 15844 8576 15896 8628
rect 17316 8576 17368 8628
rect 17776 8576 17828 8628
rect 18420 8576 18472 8628
rect 19248 8576 19300 8628
rect 8116 8483 8168 8492
rect 8116 8449 8125 8483
rect 8125 8449 8159 8483
rect 8159 8449 8168 8483
rect 8116 8440 8168 8449
rect 8300 8372 8352 8424
rect 8484 8304 8536 8356
rect 11980 8372 12032 8424
rect 12164 8415 12216 8424
rect 12164 8381 12173 8415
rect 12173 8381 12207 8415
rect 12207 8381 12216 8415
rect 12164 8372 12216 8381
rect 12808 8440 12860 8492
rect 18788 8508 18840 8560
rect 14096 8440 14148 8492
rect 12624 8372 12676 8424
rect 17776 8440 17828 8492
rect 19892 8576 19944 8628
rect 20168 8576 20220 8628
rect 20260 8508 20312 8560
rect 22008 8508 22060 8560
rect 22652 8551 22704 8560
rect 22652 8517 22661 8551
rect 22661 8517 22695 8551
rect 22695 8517 22704 8551
rect 22652 8508 22704 8517
rect 24032 8508 24084 8560
rect 14280 8415 14332 8424
rect 14280 8381 14289 8415
rect 14289 8381 14323 8415
rect 14323 8381 14332 8415
rect 14280 8372 14332 8381
rect 15108 8372 15160 8424
rect 16396 8372 16448 8424
rect 16488 8372 16540 8424
rect 11060 8304 11112 8356
rect 16764 8304 16816 8356
rect 17592 8372 17644 8424
rect 19708 8483 19760 8492
rect 19708 8449 19717 8483
rect 19717 8449 19751 8483
rect 19751 8449 19760 8483
rect 19708 8440 19760 8449
rect 18788 8415 18840 8424
rect 18788 8381 18797 8415
rect 18797 8381 18831 8415
rect 18831 8381 18840 8415
rect 18788 8372 18840 8381
rect 19248 8304 19300 8356
rect 9036 8236 9088 8288
rect 10324 8279 10376 8288
rect 10324 8245 10333 8279
rect 10333 8245 10367 8279
rect 10367 8245 10376 8279
rect 10324 8236 10376 8245
rect 13544 8279 13596 8288
rect 13544 8245 13553 8279
rect 13553 8245 13587 8279
rect 13587 8245 13596 8279
rect 13544 8236 13596 8245
rect 13820 8279 13872 8288
rect 13820 8245 13829 8279
rect 13829 8245 13863 8279
rect 13863 8245 13872 8279
rect 13820 8236 13872 8245
rect 17500 8236 17552 8288
rect 22192 8372 22244 8424
rect 22284 8372 22336 8424
rect 22744 8372 22796 8424
rect 24860 8440 24912 8492
rect 21456 8279 21508 8288
rect 21456 8245 21465 8279
rect 21465 8245 21499 8279
rect 21499 8245 21508 8279
rect 21456 8236 21508 8245
rect 22192 8236 22244 8288
rect 23388 8236 23440 8288
rect 25228 8279 25280 8288
rect 25228 8245 25237 8279
rect 25237 8245 25271 8279
rect 25271 8245 25280 8279
rect 25228 8236 25280 8245
rect 2950 8134 3002 8186
rect 3014 8134 3066 8186
rect 3078 8134 3130 8186
rect 3142 8134 3194 8186
rect 3206 8134 3258 8186
rect 12950 8134 13002 8186
rect 13014 8134 13066 8186
rect 13078 8134 13130 8186
rect 13142 8134 13194 8186
rect 13206 8134 13258 8186
rect 22950 8134 23002 8186
rect 23014 8134 23066 8186
rect 23078 8134 23130 8186
rect 23142 8134 23194 8186
rect 23206 8134 23258 8186
rect 10324 8032 10376 8084
rect 10324 7828 10376 7880
rect 8392 7760 8444 7812
rect 10876 8032 10928 8084
rect 11520 7939 11572 7948
rect 11520 7905 11529 7939
rect 11529 7905 11563 7939
rect 11563 7905 11572 7939
rect 11520 7896 11572 7905
rect 11796 8075 11848 8084
rect 11796 8041 11805 8075
rect 11805 8041 11839 8075
rect 11839 8041 11848 8075
rect 11796 8032 11848 8041
rect 16672 8032 16724 8084
rect 15568 7964 15620 8016
rect 18880 8075 18932 8084
rect 18880 8041 18889 8075
rect 18889 8041 18923 8075
rect 18923 8041 18932 8075
rect 18880 8032 18932 8041
rect 20168 8032 20220 8084
rect 20536 8032 20588 8084
rect 21088 8032 21140 8084
rect 21548 8032 21600 8084
rect 21732 7964 21784 8016
rect 12808 7896 12860 7948
rect 15016 7896 15068 7948
rect 16856 7896 16908 7948
rect 17408 7939 17460 7948
rect 17408 7905 17417 7939
rect 17417 7905 17451 7939
rect 17451 7905 17460 7939
rect 17408 7896 17460 7905
rect 18420 7896 18472 7948
rect 11980 7828 12032 7880
rect 13360 7871 13412 7880
rect 13360 7837 13369 7871
rect 13369 7837 13403 7871
rect 13403 7837 13412 7871
rect 13360 7828 13412 7837
rect 16672 7871 16724 7880
rect 16672 7837 16681 7871
rect 16681 7837 16715 7871
rect 16715 7837 16724 7871
rect 16672 7828 16724 7837
rect 18696 7828 18748 7880
rect 23204 7964 23256 8016
rect 22560 7896 22612 7948
rect 22192 7871 22244 7880
rect 22192 7837 22201 7871
rect 22201 7837 22235 7871
rect 22235 7837 22244 7871
rect 22192 7828 22244 7837
rect 9312 7692 9364 7744
rect 12348 7760 12400 7812
rect 13820 7760 13872 7812
rect 15016 7760 15068 7812
rect 18420 7760 18472 7812
rect 15568 7692 15620 7744
rect 16028 7735 16080 7744
rect 16028 7701 16037 7735
rect 16037 7701 16071 7735
rect 16071 7701 16080 7735
rect 16028 7692 16080 7701
rect 18788 7692 18840 7744
rect 22836 7692 22888 7744
rect 23388 7760 23440 7812
rect 23572 7692 23624 7744
rect 24032 7692 24084 7744
rect 7950 7590 8002 7642
rect 8014 7590 8066 7642
rect 8078 7590 8130 7642
rect 8142 7590 8194 7642
rect 8206 7590 8258 7642
rect 17950 7590 18002 7642
rect 18014 7590 18066 7642
rect 18078 7590 18130 7642
rect 18142 7590 18194 7642
rect 18206 7590 18258 7642
rect 10876 7488 10928 7540
rect 12348 7488 12400 7540
rect 12716 7488 12768 7540
rect 15476 7531 15528 7540
rect 15476 7497 15485 7531
rect 15485 7497 15519 7531
rect 15519 7497 15528 7531
rect 15476 7488 15528 7497
rect 16396 7488 16448 7540
rect 17500 7531 17552 7540
rect 17500 7497 17509 7531
rect 17509 7497 17543 7531
rect 17543 7497 17552 7531
rect 17500 7488 17552 7497
rect 17776 7488 17828 7540
rect 21916 7488 21968 7540
rect 23204 7488 23256 7540
rect 24952 7488 25004 7540
rect 9312 7463 9364 7472
rect 9312 7429 9321 7463
rect 9321 7429 9355 7463
rect 9355 7429 9364 7463
rect 9312 7420 9364 7429
rect 15108 7420 15160 7472
rect 11060 7352 11112 7404
rect 9036 7327 9088 7336
rect 9036 7293 9045 7327
rect 9045 7293 9079 7327
rect 9079 7293 9088 7327
rect 9036 7284 9088 7293
rect 12072 7395 12124 7404
rect 12072 7361 12081 7395
rect 12081 7361 12115 7395
rect 12115 7361 12124 7395
rect 12072 7352 12124 7361
rect 18144 7352 18196 7404
rect 12256 7327 12308 7336
rect 12256 7293 12265 7327
rect 12265 7293 12299 7327
rect 12299 7293 12308 7327
rect 12256 7284 12308 7293
rect 12348 7284 12400 7336
rect 13636 7327 13688 7336
rect 13636 7293 13645 7327
rect 13645 7293 13679 7327
rect 13679 7293 13688 7327
rect 13636 7284 13688 7293
rect 15568 7327 15620 7336
rect 15568 7293 15577 7327
rect 15577 7293 15611 7327
rect 15611 7293 15620 7327
rect 15568 7284 15620 7293
rect 16948 7284 17000 7336
rect 17316 7284 17368 7336
rect 17684 7327 17736 7336
rect 17684 7293 17693 7327
rect 17693 7293 17727 7327
rect 17727 7293 17736 7327
rect 17684 7284 17736 7293
rect 13360 7216 13412 7268
rect 13452 7216 13504 7268
rect 18788 7352 18840 7404
rect 25136 7463 25188 7472
rect 25136 7429 25145 7463
rect 25145 7429 25179 7463
rect 25179 7429 25188 7463
rect 25136 7420 25188 7429
rect 22468 7352 22520 7404
rect 21916 7284 21968 7336
rect 23296 7327 23348 7336
rect 23296 7293 23305 7327
rect 23305 7293 23339 7327
rect 23339 7293 23348 7327
rect 23296 7284 23348 7293
rect 22008 7216 22060 7268
rect 11980 7148 12032 7200
rect 14004 7148 14056 7200
rect 15016 7191 15068 7200
rect 15016 7157 15025 7191
rect 15025 7157 15059 7191
rect 15059 7157 15068 7191
rect 15016 7148 15068 7157
rect 15200 7148 15252 7200
rect 16120 7191 16172 7200
rect 16120 7157 16129 7191
rect 16129 7157 16163 7191
rect 16163 7157 16172 7191
rect 16120 7148 16172 7157
rect 16396 7148 16448 7200
rect 18144 7148 18196 7200
rect 21272 7148 21324 7200
rect 22100 7148 22152 7200
rect 23756 7148 23808 7200
rect 2950 7046 3002 7098
rect 3014 7046 3066 7098
rect 3078 7046 3130 7098
rect 3142 7046 3194 7098
rect 3206 7046 3258 7098
rect 12950 7046 13002 7098
rect 13014 7046 13066 7098
rect 13078 7046 13130 7098
rect 13142 7046 13194 7098
rect 13206 7046 13258 7098
rect 22950 7046 23002 7098
rect 23014 7046 23066 7098
rect 23078 7046 23130 7098
rect 23142 7046 23194 7098
rect 23206 7046 23258 7098
rect 9312 6944 9364 6996
rect 12808 6944 12860 6996
rect 15200 6987 15252 6996
rect 15200 6953 15209 6987
rect 15209 6953 15243 6987
rect 15243 6953 15252 6987
rect 15200 6944 15252 6953
rect 12716 6876 12768 6928
rect 13360 6876 13412 6928
rect 17868 6944 17920 6996
rect 22100 6944 22152 6996
rect 25228 6944 25280 6996
rect 15844 6876 15896 6928
rect 17776 6876 17828 6928
rect 21548 6919 21600 6928
rect 21548 6885 21557 6919
rect 21557 6885 21591 6919
rect 21591 6885 21600 6919
rect 21548 6876 21600 6885
rect 23388 6876 23440 6928
rect 24860 6876 24912 6928
rect 5264 6808 5316 6860
rect 10048 6808 10100 6860
rect 11612 6808 11664 6860
rect 12440 6808 12492 6860
rect 11980 6740 12032 6792
rect 16028 6808 16080 6860
rect 16948 6851 17000 6860
rect 16948 6817 16957 6851
rect 16957 6817 16991 6851
rect 16991 6817 17000 6851
rect 16948 6808 17000 6817
rect 19708 6808 19760 6860
rect 22284 6808 22336 6860
rect 22744 6808 22796 6860
rect 25044 6851 25096 6860
rect 25044 6817 25053 6851
rect 25053 6817 25087 6851
rect 25087 6817 25096 6851
rect 25044 6808 25096 6817
rect 15016 6740 15068 6792
rect 11152 6672 11204 6724
rect 15660 6715 15712 6724
rect 15660 6681 15669 6715
rect 15669 6681 15703 6715
rect 15703 6681 15712 6715
rect 15660 6672 15712 6681
rect 16028 6672 16080 6724
rect 16764 6740 16816 6792
rect 17132 6740 17184 6792
rect 2044 6604 2096 6656
rect 8760 6604 8812 6656
rect 12992 6647 13044 6656
rect 12992 6613 13001 6647
rect 13001 6613 13035 6647
rect 13035 6613 13044 6647
rect 12992 6604 13044 6613
rect 13360 6647 13412 6656
rect 13360 6613 13369 6647
rect 13369 6613 13403 6647
rect 13403 6613 13412 6647
rect 13360 6604 13412 6613
rect 13544 6604 13596 6656
rect 15292 6604 15344 6656
rect 18972 6672 19024 6724
rect 19984 6672 20036 6724
rect 24032 6647 24084 6656
rect 24032 6613 24041 6647
rect 24041 6613 24075 6647
rect 24075 6613 24084 6647
rect 24032 6604 24084 6613
rect 24584 6647 24636 6656
rect 24584 6613 24593 6647
rect 24593 6613 24627 6647
rect 24627 6613 24636 6647
rect 24584 6604 24636 6613
rect 24952 6647 25004 6656
rect 24952 6613 24961 6647
rect 24961 6613 24995 6647
rect 24995 6613 25004 6647
rect 24952 6604 25004 6613
rect 7950 6502 8002 6554
rect 8014 6502 8066 6554
rect 8078 6502 8130 6554
rect 8142 6502 8194 6554
rect 8206 6502 8258 6554
rect 17950 6502 18002 6554
rect 18014 6502 18066 6554
rect 18078 6502 18130 6554
rect 18142 6502 18194 6554
rect 18206 6502 18258 6554
rect 11152 6400 11204 6452
rect 12992 6400 13044 6452
rect 13544 6332 13596 6384
rect 13820 6332 13872 6384
rect 22100 6400 22152 6452
rect 22284 6400 22336 6452
rect 10876 6264 10928 6316
rect 11704 6307 11756 6316
rect 11704 6273 11713 6307
rect 11713 6273 11747 6307
rect 11747 6273 11756 6307
rect 11704 6264 11756 6273
rect 12256 6264 12308 6316
rect 15016 6264 15068 6316
rect 17132 6332 17184 6384
rect 18144 6332 18196 6384
rect 16120 6264 16172 6316
rect 11612 6196 11664 6248
rect 2228 6128 2280 6180
rect 12164 6128 12216 6180
rect 10232 6060 10284 6112
rect 11980 6060 12032 6112
rect 13728 6196 13780 6248
rect 13728 6060 13780 6112
rect 15200 6196 15252 6248
rect 15568 6196 15620 6248
rect 14372 6128 14424 6180
rect 16856 6307 16908 6316
rect 16856 6273 16865 6307
rect 16865 6273 16899 6307
rect 16899 6273 16908 6307
rect 16856 6264 16908 6273
rect 19340 6264 19392 6316
rect 24860 6332 24912 6384
rect 23940 6307 23992 6316
rect 23940 6273 23949 6307
rect 23949 6273 23983 6307
rect 23983 6273 23992 6307
rect 23940 6264 23992 6273
rect 17132 6239 17184 6248
rect 17132 6205 17141 6239
rect 17141 6205 17175 6239
rect 17175 6205 17184 6239
rect 17132 6196 17184 6205
rect 17684 6196 17736 6248
rect 22468 6239 22520 6248
rect 22468 6205 22477 6239
rect 22477 6205 22511 6239
rect 22511 6205 22520 6239
rect 22468 6196 22520 6205
rect 24676 6239 24728 6248
rect 24676 6205 24685 6239
rect 24685 6205 24719 6239
rect 24719 6205 24728 6239
rect 24676 6196 24728 6205
rect 19616 6128 19668 6180
rect 20352 6128 20404 6180
rect 22100 6128 22152 6180
rect 18144 6060 18196 6112
rect 18420 6060 18472 6112
rect 19984 6060 20036 6112
rect 2950 5958 3002 6010
rect 3014 5958 3066 6010
rect 3078 5958 3130 6010
rect 3142 5958 3194 6010
rect 3206 5958 3258 6010
rect 12950 5958 13002 6010
rect 13014 5958 13066 6010
rect 13078 5958 13130 6010
rect 13142 5958 13194 6010
rect 13206 5958 13258 6010
rect 22950 5958 23002 6010
rect 23014 5958 23066 6010
rect 23078 5958 23130 6010
rect 23142 5958 23194 6010
rect 23206 5958 23258 6010
rect 11704 5899 11756 5908
rect 11704 5865 11713 5899
rect 11713 5865 11747 5899
rect 11747 5865 11756 5899
rect 11704 5856 11756 5865
rect 17132 5856 17184 5908
rect 10232 5763 10284 5772
rect 10232 5729 10241 5763
rect 10241 5729 10275 5763
rect 10275 5729 10284 5763
rect 10232 5720 10284 5729
rect 11244 5720 11296 5772
rect 23940 5856 23992 5908
rect 17408 5788 17460 5840
rect 24952 5856 25004 5908
rect 19984 5763 20036 5772
rect 19984 5729 19993 5763
rect 19993 5729 20027 5763
rect 20027 5729 20036 5763
rect 19984 5720 20036 5729
rect 20260 5720 20312 5772
rect 22652 5763 22704 5772
rect 22652 5729 22661 5763
rect 22661 5729 22695 5763
rect 22695 5729 22704 5763
rect 22652 5720 22704 5729
rect 8300 5652 8352 5704
rect 9036 5652 9088 5704
rect 12716 5652 12768 5704
rect 9588 5584 9640 5636
rect 14372 5695 14424 5704
rect 14372 5661 14381 5695
rect 14381 5661 14415 5695
rect 14415 5661 14424 5695
rect 14372 5652 14424 5661
rect 15200 5652 15252 5704
rect 17592 5652 17644 5704
rect 20352 5652 20404 5704
rect 17224 5584 17276 5636
rect 17868 5584 17920 5636
rect 18696 5627 18748 5636
rect 18696 5593 18705 5627
rect 18705 5593 18739 5627
rect 18739 5593 18748 5627
rect 18696 5584 18748 5593
rect 11980 5559 12032 5568
rect 11980 5525 11989 5559
rect 11989 5525 12023 5559
rect 12023 5525 12032 5559
rect 11980 5516 12032 5525
rect 12348 5559 12400 5568
rect 12348 5525 12357 5559
rect 12357 5525 12391 5559
rect 12391 5525 12400 5559
rect 12348 5516 12400 5525
rect 14004 5516 14056 5568
rect 15108 5516 15160 5568
rect 16304 5516 16356 5568
rect 18512 5516 18564 5568
rect 20444 5584 20496 5636
rect 22284 5695 22336 5704
rect 22284 5661 22293 5695
rect 22293 5661 22327 5695
rect 22327 5661 22336 5695
rect 22284 5652 22336 5661
rect 23388 5652 23440 5704
rect 20904 5584 20956 5636
rect 19800 5516 19852 5568
rect 20076 5516 20128 5568
rect 21548 5516 21600 5568
rect 24032 5516 24084 5568
rect 24216 5516 24268 5568
rect 7950 5414 8002 5466
rect 8014 5414 8066 5466
rect 8078 5414 8130 5466
rect 8142 5414 8194 5466
rect 8206 5414 8258 5466
rect 17950 5414 18002 5466
rect 18014 5414 18066 5466
rect 18078 5414 18130 5466
rect 18142 5414 18194 5466
rect 18206 5414 18258 5466
rect 13544 5312 13596 5364
rect 10508 5244 10560 5296
rect 11152 5219 11204 5228
rect 11152 5185 11161 5219
rect 11161 5185 11195 5219
rect 11195 5185 11204 5219
rect 11152 5176 11204 5185
rect 13268 5244 13320 5296
rect 14004 5287 14056 5296
rect 14004 5253 14013 5287
rect 14013 5253 14047 5287
rect 14047 5253 14056 5287
rect 14004 5244 14056 5253
rect 15384 5244 15436 5296
rect 13728 5219 13780 5228
rect 13728 5185 13737 5219
rect 13737 5185 13771 5219
rect 13771 5185 13780 5219
rect 13728 5176 13780 5185
rect 15108 5176 15160 5228
rect 18604 5244 18656 5296
rect 24216 5312 24268 5364
rect 16856 5219 16908 5228
rect 16856 5185 16865 5219
rect 16865 5185 16899 5219
rect 16899 5185 16908 5219
rect 16856 5176 16908 5185
rect 20076 5244 20128 5296
rect 19708 5219 19760 5228
rect 19708 5185 19717 5219
rect 19717 5185 19751 5219
rect 19751 5185 19760 5219
rect 19708 5176 19760 5185
rect 10968 5108 11020 5160
rect 15844 5108 15896 5160
rect 18604 5108 18656 5160
rect 20444 5108 20496 5160
rect 23664 5176 23716 5228
rect 9496 5040 9548 5092
rect 13268 5040 13320 5092
rect 12808 4972 12860 5024
rect 15200 4972 15252 5024
rect 15476 5015 15528 5024
rect 15476 4981 15485 5015
rect 15485 4981 15519 5015
rect 15519 4981 15528 5015
rect 15476 4972 15528 4981
rect 19340 5040 19392 5092
rect 24768 5151 24820 5160
rect 24768 5117 24777 5151
rect 24777 5117 24811 5151
rect 24811 5117 24820 5151
rect 24768 5108 24820 5117
rect 18236 4972 18288 5024
rect 20720 4972 20772 5024
rect 21456 5015 21508 5024
rect 21456 4981 21465 5015
rect 21465 4981 21499 5015
rect 21499 4981 21508 5015
rect 21456 4972 21508 4981
rect 2950 4870 3002 4922
rect 3014 4870 3066 4922
rect 3078 4870 3130 4922
rect 3142 4870 3194 4922
rect 3206 4870 3258 4922
rect 12950 4870 13002 4922
rect 13014 4870 13066 4922
rect 13078 4870 13130 4922
rect 13142 4870 13194 4922
rect 13206 4870 13258 4922
rect 22950 4870 23002 4922
rect 23014 4870 23066 4922
rect 23078 4870 23130 4922
rect 23142 4870 23194 4922
rect 23206 4870 23258 4922
rect 8852 4768 8904 4820
rect 9772 4700 9824 4752
rect 12808 4768 12860 4820
rect 16672 4768 16724 4820
rect 16948 4768 17000 4820
rect 23756 4811 23808 4820
rect 23756 4777 23765 4811
rect 23765 4777 23799 4811
rect 23799 4777 23808 4811
rect 23756 4768 23808 4777
rect 8208 4632 8260 4684
rect 8484 4632 8536 4684
rect 11888 4675 11940 4684
rect 11888 4641 11897 4675
rect 11897 4641 11931 4675
rect 11931 4641 11940 4675
rect 11888 4632 11940 4641
rect 13452 4632 13504 4684
rect 14648 4700 14700 4752
rect 16488 4700 16540 4752
rect 21088 4700 21140 4752
rect 25044 4700 25096 4752
rect 14372 4632 14424 4684
rect 7104 4607 7156 4616
rect 7104 4573 7113 4607
rect 7113 4573 7147 4607
rect 7147 4573 7156 4607
rect 7104 4564 7156 4573
rect 9956 4564 10008 4616
rect 10416 4564 10468 4616
rect 16856 4632 16908 4684
rect 5356 4539 5408 4548
rect 5356 4505 5365 4539
rect 5365 4505 5399 4539
rect 5399 4505 5408 4539
rect 5356 4496 5408 4505
rect 9588 4496 9640 4548
rect 16672 4564 16724 4616
rect 18328 4632 18380 4684
rect 18788 4632 18840 4684
rect 21732 4675 21784 4684
rect 21732 4641 21741 4675
rect 21741 4641 21775 4675
rect 21775 4641 21784 4675
rect 21732 4632 21784 4641
rect 19156 4564 19208 4616
rect 20536 4564 20588 4616
rect 21364 4607 21416 4616
rect 21364 4573 21373 4607
rect 21373 4573 21407 4607
rect 21407 4573 21416 4607
rect 21364 4564 21416 4573
rect 21456 4564 21508 4616
rect 15292 4496 15344 4548
rect 15384 4539 15436 4548
rect 15384 4505 15393 4539
rect 15393 4505 15427 4539
rect 15427 4505 15436 4539
rect 15384 4496 15436 4505
rect 1492 4471 1544 4480
rect 1492 4437 1501 4471
rect 1501 4437 1535 4471
rect 1535 4437 1544 4471
rect 1492 4428 1544 4437
rect 10968 4471 11020 4480
rect 10968 4437 10977 4471
rect 10977 4437 11011 4471
rect 11011 4437 11020 4471
rect 10968 4428 11020 4437
rect 14464 4471 14516 4480
rect 14464 4437 14473 4471
rect 14473 4437 14507 4471
rect 14507 4437 14516 4471
rect 14464 4428 14516 4437
rect 15108 4428 15160 4480
rect 18328 4539 18380 4548
rect 18328 4505 18337 4539
rect 18337 4505 18371 4539
rect 18371 4505 18380 4539
rect 18328 4496 18380 4505
rect 19064 4496 19116 4548
rect 7950 4326 8002 4378
rect 8014 4326 8066 4378
rect 8078 4326 8130 4378
rect 8142 4326 8194 4378
rect 8206 4326 8258 4378
rect 17950 4326 18002 4378
rect 18014 4326 18066 4378
rect 18078 4326 18130 4378
rect 18142 4326 18194 4378
rect 18206 4326 18258 4378
rect 11152 4224 11204 4276
rect 7288 4199 7340 4208
rect 7288 4165 7297 4199
rect 7297 4165 7331 4199
rect 7331 4165 7340 4199
rect 7288 4156 7340 4165
rect 13544 4224 13596 4276
rect 21180 4224 21232 4276
rect 21364 4224 21416 4276
rect 22284 4224 22336 4276
rect 1492 4088 1544 4140
rect 1860 4088 1912 4140
rect 4068 4088 4120 4140
rect 6644 4088 6696 4140
rect 5356 3952 5408 4004
rect 2228 3927 2280 3936
rect 2228 3893 2237 3927
rect 2237 3893 2271 3927
rect 2271 3893 2280 3927
rect 2228 3884 2280 3893
rect 2872 3927 2924 3936
rect 2872 3893 2881 3927
rect 2881 3893 2915 3927
rect 2915 3893 2924 3927
rect 2872 3884 2924 3893
rect 6184 3952 6236 4004
rect 6092 3927 6144 3936
rect 6092 3893 6101 3927
rect 6101 3893 6135 3927
rect 6135 3893 6144 3927
rect 6092 3884 6144 3893
rect 6368 3884 6420 3936
rect 8392 4020 8444 4072
rect 8852 4131 8904 4140
rect 8852 4097 8861 4131
rect 8861 4097 8895 4131
rect 8895 4097 8904 4131
rect 8852 4088 8904 4097
rect 9220 4088 9272 4140
rect 8576 4020 8628 4072
rect 10416 4020 10468 4072
rect 10600 4131 10652 4140
rect 10600 4097 10609 4131
rect 10609 4097 10643 4131
rect 10643 4097 10652 4131
rect 10600 4088 10652 4097
rect 12992 4131 13044 4140
rect 12992 4097 13001 4131
rect 13001 4097 13035 4131
rect 13035 4097 13044 4131
rect 12992 4088 13044 4097
rect 15568 4156 15620 4208
rect 18420 4156 18472 4208
rect 19064 4156 19116 4208
rect 21088 4156 21140 4208
rect 12256 4020 12308 4072
rect 12808 4020 12860 4072
rect 13912 4020 13964 4072
rect 14372 4020 14424 4072
rect 15476 4020 15528 4072
rect 12072 3952 12124 4004
rect 15384 3952 15436 4004
rect 18512 4088 18564 4140
rect 21548 4131 21600 4140
rect 21548 4097 21557 4131
rect 21557 4097 21591 4131
rect 21591 4097 21600 4131
rect 21548 4088 21600 4097
rect 22100 4131 22152 4140
rect 22100 4097 22109 4131
rect 22109 4097 22143 4131
rect 22143 4097 22152 4131
rect 22100 4088 22152 4097
rect 16120 4063 16172 4072
rect 16120 4029 16129 4063
rect 16129 4029 16163 4063
rect 16163 4029 16172 4063
rect 16120 4020 16172 4029
rect 16212 4020 16264 4072
rect 18420 4020 18472 4072
rect 19248 4020 19300 4072
rect 21456 4020 21508 4072
rect 22928 4199 22980 4208
rect 22928 4165 22937 4199
rect 22937 4165 22971 4199
rect 22971 4165 22980 4199
rect 22928 4156 22980 4165
rect 22836 4088 22888 4140
rect 16856 3952 16908 4004
rect 19984 3952 20036 4004
rect 22928 3952 22980 4004
rect 7380 3884 7432 3936
rect 8668 3927 8720 3936
rect 8668 3893 8677 3927
rect 8677 3893 8711 3927
rect 8711 3893 8720 3927
rect 8668 3884 8720 3893
rect 9312 3927 9364 3936
rect 9312 3893 9321 3927
rect 9321 3893 9355 3927
rect 9355 3893 9364 3927
rect 9312 3884 9364 3893
rect 9956 3927 10008 3936
rect 9956 3893 9965 3927
rect 9965 3893 9999 3927
rect 9999 3893 10008 3927
rect 9956 3884 10008 3893
rect 11612 3927 11664 3936
rect 11612 3893 11621 3927
rect 11621 3893 11655 3927
rect 11655 3893 11664 3927
rect 11612 3884 11664 3893
rect 12716 3884 12768 3936
rect 21548 3884 21600 3936
rect 24032 3884 24084 3936
rect 2950 3782 3002 3834
rect 3014 3782 3066 3834
rect 3078 3782 3130 3834
rect 3142 3782 3194 3834
rect 3206 3782 3258 3834
rect 12950 3782 13002 3834
rect 13014 3782 13066 3834
rect 13078 3782 13130 3834
rect 13142 3782 13194 3834
rect 13206 3782 13258 3834
rect 22950 3782 23002 3834
rect 23014 3782 23066 3834
rect 23078 3782 23130 3834
rect 23142 3782 23194 3834
rect 23206 3782 23258 3834
rect 3792 3680 3844 3732
rect 6920 3680 6972 3732
rect 8668 3680 8720 3732
rect 14280 3680 14332 3732
rect 18604 3723 18656 3732
rect 18604 3689 18613 3723
rect 18613 3689 18647 3723
rect 18647 3689 18656 3723
rect 18604 3680 18656 3689
rect 19524 3680 19576 3732
rect 21732 3680 21784 3732
rect 22744 3680 22796 3732
rect 6368 3655 6420 3664
rect 6368 3621 6377 3655
rect 6377 3621 6411 3655
rect 6411 3621 6420 3655
rect 6368 3612 6420 3621
rect 6460 3612 6512 3664
rect 10140 3612 10192 3664
rect 10508 3612 10560 3664
rect 2044 3544 2096 3596
rect 2872 3544 2924 3596
rect 3700 3544 3752 3596
rect 5172 3587 5224 3596
rect 5172 3553 5181 3587
rect 5181 3553 5215 3587
rect 5215 3553 5224 3587
rect 5172 3544 5224 3553
rect 2228 3476 2280 3528
rect 4436 3519 4488 3528
rect 4436 3485 4445 3519
rect 4445 3485 4479 3519
rect 4479 3485 4488 3519
rect 4436 3476 4488 3485
rect 4896 3519 4948 3528
rect 4896 3485 4905 3519
rect 4905 3485 4939 3519
rect 4939 3485 4948 3519
rect 4896 3476 4948 3485
rect 6276 3476 6328 3528
rect 7012 3476 7064 3528
rect 7288 3519 7340 3528
rect 7288 3485 7297 3519
rect 7297 3485 7331 3519
rect 7331 3485 7340 3519
rect 7288 3476 7340 3485
rect 8484 3476 8536 3528
rect 9772 3587 9824 3596
rect 9772 3553 9781 3587
rect 9781 3553 9815 3587
rect 9815 3553 9824 3587
rect 9772 3544 9824 3553
rect 15016 3612 15068 3664
rect 17408 3612 17460 3664
rect 18328 3612 18380 3664
rect 18696 3612 18748 3664
rect 14004 3544 14056 3596
rect 15476 3544 15528 3596
rect 17684 3544 17736 3596
rect 9588 3476 9640 3528
rect 10600 3519 10652 3528
rect 10600 3485 10609 3519
rect 10609 3485 10643 3519
rect 10643 3485 10652 3519
rect 10600 3476 10652 3485
rect 12348 3476 12400 3528
rect 13912 3476 13964 3528
rect 14648 3476 14700 3528
rect 16672 3476 16724 3528
rect 16948 3476 17000 3528
rect 20812 3476 20864 3528
rect 20996 3476 21048 3528
rect 3332 3383 3384 3392
rect 3332 3349 3341 3383
rect 3341 3349 3375 3383
rect 3375 3349 3384 3383
rect 3332 3340 3384 3349
rect 7196 3340 7248 3392
rect 7748 3383 7800 3392
rect 7748 3349 7757 3383
rect 7757 3349 7791 3383
rect 7791 3349 7800 3383
rect 7748 3340 7800 3349
rect 8576 3340 8628 3392
rect 12624 3408 12676 3460
rect 17592 3408 17644 3460
rect 19156 3408 19208 3460
rect 22836 3544 22888 3596
rect 23480 3680 23532 3732
rect 24860 3655 24912 3664
rect 24860 3621 24869 3655
rect 24869 3621 24903 3655
rect 24903 3621 24912 3655
rect 24860 3612 24912 3621
rect 24400 3476 24452 3528
rect 9312 3340 9364 3392
rect 13360 3340 13412 3392
rect 17316 3340 17368 3392
rect 18880 3383 18932 3392
rect 18880 3349 18889 3383
rect 18889 3349 18923 3383
rect 18923 3349 18932 3383
rect 18880 3340 18932 3349
rect 18972 3340 19024 3392
rect 23204 3340 23256 3392
rect 7950 3238 8002 3290
rect 8014 3238 8066 3290
rect 8078 3238 8130 3290
rect 8142 3238 8194 3290
rect 8206 3238 8258 3290
rect 17950 3238 18002 3290
rect 18014 3238 18066 3290
rect 18078 3238 18130 3290
rect 18142 3238 18194 3290
rect 18206 3238 18258 3290
rect 4436 3136 4488 3188
rect 4896 3136 4948 3188
rect 8944 3136 8996 3188
rect 9312 3068 9364 3120
rect 9772 3068 9824 3120
rect 2596 3000 2648 3052
rect 3332 3000 3384 3052
rect 5080 3000 5132 3052
rect 5448 3043 5500 3052
rect 5448 3009 5457 3043
rect 5457 3009 5491 3043
rect 5491 3009 5500 3043
rect 5448 3000 5500 3009
rect 5172 2975 5224 2984
rect 5172 2941 5181 2975
rect 5181 2941 5215 2975
rect 5215 2941 5224 2975
rect 5172 2932 5224 2941
rect 7380 3043 7432 3052
rect 7380 3009 7389 3043
rect 7389 3009 7423 3043
rect 7423 3009 7432 3043
rect 7380 3000 7432 3009
rect 7748 3000 7800 3052
rect 13636 3136 13688 3188
rect 16120 3136 16172 3188
rect 16580 3068 16632 3120
rect 7656 2932 7708 2984
rect 10692 2932 10744 2984
rect 11152 3047 11204 3052
rect 11152 3013 11161 3047
rect 11161 3013 11195 3047
rect 11195 3013 11204 3047
rect 11152 3000 11204 3013
rect 11612 3000 11664 3052
rect 12532 3000 12584 3052
rect 13176 3043 13228 3052
rect 13176 3009 13185 3043
rect 13185 3009 13219 3043
rect 13219 3009 13228 3043
rect 13176 3000 13228 3009
rect 14556 3000 14608 3052
rect 17132 3000 17184 3052
rect 12164 2932 12216 2984
rect 13636 2975 13688 2984
rect 13636 2941 13645 2975
rect 13645 2941 13679 2975
rect 13679 2941 13688 2975
rect 13636 2932 13688 2941
rect 14740 2932 14792 2984
rect 15844 2932 15896 2984
rect 19248 3000 19300 3052
rect 6460 2864 6512 2916
rect 6736 2864 6788 2916
rect 8852 2864 8904 2916
rect 10324 2839 10376 2848
rect 10324 2805 10333 2839
rect 10333 2805 10367 2839
rect 10367 2805 10376 2839
rect 10324 2796 10376 2805
rect 11152 2796 11204 2848
rect 11796 2796 11848 2848
rect 15108 2864 15160 2916
rect 17316 2864 17368 2916
rect 19892 3136 19944 3188
rect 20168 3068 20220 3120
rect 21272 3179 21324 3188
rect 21272 3145 21281 3179
rect 21281 3145 21315 3179
rect 21315 3145 21324 3179
rect 21272 3136 21324 3145
rect 22192 3179 22244 3188
rect 22192 3145 22201 3179
rect 22201 3145 22235 3179
rect 22235 3145 22244 3179
rect 22192 3136 22244 3145
rect 22928 3179 22980 3188
rect 22928 3145 22937 3179
rect 22937 3145 22971 3179
rect 22971 3145 22980 3179
rect 22928 3136 22980 3145
rect 24032 3136 24084 3188
rect 23388 3068 23440 3120
rect 21364 3000 21416 3052
rect 24308 3000 24360 3052
rect 24768 3000 24820 3052
rect 21732 2932 21784 2984
rect 22468 2932 22520 2984
rect 23296 2864 23348 2916
rect 15752 2796 15804 2848
rect 16948 2796 17000 2848
rect 19892 2796 19944 2848
rect 21364 2796 21416 2848
rect 22652 2796 22704 2848
rect 2950 2694 3002 2746
rect 3014 2694 3066 2746
rect 3078 2694 3130 2746
rect 3142 2694 3194 2746
rect 3206 2694 3258 2746
rect 12950 2694 13002 2746
rect 13014 2694 13066 2746
rect 13078 2694 13130 2746
rect 13142 2694 13194 2746
rect 13206 2694 13258 2746
rect 22950 2694 23002 2746
rect 23014 2694 23066 2746
rect 23078 2694 23130 2746
rect 23142 2694 23194 2746
rect 23206 2694 23258 2746
rect 6736 2592 6788 2644
rect 10048 2592 10100 2644
rect 13820 2592 13872 2644
rect 13912 2592 13964 2644
rect 20904 2592 20956 2644
rect 21272 2635 21324 2644
rect 21272 2601 21281 2635
rect 21281 2601 21315 2635
rect 21315 2601 21324 2635
rect 21272 2592 21324 2601
rect 23848 2635 23900 2644
rect 23848 2601 23857 2635
rect 23857 2601 23891 2635
rect 23891 2601 23900 2635
rect 23848 2592 23900 2601
rect 24768 2592 24820 2644
rect 8208 2524 8260 2576
rect 5264 2456 5316 2508
rect 2872 2431 2924 2440
rect 2872 2397 2881 2431
rect 2881 2397 2915 2431
rect 2915 2397 2924 2431
rect 2872 2388 2924 2397
rect 2964 2320 3016 2372
rect 6092 2388 6144 2440
rect 7840 2388 7892 2440
rect 5908 2320 5960 2372
rect 2596 2252 2648 2304
rect 5172 2252 5224 2304
rect 7104 2295 7156 2304
rect 7104 2261 7113 2295
rect 7113 2261 7147 2295
rect 7147 2261 7156 2295
rect 7104 2252 7156 2261
rect 8392 2295 8444 2304
rect 8392 2261 8401 2295
rect 8401 2261 8435 2295
rect 8435 2261 8444 2295
rect 8392 2252 8444 2261
rect 12348 2388 12400 2440
rect 10968 2320 11020 2372
rect 13268 2363 13320 2372
rect 13268 2329 13277 2363
rect 13277 2329 13311 2363
rect 13311 2329 13320 2363
rect 13268 2320 13320 2329
rect 13820 2320 13872 2372
rect 14188 2320 14240 2372
rect 10324 2252 10376 2304
rect 14464 2431 14516 2440
rect 14464 2397 14473 2431
rect 14473 2397 14507 2431
rect 14507 2397 14516 2431
rect 14464 2388 14516 2397
rect 14372 2320 14424 2372
rect 16120 2295 16172 2304
rect 16120 2261 16129 2295
rect 16129 2261 16163 2295
rect 16163 2261 16172 2295
rect 16120 2252 16172 2261
rect 16396 2524 16448 2576
rect 17316 2499 17368 2508
rect 17316 2465 17325 2499
rect 17325 2465 17359 2499
rect 17359 2465 17368 2499
rect 17316 2456 17368 2465
rect 16764 2388 16816 2440
rect 17040 2431 17092 2440
rect 17040 2397 17049 2431
rect 17049 2397 17083 2431
rect 17083 2397 17092 2431
rect 17040 2388 17092 2397
rect 17224 2388 17276 2440
rect 18880 2431 18932 2440
rect 18880 2397 18889 2431
rect 18889 2397 18923 2431
rect 18923 2397 18932 2431
rect 18880 2388 18932 2397
rect 17500 2320 17552 2372
rect 19892 2499 19944 2508
rect 19892 2465 19901 2499
rect 19901 2465 19935 2499
rect 19935 2465 19944 2499
rect 19892 2456 19944 2465
rect 19616 2431 19668 2440
rect 19616 2397 19625 2431
rect 19625 2397 19659 2431
rect 19659 2397 19668 2431
rect 19616 2388 19668 2397
rect 21640 2524 21692 2576
rect 21548 2456 21600 2508
rect 22008 2431 22060 2440
rect 22008 2397 22017 2431
rect 22017 2397 22051 2431
rect 22051 2397 22060 2431
rect 22008 2388 22060 2397
rect 19064 2252 19116 2304
rect 22100 2320 22152 2372
rect 24768 2295 24820 2304
rect 24768 2261 24777 2295
rect 24777 2261 24811 2295
rect 24811 2261 24820 2295
rect 24768 2252 24820 2261
rect 7950 2150 8002 2202
rect 8014 2150 8066 2202
rect 8078 2150 8130 2202
rect 8142 2150 8194 2202
rect 8206 2150 8258 2202
rect 17950 2150 18002 2202
rect 18014 2150 18066 2202
rect 18078 2150 18130 2202
rect 18142 2150 18194 2202
rect 18206 2150 18258 2202
rect 8392 2048 8444 2100
rect 11336 2048 11388 2100
rect 16856 2048 16908 2100
rect 24768 2048 24820 2100
rect 2872 1980 2924 2032
rect 10876 1980 10928 2032
rect 16028 1912 16080 1964
rect 22008 1912 22060 1964
rect 10416 1844 10468 1896
rect 21272 1844 21324 1896
rect 18512 1776 18564 1828
rect 21548 1776 21600 1828
rect 5540 1708 5592 1760
rect 6092 1708 6144 1760
rect 22284 892 22336 944
rect 22468 892 22520 944
<< metal2 >>
rect 1030 56200 1086 57000
rect 2410 56200 2466 57000
rect 3790 56200 3846 57000
rect 3896 56222 4108 56250
rect 1044 53650 1072 56200
rect 2424 54126 2452 56200
rect 3804 56114 3832 56200
rect 3896 56114 3924 56222
rect 3804 56086 3924 56114
rect 3884 54188 3936 54194
rect 3884 54130 3936 54136
rect 2412 54120 2464 54126
rect 2412 54062 2464 54068
rect 2950 53884 3258 53893
rect 2950 53882 2956 53884
rect 3012 53882 3036 53884
rect 3092 53882 3116 53884
rect 3172 53882 3196 53884
rect 3252 53882 3258 53884
rect 3012 53830 3014 53882
rect 3194 53830 3196 53882
rect 2950 53828 2956 53830
rect 3012 53828 3036 53830
rect 3092 53828 3116 53830
rect 3172 53828 3196 53830
rect 3252 53828 3258 53830
rect 2950 53819 3258 53828
rect 1032 53644 1084 53650
rect 1032 53586 1084 53592
rect 3896 53242 3924 54130
rect 4080 54126 4108 56222
rect 5170 56200 5226 57000
rect 6550 56200 6606 57000
rect 6656 56222 6868 56250
rect 4068 54120 4120 54126
rect 4068 54062 4120 54068
rect 5184 53650 5212 56200
rect 6564 56114 6592 56200
rect 6656 56114 6684 56222
rect 6564 56086 6684 56114
rect 6840 54210 6868 56222
rect 7930 56200 7986 57000
rect 9310 56200 9366 57000
rect 10690 56200 10746 57000
rect 10796 56222 11008 56250
rect 7944 55214 7972 56200
rect 7852 55186 7972 55214
rect 6552 54188 6604 54194
rect 6552 54130 6604 54136
rect 6736 54188 6788 54194
rect 6840 54182 6960 54210
rect 6736 54130 6788 54136
rect 5172 53644 5224 53650
rect 5172 53586 5224 53592
rect 6564 53242 6592 54130
rect 3884 53236 3936 53242
rect 3884 53178 3936 53184
rect 6552 53236 6604 53242
rect 6552 53178 6604 53184
rect 2950 52796 3258 52805
rect 2950 52794 2956 52796
rect 3012 52794 3036 52796
rect 3092 52794 3116 52796
rect 3172 52794 3196 52796
rect 3252 52794 3258 52796
rect 3012 52742 3014 52794
rect 3194 52742 3196 52794
rect 2950 52740 2956 52742
rect 3012 52740 3036 52742
rect 3092 52740 3116 52742
rect 3172 52740 3196 52742
rect 3252 52740 3258 52742
rect 2950 52731 3258 52740
rect 6748 52154 6776 54130
rect 6932 54126 6960 54182
rect 6920 54120 6972 54126
rect 6920 54062 6972 54068
rect 7656 53576 7708 53582
rect 7656 53518 7708 53524
rect 7564 53508 7616 53514
rect 7564 53450 7616 53456
rect 7576 52578 7604 53450
rect 7668 52698 7696 53518
rect 7748 53032 7800 53038
rect 7748 52974 7800 52980
rect 7656 52692 7708 52698
rect 7656 52634 7708 52640
rect 7576 52550 7696 52578
rect 6736 52148 6788 52154
rect 6736 52090 6788 52096
rect 2950 51708 3258 51717
rect 2950 51706 2956 51708
rect 3012 51706 3036 51708
rect 3092 51706 3116 51708
rect 3172 51706 3196 51708
rect 3252 51706 3258 51708
rect 3012 51654 3014 51706
rect 3194 51654 3196 51706
rect 2950 51652 2956 51654
rect 3012 51652 3036 51654
rect 3092 51652 3116 51654
rect 3172 51652 3196 51654
rect 3252 51652 3258 51654
rect 2950 51643 3258 51652
rect 7668 51610 7696 52550
rect 7760 51610 7788 52974
rect 7852 52630 7880 55186
rect 7950 54428 8258 54437
rect 7950 54426 7956 54428
rect 8012 54426 8036 54428
rect 8092 54426 8116 54428
rect 8172 54426 8196 54428
rect 8252 54426 8258 54428
rect 8012 54374 8014 54426
rect 8194 54374 8196 54426
rect 7950 54372 7956 54374
rect 8012 54372 8036 54374
rect 8092 54372 8116 54374
rect 8172 54372 8196 54374
rect 8252 54372 8258 54374
rect 7950 54363 8258 54372
rect 8484 54120 8536 54126
rect 8484 54062 8536 54068
rect 7950 53340 8258 53349
rect 7950 53338 7956 53340
rect 8012 53338 8036 53340
rect 8092 53338 8116 53340
rect 8172 53338 8196 53340
rect 8252 53338 8258 53340
rect 8012 53286 8014 53338
rect 8194 53286 8196 53338
rect 7950 53284 7956 53286
rect 8012 53284 8036 53286
rect 8092 53284 8116 53286
rect 8172 53284 8196 53286
rect 8252 53284 8258 53286
rect 7950 53275 8258 53284
rect 7840 52624 7892 52630
rect 7840 52566 7892 52572
rect 8392 52624 8444 52630
rect 8392 52566 8444 52572
rect 7950 52252 8258 52261
rect 7950 52250 7956 52252
rect 8012 52250 8036 52252
rect 8092 52250 8116 52252
rect 8172 52250 8196 52252
rect 8252 52250 8258 52252
rect 8012 52198 8014 52250
rect 8194 52198 8196 52250
rect 7950 52196 7956 52198
rect 8012 52196 8036 52198
rect 8092 52196 8116 52198
rect 8172 52196 8196 52198
rect 8252 52196 8258 52198
rect 7950 52187 8258 52196
rect 7656 51604 7708 51610
rect 7656 51546 7708 51552
rect 7748 51604 7800 51610
rect 7748 51546 7800 51552
rect 2950 50620 3258 50629
rect 2950 50618 2956 50620
rect 3012 50618 3036 50620
rect 3092 50618 3116 50620
rect 3172 50618 3196 50620
rect 3252 50618 3258 50620
rect 3012 50566 3014 50618
rect 3194 50566 3196 50618
rect 2950 50564 2956 50566
rect 3012 50564 3036 50566
rect 3092 50564 3116 50566
rect 3172 50564 3196 50566
rect 3252 50564 3258 50566
rect 2950 50555 3258 50564
rect 2950 49532 3258 49541
rect 2950 49530 2956 49532
rect 3012 49530 3036 49532
rect 3092 49530 3116 49532
rect 3172 49530 3196 49532
rect 3252 49530 3258 49532
rect 3012 49478 3014 49530
rect 3194 49478 3196 49530
rect 2950 49476 2956 49478
rect 3012 49476 3036 49478
rect 3092 49476 3116 49478
rect 3172 49476 3196 49478
rect 3252 49476 3258 49478
rect 2950 49467 3258 49476
rect 7668 49434 7696 51546
rect 7656 49428 7708 49434
rect 7656 49370 7708 49376
rect 7760 48822 7788 51546
rect 7950 51164 8258 51173
rect 7950 51162 7956 51164
rect 8012 51162 8036 51164
rect 8092 51162 8116 51164
rect 8172 51162 8196 51164
rect 8252 51162 8258 51164
rect 8012 51110 8014 51162
rect 8194 51110 8196 51162
rect 7950 51108 7956 51110
rect 8012 51108 8036 51110
rect 8092 51108 8116 51110
rect 8172 51108 8196 51110
rect 8252 51108 8258 51110
rect 7950 51099 8258 51108
rect 7950 50076 8258 50085
rect 7950 50074 7956 50076
rect 8012 50074 8036 50076
rect 8092 50074 8116 50076
rect 8172 50074 8196 50076
rect 8252 50074 8258 50076
rect 8012 50022 8014 50074
rect 8194 50022 8196 50074
rect 7950 50020 7956 50022
rect 8012 50020 8036 50022
rect 8092 50020 8116 50022
rect 8172 50020 8196 50022
rect 8252 50020 8258 50022
rect 7950 50011 8258 50020
rect 8300 49088 8352 49094
rect 8300 49030 8352 49036
rect 7950 48988 8258 48997
rect 7950 48986 7956 48988
rect 8012 48986 8036 48988
rect 8092 48986 8116 48988
rect 8172 48986 8196 48988
rect 8252 48986 8258 48988
rect 8012 48934 8014 48986
rect 8194 48934 8196 48986
rect 7950 48932 7956 48934
rect 8012 48932 8036 48934
rect 8092 48932 8116 48934
rect 8172 48932 8196 48934
rect 8252 48932 8258 48934
rect 7950 48923 8258 48932
rect 7748 48816 7800 48822
rect 7748 48758 7800 48764
rect 7748 48680 7800 48686
rect 7748 48622 7800 48628
rect 2950 48444 3258 48453
rect 2950 48442 2956 48444
rect 3012 48442 3036 48444
rect 3092 48442 3116 48444
rect 3172 48442 3196 48444
rect 3252 48442 3258 48444
rect 3012 48390 3014 48442
rect 3194 48390 3196 48442
rect 2950 48388 2956 48390
rect 3012 48388 3036 48390
rect 3092 48388 3116 48390
rect 3172 48388 3196 48390
rect 3252 48388 3258 48390
rect 2950 48379 3258 48388
rect 2950 47356 3258 47365
rect 2950 47354 2956 47356
rect 3012 47354 3036 47356
rect 3092 47354 3116 47356
rect 3172 47354 3196 47356
rect 3252 47354 3258 47356
rect 3012 47302 3014 47354
rect 3194 47302 3196 47354
rect 2950 47300 2956 47302
rect 3012 47300 3036 47302
rect 3092 47300 3116 47302
rect 3172 47300 3196 47302
rect 3252 47300 3258 47302
rect 2950 47291 3258 47300
rect 2950 46268 3258 46277
rect 2950 46266 2956 46268
rect 3012 46266 3036 46268
rect 3092 46266 3116 46268
rect 3172 46266 3196 46268
rect 3252 46266 3258 46268
rect 3012 46214 3014 46266
rect 3194 46214 3196 46266
rect 2950 46212 2956 46214
rect 3012 46212 3036 46214
rect 3092 46212 3116 46214
rect 3172 46212 3196 46214
rect 3252 46212 3258 46214
rect 2950 46203 3258 46212
rect 2950 45180 3258 45189
rect 2950 45178 2956 45180
rect 3012 45178 3036 45180
rect 3092 45178 3116 45180
rect 3172 45178 3196 45180
rect 3252 45178 3258 45180
rect 3012 45126 3014 45178
rect 3194 45126 3196 45178
rect 2950 45124 2956 45126
rect 3012 45124 3036 45126
rect 3092 45124 3116 45126
rect 3172 45124 3196 45126
rect 3252 45124 3258 45126
rect 2950 45115 3258 45124
rect 2950 44092 3258 44101
rect 2950 44090 2956 44092
rect 3012 44090 3036 44092
rect 3092 44090 3116 44092
rect 3172 44090 3196 44092
rect 3252 44090 3258 44092
rect 3012 44038 3014 44090
rect 3194 44038 3196 44090
rect 2950 44036 2956 44038
rect 3012 44036 3036 44038
rect 3092 44036 3116 44038
rect 3172 44036 3196 44038
rect 3252 44036 3258 44038
rect 2950 44027 3258 44036
rect 2950 43004 3258 43013
rect 2950 43002 2956 43004
rect 3012 43002 3036 43004
rect 3092 43002 3116 43004
rect 3172 43002 3196 43004
rect 3252 43002 3258 43004
rect 3012 42950 3014 43002
rect 3194 42950 3196 43002
rect 2950 42948 2956 42950
rect 3012 42948 3036 42950
rect 3092 42948 3116 42950
rect 3172 42948 3196 42950
rect 3252 42948 3258 42950
rect 2950 42939 3258 42948
rect 2950 41916 3258 41925
rect 2950 41914 2956 41916
rect 3012 41914 3036 41916
rect 3092 41914 3116 41916
rect 3172 41914 3196 41916
rect 3252 41914 3258 41916
rect 3012 41862 3014 41914
rect 3194 41862 3196 41914
rect 2950 41860 2956 41862
rect 3012 41860 3036 41862
rect 3092 41860 3116 41862
rect 3172 41860 3196 41862
rect 3252 41860 3258 41862
rect 2950 41851 3258 41860
rect 2950 40828 3258 40837
rect 2950 40826 2956 40828
rect 3012 40826 3036 40828
rect 3092 40826 3116 40828
rect 3172 40826 3196 40828
rect 3252 40826 3258 40828
rect 3012 40774 3014 40826
rect 3194 40774 3196 40826
rect 2950 40772 2956 40774
rect 3012 40772 3036 40774
rect 3092 40772 3116 40774
rect 3172 40772 3196 40774
rect 3252 40772 3258 40774
rect 2950 40763 3258 40772
rect 2950 39740 3258 39749
rect 2950 39738 2956 39740
rect 3012 39738 3036 39740
rect 3092 39738 3116 39740
rect 3172 39738 3196 39740
rect 3252 39738 3258 39740
rect 3012 39686 3014 39738
rect 3194 39686 3196 39738
rect 2950 39684 2956 39686
rect 3012 39684 3036 39686
rect 3092 39684 3116 39686
rect 3172 39684 3196 39686
rect 3252 39684 3258 39686
rect 2950 39675 3258 39684
rect 7760 39642 7788 48622
rect 8312 48278 8340 49030
rect 8404 48686 8432 52566
rect 8496 51610 8524 54062
rect 8484 51604 8536 51610
rect 8484 51546 8536 51552
rect 8496 51406 8524 51546
rect 8484 51400 8536 51406
rect 8484 51342 8536 51348
rect 8496 49366 8524 51342
rect 9128 49428 9180 49434
rect 9128 49370 9180 49376
rect 8484 49360 8536 49366
rect 8484 49302 8536 49308
rect 8760 49292 8812 49298
rect 8760 49234 8812 49240
rect 8772 49094 8800 49234
rect 8760 49088 8812 49094
rect 8760 49030 8812 49036
rect 8392 48680 8444 48686
rect 8392 48622 8444 48628
rect 8300 48272 8352 48278
rect 8300 48214 8352 48220
rect 7950 47900 8258 47909
rect 7950 47898 7956 47900
rect 8012 47898 8036 47900
rect 8092 47898 8116 47900
rect 8172 47898 8196 47900
rect 8252 47898 8258 47900
rect 8012 47846 8014 47898
rect 8194 47846 8196 47898
rect 7950 47844 7956 47846
rect 8012 47844 8036 47846
rect 8092 47844 8116 47846
rect 8172 47844 8196 47846
rect 8252 47844 8258 47846
rect 7950 47835 8258 47844
rect 7950 46812 8258 46821
rect 7950 46810 7956 46812
rect 8012 46810 8036 46812
rect 8092 46810 8116 46812
rect 8172 46810 8196 46812
rect 8252 46810 8258 46812
rect 8012 46758 8014 46810
rect 8194 46758 8196 46810
rect 7950 46756 7956 46758
rect 8012 46756 8036 46758
rect 8092 46756 8116 46758
rect 8172 46756 8196 46758
rect 8252 46756 8258 46758
rect 7950 46747 8258 46756
rect 8772 46510 8800 49030
rect 9140 48142 9168 49370
rect 9128 48136 9180 48142
rect 9128 48078 9180 48084
rect 9036 47524 9088 47530
rect 9036 47466 9088 47472
rect 8760 46504 8812 46510
rect 8760 46446 8812 46452
rect 7950 45724 8258 45733
rect 7950 45722 7956 45724
rect 8012 45722 8036 45724
rect 8092 45722 8116 45724
rect 8172 45722 8196 45724
rect 8252 45722 8258 45724
rect 8012 45670 8014 45722
rect 8194 45670 8196 45722
rect 7950 45668 7956 45670
rect 8012 45668 8036 45670
rect 8092 45668 8116 45670
rect 8172 45668 8196 45670
rect 8252 45668 8258 45670
rect 7950 45659 8258 45668
rect 8944 45416 8996 45422
rect 8944 45358 8996 45364
rect 7950 44636 8258 44645
rect 7950 44634 7956 44636
rect 8012 44634 8036 44636
rect 8092 44634 8116 44636
rect 8172 44634 8196 44636
rect 8252 44634 8258 44636
rect 8012 44582 8014 44634
rect 8194 44582 8196 44634
rect 7950 44580 7956 44582
rect 8012 44580 8036 44582
rect 8092 44580 8116 44582
rect 8172 44580 8196 44582
rect 8252 44580 8258 44582
rect 7950 44571 8258 44580
rect 7950 43548 8258 43557
rect 7950 43546 7956 43548
rect 8012 43546 8036 43548
rect 8092 43546 8116 43548
rect 8172 43546 8196 43548
rect 8252 43546 8258 43548
rect 8012 43494 8014 43546
rect 8194 43494 8196 43546
rect 7950 43492 7956 43494
rect 8012 43492 8036 43494
rect 8092 43492 8116 43494
rect 8172 43492 8196 43494
rect 8252 43492 8258 43494
rect 7950 43483 8258 43492
rect 7950 42460 8258 42469
rect 7950 42458 7956 42460
rect 8012 42458 8036 42460
rect 8092 42458 8116 42460
rect 8172 42458 8196 42460
rect 8252 42458 8258 42460
rect 8012 42406 8014 42458
rect 8194 42406 8196 42458
rect 7950 42404 7956 42406
rect 8012 42404 8036 42406
rect 8092 42404 8116 42406
rect 8172 42404 8196 42406
rect 8252 42404 8258 42406
rect 7950 42395 8258 42404
rect 7950 41372 8258 41381
rect 7950 41370 7956 41372
rect 8012 41370 8036 41372
rect 8092 41370 8116 41372
rect 8172 41370 8196 41372
rect 8252 41370 8258 41372
rect 8012 41318 8014 41370
rect 8194 41318 8196 41370
rect 7950 41316 7956 41318
rect 8012 41316 8036 41318
rect 8092 41316 8116 41318
rect 8172 41316 8196 41318
rect 8252 41316 8258 41318
rect 7950 41307 8258 41316
rect 7950 40284 8258 40293
rect 7950 40282 7956 40284
rect 8012 40282 8036 40284
rect 8092 40282 8116 40284
rect 8172 40282 8196 40284
rect 8252 40282 8258 40284
rect 8012 40230 8014 40282
rect 8194 40230 8196 40282
rect 7950 40228 7956 40230
rect 8012 40228 8036 40230
rect 8092 40228 8116 40230
rect 8172 40228 8196 40230
rect 8252 40228 8258 40230
rect 7950 40219 8258 40228
rect 7748 39636 7800 39642
rect 7748 39578 7800 39584
rect 7950 39196 8258 39205
rect 7950 39194 7956 39196
rect 8012 39194 8036 39196
rect 8092 39194 8116 39196
rect 8172 39194 8196 39196
rect 8252 39194 8258 39196
rect 8012 39142 8014 39194
rect 8194 39142 8196 39194
rect 7950 39140 7956 39142
rect 8012 39140 8036 39142
rect 8092 39140 8116 39142
rect 8172 39140 8196 39142
rect 8252 39140 8258 39142
rect 7950 39131 8258 39140
rect 2950 38652 3258 38661
rect 2950 38650 2956 38652
rect 3012 38650 3036 38652
rect 3092 38650 3116 38652
rect 3172 38650 3196 38652
rect 3252 38650 3258 38652
rect 3012 38598 3014 38650
rect 3194 38598 3196 38650
rect 2950 38596 2956 38598
rect 3012 38596 3036 38598
rect 3092 38596 3116 38598
rect 3172 38596 3196 38598
rect 3252 38596 3258 38598
rect 2950 38587 3258 38596
rect 7950 38108 8258 38117
rect 7950 38106 7956 38108
rect 8012 38106 8036 38108
rect 8092 38106 8116 38108
rect 8172 38106 8196 38108
rect 8252 38106 8258 38108
rect 8012 38054 8014 38106
rect 8194 38054 8196 38106
rect 7950 38052 7956 38054
rect 8012 38052 8036 38054
rect 8092 38052 8116 38054
rect 8172 38052 8196 38054
rect 8252 38052 8258 38054
rect 7950 38043 8258 38052
rect 2950 37564 3258 37573
rect 2950 37562 2956 37564
rect 3012 37562 3036 37564
rect 3092 37562 3116 37564
rect 3172 37562 3196 37564
rect 3252 37562 3258 37564
rect 3012 37510 3014 37562
rect 3194 37510 3196 37562
rect 2950 37508 2956 37510
rect 3012 37508 3036 37510
rect 3092 37508 3116 37510
rect 3172 37508 3196 37510
rect 3252 37508 3258 37510
rect 2950 37499 3258 37508
rect 7950 37020 8258 37029
rect 7950 37018 7956 37020
rect 8012 37018 8036 37020
rect 8092 37018 8116 37020
rect 8172 37018 8196 37020
rect 8252 37018 8258 37020
rect 8012 36966 8014 37018
rect 8194 36966 8196 37018
rect 7950 36964 7956 36966
rect 8012 36964 8036 36966
rect 8092 36964 8116 36966
rect 8172 36964 8196 36966
rect 8252 36964 8258 36966
rect 7950 36955 8258 36964
rect 2950 36476 3258 36485
rect 2950 36474 2956 36476
rect 3012 36474 3036 36476
rect 3092 36474 3116 36476
rect 3172 36474 3196 36476
rect 3252 36474 3258 36476
rect 3012 36422 3014 36474
rect 3194 36422 3196 36474
rect 2950 36420 2956 36422
rect 3012 36420 3036 36422
rect 3092 36420 3116 36422
rect 3172 36420 3196 36422
rect 3252 36420 3258 36422
rect 2950 36411 3258 36420
rect 7950 35932 8258 35941
rect 7950 35930 7956 35932
rect 8012 35930 8036 35932
rect 8092 35930 8116 35932
rect 8172 35930 8196 35932
rect 8252 35930 8258 35932
rect 8012 35878 8014 35930
rect 8194 35878 8196 35930
rect 7950 35876 7956 35878
rect 8012 35876 8036 35878
rect 8092 35876 8116 35878
rect 8172 35876 8196 35878
rect 8252 35876 8258 35878
rect 7950 35867 8258 35876
rect 2950 35388 3258 35397
rect 2950 35386 2956 35388
rect 3012 35386 3036 35388
rect 3092 35386 3116 35388
rect 3172 35386 3196 35388
rect 3252 35386 3258 35388
rect 3012 35334 3014 35386
rect 3194 35334 3196 35386
rect 2950 35332 2956 35334
rect 3012 35332 3036 35334
rect 3092 35332 3116 35334
rect 3172 35332 3196 35334
rect 3252 35332 3258 35334
rect 2950 35323 3258 35332
rect 7950 34844 8258 34853
rect 7950 34842 7956 34844
rect 8012 34842 8036 34844
rect 8092 34842 8116 34844
rect 8172 34842 8196 34844
rect 8252 34842 8258 34844
rect 8012 34790 8014 34842
rect 8194 34790 8196 34842
rect 7950 34788 7956 34790
rect 8012 34788 8036 34790
rect 8092 34788 8116 34790
rect 8172 34788 8196 34790
rect 8252 34788 8258 34790
rect 7950 34779 8258 34788
rect 2950 34300 3258 34309
rect 2950 34298 2956 34300
rect 3012 34298 3036 34300
rect 3092 34298 3116 34300
rect 3172 34298 3196 34300
rect 3252 34298 3258 34300
rect 3012 34246 3014 34298
rect 3194 34246 3196 34298
rect 2950 34244 2956 34246
rect 3012 34244 3036 34246
rect 3092 34244 3116 34246
rect 3172 34244 3196 34246
rect 3252 34244 3258 34246
rect 2950 34235 3258 34244
rect 7950 33756 8258 33765
rect 7950 33754 7956 33756
rect 8012 33754 8036 33756
rect 8092 33754 8116 33756
rect 8172 33754 8196 33756
rect 8252 33754 8258 33756
rect 8012 33702 8014 33754
rect 8194 33702 8196 33754
rect 7950 33700 7956 33702
rect 8012 33700 8036 33702
rect 8092 33700 8116 33702
rect 8172 33700 8196 33702
rect 8252 33700 8258 33702
rect 7950 33691 8258 33700
rect 2950 33212 3258 33221
rect 2950 33210 2956 33212
rect 3012 33210 3036 33212
rect 3092 33210 3116 33212
rect 3172 33210 3196 33212
rect 3252 33210 3258 33212
rect 3012 33158 3014 33210
rect 3194 33158 3196 33210
rect 2950 33156 2956 33158
rect 3012 33156 3036 33158
rect 3092 33156 3116 33158
rect 3172 33156 3196 33158
rect 3252 33156 3258 33158
rect 2950 33147 3258 33156
rect 7950 32668 8258 32677
rect 7950 32666 7956 32668
rect 8012 32666 8036 32668
rect 8092 32666 8116 32668
rect 8172 32666 8196 32668
rect 8252 32666 8258 32668
rect 8012 32614 8014 32666
rect 8194 32614 8196 32666
rect 7950 32612 7956 32614
rect 8012 32612 8036 32614
rect 8092 32612 8116 32614
rect 8172 32612 8196 32614
rect 8252 32612 8258 32614
rect 7950 32603 8258 32612
rect 8956 32570 8984 45358
rect 9048 36378 9076 47466
rect 9140 46714 9168 48078
rect 9324 47598 9352 56200
rect 10704 56114 10732 56200
rect 10796 56114 10824 56222
rect 10704 56086 10824 56114
rect 10980 55214 11008 56222
rect 12070 56200 12126 57000
rect 13450 56200 13506 57000
rect 14830 56200 14886 57000
rect 16210 56200 16266 57000
rect 16316 56222 16528 56250
rect 10888 55186 11008 55214
rect 9588 53100 9640 53106
rect 9588 53042 9640 53048
rect 9496 52488 9548 52494
rect 9496 52430 9548 52436
rect 9312 47592 9364 47598
rect 9312 47534 9364 47540
rect 9508 47190 9536 52430
rect 9600 49434 9628 53042
rect 10324 52012 10376 52018
rect 10324 51954 10376 51960
rect 9588 49428 9640 49434
rect 9588 49370 9640 49376
rect 9600 48346 9628 49370
rect 9680 49156 9732 49162
rect 9680 49098 9732 49104
rect 9588 48340 9640 48346
rect 9588 48282 9640 48288
rect 9600 47734 9628 48282
rect 9588 47728 9640 47734
rect 9588 47670 9640 47676
rect 9496 47184 9548 47190
rect 9496 47126 9548 47132
rect 9128 46708 9180 46714
rect 9128 46650 9180 46656
rect 9220 46368 9272 46374
rect 9220 46310 9272 46316
rect 9232 43246 9260 46310
rect 9508 45558 9536 47126
rect 9692 46646 9720 49098
rect 9680 46640 9732 46646
rect 9680 46582 9732 46588
rect 9692 46374 9720 46582
rect 9680 46368 9732 46374
rect 9680 46310 9732 46316
rect 10336 46034 10364 51954
rect 10692 47252 10744 47258
rect 10692 47194 10744 47200
rect 10600 46504 10652 46510
rect 10600 46446 10652 46452
rect 10324 46028 10376 46034
rect 10324 45970 10376 45976
rect 10416 45960 10468 45966
rect 10416 45902 10468 45908
rect 9496 45552 9548 45558
rect 9496 45494 9548 45500
rect 9956 44872 10008 44878
rect 9956 44814 10008 44820
rect 9968 43450 9996 44814
rect 9956 43444 10008 43450
rect 9956 43386 10008 43392
rect 9220 43240 9272 43246
rect 9220 43182 9272 43188
rect 9772 39432 9824 39438
rect 9772 39374 9824 39380
rect 9680 36712 9732 36718
rect 9680 36654 9732 36660
rect 9036 36372 9088 36378
rect 9036 36314 9088 36320
rect 9220 36168 9272 36174
rect 9220 36110 9272 36116
rect 8944 32564 8996 32570
rect 8944 32506 8996 32512
rect 8668 32428 8720 32434
rect 8668 32370 8720 32376
rect 2950 32124 3258 32133
rect 2950 32122 2956 32124
rect 3012 32122 3036 32124
rect 3092 32122 3116 32124
rect 3172 32122 3196 32124
rect 3252 32122 3258 32124
rect 3012 32070 3014 32122
rect 3194 32070 3196 32122
rect 2950 32068 2956 32070
rect 3012 32068 3036 32070
rect 3092 32068 3116 32070
rect 3172 32068 3196 32070
rect 3252 32068 3258 32070
rect 2950 32059 3258 32068
rect 7950 31580 8258 31589
rect 7950 31578 7956 31580
rect 8012 31578 8036 31580
rect 8092 31578 8116 31580
rect 8172 31578 8196 31580
rect 8252 31578 8258 31580
rect 8012 31526 8014 31578
rect 8194 31526 8196 31578
rect 7950 31524 7956 31526
rect 8012 31524 8036 31526
rect 8092 31524 8116 31526
rect 8172 31524 8196 31526
rect 8252 31524 8258 31526
rect 7950 31515 8258 31524
rect 2950 31036 3258 31045
rect 2950 31034 2956 31036
rect 3012 31034 3036 31036
rect 3092 31034 3116 31036
rect 3172 31034 3196 31036
rect 3252 31034 3258 31036
rect 3012 30982 3014 31034
rect 3194 30982 3196 31034
rect 2950 30980 2956 30982
rect 3012 30980 3036 30982
rect 3092 30980 3116 30982
rect 3172 30980 3196 30982
rect 3252 30980 3258 30982
rect 2950 30971 3258 30980
rect 7950 30492 8258 30501
rect 7950 30490 7956 30492
rect 8012 30490 8036 30492
rect 8092 30490 8116 30492
rect 8172 30490 8196 30492
rect 8252 30490 8258 30492
rect 8012 30438 8014 30490
rect 8194 30438 8196 30490
rect 7950 30436 7956 30438
rect 8012 30436 8036 30438
rect 8092 30436 8116 30438
rect 8172 30436 8196 30438
rect 8252 30436 8258 30438
rect 7950 30427 8258 30436
rect 2950 29948 3258 29957
rect 2950 29946 2956 29948
rect 3012 29946 3036 29948
rect 3092 29946 3116 29948
rect 3172 29946 3196 29948
rect 3252 29946 3258 29948
rect 3012 29894 3014 29946
rect 3194 29894 3196 29946
rect 2950 29892 2956 29894
rect 3012 29892 3036 29894
rect 3092 29892 3116 29894
rect 3172 29892 3196 29894
rect 3252 29892 3258 29894
rect 2950 29883 3258 29892
rect 7950 29404 8258 29413
rect 7950 29402 7956 29404
rect 8012 29402 8036 29404
rect 8092 29402 8116 29404
rect 8172 29402 8196 29404
rect 8252 29402 8258 29404
rect 8012 29350 8014 29402
rect 8194 29350 8196 29402
rect 7950 29348 7956 29350
rect 8012 29348 8036 29350
rect 8092 29348 8116 29350
rect 8172 29348 8196 29350
rect 8252 29348 8258 29350
rect 7950 29339 8258 29348
rect 2950 28860 3258 28869
rect 2950 28858 2956 28860
rect 3012 28858 3036 28860
rect 3092 28858 3116 28860
rect 3172 28858 3196 28860
rect 3252 28858 3258 28860
rect 3012 28806 3014 28858
rect 3194 28806 3196 28858
rect 2950 28804 2956 28806
rect 3012 28804 3036 28806
rect 3092 28804 3116 28806
rect 3172 28804 3196 28806
rect 3252 28804 3258 28806
rect 2950 28795 3258 28804
rect 7950 28316 8258 28325
rect 7950 28314 7956 28316
rect 8012 28314 8036 28316
rect 8092 28314 8116 28316
rect 8172 28314 8196 28316
rect 8252 28314 8258 28316
rect 8012 28262 8014 28314
rect 8194 28262 8196 28314
rect 7950 28260 7956 28262
rect 8012 28260 8036 28262
rect 8092 28260 8116 28262
rect 8172 28260 8196 28262
rect 8252 28260 8258 28262
rect 7950 28251 8258 28260
rect 2950 27772 3258 27781
rect 2950 27770 2956 27772
rect 3012 27770 3036 27772
rect 3092 27770 3116 27772
rect 3172 27770 3196 27772
rect 3252 27770 3258 27772
rect 3012 27718 3014 27770
rect 3194 27718 3196 27770
rect 2950 27716 2956 27718
rect 3012 27716 3036 27718
rect 3092 27716 3116 27718
rect 3172 27716 3196 27718
rect 3252 27716 3258 27718
rect 2950 27707 3258 27716
rect 7950 27228 8258 27237
rect 7950 27226 7956 27228
rect 8012 27226 8036 27228
rect 8092 27226 8116 27228
rect 8172 27226 8196 27228
rect 8252 27226 8258 27228
rect 8012 27174 8014 27226
rect 8194 27174 8196 27226
rect 7950 27172 7956 27174
rect 8012 27172 8036 27174
rect 8092 27172 8116 27174
rect 8172 27172 8196 27174
rect 8252 27172 8258 27174
rect 7950 27163 8258 27172
rect 2950 26684 3258 26693
rect 2950 26682 2956 26684
rect 3012 26682 3036 26684
rect 3092 26682 3116 26684
rect 3172 26682 3196 26684
rect 3252 26682 3258 26684
rect 3012 26630 3014 26682
rect 3194 26630 3196 26682
rect 2950 26628 2956 26630
rect 3012 26628 3036 26630
rect 3092 26628 3116 26630
rect 3172 26628 3196 26630
rect 3252 26628 3258 26630
rect 2950 26619 3258 26628
rect 7950 26140 8258 26149
rect 7950 26138 7956 26140
rect 8012 26138 8036 26140
rect 8092 26138 8116 26140
rect 8172 26138 8196 26140
rect 8252 26138 8258 26140
rect 8012 26086 8014 26138
rect 8194 26086 8196 26138
rect 7950 26084 7956 26086
rect 8012 26084 8036 26086
rect 8092 26084 8116 26086
rect 8172 26084 8196 26086
rect 8252 26084 8258 26086
rect 7950 26075 8258 26084
rect 2950 25596 3258 25605
rect 2950 25594 2956 25596
rect 3012 25594 3036 25596
rect 3092 25594 3116 25596
rect 3172 25594 3196 25596
rect 3252 25594 3258 25596
rect 3012 25542 3014 25594
rect 3194 25542 3196 25594
rect 2950 25540 2956 25542
rect 3012 25540 3036 25542
rect 3092 25540 3116 25542
rect 3172 25540 3196 25542
rect 3252 25540 3258 25542
rect 2950 25531 3258 25540
rect 7950 25052 8258 25061
rect 7950 25050 7956 25052
rect 8012 25050 8036 25052
rect 8092 25050 8116 25052
rect 8172 25050 8196 25052
rect 8252 25050 8258 25052
rect 8012 24998 8014 25050
rect 8194 24998 8196 25050
rect 7950 24996 7956 24998
rect 8012 24996 8036 24998
rect 8092 24996 8116 24998
rect 8172 24996 8196 24998
rect 8252 24996 8258 24998
rect 7950 24987 8258 24996
rect 8576 24744 8628 24750
rect 8576 24686 8628 24692
rect 8392 24676 8444 24682
rect 8392 24618 8444 24624
rect 2950 24508 3258 24517
rect 2950 24506 2956 24508
rect 3012 24506 3036 24508
rect 3092 24506 3116 24508
rect 3172 24506 3196 24508
rect 3252 24506 3258 24508
rect 3012 24454 3014 24506
rect 3194 24454 3196 24506
rect 2950 24452 2956 24454
rect 3012 24452 3036 24454
rect 3092 24452 3116 24454
rect 3172 24452 3196 24454
rect 3252 24452 3258 24454
rect 2950 24443 3258 24452
rect 7748 24268 7800 24274
rect 7748 24210 7800 24216
rect 7760 23730 7788 24210
rect 7950 23964 8258 23973
rect 7950 23962 7956 23964
rect 8012 23962 8036 23964
rect 8092 23962 8116 23964
rect 8172 23962 8196 23964
rect 8252 23962 8258 23964
rect 8012 23910 8014 23962
rect 8194 23910 8196 23962
rect 7950 23908 7956 23910
rect 8012 23908 8036 23910
rect 8092 23908 8116 23910
rect 8172 23908 8196 23910
rect 8252 23908 8258 23910
rect 7950 23899 8258 23908
rect 7748 23724 7800 23730
rect 7748 23666 7800 23672
rect 2950 23420 3258 23429
rect 2950 23418 2956 23420
rect 3012 23418 3036 23420
rect 3092 23418 3116 23420
rect 3172 23418 3196 23420
rect 3252 23418 3258 23420
rect 3012 23366 3014 23418
rect 3194 23366 3196 23418
rect 2950 23364 2956 23366
rect 3012 23364 3036 23366
rect 3092 23364 3116 23366
rect 3172 23364 3196 23366
rect 3252 23364 3258 23366
rect 2950 23355 3258 23364
rect 7760 22642 7788 23666
rect 7950 22876 8258 22885
rect 7950 22874 7956 22876
rect 8012 22874 8036 22876
rect 8092 22874 8116 22876
rect 8172 22874 8196 22876
rect 8252 22874 8258 22876
rect 8012 22822 8014 22874
rect 8194 22822 8196 22874
rect 7950 22820 7956 22822
rect 8012 22820 8036 22822
rect 8092 22820 8116 22822
rect 8172 22820 8196 22822
rect 8252 22820 8258 22822
rect 7950 22811 8258 22820
rect 7748 22636 7800 22642
rect 7748 22578 7800 22584
rect 7288 22432 7340 22438
rect 7288 22374 7340 22380
rect 2950 22332 3258 22341
rect 2950 22330 2956 22332
rect 3012 22330 3036 22332
rect 3092 22330 3116 22332
rect 3172 22330 3196 22332
rect 3252 22330 3258 22332
rect 3012 22278 3014 22330
rect 3194 22278 3196 22330
rect 2950 22276 2956 22278
rect 3012 22276 3036 22278
rect 3092 22276 3116 22278
rect 3172 22276 3196 22278
rect 3252 22276 3258 22278
rect 2950 22267 3258 22276
rect 6276 21888 6328 21894
rect 6276 21830 6328 21836
rect 2950 21244 3258 21253
rect 2950 21242 2956 21244
rect 3012 21242 3036 21244
rect 3092 21242 3116 21244
rect 3172 21242 3196 21244
rect 3252 21242 3258 21244
rect 3012 21190 3014 21242
rect 3194 21190 3196 21242
rect 2950 21188 2956 21190
rect 3012 21188 3036 21190
rect 3092 21188 3116 21190
rect 3172 21188 3196 21190
rect 3252 21188 3258 21190
rect 2950 21179 3258 21188
rect 5264 21072 5316 21078
rect 5264 21014 5316 21020
rect 2950 20156 3258 20165
rect 2950 20154 2956 20156
rect 3012 20154 3036 20156
rect 3092 20154 3116 20156
rect 3172 20154 3196 20156
rect 3252 20154 3258 20156
rect 3012 20102 3014 20154
rect 3194 20102 3196 20154
rect 2950 20100 2956 20102
rect 3012 20100 3036 20102
rect 3092 20100 3116 20102
rect 3172 20100 3196 20102
rect 3252 20100 3258 20102
rect 2950 20091 3258 20100
rect 3516 19168 3568 19174
rect 3516 19110 3568 19116
rect 2950 19068 3258 19077
rect 2950 19066 2956 19068
rect 3012 19066 3036 19068
rect 3092 19066 3116 19068
rect 3172 19066 3196 19068
rect 3252 19066 3258 19068
rect 3012 19014 3014 19066
rect 3194 19014 3196 19066
rect 2950 19012 2956 19014
rect 3012 19012 3036 19014
rect 3092 19012 3116 19014
rect 3172 19012 3196 19014
rect 3252 19012 3258 19014
rect 2950 19003 3258 19012
rect 2950 17980 3258 17989
rect 2950 17978 2956 17980
rect 3012 17978 3036 17980
rect 3092 17978 3116 17980
rect 3172 17978 3196 17980
rect 3252 17978 3258 17980
rect 3012 17926 3014 17978
rect 3194 17926 3196 17978
rect 2950 17924 2956 17926
rect 3012 17924 3036 17926
rect 3092 17924 3116 17926
rect 3172 17924 3196 17926
rect 3252 17924 3258 17926
rect 2950 17915 3258 17924
rect 2950 16892 3258 16901
rect 2950 16890 2956 16892
rect 3012 16890 3036 16892
rect 3092 16890 3116 16892
rect 3172 16890 3196 16892
rect 3252 16890 3258 16892
rect 3012 16838 3014 16890
rect 3194 16838 3196 16890
rect 2950 16836 2956 16838
rect 3012 16836 3036 16838
rect 3092 16836 3116 16838
rect 3172 16836 3196 16838
rect 3252 16836 3258 16838
rect 2950 16827 3258 16836
rect 2950 15804 3258 15813
rect 2950 15802 2956 15804
rect 3012 15802 3036 15804
rect 3092 15802 3116 15804
rect 3172 15802 3196 15804
rect 3252 15802 3258 15804
rect 3012 15750 3014 15802
rect 3194 15750 3196 15802
rect 2950 15748 2956 15750
rect 3012 15748 3036 15750
rect 3092 15748 3116 15750
rect 3172 15748 3196 15750
rect 3252 15748 3258 15750
rect 2950 15739 3258 15748
rect 3424 15020 3476 15026
rect 3424 14962 3476 14968
rect 2950 14716 3258 14725
rect 2950 14714 2956 14716
rect 3012 14714 3036 14716
rect 3092 14714 3116 14716
rect 3172 14714 3196 14716
rect 3252 14714 3258 14716
rect 3012 14662 3014 14714
rect 3194 14662 3196 14714
rect 2950 14660 2956 14662
rect 3012 14660 3036 14662
rect 3092 14660 3116 14662
rect 3172 14660 3196 14662
rect 3252 14660 3258 14662
rect 2950 14651 3258 14660
rect 2950 13628 3258 13637
rect 2950 13626 2956 13628
rect 3012 13626 3036 13628
rect 3092 13626 3116 13628
rect 3172 13626 3196 13628
rect 3252 13626 3258 13628
rect 3012 13574 3014 13626
rect 3194 13574 3196 13626
rect 2950 13572 2956 13574
rect 3012 13572 3036 13574
rect 3092 13572 3116 13574
rect 3172 13572 3196 13574
rect 3252 13572 3258 13574
rect 2950 13563 3258 13572
rect 2950 12540 3258 12549
rect 2950 12538 2956 12540
rect 3012 12538 3036 12540
rect 3092 12538 3116 12540
rect 3172 12538 3196 12540
rect 3252 12538 3258 12540
rect 3012 12486 3014 12538
rect 3194 12486 3196 12538
rect 2950 12484 2956 12486
rect 3012 12484 3036 12486
rect 3092 12484 3116 12486
rect 3172 12484 3196 12486
rect 3252 12484 3258 12486
rect 2950 12475 3258 12484
rect 2950 11452 3258 11461
rect 2950 11450 2956 11452
rect 3012 11450 3036 11452
rect 3092 11450 3116 11452
rect 3172 11450 3196 11452
rect 3252 11450 3258 11452
rect 3012 11398 3014 11450
rect 3194 11398 3196 11450
rect 2950 11396 2956 11398
rect 3012 11396 3036 11398
rect 3092 11396 3116 11398
rect 3172 11396 3196 11398
rect 3252 11396 3258 11398
rect 2950 11387 3258 11396
rect 2950 10364 3258 10373
rect 2950 10362 2956 10364
rect 3012 10362 3036 10364
rect 3092 10362 3116 10364
rect 3172 10362 3196 10364
rect 3252 10362 3258 10364
rect 3012 10310 3014 10362
rect 3194 10310 3196 10362
rect 2950 10308 2956 10310
rect 3012 10308 3036 10310
rect 3092 10308 3116 10310
rect 3172 10308 3196 10310
rect 3252 10308 3258 10310
rect 2950 10299 3258 10308
rect 3332 9648 3384 9654
rect 3332 9590 3384 9596
rect 2950 9276 3258 9285
rect 2950 9274 2956 9276
rect 3012 9274 3036 9276
rect 3092 9274 3116 9276
rect 3172 9274 3196 9276
rect 3252 9274 3258 9276
rect 3012 9222 3014 9274
rect 3194 9222 3196 9274
rect 2950 9220 2956 9222
rect 3012 9220 3036 9222
rect 3092 9220 3116 9222
rect 3172 9220 3196 9222
rect 3252 9220 3258 9222
rect 2950 9211 3258 9220
rect 3344 8809 3372 9590
rect 3330 8800 3386 8809
rect 3330 8735 3386 8744
rect 2950 8188 3258 8197
rect 2950 8186 2956 8188
rect 3012 8186 3036 8188
rect 3092 8186 3116 8188
rect 3172 8186 3196 8188
rect 3252 8186 3258 8188
rect 3012 8134 3014 8186
rect 3194 8134 3196 8186
rect 2950 8132 2956 8134
rect 3012 8132 3036 8134
rect 3092 8132 3116 8134
rect 3172 8132 3196 8134
rect 3252 8132 3258 8134
rect 2950 8123 3258 8132
rect 2950 7100 3258 7109
rect 2950 7098 2956 7100
rect 3012 7098 3036 7100
rect 3092 7098 3116 7100
rect 3172 7098 3196 7100
rect 3252 7098 3258 7100
rect 3012 7046 3014 7098
rect 3194 7046 3196 7098
rect 2950 7044 2956 7046
rect 3012 7044 3036 7046
rect 3092 7044 3116 7046
rect 3172 7044 3196 7046
rect 3252 7044 3258 7046
rect 2950 7035 3258 7044
rect 2044 6656 2096 6662
rect 2044 6598 2096 6604
rect 1492 4480 1544 4486
rect 1492 4422 1544 4428
rect 1504 4146 1532 4422
rect 1492 4140 1544 4146
rect 1492 4082 1544 4088
rect 1860 4140 1912 4146
rect 1860 4082 1912 4088
rect 1504 800 1532 4082
rect 1872 800 1900 4082
rect 2056 3602 2084 6598
rect 2228 6180 2280 6186
rect 2228 6122 2280 6128
rect 2240 3942 2268 6122
rect 2950 6012 3258 6021
rect 2950 6010 2956 6012
rect 3012 6010 3036 6012
rect 3092 6010 3116 6012
rect 3172 6010 3196 6012
rect 3252 6010 3258 6012
rect 3012 5958 3014 6010
rect 3194 5958 3196 6010
rect 2950 5956 2956 5958
rect 3012 5956 3036 5958
rect 3092 5956 3116 5958
rect 3172 5956 3196 5958
rect 3252 5956 3258 5958
rect 2950 5947 3258 5956
rect 2950 4924 3258 4933
rect 2950 4922 2956 4924
rect 3012 4922 3036 4924
rect 3092 4922 3116 4924
rect 3172 4922 3196 4924
rect 3252 4922 3258 4924
rect 3012 4870 3014 4922
rect 3194 4870 3196 4922
rect 2950 4868 2956 4870
rect 3012 4868 3036 4870
rect 3092 4868 3116 4870
rect 3172 4868 3196 4870
rect 3252 4868 3258 4870
rect 2950 4859 3258 4868
rect 2228 3936 2280 3942
rect 2228 3878 2280 3884
rect 2872 3936 2924 3942
rect 2872 3878 2924 3884
rect 2884 3602 2912 3878
rect 2950 3836 3258 3845
rect 2950 3834 2956 3836
rect 3012 3834 3036 3836
rect 3092 3834 3116 3836
rect 3172 3834 3196 3836
rect 3252 3834 3258 3836
rect 3012 3782 3014 3834
rect 3194 3782 3196 3834
rect 2950 3780 2956 3782
rect 3012 3780 3036 3782
rect 3092 3780 3116 3782
rect 3172 3780 3196 3782
rect 3252 3780 3258 3782
rect 2950 3771 3258 3780
rect 2044 3596 2096 3602
rect 2044 3538 2096 3544
rect 2872 3596 2924 3602
rect 2872 3538 2924 3544
rect 2228 3528 2280 3534
rect 2228 3470 2280 3476
rect 2240 800 2268 3470
rect 3332 3392 3384 3398
rect 3332 3334 3384 3340
rect 3344 3058 3372 3334
rect 2596 3052 2648 3058
rect 2596 2994 2648 3000
rect 3332 3052 3384 3058
rect 3332 2994 3384 3000
rect 2608 2310 2636 2994
rect 2950 2748 3258 2757
rect 2950 2746 2956 2748
rect 3012 2746 3036 2748
rect 3092 2746 3116 2748
rect 3172 2746 3196 2748
rect 3252 2746 3258 2748
rect 3012 2694 3014 2746
rect 3194 2694 3196 2746
rect 2950 2692 2956 2694
rect 3012 2692 3036 2694
rect 3092 2692 3116 2694
rect 3172 2692 3196 2694
rect 3252 2692 3258 2694
rect 2950 2683 3258 2692
rect 2872 2440 2924 2446
rect 2872 2382 2924 2388
rect 2596 2304 2648 2310
rect 2596 2246 2648 2252
rect 2608 800 2636 2246
rect 2884 2038 2912 2382
rect 2964 2372 3016 2378
rect 2964 2314 3016 2320
rect 2872 2032 2924 2038
rect 2872 1974 2924 1980
rect 2976 800 3004 2314
rect 3344 800 3372 2994
rect 3436 1873 3464 14962
rect 3528 6497 3556 19110
rect 5172 18080 5224 18086
rect 5172 18022 5224 18028
rect 3792 17536 3844 17542
rect 3792 17478 3844 17484
rect 3514 6488 3570 6497
rect 3514 6423 3570 6432
rect 3804 3738 3832 17478
rect 5080 12164 5132 12170
rect 5080 12106 5132 12112
rect 3976 9716 4028 9722
rect 3976 9658 4028 9664
rect 3988 4185 4016 9658
rect 3974 4176 4030 4185
rect 3974 4111 4030 4120
rect 4068 4140 4120 4146
rect 4068 4082 4120 4088
rect 3792 3732 3844 3738
rect 3792 3674 3844 3680
rect 3700 3596 3752 3602
rect 3700 3538 3752 3544
rect 3422 1864 3478 1873
rect 3422 1799 3478 1808
rect 3712 800 3740 3538
rect 4080 800 4108 4082
rect 4436 3528 4488 3534
rect 4436 3470 4488 3476
rect 4896 3528 4948 3534
rect 4896 3470 4948 3476
rect 4448 3194 4476 3470
rect 4908 3194 4936 3470
rect 4436 3188 4488 3194
rect 4436 3130 4488 3136
rect 4896 3188 4948 3194
rect 4896 3130 4948 3136
rect 4448 800 4476 3130
rect 4908 2774 4936 3130
rect 5092 3058 5120 12106
rect 5184 3602 5212 18022
rect 5276 15026 5304 21014
rect 6184 16516 6236 16522
rect 6184 16458 6236 16464
rect 5448 16244 5500 16250
rect 5448 16186 5500 16192
rect 5264 15020 5316 15026
rect 5264 14962 5316 14968
rect 5264 6860 5316 6866
rect 5264 6802 5316 6808
rect 5172 3596 5224 3602
rect 5172 3538 5224 3544
rect 5080 3052 5132 3058
rect 5080 2994 5132 3000
rect 5172 2984 5224 2990
rect 5172 2926 5224 2932
rect 4816 2746 4936 2774
rect 4816 800 4844 2746
rect 5184 2310 5212 2926
rect 5276 2514 5304 6802
rect 5356 4548 5408 4554
rect 5356 4490 5408 4496
rect 5368 4010 5396 4490
rect 5356 4004 5408 4010
rect 5356 3946 5408 3952
rect 5460 3058 5488 16186
rect 6196 15162 6224 16458
rect 6184 15156 6236 15162
rect 6184 15098 6236 15104
rect 6184 13252 6236 13258
rect 6184 13194 6236 13200
rect 6196 4010 6224 13194
rect 6288 9654 6316 21830
rect 7196 20256 7248 20262
rect 7196 20198 7248 20204
rect 6736 19916 6788 19922
rect 6736 19858 6788 19864
rect 6748 19802 6776 19858
rect 6748 19774 6868 19802
rect 6840 19378 6868 19774
rect 7012 19712 7064 19718
rect 7012 19654 7064 19660
rect 6828 19372 6880 19378
rect 6828 19314 6880 19320
rect 6840 18834 6868 19314
rect 6828 18828 6880 18834
rect 6828 18770 6880 18776
rect 6840 16658 6868 18770
rect 6828 16652 6880 16658
rect 6828 16594 6880 16600
rect 6840 16130 6868 16594
rect 6840 16114 6960 16130
rect 6840 16108 6972 16114
rect 6840 16102 6920 16108
rect 6920 16050 6972 16056
rect 6368 15496 6420 15502
rect 6368 15438 6420 15444
rect 6380 14958 6408 15438
rect 6368 14952 6420 14958
rect 6368 14894 6420 14900
rect 6380 13938 6408 14894
rect 6368 13932 6420 13938
rect 6368 13874 6420 13880
rect 7024 13394 7052 19654
rect 7208 18834 7236 20198
rect 7300 19718 7328 22374
rect 7564 22094 7616 22098
rect 7760 22094 7788 22578
rect 7564 22092 7788 22094
rect 7616 22066 7788 22092
rect 7564 22034 7616 22040
rect 7576 21486 7604 22034
rect 8208 22024 8260 22030
rect 8208 21966 8260 21972
rect 8220 21876 8248 21966
rect 8220 21848 8340 21876
rect 7950 21788 8258 21797
rect 7950 21786 7956 21788
rect 8012 21786 8036 21788
rect 8092 21786 8116 21788
rect 8172 21786 8196 21788
rect 8252 21786 8258 21788
rect 8012 21734 8014 21786
rect 8194 21734 8196 21786
rect 7950 21732 7956 21734
rect 8012 21732 8036 21734
rect 8092 21732 8116 21734
rect 8172 21732 8196 21734
rect 8252 21732 8258 21734
rect 7950 21723 8258 21732
rect 8312 21622 8340 21848
rect 8300 21616 8352 21622
rect 8300 21558 8352 21564
rect 7564 21480 7616 21486
rect 7564 21422 7616 21428
rect 7288 19712 7340 19718
rect 7288 19654 7340 19660
rect 7576 19514 7604 21422
rect 8312 20806 8340 21558
rect 8300 20800 8352 20806
rect 8300 20742 8352 20748
rect 7950 20700 8258 20709
rect 7950 20698 7956 20700
rect 8012 20698 8036 20700
rect 8092 20698 8116 20700
rect 8172 20698 8196 20700
rect 8252 20698 8258 20700
rect 8012 20646 8014 20698
rect 8194 20646 8196 20698
rect 7950 20644 7956 20646
rect 8012 20644 8036 20646
rect 8092 20644 8116 20646
rect 8172 20644 8196 20646
rect 8252 20644 8258 20646
rect 7950 20635 8258 20644
rect 8300 20460 8352 20466
rect 8300 20402 8352 20408
rect 7656 20324 7708 20330
rect 7656 20266 7708 20272
rect 7564 19508 7616 19514
rect 7564 19450 7616 19456
rect 7196 18828 7248 18834
rect 7196 18770 7248 18776
rect 7380 18624 7432 18630
rect 7380 18566 7432 18572
rect 7104 14000 7156 14006
rect 7104 13942 7156 13948
rect 7012 13388 7064 13394
rect 7012 13330 7064 13336
rect 7116 12850 7144 13942
rect 7392 13530 7420 18566
rect 7668 17202 7696 20266
rect 8312 19718 8340 20402
rect 8404 19938 8432 24618
rect 8484 22976 8536 22982
rect 8484 22918 8536 22924
rect 8496 22710 8524 22918
rect 8484 22704 8536 22710
rect 8484 22646 8536 22652
rect 8588 22094 8616 24686
rect 8496 22066 8616 22094
rect 8496 21894 8524 22066
rect 8484 21888 8536 21894
rect 8484 21830 8536 21836
rect 8496 20942 8524 21830
rect 8576 21480 8628 21486
rect 8576 21422 8628 21428
rect 8588 21146 8616 21422
rect 8576 21140 8628 21146
rect 8576 21082 8628 21088
rect 8484 20936 8536 20942
rect 8484 20878 8536 20884
rect 8484 20800 8536 20806
rect 8484 20742 8536 20748
rect 8496 20058 8524 20742
rect 8484 20052 8536 20058
rect 8484 19994 8536 20000
rect 8404 19910 8616 19938
rect 8484 19780 8536 19786
rect 8484 19722 8536 19728
rect 8300 19712 8352 19718
rect 8300 19654 8352 19660
rect 8392 19712 8444 19718
rect 8392 19654 8444 19660
rect 7950 19612 8258 19621
rect 7950 19610 7956 19612
rect 8012 19610 8036 19612
rect 8092 19610 8116 19612
rect 8172 19610 8196 19612
rect 8252 19610 8258 19612
rect 8012 19558 8014 19610
rect 8194 19558 8196 19610
rect 7950 19556 7956 19558
rect 8012 19556 8036 19558
rect 8092 19556 8116 19558
rect 8172 19556 8196 19558
rect 8252 19556 8258 19558
rect 7950 19547 8258 19556
rect 8312 18834 8340 19654
rect 8300 18828 8352 18834
rect 8300 18770 8352 18776
rect 8404 18766 8432 19654
rect 8392 18760 8444 18766
rect 8392 18702 8444 18708
rect 8496 18630 8524 19722
rect 8484 18624 8536 18630
rect 8484 18566 8536 18572
rect 7950 18524 8258 18533
rect 7950 18522 7956 18524
rect 8012 18522 8036 18524
rect 8092 18522 8116 18524
rect 8172 18522 8196 18524
rect 8252 18522 8258 18524
rect 8012 18470 8014 18522
rect 8194 18470 8196 18522
rect 7950 18468 7956 18470
rect 8012 18468 8036 18470
rect 8092 18468 8116 18470
rect 8172 18468 8196 18470
rect 8252 18468 8258 18470
rect 7950 18459 8258 18468
rect 8300 18284 8352 18290
rect 8300 18226 8352 18232
rect 7748 18148 7800 18154
rect 7748 18090 7800 18096
rect 7656 17196 7708 17202
rect 7656 17138 7708 17144
rect 7668 16794 7696 17138
rect 7656 16788 7708 16794
rect 7656 16730 7708 16736
rect 7472 16652 7524 16658
rect 7472 16594 7524 16600
rect 7380 13524 7432 13530
rect 7380 13466 7432 13472
rect 7380 13184 7432 13190
rect 7380 13126 7432 13132
rect 7392 12986 7420 13126
rect 7380 12980 7432 12986
rect 7380 12922 7432 12928
rect 7104 12844 7156 12850
rect 7104 12786 7156 12792
rect 6920 12096 6972 12102
rect 6920 12038 6972 12044
rect 6276 9648 6328 9654
rect 6276 9590 6328 9596
rect 6644 4140 6696 4146
rect 6644 4082 6696 4088
rect 6184 4004 6236 4010
rect 6184 3946 6236 3952
rect 6092 3936 6144 3942
rect 6092 3878 6144 3884
rect 6368 3936 6420 3942
rect 6368 3878 6420 3884
rect 5448 3052 5500 3058
rect 5448 2994 5500 3000
rect 5264 2508 5316 2514
rect 5264 2450 5316 2456
rect 6104 2446 6132 3878
rect 6380 3670 6408 3878
rect 6368 3664 6420 3670
rect 6368 3606 6420 3612
rect 6460 3664 6512 3670
rect 6460 3606 6512 3612
rect 6276 3528 6328 3534
rect 6276 3470 6328 3476
rect 6092 2440 6144 2446
rect 6092 2382 6144 2388
rect 5908 2372 5960 2378
rect 5908 2314 5960 2320
rect 5172 2304 5224 2310
rect 5172 2246 5224 2252
rect 5184 800 5212 2246
rect 5540 1760 5592 1766
rect 5540 1702 5592 1708
rect 5552 800 5580 1702
rect 5920 800 5948 2314
rect 6104 1766 6132 2382
rect 6092 1760 6144 1766
rect 6092 1702 6144 1708
rect 6288 800 6316 3470
rect 6472 2922 6500 3606
rect 6460 2916 6512 2922
rect 6460 2858 6512 2864
rect 6656 800 6684 4082
rect 6932 3738 6960 12038
rect 7116 9518 7144 12786
rect 7484 12442 7512 16594
rect 7760 15706 7788 18090
rect 7840 17536 7892 17542
rect 7840 17478 7892 17484
rect 7852 17338 7880 17478
rect 7950 17436 8258 17445
rect 7950 17434 7956 17436
rect 8012 17434 8036 17436
rect 8092 17434 8116 17436
rect 8172 17434 8196 17436
rect 8252 17434 8258 17436
rect 8012 17382 8014 17434
rect 8194 17382 8196 17434
rect 7950 17380 7956 17382
rect 8012 17380 8036 17382
rect 8092 17380 8116 17382
rect 8172 17380 8196 17382
rect 8252 17380 8258 17382
rect 7950 17371 8258 17380
rect 7840 17332 7892 17338
rect 7840 17274 7892 17280
rect 7840 16992 7892 16998
rect 7840 16934 7892 16940
rect 7852 16182 7880 16934
rect 7950 16348 8258 16357
rect 7950 16346 7956 16348
rect 8012 16346 8036 16348
rect 8092 16346 8116 16348
rect 8172 16346 8196 16348
rect 8252 16346 8258 16348
rect 8012 16294 8014 16346
rect 8194 16294 8196 16346
rect 7950 16292 7956 16294
rect 8012 16292 8036 16294
rect 8092 16292 8116 16294
rect 8172 16292 8196 16294
rect 8252 16292 8258 16294
rect 7950 16283 8258 16292
rect 7840 16176 7892 16182
rect 7840 16118 7892 16124
rect 7748 15700 7800 15706
rect 7748 15642 7800 15648
rect 7564 15020 7616 15026
rect 7564 14962 7616 14968
rect 7576 14482 7604 14962
rect 7564 14476 7616 14482
rect 7564 14418 7616 14424
rect 7576 13870 7604 14418
rect 7760 14414 7788 15642
rect 7950 15260 8258 15269
rect 7950 15258 7956 15260
rect 8012 15258 8036 15260
rect 8092 15258 8116 15260
rect 8172 15258 8196 15260
rect 8252 15258 8258 15260
rect 8012 15206 8014 15258
rect 8194 15206 8196 15258
rect 7950 15204 7956 15206
rect 8012 15204 8036 15206
rect 8092 15204 8116 15206
rect 8172 15204 8196 15206
rect 8252 15204 8258 15206
rect 7950 15195 8258 15204
rect 7748 14408 7800 14414
rect 7748 14350 7800 14356
rect 7950 14172 8258 14181
rect 7950 14170 7956 14172
rect 8012 14170 8036 14172
rect 8092 14170 8116 14172
rect 8172 14170 8196 14172
rect 8252 14170 8258 14172
rect 8012 14118 8014 14170
rect 8194 14118 8196 14170
rect 7950 14116 7956 14118
rect 8012 14116 8036 14118
rect 8092 14116 8116 14118
rect 8172 14116 8196 14118
rect 8252 14116 8258 14118
rect 7950 14107 8258 14116
rect 8312 14074 8340 18226
rect 8392 18216 8444 18222
rect 8392 18158 8444 18164
rect 8300 14068 8352 14074
rect 8300 14010 8352 14016
rect 7564 13864 7616 13870
rect 7564 13806 7616 13812
rect 7950 13084 8258 13093
rect 7950 13082 7956 13084
rect 8012 13082 8036 13084
rect 8092 13082 8116 13084
rect 8172 13082 8196 13084
rect 8252 13082 8258 13084
rect 8012 13030 8014 13082
rect 8194 13030 8196 13082
rect 7950 13028 7956 13030
rect 8012 13028 8036 13030
rect 8092 13028 8116 13030
rect 8172 13028 8196 13030
rect 8252 13028 8258 13030
rect 7950 13019 8258 13028
rect 8404 12986 8432 18158
rect 8392 12980 8444 12986
rect 8392 12922 8444 12928
rect 7656 12640 7708 12646
rect 7656 12582 7708 12588
rect 7472 12436 7524 12442
rect 7472 12378 7524 12384
rect 7196 11552 7248 11558
rect 7196 11494 7248 11500
rect 7104 9512 7156 9518
rect 7104 9454 7156 9460
rect 7104 9376 7156 9382
rect 7104 9318 7156 9324
rect 7116 4622 7144 9318
rect 7104 4616 7156 4622
rect 7104 4558 7156 4564
rect 6920 3732 6972 3738
rect 6920 3674 6972 3680
rect 7012 3528 7064 3534
rect 7012 3470 7064 3476
rect 6736 2916 6788 2922
rect 6736 2858 6788 2864
rect 6748 2650 6776 2858
rect 6736 2644 6788 2650
rect 6736 2586 6788 2592
rect 7024 800 7052 3470
rect 7208 3398 7236 11494
rect 7288 4208 7340 4214
rect 7288 4150 7340 4156
rect 7300 3534 7328 4150
rect 7380 3936 7432 3942
rect 7380 3878 7432 3884
rect 7288 3528 7340 3534
rect 7288 3470 7340 3476
rect 7196 3392 7248 3398
rect 7196 3334 7248 3340
rect 7392 3058 7420 3878
rect 7380 3052 7432 3058
rect 7380 2994 7432 3000
rect 7102 2408 7158 2417
rect 7102 2343 7158 2352
rect 7116 2310 7144 2343
rect 7104 2304 7156 2310
rect 7104 2246 7156 2252
rect 7392 800 7420 2994
rect 7668 2990 7696 12582
rect 8496 12306 8524 18566
rect 8588 17270 8616 19910
rect 8680 18426 8708 32370
rect 9128 29640 9180 29646
rect 9128 29582 9180 29588
rect 9140 28626 9168 29582
rect 9128 28620 9180 28626
rect 9128 28562 9180 28568
rect 9128 27464 9180 27470
rect 9128 27406 9180 27412
rect 9140 26450 9168 27406
rect 9128 26444 9180 26450
rect 9128 26386 9180 26392
rect 9232 24698 9260 36110
rect 9692 33658 9720 36654
rect 9680 33652 9732 33658
rect 9680 33594 9732 33600
rect 9312 32904 9364 32910
rect 9312 32846 9364 32852
rect 9140 24670 9260 24698
rect 9140 24614 9168 24670
rect 9128 24608 9180 24614
rect 9128 24550 9180 24556
rect 9220 24200 9272 24206
rect 9220 24142 9272 24148
rect 8944 24132 8996 24138
rect 8944 24074 8996 24080
rect 8956 23798 8984 24074
rect 8944 23792 8996 23798
rect 8944 23734 8996 23740
rect 8956 22710 8984 23734
rect 9128 23044 9180 23050
rect 9128 22986 9180 22992
rect 8944 22704 8996 22710
rect 8944 22646 8996 22652
rect 9036 20460 9088 20466
rect 9036 20402 9088 20408
rect 8760 18760 8812 18766
rect 8760 18702 8812 18708
rect 8668 18420 8720 18426
rect 8668 18362 8720 18368
rect 8772 17882 8800 18702
rect 8760 17876 8812 17882
rect 8760 17818 8812 17824
rect 8576 17264 8628 17270
rect 8576 17206 8628 17212
rect 8772 16794 8800 17818
rect 8852 16992 8904 16998
rect 8852 16934 8904 16940
rect 8760 16788 8812 16794
rect 8760 16730 8812 16736
rect 8772 15706 8800 16730
rect 8760 15700 8812 15706
rect 8760 15642 8812 15648
rect 8772 15434 8800 15642
rect 8760 15428 8812 15434
rect 8760 15370 8812 15376
rect 8772 15094 8800 15370
rect 8760 15088 8812 15094
rect 8760 15030 8812 15036
rect 8576 14952 8628 14958
rect 8576 14894 8628 14900
rect 8588 14618 8616 14894
rect 8576 14612 8628 14618
rect 8576 14554 8628 14560
rect 8772 14006 8800 15030
rect 8864 14498 8892 16934
rect 9048 14618 9076 20402
rect 9140 19990 9168 22986
rect 9128 19984 9180 19990
rect 9128 19926 9180 19932
rect 9128 19848 9180 19854
rect 9128 19790 9180 19796
rect 9140 19514 9168 19790
rect 9128 19508 9180 19514
rect 9128 19450 9180 19456
rect 9140 18222 9168 19450
rect 9128 18216 9180 18222
rect 9128 18158 9180 18164
rect 9232 17202 9260 24142
rect 9324 20602 9352 32846
rect 9784 30122 9812 39374
rect 10232 33516 10284 33522
rect 10232 33458 10284 33464
rect 10244 30190 10272 33458
rect 10428 33114 10456 45902
rect 10612 45082 10640 46446
rect 10600 45076 10652 45082
rect 10600 45018 10652 45024
rect 10704 44878 10732 47194
rect 10888 45422 10916 55186
rect 10968 49360 11020 49366
rect 10968 49302 11020 49308
rect 10980 47258 11008 49302
rect 10968 47252 11020 47258
rect 10968 47194 11020 47200
rect 10980 47002 11008 47194
rect 11520 47116 11572 47122
rect 11520 47058 11572 47064
rect 10980 46986 11100 47002
rect 10968 46980 11100 46986
rect 11020 46974 11100 46980
rect 10968 46922 11020 46928
rect 10968 46368 11020 46374
rect 10968 46310 11020 46316
rect 10876 45416 10928 45422
rect 10876 45358 10928 45364
rect 10692 44872 10744 44878
rect 10692 44814 10744 44820
rect 10980 44146 11008 46310
rect 11072 44878 11100 46974
rect 11152 46436 11204 46442
rect 11152 46378 11204 46384
rect 11060 44872 11112 44878
rect 11060 44814 11112 44820
rect 10980 44118 11100 44146
rect 11072 43178 11100 44118
rect 11164 43314 11192 46378
rect 11532 46034 11560 47058
rect 12084 46034 12112 56200
rect 13464 54194 13492 56200
rect 14844 54194 14872 56200
rect 16224 56114 16252 56200
rect 16316 56114 16344 56222
rect 16224 56086 16344 56114
rect 16500 54210 16528 56222
rect 17590 56200 17646 57000
rect 18970 56200 19026 57000
rect 20350 56200 20406 57000
rect 21730 56200 21786 57000
rect 22756 56222 23060 56250
rect 16500 54194 16620 54210
rect 17604 54194 17632 56200
rect 17950 54428 18258 54437
rect 17950 54426 17956 54428
rect 18012 54426 18036 54428
rect 18092 54426 18116 54428
rect 18172 54426 18196 54428
rect 18252 54426 18258 54428
rect 18012 54374 18014 54426
rect 18194 54374 18196 54426
rect 17950 54372 17956 54374
rect 18012 54372 18036 54374
rect 18092 54372 18116 54374
rect 18172 54372 18196 54374
rect 18252 54372 18258 54374
rect 17950 54363 18258 54372
rect 18984 54330 19012 56200
rect 18972 54324 19024 54330
rect 18972 54266 19024 54272
rect 13452 54188 13504 54194
rect 13452 54130 13504 54136
rect 14832 54188 14884 54194
rect 16500 54188 16632 54194
rect 16500 54182 16580 54188
rect 14832 54130 14884 54136
rect 16580 54130 16632 54136
rect 17592 54188 17644 54194
rect 17592 54130 17644 54136
rect 18984 54126 19012 54266
rect 18972 54120 19024 54126
rect 18972 54062 19024 54068
rect 18788 54052 18840 54058
rect 18788 53994 18840 54000
rect 12624 53984 12676 53990
rect 12624 53926 12676 53932
rect 14924 53984 14976 53990
rect 14924 53926 14976 53932
rect 15476 53984 15528 53990
rect 15476 53926 15528 53932
rect 17132 53984 17184 53990
rect 17132 53926 17184 53932
rect 12348 48544 12400 48550
rect 12348 48486 12400 48492
rect 12360 47734 12388 48486
rect 12348 47728 12400 47734
rect 12348 47670 12400 47676
rect 12636 47666 12664 53926
rect 12950 53884 13258 53893
rect 12950 53882 12956 53884
rect 13012 53882 13036 53884
rect 13092 53882 13116 53884
rect 13172 53882 13196 53884
rect 13252 53882 13258 53884
rect 13012 53830 13014 53882
rect 13194 53830 13196 53882
rect 12950 53828 12956 53830
rect 13012 53828 13036 53830
rect 13092 53828 13116 53830
rect 13172 53828 13196 53830
rect 13252 53828 13258 53830
rect 12950 53819 13258 53828
rect 12950 52796 13258 52805
rect 12950 52794 12956 52796
rect 13012 52794 13036 52796
rect 13092 52794 13116 52796
rect 13172 52794 13196 52796
rect 13252 52794 13258 52796
rect 13012 52742 13014 52794
rect 13194 52742 13196 52794
rect 12950 52740 12956 52742
rect 13012 52740 13036 52742
rect 13092 52740 13116 52742
rect 13172 52740 13196 52742
rect 13252 52740 13258 52742
rect 12950 52731 13258 52740
rect 12950 51708 13258 51717
rect 12950 51706 12956 51708
rect 13012 51706 13036 51708
rect 13092 51706 13116 51708
rect 13172 51706 13196 51708
rect 13252 51706 13258 51708
rect 13012 51654 13014 51706
rect 13194 51654 13196 51706
rect 12950 51652 12956 51654
rect 13012 51652 13036 51654
rect 13092 51652 13116 51654
rect 13172 51652 13196 51654
rect 13252 51652 13258 51654
rect 12950 51643 13258 51652
rect 12950 50620 13258 50629
rect 12950 50618 12956 50620
rect 13012 50618 13036 50620
rect 13092 50618 13116 50620
rect 13172 50618 13196 50620
rect 13252 50618 13258 50620
rect 13012 50566 13014 50618
rect 13194 50566 13196 50618
rect 12950 50564 12956 50566
rect 13012 50564 13036 50566
rect 13092 50564 13116 50566
rect 13172 50564 13196 50566
rect 13252 50564 13258 50566
rect 12950 50555 13258 50564
rect 12950 49532 13258 49541
rect 12950 49530 12956 49532
rect 13012 49530 13036 49532
rect 13092 49530 13116 49532
rect 13172 49530 13196 49532
rect 13252 49530 13258 49532
rect 13012 49478 13014 49530
rect 13194 49478 13196 49530
rect 12950 49476 12956 49478
rect 13012 49476 13036 49478
rect 13092 49476 13116 49478
rect 13172 49476 13196 49478
rect 13252 49476 13258 49478
rect 12950 49467 13258 49476
rect 12950 48444 13258 48453
rect 12950 48442 12956 48444
rect 13012 48442 13036 48444
rect 13092 48442 13116 48444
rect 13172 48442 13196 48444
rect 13252 48442 13258 48444
rect 13012 48390 13014 48442
rect 13194 48390 13196 48442
rect 12950 48388 12956 48390
rect 13012 48388 13036 48390
rect 13092 48388 13116 48390
rect 13172 48388 13196 48390
rect 13252 48388 13258 48390
rect 12950 48379 13258 48388
rect 14464 48000 14516 48006
rect 14464 47942 14516 47948
rect 12624 47660 12676 47666
rect 12624 47602 12676 47608
rect 12950 47356 13258 47365
rect 12950 47354 12956 47356
rect 13012 47354 13036 47356
rect 13092 47354 13116 47356
rect 13172 47354 13196 47356
rect 13252 47354 13258 47356
rect 13012 47302 13014 47354
rect 13194 47302 13196 47354
rect 12950 47300 12956 47302
rect 13012 47300 13036 47302
rect 13092 47300 13116 47302
rect 13172 47300 13196 47302
rect 13252 47300 13258 47302
rect 12950 47291 13258 47300
rect 14188 47048 14240 47054
rect 14188 46990 14240 46996
rect 12950 46268 13258 46277
rect 12950 46266 12956 46268
rect 13012 46266 13036 46268
rect 13092 46266 13116 46268
rect 13172 46266 13196 46268
rect 13252 46266 13258 46268
rect 13012 46214 13014 46266
rect 13194 46214 13196 46266
rect 12950 46212 12956 46214
rect 13012 46212 13036 46214
rect 13092 46212 13116 46214
rect 13172 46212 13196 46214
rect 13252 46212 13258 46214
rect 12950 46203 13258 46212
rect 14200 46034 14228 46990
rect 14476 46986 14504 47942
rect 14832 47592 14884 47598
rect 14832 47534 14884 47540
rect 14280 46980 14332 46986
rect 14280 46922 14332 46928
rect 14464 46980 14516 46986
rect 14464 46922 14516 46928
rect 14292 46646 14320 46922
rect 14280 46640 14332 46646
rect 14280 46582 14332 46588
rect 11520 46028 11572 46034
rect 11520 45970 11572 45976
rect 12072 46028 12124 46034
rect 12072 45970 12124 45976
rect 14188 46028 14240 46034
rect 14188 45970 14240 45976
rect 11532 45082 11560 45970
rect 12950 45180 13258 45189
rect 12950 45178 12956 45180
rect 13012 45178 13036 45180
rect 13092 45178 13116 45180
rect 13172 45178 13196 45180
rect 13252 45178 13258 45180
rect 13012 45126 13014 45178
rect 13194 45126 13196 45178
rect 12950 45124 12956 45126
rect 13012 45124 13036 45126
rect 13092 45124 13116 45126
rect 13172 45124 13196 45126
rect 13252 45124 13258 45126
rect 12950 45115 13258 45124
rect 11336 45076 11388 45082
rect 11336 45018 11388 45024
rect 11520 45076 11572 45082
rect 11520 45018 11572 45024
rect 11152 43308 11204 43314
rect 11152 43250 11204 43256
rect 11060 43172 11112 43178
rect 11060 43114 11112 43120
rect 11348 40050 11376 45018
rect 12950 44092 13258 44101
rect 12950 44090 12956 44092
rect 13012 44090 13036 44092
rect 13092 44090 13116 44092
rect 13172 44090 13196 44092
rect 13252 44090 13258 44092
rect 13012 44038 13014 44090
rect 13194 44038 13196 44090
rect 12950 44036 12956 44038
rect 13012 44036 13036 44038
rect 13092 44036 13116 44038
rect 13172 44036 13196 44038
rect 13252 44036 13258 44038
rect 12950 44027 13258 44036
rect 11704 43308 11756 43314
rect 11704 43250 11756 43256
rect 11612 43104 11664 43110
rect 11612 43046 11664 43052
rect 11336 40044 11388 40050
rect 11336 39986 11388 39992
rect 11348 36922 11376 39986
rect 11336 36916 11388 36922
rect 11336 36858 11388 36864
rect 11244 36848 11296 36854
rect 11244 36790 11296 36796
rect 10416 33108 10468 33114
rect 10416 33050 10468 33056
rect 11256 30326 11284 36790
rect 11624 36582 11652 43046
rect 11716 36922 11744 43250
rect 12348 43240 12400 43246
rect 12348 43182 12400 43188
rect 12360 40186 12388 43182
rect 12950 43004 13258 43013
rect 12950 43002 12956 43004
rect 13012 43002 13036 43004
rect 13092 43002 13116 43004
rect 13172 43002 13196 43004
rect 13252 43002 13258 43004
rect 13012 42950 13014 43002
rect 13194 42950 13196 43002
rect 12950 42948 12956 42950
rect 13012 42948 13036 42950
rect 13092 42948 13116 42950
rect 13172 42948 13196 42950
rect 13252 42948 13258 42950
rect 12950 42939 13258 42948
rect 12950 41916 13258 41925
rect 12950 41914 12956 41916
rect 13012 41914 13036 41916
rect 13092 41914 13116 41916
rect 13172 41914 13196 41916
rect 13252 41914 13258 41916
rect 13012 41862 13014 41914
rect 13194 41862 13196 41914
rect 12950 41860 12956 41862
rect 13012 41860 13036 41862
rect 13092 41860 13116 41862
rect 13172 41860 13196 41862
rect 13252 41860 13258 41862
rect 12950 41851 13258 41860
rect 14844 41414 14872 47534
rect 14936 47122 14964 53926
rect 14924 47116 14976 47122
rect 14924 47058 14976 47064
rect 15488 46510 15516 53926
rect 16948 52488 17000 52494
rect 16948 52430 17000 52436
rect 16028 50516 16080 50522
rect 16028 50458 16080 50464
rect 15476 46504 15528 46510
rect 15476 46446 15528 46452
rect 15752 45076 15804 45082
rect 15752 45018 15804 45024
rect 14844 41386 14964 41414
rect 12950 40828 13258 40837
rect 12950 40826 12956 40828
rect 13012 40826 13036 40828
rect 13092 40826 13116 40828
rect 13172 40826 13196 40828
rect 13252 40826 13258 40828
rect 13012 40774 13014 40826
rect 13194 40774 13196 40826
rect 12950 40772 12956 40774
rect 13012 40772 13036 40774
rect 13092 40772 13116 40774
rect 13172 40772 13196 40774
rect 13252 40772 13258 40774
rect 12950 40763 13258 40772
rect 12348 40180 12400 40186
rect 12348 40122 12400 40128
rect 12950 39740 13258 39749
rect 12950 39738 12956 39740
rect 13012 39738 13036 39740
rect 13092 39738 13116 39740
rect 13172 39738 13196 39740
rect 13252 39738 13258 39740
rect 13012 39686 13014 39738
rect 13194 39686 13196 39738
rect 12950 39684 12956 39686
rect 13012 39684 13036 39686
rect 13092 39684 13116 39686
rect 13172 39684 13196 39686
rect 13252 39684 13258 39686
rect 12950 39675 13258 39684
rect 12950 38652 13258 38661
rect 12950 38650 12956 38652
rect 13012 38650 13036 38652
rect 13092 38650 13116 38652
rect 13172 38650 13196 38652
rect 13252 38650 13258 38652
rect 13012 38598 13014 38650
rect 13194 38598 13196 38650
rect 12950 38596 12956 38598
rect 13012 38596 13036 38598
rect 13092 38596 13116 38598
rect 13172 38596 13196 38598
rect 13252 38596 13258 38598
rect 12950 38587 13258 38596
rect 12950 37564 13258 37573
rect 12950 37562 12956 37564
rect 13012 37562 13036 37564
rect 13092 37562 13116 37564
rect 13172 37562 13196 37564
rect 13252 37562 13258 37564
rect 13012 37510 13014 37562
rect 13194 37510 13196 37562
rect 12950 37508 12956 37510
rect 13012 37508 13036 37510
rect 13092 37508 13116 37510
rect 13172 37508 13196 37510
rect 13252 37508 13258 37510
rect 12950 37499 13258 37508
rect 11704 36916 11756 36922
rect 11704 36858 11756 36864
rect 11612 36576 11664 36582
rect 11612 36518 11664 36524
rect 11624 34678 11652 36518
rect 12950 36476 13258 36485
rect 12950 36474 12956 36476
rect 13012 36474 13036 36476
rect 13092 36474 13116 36476
rect 13172 36474 13196 36476
rect 13252 36474 13258 36476
rect 13012 36422 13014 36474
rect 13194 36422 13196 36474
rect 12950 36420 12956 36422
rect 13012 36420 13036 36422
rect 13092 36420 13116 36422
rect 13172 36420 13196 36422
rect 13252 36420 13258 36422
rect 12950 36411 13258 36420
rect 12950 35388 13258 35397
rect 12950 35386 12956 35388
rect 13012 35386 13036 35388
rect 13092 35386 13116 35388
rect 13172 35386 13196 35388
rect 13252 35386 13258 35388
rect 13012 35334 13014 35386
rect 13194 35334 13196 35386
rect 12950 35332 12956 35334
rect 13012 35332 13036 35334
rect 13092 35332 13116 35334
rect 13172 35332 13196 35334
rect 13252 35332 13258 35334
rect 12950 35323 13258 35332
rect 11612 34672 11664 34678
rect 11612 34614 11664 34620
rect 12950 34300 13258 34309
rect 12950 34298 12956 34300
rect 13012 34298 13036 34300
rect 13092 34298 13116 34300
rect 13172 34298 13196 34300
rect 13252 34298 13258 34300
rect 13012 34246 13014 34298
rect 13194 34246 13196 34298
rect 12950 34244 12956 34246
rect 13012 34244 13036 34246
rect 13092 34244 13116 34246
rect 13172 34244 13196 34246
rect 13252 34244 13258 34246
rect 12950 34235 13258 34244
rect 12950 33212 13258 33221
rect 12950 33210 12956 33212
rect 13012 33210 13036 33212
rect 13092 33210 13116 33212
rect 13172 33210 13196 33212
rect 13252 33210 13258 33212
rect 13012 33158 13014 33210
rect 13194 33158 13196 33210
rect 12950 33156 12956 33158
rect 13012 33156 13036 33158
rect 13092 33156 13116 33158
rect 13172 33156 13196 33158
rect 13252 33156 13258 33158
rect 12950 33147 13258 33156
rect 13452 32224 13504 32230
rect 13452 32166 13504 32172
rect 12950 32124 13258 32133
rect 12950 32122 12956 32124
rect 13012 32122 13036 32124
rect 13092 32122 13116 32124
rect 13172 32122 13196 32124
rect 13252 32122 13258 32124
rect 13012 32070 13014 32122
rect 13194 32070 13196 32122
rect 12950 32068 12956 32070
rect 13012 32068 13036 32070
rect 13092 32068 13116 32070
rect 13172 32068 13196 32070
rect 13252 32068 13258 32070
rect 12950 32059 13258 32068
rect 13360 31952 13412 31958
rect 13360 31894 13412 31900
rect 11520 31816 11572 31822
rect 11520 31758 11572 31764
rect 11244 30320 11296 30326
rect 11244 30262 11296 30268
rect 10324 30252 10376 30258
rect 10324 30194 10376 30200
rect 10232 30184 10284 30190
rect 10232 30126 10284 30132
rect 9772 30116 9824 30122
rect 9772 30058 9824 30064
rect 10048 30116 10100 30122
rect 10048 30058 10100 30064
rect 9588 29504 9640 29510
rect 9588 29446 9640 29452
rect 9496 29028 9548 29034
rect 9496 28970 9548 28976
rect 9404 28620 9456 28626
rect 9404 28562 9456 28568
rect 9416 26994 9444 28562
rect 9404 26988 9456 26994
rect 9404 26930 9456 26936
rect 9508 26450 9536 28970
rect 9496 26444 9548 26450
rect 9496 26386 9548 26392
rect 9600 25362 9628 29446
rect 9772 28484 9824 28490
rect 9772 28426 9824 28432
rect 9784 28218 9812 28426
rect 9772 28212 9824 28218
rect 9772 28154 9824 28160
rect 9680 26784 9732 26790
rect 9680 26726 9732 26732
rect 9588 25356 9640 25362
rect 9588 25298 9640 25304
rect 9404 24404 9456 24410
rect 9600 24392 9628 25298
rect 9456 24364 9628 24392
rect 9404 24346 9456 24352
rect 9404 22228 9456 22234
rect 9404 22170 9456 22176
rect 9416 21418 9444 22170
rect 9508 22166 9536 24364
rect 9692 24070 9720 26726
rect 9772 24880 9824 24886
rect 9772 24822 9824 24828
rect 9680 24064 9732 24070
rect 9680 24006 9732 24012
rect 9496 22160 9548 22166
rect 9496 22102 9548 22108
rect 9496 21888 9548 21894
rect 9496 21830 9548 21836
rect 9404 21412 9456 21418
rect 9404 21354 9456 21360
rect 9312 20596 9364 20602
rect 9312 20538 9364 20544
rect 9312 19508 9364 19514
rect 9416 19496 9444 21354
rect 9508 20942 9536 21830
rect 9784 21690 9812 24822
rect 9864 22772 9916 22778
rect 9864 22714 9916 22720
rect 9876 22098 9904 22714
rect 9956 22432 10008 22438
rect 9956 22374 10008 22380
rect 9968 22234 9996 22374
rect 9956 22228 10008 22234
rect 9956 22170 10008 22176
rect 9864 22092 9916 22098
rect 9864 22034 9916 22040
rect 9772 21684 9824 21690
rect 9772 21626 9824 21632
rect 9876 21622 9904 22034
rect 10060 21894 10088 30058
rect 10244 29510 10272 30126
rect 10232 29504 10284 29510
rect 10232 29446 10284 29452
rect 10232 28756 10284 28762
rect 10232 28698 10284 28704
rect 10140 28416 10192 28422
rect 10140 28358 10192 28364
rect 10152 27062 10180 28358
rect 10244 27946 10272 28698
rect 10232 27940 10284 27946
rect 10232 27882 10284 27888
rect 10140 27056 10192 27062
rect 10140 26998 10192 27004
rect 10152 26450 10180 26998
rect 10244 26926 10272 27882
rect 10232 26920 10284 26926
rect 10232 26862 10284 26868
rect 10140 26444 10192 26450
rect 10140 26386 10192 26392
rect 10152 26314 10180 26386
rect 10140 26308 10192 26314
rect 10140 26250 10192 26256
rect 10140 24064 10192 24070
rect 10140 24006 10192 24012
rect 10152 23866 10180 24006
rect 10140 23860 10192 23866
rect 10140 23802 10192 23808
rect 10244 23746 10272 26862
rect 10336 25498 10364 30194
rect 11256 29850 11284 30262
rect 11244 29844 11296 29850
rect 11244 29786 11296 29792
rect 11256 29578 11284 29786
rect 11532 29714 11560 31758
rect 12950 31036 13258 31045
rect 12950 31034 12956 31036
rect 13012 31034 13036 31036
rect 13092 31034 13116 31036
rect 13172 31034 13196 31036
rect 13252 31034 13258 31036
rect 13012 30982 13014 31034
rect 13194 30982 13196 31034
rect 12950 30980 12956 30982
rect 13012 30980 13036 30982
rect 13092 30980 13116 30982
rect 13172 30980 13196 30982
rect 13252 30980 13258 30982
rect 12950 30971 13258 30980
rect 12532 30048 12584 30054
rect 12532 29990 12584 29996
rect 12544 29714 12572 29990
rect 12950 29948 13258 29957
rect 12950 29946 12956 29948
rect 13012 29946 13036 29948
rect 13092 29946 13116 29948
rect 13172 29946 13196 29948
rect 13252 29946 13258 29948
rect 13012 29894 13014 29946
rect 13194 29894 13196 29946
rect 12950 29892 12956 29894
rect 13012 29892 13036 29894
rect 13092 29892 13116 29894
rect 13172 29892 13196 29894
rect 13252 29892 13258 29894
rect 12950 29883 13258 29892
rect 11520 29708 11572 29714
rect 11520 29650 11572 29656
rect 12532 29708 12584 29714
rect 12532 29650 12584 29656
rect 11244 29572 11296 29578
rect 11244 29514 11296 29520
rect 10784 29164 10836 29170
rect 10784 29106 10836 29112
rect 10692 26308 10744 26314
rect 10692 26250 10744 26256
rect 10324 25492 10376 25498
rect 10324 25434 10376 25440
rect 10324 25152 10376 25158
rect 10324 25094 10376 25100
rect 10152 23718 10272 23746
rect 10152 22094 10180 23718
rect 10232 23520 10284 23526
rect 10232 23462 10284 23468
rect 10244 22778 10272 23462
rect 10232 22772 10284 22778
rect 10232 22714 10284 22720
rect 10152 22066 10272 22094
rect 10048 21888 10100 21894
rect 10048 21830 10100 21836
rect 9864 21616 9916 21622
rect 9864 21558 9916 21564
rect 9588 21480 9640 21486
rect 9588 21422 9640 21428
rect 9496 20936 9548 20942
rect 9496 20878 9548 20884
rect 9496 19712 9548 19718
rect 9496 19654 9548 19660
rect 9508 19514 9536 19654
rect 9364 19468 9444 19496
rect 9496 19508 9548 19514
rect 9312 19450 9364 19456
rect 9496 19450 9548 19456
rect 9220 17196 9272 17202
rect 9220 17138 9272 17144
rect 9324 17066 9352 19450
rect 9496 18624 9548 18630
rect 9496 18566 9548 18572
rect 9404 18216 9456 18222
rect 9404 18158 9456 18164
rect 9416 17746 9444 18158
rect 9404 17740 9456 17746
rect 9404 17682 9456 17688
rect 9508 17338 9536 18566
rect 9600 18426 9628 21422
rect 10244 21010 10272 22066
rect 10232 21004 10284 21010
rect 10232 20946 10284 20952
rect 10232 20800 10284 20806
rect 10232 20742 10284 20748
rect 10140 20528 10192 20534
rect 10140 20470 10192 20476
rect 9864 20052 9916 20058
rect 9864 19994 9916 20000
rect 9876 19786 9904 19994
rect 9864 19780 9916 19786
rect 9864 19722 9916 19728
rect 9680 19712 9732 19718
rect 9680 19654 9732 19660
rect 9588 18420 9640 18426
rect 9588 18362 9640 18368
rect 9496 17332 9548 17338
rect 9496 17274 9548 17280
rect 9312 17060 9364 17066
rect 9312 17002 9364 17008
rect 9588 16788 9640 16794
rect 9588 16730 9640 16736
rect 9600 16182 9628 16730
rect 9692 16658 9720 19654
rect 9772 19304 9824 19310
rect 9772 19246 9824 19252
rect 9784 17542 9812 19246
rect 9876 18358 9904 19722
rect 9864 18352 9916 18358
rect 9864 18294 9916 18300
rect 9772 17536 9824 17542
rect 9772 17478 9824 17484
rect 9680 16652 9732 16658
rect 9680 16594 9732 16600
rect 9588 16176 9640 16182
rect 9588 16118 9640 16124
rect 9588 16040 9640 16046
rect 9588 15982 9640 15988
rect 9312 15700 9364 15706
rect 9312 15642 9364 15648
rect 9036 14612 9088 14618
rect 9036 14554 9088 14560
rect 8864 14470 9076 14498
rect 8944 14408 8996 14414
rect 8944 14350 8996 14356
rect 8760 14000 8812 14006
rect 8760 13942 8812 13948
rect 8772 13258 8800 13942
rect 8760 13252 8812 13258
rect 8760 13194 8812 13200
rect 8772 12918 8800 13194
rect 8760 12912 8812 12918
rect 8760 12854 8812 12860
rect 8576 12708 8628 12714
rect 8576 12650 8628 12656
rect 8484 12300 8536 12306
rect 8484 12242 8536 12248
rect 7950 11996 8258 12005
rect 7950 11994 7956 11996
rect 8012 11994 8036 11996
rect 8092 11994 8116 11996
rect 8172 11994 8196 11996
rect 8252 11994 8258 11996
rect 8012 11942 8014 11994
rect 8194 11942 8196 11994
rect 7950 11940 7956 11942
rect 8012 11940 8036 11942
rect 8092 11940 8116 11942
rect 8172 11940 8196 11942
rect 8252 11940 8258 11942
rect 7950 11931 8258 11940
rect 8588 11354 8616 12650
rect 8760 12096 8812 12102
rect 8760 12038 8812 12044
rect 8772 11762 8800 12038
rect 8760 11756 8812 11762
rect 8760 11698 8812 11704
rect 8576 11348 8628 11354
rect 8576 11290 8628 11296
rect 7950 10908 8258 10917
rect 7950 10906 7956 10908
rect 8012 10906 8036 10908
rect 8092 10906 8116 10908
rect 8172 10906 8196 10908
rect 8252 10906 8258 10908
rect 8012 10854 8014 10906
rect 8194 10854 8196 10906
rect 7950 10852 7956 10854
rect 8012 10852 8036 10854
rect 8092 10852 8116 10854
rect 8172 10852 8196 10854
rect 8252 10852 8258 10854
rect 7950 10843 8258 10852
rect 8390 10024 8446 10033
rect 8390 9959 8446 9968
rect 8404 9926 8432 9959
rect 8392 9920 8444 9926
rect 8392 9862 8444 9868
rect 7950 9820 8258 9829
rect 7950 9818 7956 9820
rect 8012 9818 8036 9820
rect 8092 9818 8116 9820
rect 8172 9818 8196 9820
rect 8252 9818 8258 9820
rect 8012 9766 8014 9818
rect 8194 9766 8196 9818
rect 7950 9764 7956 9766
rect 8012 9764 8036 9766
rect 8092 9764 8116 9766
rect 8172 9764 8196 9766
rect 8252 9764 8258 9766
rect 7950 9755 8258 9764
rect 8208 9512 8260 9518
rect 8208 9454 8260 9460
rect 8220 8820 8248 9454
rect 8220 8792 8340 8820
rect 7950 8732 8258 8741
rect 7950 8730 7956 8732
rect 8012 8730 8036 8732
rect 8092 8730 8116 8732
rect 8172 8730 8196 8732
rect 8252 8730 8258 8732
rect 8012 8678 8014 8730
rect 8194 8678 8196 8730
rect 7950 8676 7956 8678
rect 8012 8676 8036 8678
rect 8092 8676 8116 8678
rect 8172 8676 8196 8678
rect 8252 8676 8258 8678
rect 7950 8667 8258 8676
rect 8114 8528 8170 8537
rect 8114 8463 8116 8472
rect 8168 8463 8170 8472
rect 8116 8434 8168 8440
rect 8312 8430 8340 8792
rect 8300 8424 8352 8430
rect 8300 8366 8352 8372
rect 8484 8356 8536 8362
rect 8484 8298 8536 8304
rect 8392 7812 8444 7818
rect 8392 7754 8444 7760
rect 7950 7644 8258 7653
rect 7950 7642 7956 7644
rect 8012 7642 8036 7644
rect 8092 7642 8116 7644
rect 8172 7642 8196 7644
rect 8252 7642 8258 7644
rect 8012 7590 8014 7642
rect 8194 7590 8196 7642
rect 7950 7588 7956 7590
rect 8012 7588 8036 7590
rect 8092 7588 8116 7590
rect 8172 7588 8196 7590
rect 8252 7588 8258 7590
rect 7950 7579 8258 7588
rect 7950 6556 8258 6565
rect 7950 6554 7956 6556
rect 8012 6554 8036 6556
rect 8092 6554 8116 6556
rect 8172 6554 8196 6556
rect 8252 6554 8258 6556
rect 8012 6502 8014 6554
rect 8194 6502 8196 6554
rect 7950 6500 7956 6502
rect 8012 6500 8036 6502
rect 8092 6500 8116 6502
rect 8172 6500 8196 6502
rect 8252 6500 8258 6502
rect 7950 6491 8258 6500
rect 8300 5704 8352 5710
rect 8300 5646 8352 5652
rect 7950 5468 8258 5477
rect 7950 5466 7956 5468
rect 8012 5466 8036 5468
rect 8092 5466 8116 5468
rect 8172 5466 8196 5468
rect 8252 5466 8258 5468
rect 8012 5414 8014 5466
rect 8194 5414 8196 5466
rect 7950 5412 7956 5414
rect 8012 5412 8036 5414
rect 8092 5412 8116 5414
rect 8172 5412 8196 5414
rect 8252 5412 8258 5414
rect 7950 5403 8258 5412
rect 8312 5250 8340 5646
rect 8220 5222 8340 5250
rect 8220 4690 8248 5222
rect 8208 4684 8260 4690
rect 8208 4626 8260 4632
rect 7950 4380 8258 4389
rect 7950 4378 7956 4380
rect 8012 4378 8036 4380
rect 8092 4378 8116 4380
rect 8172 4378 8196 4380
rect 8252 4378 8258 4380
rect 8012 4326 8014 4378
rect 8194 4326 8196 4378
rect 7950 4324 7956 4326
rect 8012 4324 8036 4326
rect 8092 4324 8116 4326
rect 8172 4324 8196 4326
rect 8252 4324 8258 4326
rect 7950 4315 8258 4324
rect 8404 4078 8432 7754
rect 8496 4690 8524 8298
rect 8772 6662 8800 11698
rect 8956 10742 8984 14350
rect 9048 12102 9076 14470
rect 9220 13320 9272 13326
rect 9220 13262 9272 13268
rect 9128 13184 9180 13190
rect 9128 13126 9180 13132
rect 9140 12238 9168 13126
rect 9128 12232 9180 12238
rect 9128 12174 9180 12180
rect 9036 12096 9088 12102
rect 9036 12038 9088 12044
rect 9128 12096 9180 12102
rect 9128 12038 9180 12044
rect 9140 11558 9168 12038
rect 9128 11552 9180 11558
rect 9128 11494 9180 11500
rect 8944 10736 8996 10742
rect 8944 10678 8996 10684
rect 9232 10674 9260 13262
rect 9220 10668 9272 10674
rect 9220 10610 9272 10616
rect 8944 10600 8996 10606
rect 9232 10554 9260 10610
rect 8944 10542 8996 10548
rect 8852 8832 8904 8838
rect 8852 8774 8904 8780
rect 8864 8566 8892 8774
rect 8852 8560 8904 8566
rect 8852 8502 8904 8508
rect 8760 6656 8812 6662
rect 8760 6598 8812 6604
rect 8852 4820 8904 4826
rect 8852 4762 8904 4768
rect 8484 4684 8536 4690
rect 8484 4626 8536 4632
rect 8864 4146 8892 4762
rect 8852 4140 8904 4146
rect 8852 4082 8904 4088
rect 8392 4072 8444 4078
rect 8392 4014 8444 4020
rect 8576 4072 8628 4078
rect 8576 4014 8628 4020
rect 8484 3528 8536 3534
rect 8484 3470 8536 3476
rect 7748 3392 7800 3398
rect 7748 3334 7800 3340
rect 7760 3058 7788 3334
rect 7950 3292 8258 3301
rect 7950 3290 7956 3292
rect 8012 3290 8036 3292
rect 8092 3290 8116 3292
rect 8172 3290 8196 3292
rect 8252 3290 8258 3292
rect 8012 3238 8014 3290
rect 8194 3238 8196 3290
rect 7950 3236 7956 3238
rect 8012 3236 8036 3238
rect 8092 3236 8116 3238
rect 8172 3236 8196 3238
rect 8252 3236 8258 3238
rect 7950 3227 8258 3236
rect 7748 3052 7800 3058
rect 7748 2994 7800 3000
rect 7656 2984 7708 2990
rect 7656 2926 7708 2932
rect 7760 800 7788 2994
rect 8208 2576 8260 2582
rect 8206 2544 8208 2553
rect 8260 2544 8262 2553
rect 8206 2479 8262 2488
rect 7840 2440 7892 2446
rect 7840 2382 7892 2388
rect 1490 0 1546 800
rect 1858 0 1914 800
rect 2226 0 2282 800
rect 2594 0 2650 800
rect 2962 0 3018 800
rect 3330 0 3386 800
rect 3698 0 3754 800
rect 4066 0 4122 800
rect 4434 0 4490 800
rect 4802 0 4858 800
rect 5170 0 5226 800
rect 5538 0 5594 800
rect 5906 0 5962 800
rect 6274 0 6330 800
rect 6642 0 6698 800
rect 7010 0 7066 800
rect 7378 0 7434 800
rect 7746 0 7802 800
rect 7852 762 7880 2382
rect 8392 2304 8444 2310
rect 8392 2246 8444 2252
rect 7950 2204 8258 2213
rect 7950 2202 7956 2204
rect 8012 2202 8036 2204
rect 8092 2202 8116 2204
rect 8172 2202 8196 2204
rect 8252 2202 8258 2204
rect 8012 2150 8014 2202
rect 8194 2150 8196 2202
rect 7950 2148 7956 2150
rect 8012 2148 8036 2150
rect 8092 2148 8116 2150
rect 8172 2148 8196 2150
rect 8252 2148 8258 2150
rect 7950 2139 8258 2148
rect 8404 2106 8432 2246
rect 8392 2100 8444 2106
rect 8392 2042 8444 2048
rect 8036 870 8156 898
rect 8036 762 8064 870
rect 8128 800 8156 870
rect 8496 800 8524 3470
rect 8588 3398 8616 4014
rect 8668 3936 8720 3942
rect 8668 3878 8720 3884
rect 8680 3738 8708 3878
rect 8668 3732 8720 3738
rect 8668 3674 8720 3680
rect 8576 3392 8628 3398
rect 8576 3334 8628 3340
rect 8956 3194 8984 10542
rect 9140 10526 9260 10554
rect 9140 10130 9168 10526
rect 9128 10124 9180 10130
rect 9128 10066 9180 10072
rect 9324 9722 9352 15642
rect 9404 15564 9456 15570
rect 9404 15506 9456 15512
rect 9416 13870 9444 15506
rect 9600 14414 9628 15982
rect 9956 15496 10008 15502
rect 9956 15438 10008 15444
rect 9680 15020 9732 15026
rect 9680 14962 9732 14968
rect 9692 14482 9720 14962
rect 9968 14822 9996 15438
rect 10152 14890 10180 20470
rect 10244 19394 10272 20742
rect 10336 19514 10364 25094
rect 10508 24132 10560 24138
rect 10508 24074 10560 24080
rect 10416 21480 10468 21486
rect 10416 21422 10468 21428
rect 10324 19508 10376 19514
rect 10324 19450 10376 19456
rect 10244 19378 10364 19394
rect 10244 19372 10376 19378
rect 10244 19366 10324 19372
rect 10324 19314 10376 19320
rect 10336 16266 10364 19314
rect 10428 16454 10456 21422
rect 10520 19242 10548 24074
rect 10600 23656 10652 23662
rect 10600 23598 10652 23604
rect 10612 23118 10640 23598
rect 10600 23112 10652 23118
rect 10600 23054 10652 23060
rect 10612 22710 10640 23054
rect 10600 22704 10652 22710
rect 10600 22646 10652 22652
rect 10600 21888 10652 21894
rect 10600 21830 10652 21836
rect 10508 19236 10560 19242
rect 10508 19178 10560 19184
rect 10612 16590 10640 21830
rect 10704 21146 10732 26250
rect 10692 21140 10744 21146
rect 10692 21082 10744 21088
rect 10796 18986 10824 29106
rect 11532 28626 11560 29650
rect 11796 29572 11848 29578
rect 11796 29514 11848 29520
rect 11520 28620 11572 28626
rect 11520 28562 11572 28568
rect 11808 28218 11836 29514
rect 12164 29028 12216 29034
rect 12164 28970 12216 28976
rect 11980 28416 12032 28422
rect 11980 28358 12032 28364
rect 11796 28212 11848 28218
rect 11796 28154 11848 28160
rect 11992 28150 12020 28358
rect 11980 28144 12032 28150
rect 11980 28086 12032 28092
rect 11152 28076 11204 28082
rect 11152 28018 11204 28024
rect 11164 26790 11192 28018
rect 11992 27606 12020 28086
rect 11980 27600 12032 27606
rect 11980 27542 12032 27548
rect 12072 27464 12124 27470
rect 12072 27406 12124 27412
rect 11336 27328 11388 27334
rect 11336 27270 11388 27276
rect 11348 26926 11376 27270
rect 11520 26988 11572 26994
rect 11520 26930 11572 26936
rect 11336 26920 11388 26926
rect 11336 26862 11388 26868
rect 11152 26784 11204 26790
rect 11152 26726 11204 26732
rect 11164 26450 11192 26726
rect 11152 26444 11204 26450
rect 11152 26386 11204 26392
rect 11244 26376 11296 26382
rect 11244 26318 11296 26324
rect 11152 25696 11204 25702
rect 11152 25638 11204 25644
rect 11060 25152 11112 25158
rect 11060 25094 11112 25100
rect 10876 24948 10928 24954
rect 10876 24890 10928 24896
rect 10888 24614 10916 24890
rect 10968 24744 11020 24750
rect 10968 24686 11020 24692
rect 10876 24608 10928 24614
rect 10876 24550 10928 24556
rect 10888 23186 10916 24550
rect 10980 23322 11008 24686
rect 10968 23316 11020 23322
rect 10968 23258 11020 23264
rect 10876 23180 10928 23186
rect 10876 23122 10928 23128
rect 10968 20800 11020 20806
rect 10968 20742 11020 20748
rect 10980 20058 11008 20742
rect 10968 20052 11020 20058
rect 10968 19994 11020 20000
rect 10980 19718 11008 19994
rect 10968 19712 11020 19718
rect 10968 19654 11020 19660
rect 10968 19236 11020 19242
rect 10968 19178 11020 19184
rect 10704 18958 10824 18986
rect 10704 17882 10732 18958
rect 10980 18766 11008 19178
rect 10784 18760 10836 18766
rect 10784 18702 10836 18708
rect 10968 18760 11020 18766
rect 10968 18702 11020 18708
rect 10692 17876 10744 17882
rect 10692 17818 10744 17824
rect 10600 16584 10652 16590
rect 10600 16526 10652 16532
rect 10416 16448 10468 16454
rect 10416 16390 10468 16396
rect 10692 16448 10744 16454
rect 10692 16390 10744 16396
rect 10336 16238 10456 16266
rect 10230 15464 10286 15473
rect 10230 15399 10232 15408
rect 10284 15399 10286 15408
rect 10232 15370 10284 15376
rect 10244 15094 10272 15370
rect 10232 15088 10284 15094
rect 10232 15030 10284 15036
rect 10140 14884 10192 14890
rect 10140 14826 10192 14832
rect 9956 14816 10008 14822
rect 9956 14758 10008 14764
rect 10324 14816 10376 14822
rect 10324 14758 10376 14764
rect 9968 14482 9996 14758
rect 9680 14476 9732 14482
rect 9680 14418 9732 14424
rect 9956 14476 10008 14482
rect 9956 14418 10008 14424
rect 9588 14408 9640 14414
rect 9588 14350 9640 14356
rect 9496 14272 9548 14278
rect 9496 14214 9548 14220
rect 9588 14272 9640 14278
rect 9588 14214 9640 14220
rect 10232 14272 10284 14278
rect 10232 14214 10284 14220
rect 9508 14074 9536 14214
rect 9496 14068 9548 14074
rect 9496 14010 9548 14016
rect 9404 13864 9456 13870
rect 9404 13806 9456 13812
rect 9416 12850 9444 13806
rect 9496 13728 9548 13734
rect 9496 13670 9548 13676
rect 9404 12844 9456 12850
rect 9404 12786 9456 12792
rect 9416 12714 9444 12786
rect 9404 12708 9456 12714
rect 9404 12650 9456 12656
rect 9508 11694 9536 13670
rect 9600 11830 9628 14214
rect 10140 14000 10192 14006
rect 10140 13942 10192 13948
rect 9772 13932 9824 13938
rect 9772 13874 9824 13880
rect 9680 12708 9732 12714
rect 9680 12650 9732 12656
rect 9692 11898 9720 12650
rect 9784 12442 9812 13874
rect 9772 12436 9824 12442
rect 9772 12378 9824 12384
rect 10152 11898 10180 13942
rect 9680 11892 9732 11898
rect 9680 11834 9732 11840
rect 10140 11892 10192 11898
rect 10140 11834 10192 11840
rect 9588 11824 9640 11830
rect 9588 11766 9640 11772
rect 9496 11688 9548 11694
rect 9496 11630 9548 11636
rect 9956 11688 10008 11694
rect 9956 11630 10008 11636
rect 9404 11620 9456 11626
rect 9404 11562 9456 11568
rect 9416 10130 9444 11562
rect 9496 11212 9548 11218
rect 9496 11154 9548 11160
rect 9404 10124 9456 10130
rect 9404 10066 9456 10072
rect 9312 9716 9364 9722
rect 9312 9658 9364 9664
rect 9036 8288 9088 8294
rect 9036 8230 9088 8236
rect 9048 7342 9076 8230
rect 9312 7744 9364 7750
rect 9312 7686 9364 7692
rect 9324 7478 9352 7686
rect 9312 7472 9364 7478
rect 9312 7414 9364 7420
rect 9036 7336 9088 7342
rect 9036 7278 9088 7284
rect 9048 5710 9076 7278
rect 9312 6996 9364 7002
rect 9312 6938 9364 6944
rect 9036 5704 9088 5710
rect 9036 5646 9088 5652
rect 9220 4140 9272 4146
rect 9220 4082 9272 4088
rect 8944 3188 8996 3194
rect 8944 3130 8996 3136
rect 8852 2916 8904 2922
rect 8852 2858 8904 2864
rect 8864 800 8892 2858
rect 9232 800 9260 4082
rect 9324 3942 9352 6938
rect 9508 5098 9536 11154
rect 9680 9988 9732 9994
rect 9680 9930 9732 9936
rect 9692 9178 9720 9930
rect 9968 9518 9996 11630
rect 10048 11212 10100 11218
rect 10048 11154 10100 11160
rect 9956 9512 10008 9518
rect 9956 9454 10008 9460
rect 9772 9444 9824 9450
rect 9772 9386 9824 9392
rect 9680 9172 9732 9178
rect 9680 9114 9732 9120
rect 9588 5636 9640 5642
rect 9588 5578 9640 5584
rect 9496 5092 9548 5098
rect 9496 5034 9548 5040
rect 9600 4554 9628 5578
rect 9784 4758 9812 9386
rect 10060 9330 10088 11154
rect 9968 9302 10088 9330
rect 9968 6746 9996 9302
rect 10244 8480 10272 14214
rect 10336 13258 10364 14758
rect 10324 13252 10376 13258
rect 10324 13194 10376 13200
rect 10428 12434 10456 16238
rect 10508 13252 10560 13258
rect 10508 13194 10560 13200
rect 10060 8452 10272 8480
rect 10336 12406 10456 12434
rect 10060 6866 10088 8452
rect 10336 8378 10364 12406
rect 10520 10742 10548 13194
rect 10508 10736 10560 10742
rect 10508 10678 10560 10684
rect 10520 10062 10548 10678
rect 10508 10056 10560 10062
rect 10508 9998 10560 10004
rect 10416 9920 10468 9926
rect 10416 9862 10468 9868
rect 10428 8974 10456 9862
rect 10520 9722 10548 9998
rect 10508 9716 10560 9722
rect 10508 9658 10560 9664
rect 10600 9512 10652 9518
rect 10600 9454 10652 9460
rect 10416 8968 10468 8974
rect 10416 8910 10468 8916
rect 10612 8634 10640 9454
rect 10600 8628 10652 8634
rect 10600 8570 10652 8576
rect 10416 8560 10468 8566
rect 10416 8502 10468 8508
rect 10152 8350 10364 8378
rect 10048 6860 10100 6866
rect 10048 6802 10100 6808
rect 9968 6718 10088 6746
rect 9772 4752 9824 4758
rect 9772 4694 9824 4700
rect 9956 4616 10008 4622
rect 9770 4584 9826 4593
rect 9588 4548 9640 4554
rect 9956 4558 10008 4564
rect 9770 4519 9826 4528
rect 9588 4490 9640 4496
rect 9312 3936 9364 3942
rect 9312 3878 9364 3884
rect 9784 3602 9812 4519
rect 9968 3942 9996 4558
rect 9956 3936 10008 3942
rect 9956 3878 10008 3884
rect 9772 3596 9824 3602
rect 9772 3538 9824 3544
rect 9588 3528 9640 3534
rect 9588 3470 9640 3476
rect 9312 3392 9364 3398
rect 9312 3334 9364 3340
rect 9324 3126 9352 3334
rect 9312 3120 9364 3126
rect 9312 3062 9364 3068
rect 9600 800 9628 3470
rect 9772 3120 9824 3126
rect 9770 3088 9772 3097
rect 9824 3088 9826 3097
rect 9770 3023 9826 3032
rect 9968 800 9996 3878
rect 10060 2650 10088 6718
rect 10152 3670 10180 8350
rect 10324 8288 10376 8294
rect 10324 8230 10376 8236
rect 10336 8090 10364 8230
rect 10324 8084 10376 8090
rect 10324 8026 10376 8032
rect 10336 7886 10364 8026
rect 10324 7880 10376 7886
rect 10324 7822 10376 7828
rect 10428 7528 10456 8502
rect 10704 7562 10732 16390
rect 10796 12434 10824 18702
rect 10876 17876 10928 17882
rect 10876 17818 10928 17824
rect 10888 17678 10916 17818
rect 11072 17814 11100 25094
rect 11164 24886 11192 25638
rect 11152 24880 11204 24886
rect 11152 24822 11204 24828
rect 11256 24818 11284 26318
rect 11532 25906 11560 26930
rect 12084 26586 12112 27406
rect 12072 26580 12124 26586
rect 12072 26522 12124 26528
rect 11520 25900 11572 25906
rect 11520 25842 11572 25848
rect 11244 24812 11296 24818
rect 11244 24754 11296 24760
rect 11152 24744 11204 24750
rect 11152 24686 11204 24692
rect 11164 24070 11192 24686
rect 11336 24132 11388 24138
rect 11336 24074 11388 24080
rect 11152 24064 11204 24070
rect 11152 24006 11204 24012
rect 11164 21486 11192 24006
rect 11348 23526 11376 24074
rect 11336 23520 11388 23526
rect 11336 23462 11388 23468
rect 11244 21888 11296 21894
rect 11244 21830 11296 21836
rect 11152 21480 11204 21486
rect 11152 21422 11204 21428
rect 11164 21010 11192 21422
rect 11152 21004 11204 21010
rect 11152 20946 11204 20952
rect 11152 19304 11204 19310
rect 11152 19246 11204 19252
rect 11164 18358 11192 19246
rect 11256 18698 11284 21830
rect 11428 20868 11480 20874
rect 11428 20810 11480 20816
rect 11440 20602 11468 20810
rect 11428 20596 11480 20602
rect 11428 20538 11480 20544
rect 11336 19168 11388 19174
rect 11336 19110 11388 19116
rect 11348 18970 11376 19110
rect 11336 18964 11388 18970
rect 11336 18906 11388 18912
rect 11532 18834 11560 25842
rect 11704 25696 11756 25702
rect 11704 25638 11756 25644
rect 11716 22030 11744 25638
rect 12084 25362 12112 26522
rect 12072 25356 12124 25362
rect 12072 25298 12124 25304
rect 12176 25226 12204 28970
rect 12440 28960 12492 28966
rect 12440 28902 12492 28908
rect 12452 28626 12480 28902
rect 12440 28620 12492 28626
rect 12440 28562 12492 28568
rect 12544 27588 12572 29650
rect 13372 29306 13400 31894
rect 13464 29306 13492 32166
rect 14280 31748 14332 31754
rect 14280 31690 14332 31696
rect 13912 31136 13964 31142
rect 13912 31078 13964 31084
rect 13728 30048 13780 30054
rect 13728 29990 13780 29996
rect 13544 29504 13596 29510
rect 13544 29446 13596 29452
rect 13360 29300 13412 29306
rect 13360 29242 13412 29248
rect 13452 29300 13504 29306
rect 13452 29242 13504 29248
rect 12624 29164 12676 29170
rect 12624 29106 12676 29112
rect 12360 27560 12572 27588
rect 12256 27124 12308 27130
rect 12256 27066 12308 27072
rect 12268 26790 12296 27066
rect 12360 26926 12388 27560
rect 12636 27520 12664 29106
rect 12950 28860 13258 28869
rect 12950 28858 12956 28860
rect 13012 28858 13036 28860
rect 13092 28858 13116 28860
rect 13172 28858 13196 28860
rect 13252 28858 13258 28860
rect 13012 28806 13014 28858
rect 13194 28806 13196 28858
rect 12950 28804 12956 28806
rect 13012 28804 13036 28806
rect 13092 28804 13116 28806
rect 13172 28804 13196 28806
rect 13252 28804 13258 28806
rect 12950 28795 13258 28804
rect 13556 28694 13584 29446
rect 13740 29170 13768 29990
rect 13728 29164 13780 29170
rect 13728 29106 13780 29112
rect 13924 29102 13952 31078
rect 14292 30666 14320 31690
rect 14280 30660 14332 30666
rect 14280 30602 14332 30608
rect 14372 30252 14424 30258
rect 14372 30194 14424 30200
rect 14384 29850 14412 30194
rect 14556 30048 14608 30054
rect 14556 29990 14608 29996
rect 14372 29844 14424 29850
rect 14372 29786 14424 29792
rect 14568 29306 14596 29990
rect 14832 29572 14884 29578
rect 14832 29514 14884 29520
rect 14556 29300 14608 29306
rect 14556 29242 14608 29248
rect 13912 29096 13964 29102
rect 13912 29038 13964 29044
rect 13636 29028 13688 29034
rect 13636 28970 13688 28976
rect 13544 28688 13596 28694
rect 13544 28630 13596 28636
rect 13084 28552 13136 28558
rect 13084 28494 13136 28500
rect 13096 28218 13124 28494
rect 13452 28416 13504 28422
rect 13452 28358 13504 28364
rect 12716 28212 12768 28218
rect 12716 28154 12768 28160
rect 13084 28212 13136 28218
rect 13084 28154 13136 28160
rect 12452 27492 12664 27520
rect 12348 26920 12400 26926
rect 12348 26862 12400 26868
rect 12256 26784 12308 26790
rect 12256 26726 12308 26732
rect 12360 25906 12388 26862
rect 12348 25900 12400 25906
rect 12348 25842 12400 25848
rect 12256 25288 12308 25294
rect 12256 25230 12308 25236
rect 12164 25220 12216 25226
rect 12164 25162 12216 25168
rect 12072 25152 12124 25158
rect 12072 25094 12124 25100
rect 11888 23588 11940 23594
rect 11888 23530 11940 23536
rect 11796 22636 11848 22642
rect 11796 22578 11848 22584
rect 11704 22024 11756 22030
rect 11704 21966 11756 21972
rect 11612 21888 11664 21894
rect 11612 21830 11664 21836
rect 11520 18828 11572 18834
rect 11520 18770 11572 18776
rect 11244 18692 11296 18698
rect 11244 18634 11296 18640
rect 11520 18420 11572 18426
rect 11520 18362 11572 18368
rect 11152 18352 11204 18358
rect 11152 18294 11204 18300
rect 11164 17898 11192 18294
rect 11532 18086 11560 18362
rect 11520 18080 11572 18086
rect 11520 18022 11572 18028
rect 11164 17882 11284 17898
rect 11164 17876 11296 17882
rect 11164 17870 11244 17876
rect 11060 17808 11112 17814
rect 11060 17750 11112 17756
rect 10876 17672 10928 17678
rect 11060 17672 11112 17678
rect 10876 17614 10928 17620
rect 10980 17632 11060 17660
rect 10980 16454 11008 17632
rect 11060 17614 11112 17620
rect 11164 17066 11192 17870
rect 11244 17818 11296 17824
rect 11336 17808 11388 17814
rect 11336 17750 11388 17756
rect 11244 17604 11296 17610
rect 11244 17546 11296 17552
rect 11152 17060 11204 17066
rect 11152 17002 11204 17008
rect 11164 16794 11192 17002
rect 11152 16788 11204 16794
rect 11152 16730 11204 16736
rect 11256 16658 11284 17546
rect 11244 16652 11296 16658
rect 11244 16594 11296 16600
rect 11060 16584 11112 16590
rect 11060 16526 11112 16532
rect 10968 16448 11020 16454
rect 10968 16390 11020 16396
rect 11072 16250 11100 16526
rect 11060 16244 11112 16250
rect 11060 16186 11112 16192
rect 11256 15570 11284 16594
rect 11244 15564 11296 15570
rect 11244 15506 11296 15512
rect 11348 15162 11376 17750
rect 11520 17536 11572 17542
rect 11520 17478 11572 17484
rect 11532 16182 11560 17478
rect 11624 17338 11652 21830
rect 11808 21536 11836 22578
rect 11900 21706 11928 23530
rect 12084 22094 12112 25094
rect 12268 24954 12296 25230
rect 12256 24948 12308 24954
rect 12256 24890 12308 24896
rect 12348 24744 12400 24750
rect 12348 24686 12400 24692
rect 12360 24410 12388 24686
rect 12348 24404 12400 24410
rect 12348 24346 12400 24352
rect 12348 22976 12400 22982
rect 12348 22918 12400 22924
rect 11992 22066 12112 22094
rect 11992 22030 12020 22066
rect 11980 22024 12032 22030
rect 11980 21966 12032 21972
rect 11900 21678 12112 21706
rect 11808 21508 12020 21536
rect 11796 21412 11848 21418
rect 11796 21354 11848 21360
rect 11704 20460 11756 20466
rect 11704 20402 11756 20408
rect 11716 19922 11744 20402
rect 11704 19916 11756 19922
rect 11704 19858 11756 19864
rect 11704 18624 11756 18630
rect 11704 18566 11756 18572
rect 11716 18426 11744 18566
rect 11704 18420 11756 18426
rect 11704 18362 11756 18368
rect 11612 17332 11664 17338
rect 11612 17274 11664 17280
rect 11704 17196 11756 17202
rect 11704 17138 11756 17144
rect 11612 16244 11664 16250
rect 11612 16186 11664 16192
rect 11520 16176 11572 16182
rect 11520 16118 11572 16124
rect 11624 16114 11652 16186
rect 11612 16108 11664 16114
rect 11612 16050 11664 16056
rect 11336 15156 11388 15162
rect 11336 15098 11388 15104
rect 10968 15020 11020 15026
rect 10968 14962 11020 14968
rect 10980 14278 11008 14962
rect 11348 14414 11376 15098
rect 11520 15088 11572 15094
rect 11520 15030 11572 15036
rect 11428 14884 11480 14890
rect 11428 14826 11480 14832
rect 11336 14408 11388 14414
rect 11336 14350 11388 14356
rect 10968 14272 11020 14278
rect 10968 14214 11020 14220
rect 11348 13326 11376 14350
rect 11336 13320 11388 13326
rect 11336 13262 11388 13268
rect 11060 13184 11112 13190
rect 11060 13126 11112 13132
rect 10796 12406 10916 12434
rect 10784 12300 10836 12306
rect 10784 12242 10836 12248
rect 10796 11694 10824 12242
rect 10888 12170 10916 12406
rect 10876 12164 10928 12170
rect 10876 12106 10928 12112
rect 11072 11898 11100 13126
rect 11440 12442 11468 14826
rect 11428 12436 11480 12442
rect 11428 12378 11480 12384
rect 11532 11898 11560 15030
rect 11716 14618 11744 17138
rect 11704 14612 11756 14618
rect 11704 14554 11756 14560
rect 11704 13388 11756 13394
rect 11704 13330 11756 13336
rect 11612 12776 11664 12782
rect 11612 12718 11664 12724
rect 11624 12646 11652 12718
rect 11612 12640 11664 12646
rect 11612 12582 11664 12588
rect 11060 11892 11112 11898
rect 11060 11834 11112 11840
rect 11520 11892 11572 11898
rect 11520 11834 11572 11840
rect 11072 11694 11100 11834
rect 11624 11778 11652 12582
rect 11428 11756 11480 11762
rect 11428 11698 11480 11704
rect 11532 11750 11652 11778
rect 10784 11688 10836 11694
rect 10784 11630 10836 11636
rect 11060 11688 11112 11694
rect 11060 11630 11112 11636
rect 10796 11354 10824 11630
rect 11244 11552 11296 11558
rect 11244 11494 11296 11500
rect 10784 11348 10836 11354
rect 10784 11290 10836 11296
rect 10796 11082 10824 11290
rect 10876 11144 10928 11150
rect 10876 11086 10928 11092
rect 10784 11076 10836 11082
rect 10784 11018 10836 11024
rect 10796 10810 10824 11018
rect 10784 10804 10836 10810
rect 10784 10746 10836 10752
rect 10888 10713 10916 11086
rect 11256 10849 11284 11494
rect 11336 11008 11388 11014
rect 11336 10950 11388 10956
rect 11242 10840 11298 10849
rect 11242 10775 11298 10784
rect 10874 10704 10930 10713
rect 10874 10639 10930 10648
rect 11348 10130 11376 10950
rect 11440 10810 11468 11698
rect 11428 10804 11480 10810
rect 11428 10746 11480 10752
rect 11060 10124 11112 10130
rect 11060 10066 11112 10072
rect 11336 10124 11388 10130
rect 11336 10066 11388 10072
rect 11072 9382 11100 10066
rect 11532 9654 11560 11750
rect 11520 9648 11572 9654
rect 11520 9590 11572 9596
rect 11716 9586 11744 13330
rect 11808 11218 11836 21354
rect 11992 16998 12020 21508
rect 12084 17610 12112 21678
rect 12360 19854 12388 22918
rect 12452 22234 12480 27492
rect 12728 27402 12756 28154
rect 13464 28082 13492 28358
rect 13452 28076 13504 28082
rect 13452 28018 13504 28024
rect 12808 27872 12860 27878
rect 12808 27814 12860 27820
rect 12716 27396 12768 27402
rect 12716 27338 12768 27344
rect 12728 26790 12756 27338
rect 12716 26784 12768 26790
rect 12716 26726 12768 26732
rect 12532 26308 12584 26314
rect 12532 26250 12584 26256
rect 12440 22228 12492 22234
rect 12440 22170 12492 22176
rect 12440 22092 12492 22098
rect 12440 22034 12492 22040
rect 12348 19848 12400 19854
rect 12348 19790 12400 19796
rect 12452 17814 12480 22034
rect 12544 21894 12572 26250
rect 12728 25974 12756 26726
rect 12820 26382 12848 27814
rect 12950 27772 13258 27781
rect 12950 27770 12956 27772
rect 13012 27770 13036 27772
rect 13092 27770 13116 27772
rect 13172 27770 13196 27772
rect 13252 27770 13258 27772
rect 13012 27718 13014 27770
rect 13194 27718 13196 27770
rect 12950 27716 12956 27718
rect 13012 27716 13036 27718
rect 13092 27716 13116 27718
rect 13172 27716 13196 27718
rect 13252 27716 13258 27718
rect 12950 27707 13258 27716
rect 12950 26684 13258 26693
rect 12950 26682 12956 26684
rect 13012 26682 13036 26684
rect 13092 26682 13116 26684
rect 13172 26682 13196 26684
rect 13252 26682 13258 26684
rect 13012 26630 13014 26682
rect 13194 26630 13196 26682
rect 12950 26628 12956 26630
rect 13012 26628 13036 26630
rect 13092 26628 13116 26630
rect 13172 26628 13196 26630
rect 13252 26628 13258 26630
rect 12950 26619 13258 26628
rect 12900 26512 12952 26518
rect 12900 26454 12952 26460
rect 12808 26376 12860 26382
rect 12808 26318 12860 26324
rect 12912 26042 12940 26454
rect 13464 26450 13492 28018
rect 13452 26444 13504 26450
rect 13452 26386 13504 26392
rect 13648 26314 13676 28970
rect 13924 28762 13952 29038
rect 13912 28756 13964 28762
rect 13912 28698 13964 28704
rect 14740 28416 14792 28422
rect 14740 28358 14792 28364
rect 14752 28218 14780 28358
rect 14844 28218 14872 29514
rect 14936 29238 14964 41386
rect 15476 31408 15528 31414
rect 15476 31350 15528 31356
rect 15488 31142 15516 31350
rect 15476 31136 15528 31142
rect 15476 31078 15528 31084
rect 15488 30734 15516 31078
rect 15476 30728 15528 30734
rect 15476 30670 15528 30676
rect 15108 30660 15160 30666
rect 15108 30602 15160 30608
rect 15120 29714 15148 30602
rect 15108 29708 15160 29714
rect 15108 29650 15160 29656
rect 15488 29510 15516 30670
rect 15200 29504 15252 29510
rect 15200 29446 15252 29452
rect 15476 29504 15528 29510
rect 15476 29446 15528 29452
rect 14924 29232 14976 29238
rect 14924 29174 14976 29180
rect 15212 28948 15240 29446
rect 15764 29170 15792 45018
rect 16040 31754 16068 50458
rect 16120 46980 16172 46986
rect 16120 46922 16172 46928
rect 16132 35834 16160 46922
rect 16304 46504 16356 46510
rect 16304 46446 16356 46452
rect 16120 35828 16172 35834
rect 16120 35770 16172 35776
rect 16316 35698 16344 46446
rect 16856 41472 16908 41478
rect 16856 41414 16908 41420
rect 16960 41414 16988 52430
rect 17144 45898 17172 53926
rect 17950 53340 18258 53349
rect 17950 53338 17956 53340
rect 18012 53338 18036 53340
rect 18092 53338 18116 53340
rect 18172 53338 18196 53340
rect 18252 53338 18258 53340
rect 18012 53286 18014 53338
rect 18194 53286 18196 53338
rect 17950 53284 17956 53286
rect 18012 53284 18036 53286
rect 18092 53284 18116 53286
rect 18172 53284 18196 53286
rect 18252 53284 18258 53286
rect 17950 53275 18258 53284
rect 17950 52252 18258 52261
rect 17950 52250 17956 52252
rect 18012 52250 18036 52252
rect 18092 52250 18116 52252
rect 18172 52250 18196 52252
rect 18252 52250 18258 52252
rect 18012 52198 18014 52250
rect 18194 52198 18196 52250
rect 17950 52196 17956 52198
rect 18012 52196 18036 52198
rect 18092 52196 18116 52198
rect 18172 52196 18196 52198
rect 18252 52196 18258 52198
rect 17950 52187 18258 52196
rect 17950 51164 18258 51173
rect 17950 51162 17956 51164
rect 18012 51162 18036 51164
rect 18092 51162 18116 51164
rect 18172 51162 18196 51164
rect 18252 51162 18258 51164
rect 18012 51110 18014 51162
rect 18194 51110 18196 51162
rect 17950 51108 17956 51110
rect 18012 51108 18036 51110
rect 18092 51108 18116 51110
rect 18172 51108 18196 51110
rect 18252 51108 18258 51110
rect 17950 51099 18258 51108
rect 17224 50448 17276 50454
rect 17224 50390 17276 50396
rect 17132 45892 17184 45898
rect 17132 45834 17184 45840
rect 17236 45554 17264 50390
rect 17950 50076 18258 50085
rect 17950 50074 17956 50076
rect 18012 50074 18036 50076
rect 18092 50074 18116 50076
rect 18172 50074 18196 50076
rect 18252 50074 18258 50076
rect 18012 50022 18014 50074
rect 18194 50022 18196 50074
rect 17950 50020 17956 50022
rect 18012 50020 18036 50022
rect 18092 50020 18116 50022
rect 18172 50020 18196 50022
rect 18252 50020 18258 50022
rect 17950 50011 18258 50020
rect 17950 48988 18258 48997
rect 17950 48986 17956 48988
rect 18012 48986 18036 48988
rect 18092 48986 18116 48988
rect 18172 48986 18196 48988
rect 18252 48986 18258 48988
rect 18012 48934 18014 48986
rect 18194 48934 18196 48986
rect 17950 48932 17956 48934
rect 18012 48932 18036 48934
rect 18092 48932 18116 48934
rect 18172 48932 18196 48934
rect 18252 48932 18258 48934
rect 17950 48923 18258 48932
rect 17592 48000 17644 48006
rect 17592 47942 17644 47948
rect 17500 45892 17552 45898
rect 17500 45834 17552 45840
rect 17144 45526 17264 45554
rect 16672 38344 16724 38350
rect 16672 38286 16724 38292
rect 16304 35692 16356 35698
rect 16304 35634 16356 35640
rect 16580 34468 16632 34474
rect 16580 34410 16632 34416
rect 16592 33862 16620 34410
rect 16580 33856 16632 33862
rect 16580 33798 16632 33804
rect 15948 31726 16068 31754
rect 15844 30252 15896 30258
rect 15844 30194 15896 30200
rect 15384 29164 15436 29170
rect 15384 29106 15436 29112
rect 15752 29164 15804 29170
rect 15752 29106 15804 29112
rect 15120 28920 15240 28948
rect 15120 28694 15148 28920
rect 15108 28688 15160 28694
rect 15108 28630 15160 28636
rect 14740 28212 14792 28218
rect 14740 28154 14792 28160
rect 14832 28212 14884 28218
rect 14832 28154 14884 28160
rect 14832 27940 14884 27946
rect 14832 27882 14884 27888
rect 14004 27872 14056 27878
rect 14004 27814 14056 27820
rect 14016 26926 14044 27814
rect 14648 27668 14700 27674
rect 14648 27610 14700 27616
rect 14660 27062 14688 27610
rect 14648 27056 14700 27062
rect 14648 26998 14700 27004
rect 14004 26920 14056 26926
rect 14004 26862 14056 26868
rect 14096 26852 14148 26858
rect 14096 26794 14148 26800
rect 14004 26580 14056 26586
rect 14004 26522 14056 26528
rect 13636 26308 13688 26314
rect 13636 26250 13688 26256
rect 12900 26036 12952 26042
rect 12900 25978 12952 25984
rect 12716 25968 12768 25974
rect 12768 25916 12848 25922
rect 12716 25910 12848 25916
rect 12728 25894 12848 25910
rect 12624 25832 12676 25838
rect 12624 25774 12676 25780
rect 12716 25832 12768 25838
rect 12716 25774 12768 25780
rect 12636 25498 12664 25774
rect 12624 25492 12676 25498
rect 12624 25434 12676 25440
rect 12728 25362 12756 25774
rect 12716 25356 12768 25362
rect 12716 25298 12768 25304
rect 12820 25242 12848 25894
rect 14016 25838 14044 26522
rect 14004 25832 14056 25838
rect 14004 25774 14056 25780
rect 14108 25702 14136 26794
rect 14280 26784 14332 26790
rect 14280 26726 14332 26732
rect 14372 26784 14424 26790
rect 14372 26726 14424 26732
rect 14292 26382 14320 26726
rect 14280 26376 14332 26382
rect 14280 26318 14332 26324
rect 14096 25696 14148 25702
rect 14096 25638 14148 25644
rect 12950 25596 13258 25605
rect 12950 25594 12956 25596
rect 13012 25594 13036 25596
rect 13092 25594 13116 25596
rect 13172 25594 13196 25596
rect 13252 25594 13258 25596
rect 13012 25542 13014 25594
rect 13194 25542 13196 25594
rect 12950 25540 12956 25542
rect 13012 25540 13036 25542
rect 13092 25540 13116 25542
rect 13172 25540 13196 25542
rect 13252 25540 13258 25542
rect 12950 25531 13258 25540
rect 12728 25214 12848 25242
rect 13452 25288 13504 25294
rect 13452 25230 13504 25236
rect 12728 24886 12756 25214
rect 12716 24880 12768 24886
rect 12716 24822 12768 24828
rect 12728 24410 12756 24822
rect 13464 24614 13492 25230
rect 13452 24608 13504 24614
rect 13452 24550 13504 24556
rect 13544 24608 13596 24614
rect 13544 24550 13596 24556
rect 14004 24608 14056 24614
rect 14004 24550 14056 24556
rect 12950 24508 13258 24517
rect 12950 24506 12956 24508
rect 13012 24506 13036 24508
rect 13092 24506 13116 24508
rect 13172 24506 13196 24508
rect 13252 24506 13258 24508
rect 13012 24454 13014 24506
rect 13194 24454 13196 24506
rect 12950 24452 12956 24454
rect 13012 24452 13036 24454
rect 13092 24452 13116 24454
rect 13172 24452 13196 24454
rect 13252 24452 13258 24454
rect 12950 24443 13258 24452
rect 12716 24404 12768 24410
rect 12716 24346 12768 24352
rect 12728 23866 12756 24346
rect 12716 23860 12768 23866
rect 12716 23802 12768 23808
rect 12624 23724 12676 23730
rect 12624 23666 12676 23672
rect 12532 21888 12584 21894
rect 12532 21830 12584 21836
rect 12636 21570 12664 23666
rect 12728 23526 12756 23802
rect 13464 23662 13492 24550
rect 13452 23656 13504 23662
rect 13452 23598 13504 23604
rect 12716 23520 12768 23526
rect 12716 23462 12768 23468
rect 12950 23420 13258 23429
rect 12950 23418 12956 23420
rect 13012 23418 13036 23420
rect 13092 23418 13116 23420
rect 13172 23418 13196 23420
rect 13252 23418 13258 23420
rect 13012 23366 13014 23418
rect 13194 23366 13196 23418
rect 12950 23364 12956 23366
rect 13012 23364 13036 23366
rect 13092 23364 13116 23366
rect 13172 23364 13196 23366
rect 13252 23364 13258 23366
rect 12950 23355 13258 23364
rect 13556 22522 13584 24550
rect 13372 22506 13584 22522
rect 13728 22568 13780 22574
rect 13728 22510 13780 22516
rect 13360 22500 13584 22506
rect 13412 22494 13584 22500
rect 13360 22442 13412 22448
rect 12808 22432 12860 22438
rect 12808 22374 12860 22380
rect 12716 22228 12768 22234
rect 12716 22170 12768 22176
rect 12544 21542 12664 21570
rect 12728 21554 12756 22170
rect 12820 22098 12848 22374
rect 12950 22332 13258 22341
rect 12950 22330 12956 22332
rect 13012 22330 13036 22332
rect 13092 22330 13116 22332
rect 13172 22330 13196 22332
rect 13252 22330 13258 22332
rect 13012 22278 13014 22330
rect 13194 22278 13196 22330
rect 12950 22276 12956 22278
rect 13012 22276 13036 22278
rect 13092 22276 13116 22278
rect 13172 22276 13196 22278
rect 13252 22276 13258 22278
rect 12950 22267 13258 22276
rect 13740 22234 13768 22510
rect 13728 22228 13780 22234
rect 13728 22170 13780 22176
rect 12808 22092 12860 22098
rect 14016 22094 14044 24550
rect 14108 24206 14136 25638
rect 14384 24818 14412 26726
rect 14660 26450 14688 26998
rect 14740 26988 14792 26994
rect 14740 26930 14792 26936
rect 14648 26444 14700 26450
rect 14648 26386 14700 26392
rect 14464 26240 14516 26246
rect 14464 26182 14516 26188
rect 14372 24812 14424 24818
rect 14372 24754 14424 24760
rect 14096 24200 14148 24206
rect 14096 24142 14148 24148
rect 14476 23866 14504 26182
rect 14464 23860 14516 23866
rect 14464 23802 14516 23808
rect 14648 23520 14700 23526
rect 14648 23462 14700 23468
rect 14464 22568 14516 22574
rect 14464 22510 14516 22516
rect 12808 22034 12860 22040
rect 13832 22066 14044 22094
rect 13360 21956 13412 21962
rect 13360 21898 13412 21904
rect 12716 21548 12768 21554
rect 12544 18766 12572 21542
rect 12768 21508 12848 21536
rect 12716 21490 12768 21496
rect 12624 21480 12676 21486
rect 12624 21422 12676 21428
rect 12636 20398 12664 21422
rect 12716 21344 12768 21350
rect 12716 21286 12768 21292
rect 12728 20534 12756 21286
rect 12820 21146 12848 21508
rect 12950 21244 13258 21253
rect 12950 21242 12956 21244
rect 13012 21242 13036 21244
rect 13092 21242 13116 21244
rect 13172 21242 13196 21244
rect 13252 21242 13258 21244
rect 13012 21190 13014 21242
rect 13194 21190 13196 21242
rect 12950 21188 12956 21190
rect 13012 21188 13036 21190
rect 13092 21188 13116 21190
rect 13172 21188 13196 21190
rect 13252 21188 13258 21190
rect 12950 21179 13258 21188
rect 12808 21140 12860 21146
rect 12808 21082 12860 21088
rect 13372 21010 13400 21898
rect 13636 21616 13688 21622
rect 13636 21558 13688 21564
rect 13544 21140 13596 21146
rect 13544 21082 13596 21088
rect 13360 21004 13412 21010
rect 13360 20946 13412 20952
rect 13360 20868 13412 20874
rect 13360 20810 13412 20816
rect 13372 20534 13400 20810
rect 13556 20618 13584 21082
rect 13648 20874 13676 21558
rect 13832 21486 13860 22066
rect 13820 21480 13872 21486
rect 13820 21422 13872 21428
rect 14096 21480 14148 21486
rect 14096 21422 14148 21428
rect 13636 20868 13688 20874
rect 13636 20810 13688 20816
rect 14108 20806 14136 21422
rect 14096 20800 14148 20806
rect 14096 20742 14148 20748
rect 13556 20590 13768 20618
rect 12716 20528 12768 20534
rect 12716 20470 12768 20476
rect 13360 20528 13412 20534
rect 13360 20470 13412 20476
rect 12624 20392 12676 20398
rect 12624 20334 12676 20340
rect 12636 19854 12664 20334
rect 12950 20156 13258 20165
rect 12950 20154 12956 20156
rect 13012 20154 13036 20156
rect 13092 20154 13116 20156
rect 13172 20154 13196 20156
rect 13252 20154 13258 20156
rect 13012 20102 13014 20154
rect 13194 20102 13196 20154
rect 12950 20100 12956 20102
rect 13012 20100 13036 20102
rect 13092 20100 13116 20102
rect 13172 20100 13196 20102
rect 13252 20100 13258 20102
rect 12950 20091 13258 20100
rect 12624 19848 12676 19854
rect 12624 19790 12676 19796
rect 12636 19446 12664 19790
rect 13372 19718 13400 20470
rect 13544 20392 13596 20398
rect 13544 20334 13596 20340
rect 13084 19712 13136 19718
rect 13084 19654 13136 19660
rect 13360 19712 13412 19718
rect 13360 19654 13412 19660
rect 12716 19508 12768 19514
rect 12716 19450 12768 19456
rect 12808 19508 12860 19514
rect 12808 19450 12860 19456
rect 12624 19440 12676 19446
rect 12624 19382 12676 19388
rect 12532 18760 12584 18766
rect 12532 18702 12584 18708
rect 12636 18698 12664 19382
rect 12624 18692 12676 18698
rect 12624 18634 12676 18640
rect 12532 18080 12584 18086
rect 12532 18022 12584 18028
rect 12164 17808 12216 17814
rect 12164 17750 12216 17756
rect 12440 17808 12492 17814
rect 12440 17750 12492 17756
rect 12176 17610 12204 17750
rect 12072 17604 12124 17610
rect 12072 17546 12124 17552
rect 12164 17604 12216 17610
rect 12164 17546 12216 17552
rect 12256 17264 12308 17270
rect 12256 17206 12308 17212
rect 12072 17196 12124 17202
rect 12072 17138 12124 17144
rect 11980 16992 12032 16998
rect 11980 16934 12032 16940
rect 11980 15564 12032 15570
rect 11980 15506 12032 15512
rect 11992 14482 12020 15506
rect 11980 14476 12032 14482
rect 11980 14418 12032 14424
rect 11992 13802 12020 14418
rect 11980 13796 12032 13802
rect 11980 13738 12032 13744
rect 11888 13728 11940 13734
rect 11888 13670 11940 13676
rect 11900 12345 11928 13670
rect 11980 12844 12032 12850
rect 11980 12786 12032 12792
rect 11886 12336 11942 12345
rect 11886 12271 11942 12280
rect 11888 11688 11940 11694
rect 11888 11630 11940 11636
rect 11900 11218 11928 11630
rect 11796 11212 11848 11218
rect 11796 11154 11848 11160
rect 11888 11212 11940 11218
rect 11888 11154 11940 11160
rect 11808 10810 11836 11154
rect 11796 10804 11848 10810
rect 11796 10746 11848 10752
rect 11888 9920 11940 9926
rect 11888 9862 11940 9868
rect 11704 9580 11756 9586
rect 11704 9522 11756 9528
rect 11060 9376 11112 9382
rect 11060 9318 11112 9324
rect 11072 8362 11100 9318
rect 11244 8968 11296 8974
rect 11244 8910 11296 8916
rect 11060 8356 11112 8362
rect 11060 8298 11112 8304
rect 10876 8084 10928 8090
rect 10876 8026 10928 8032
rect 10704 7534 10824 7562
rect 10888 7546 10916 8026
rect 10336 7500 10456 7528
rect 10232 6112 10284 6118
rect 10232 6054 10284 6060
rect 10244 5778 10272 6054
rect 10232 5772 10284 5778
rect 10232 5714 10284 5720
rect 10140 3664 10192 3670
rect 10140 3606 10192 3612
rect 10336 2854 10364 7500
rect 10414 6760 10470 6769
rect 10414 6695 10470 6704
rect 10428 4622 10456 6695
rect 10598 6216 10654 6225
rect 10598 6151 10654 6160
rect 10508 5296 10560 5302
rect 10508 5238 10560 5244
rect 10416 4616 10468 4622
rect 10416 4558 10468 4564
rect 10416 4072 10468 4078
rect 10416 4014 10468 4020
rect 10324 2848 10376 2854
rect 10324 2790 10376 2796
rect 10048 2644 10100 2650
rect 10048 2586 10100 2592
rect 10324 2304 10376 2310
rect 10324 2246 10376 2252
rect 10336 800 10364 2246
rect 10428 1902 10456 4014
rect 10520 3670 10548 5238
rect 10612 4146 10640 6151
rect 10600 4140 10652 4146
rect 10600 4082 10652 4088
rect 10508 3664 10560 3670
rect 10508 3606 10560 3612
rect 10600 3528 10652 3534
rect 10598 3496 10600 3505
rect 10652 3496 10654 3505
rect 10598 3431 10654 3440
rect 10692 2984 10744 2990
rect 10692 2926 10744 2932
rect 10416 1896 10468 1902
rect 10416 1838 10468 1844
rect 10704 800 10732 2926
rect 10796 2774 10824 7534
rect 10876 7540 10928 7546
rect 10876 7482 10928 7488
rect 10888 6322 10916 7482
rect 11072 7410 11100 8298
rect 11060 7404 11112 7410
rect 11060 7346 11112 7352
rect 11152 6724 11204 6730
rect 11152 6666 11204 6672
rect 11164 6458 11192 6666
rect 11152 6452 11204 6458
rect 11152 6394 11204 6400
rect 10876 6316 10928 6322
rect 10876 6258 10928 6264
rect 11256 5778 11284 8910
rect 11428 8900 11480 8906
rect 11428 8842 11480 8848
rect 11440 5930 11468 8842
rect 11518 7984 11574 7993
rect 11518 7919 11520 7928
rect 11572 7919 11574 7928
rect 11520 7890 11572 7896
rect 11612 6860 11664 6866
rect 11716 6848 11744 9522
rect 11900 8974 11928 9862
rect 11992 9110 12020 12786
rect 12084 12442 12112 17138
rect 12164 17128 12216 17134
rect 12164 17070 12216 17076
rect 12072 12436 12124 12442
rect 12072 12378 12124 12384
rect 12070 12336 12126 12345
rect 12070 12271 12072 12280
rect 12124 12271 12126 12280
rect 12072 12242 12124 12248
rect 12084 11694 12112 12242
rect 12176 11898 12204 17070
rect 12268 14074 12296 17206
rect 12348 17060 12400 17066
rect 12348 17002 12400 17008
rect 12360 16658 12388 17002
rect 12440 16788 12492 16794
rect 12440 16730 12492 16736
rect 12348 16652 12400 16658
rect 12348 16594 12400 16600
rect 12452 16454 12480 16730
rect 12440 16448 12492 16454
rect 12440 16390 12492 16396
rect 12440 16176 12492 16182
rect 12440 16118 12492 16124
rect 12452 15910 12480 16118
rect 12440 15904 12492 15910
rect 12440 15846 12492 15852
rect 12452 15570 12480 15846
rect 12440 15564 12492 15570
rect 12440 15506 12492 15512
rect 12348 14544 12400 14550
rect 12348 14486 12400 14492
rect 12256 14068 12308 14074
rect 12256 14010 12308 14016
rect 12360 13546 12388 14486
rect 12544 14464 12572 18022
rect 12636 16250 12664 18634
rect 12728 18426 12756 19450
rect 12716 18420 12768 18426
rect 12716 18362 12768 18368
rect 12820 17678 12848 19450
rect 13096 19446 13124 19654
rect 13084 19440 13136 19446
rect 13084 19382 13136 19388
rect 12950 19068 13258 19077
rect 12950 19066 12956 19068
rect 13012 19066 13036 19068
rect 13092 19066 13116 19068
rect 13172 19066 13196 19068
rect 13252 19066 13258 19068
rect 13012 19014 13014 19066
rect 13194 19014 13196 19066
rect 12950 19012 12956 19014
rect 13012 19012 13036 19014
rect 13092 19012 13116 19014
rect 13172 19012 13196 19014
rect 13252 19012 13258 19014
rect 12950 19003 13258 19012
rect 13452 18624 13504 18630
rect 13452 18566 13504 18572
rect 12950 17980 13258 17989
rect 12950 17978 12956 17980
rect 13012 17978 13036 17980
rect 13092 17978 13116 17980
rect 13172 17978 13196 17980
rect 13252 17978 13258 17980
rect 13012 17926 13014 17978
rect 13194 17926 13196 17978
rect 12950 17924 12956 17926
rect 13012 17924 13036 17926
rect 13092 17924 13116 17926
rect 13172 17924 13196 17926
rect 13252 17924 13258 17926
rect 12950 17915 13258 17924
rect 13464 17882 13492 18566
rect 13452 17876 13504 17882
rect 13452 17818 13504 17824
rect 12808 17672 12860 17678
rect 12808 17614 12860 17620
rect 12624 16244 12676 16250
rect 12624 16186 12676 16192
rect 12820 15570 12848 17614
rect 13452 17536 13504 17542
rect 13452 17478 13504 17484
rect 13360 17128 13412 17134
rect 13360 17070 13412 17076
rect 12950 16892 13258 16901
rect 12950 16890 12956 16892
rect 13012 16890 13036 16892
rect 13092 16890 13116 16892
rect 13172 16890 13196 16892
rect 13252 16890 13258 16892
rect 13012 16838 13014 16890
rect 13194 16838 13196 16890
rect 12950 16836 12956 16838
rect 13012 16836 13036 16838
rect 13092 16836 13116 16838
rect 13172 16836 13196 16838
rect 13252 16836 13258 16838
rect 12950 16827 13258 16836
rect 13372 16658 13400 17070
rect 13360 16652 13412 16658
rect 13360 16594 13412 16600
rect 13464 16046 13492 17478
rect 13556 17270 13584 20334
rect 13636 18624 13688 18630
rect 13636 18566 13688 18572
rect 13648 18426 13676 18566
rect 13636 18420 13688 18426
rect 13636 18362 13688 18368
rect 13636 18284 13688 18290
rect 13636 18226 13688 18232
rect 13544 17264 13596 17270
rect 13544 17206 13596 17212
rect 13544 16652 13596 16658
rect 13648 16640 13676 18226
rect 13740 17134 13768 20590
rect 13912 19440 13964 19446
rect 13912 19382 13964 19388
rect 13924 18290 13952 19382
rect 14096 19236 14148 19242
rect 14096 19178 14148 19184
rect 14108 18902 14136 19178
rect 14372 19168 14424 19174
rect 14372 19110 14424 19116
rect 14096 18896 14148 18902
rect 14096 18838 14148 18844
rect 14004 18624 14056 18630
rect 14004 18566 14056 18572
rect 13912 18284 13964 18290
rect 13912 18226 13964 18232
rect 13820 18148 13872 18154
rect 13820 18090 13872 18096
rect 13832 17814 13860 18090
rect 13820 17808 13872 17814
rect 13820 17750 13872 17756
rect 14016 17610 14044 18566
rect 14004 17604 14056 17610
rect 14004 17546 14056 17552
rect 13912 17536 13964 17542
rect 13912 17478 13964 17484
rect 13924 17338 13952 17478
rect 13912 17332 13964 17338
rect 13912 17274 13964 17280
rect 14016 17218 14044 17546
rect 13924 17190 14044 17218
rect 13728 17128 13780 17134
rect 13728 17070 13780 17076
rect 13648 16612 13768 16640
rect 13544 16594 13596 16600
rect 13556 16561 13584 16594
rect 13542 16552 13598 16561
rect 13542 16487 13598 16496
rect 13636 16516 13688 16522
rect 13636 16458 13688 16464
rect 13452 16040 13504 16046
rect 13452 15982 13504 15988
rect 13452 15904 13504 15910
rect 13452 15846 13504 15852
rect 12950 15804 13258 15813
rect 12950 15802 12956 15804
rect 13012 15802 13036 15804
rect 13092 15802 13116 15804
rect 13172 15802 13196 15804
rect 13252 15802 13258 15804
rect 13012 15750 13014 15802
rect 13194 15750 13196 15802
rect 12950 15748 12956 15750
rect 13012 15748 13036 15750
rect 13092 15748 13116 15750
rect 13172 15748 13196 15750
rect 13252 15748 13258 15750
rect 12950 15739 13258 15748
rect 12808 15564 12860 15570
rect 12808 15506 12860 15512
rect 12716 15360 12768 15366
rect 12716 15302 12768 15308
rect 13360 15360 13412 15366
rect 13360 15302 13412 15308
rect 12728 15162 12756 15302
rect 12716 15156 12768 15162
rect 12716 15098 12768 15104
rect 12624 15088 12676 15094
rect 12624 15030 12676 15036
rect 12268 13518 12388 13546
rect 12452 14436 12572 14464
rect 12164 11892 12216 11898
rect 12164 11834 12216 11840
rect 12268 11762 12296 13518
rect 12348 12640 12400 12646
rect 12348 12582 12400 12588
rect 12256 11756 12308 11762
rect 12256 11698 12308 11704
rect 12072 11688 12124 11694
rect 12072 11630 12124 11636
rect 12256 10804 12308 10810
rect 12256 10746 12308 10752
rect 12268 9738 12296 10746
rect 12360 10169 12388 12582
rect 12452 12306 12480 14436
rect 12532 14340 12584 14346
rect 12532 14282 12584 14288
rect 12440 12300 12492 12306
rect 12440 12242 12492 12248
rect 12440 12164 12492 12170
rect 12440 12106 12492 12112
rect 12452 11937 12480 12106
rect 12438 11928 12494 11937
rect 12438 11863 12494 11872
rect 12440 11756 12492 11762
rect 12440 11698 12492 11704
rect 12452 10198 12480 11698
rect 12544 10810 12572 14282
rect 12636 14006 12664 15030
rect 13372 14906 13400 15302
rect 13464 15026 13492 15846
rect 13452 15020 13504 15026
rect 13452 14962 13504 14968
rect 13542 14920 13598 14929
rect 13372 14890 13492 14906
rect 13372 14884 13504 14890
rect 13372 14878 13452 14884
rect 13542 14855 13598 14864
rect 13452 14826 13504 14832
rect 12950 14716 13258 14725
rect 12950 14714 12956 14716
rect 13012 14714 13036 14716
rect 13092 14714 13116 14716
rect 13172 14714 13196 14716
rect 13252 14714 13258 14716
rect 13012 14662 13014 14714
rect 13194 14662 13196 14714
rect 12950 14660 12956 14662
rect 13012 14660 13036 14662
rect 13092 14660 13116 14662
rect 13172 14660 13196 14662
rect 13252 14660 13258 14662
rect 12950 14651 13258 14660
rect 13464 14482 13492 14826
rect 13556 14822 13584 14855
rect 13544 14816 13596 14822
rect 13544 14758 13596 14764
rect 13452 14476 13504 14482
rect 13452 14418 13504 14424
rect 13556 14346 13584 14758
rect 13544 14340 13596 14346
rect 13544 14282 13596 14288
rect 12716 14272 12768 14278
rect 12716 14214 12768 14220
rect 12808 14272 12860 14278
rect 12808 14214 12860 14220
rect 12624 14000 12676 14006
rect 12624 13942 12676 13948
rect 12624 12912 12676 12918
rect 12624 12854 12676 12860
rect 12636 11354 12664 12854
rect 12624 11348 12676 11354
rect 12624 11290 12676 11296
rect 12624 11076 12676 11082
rect 12624 11018 12676 11024
rect 12532 10804 12584 10810
rect 12532 10746 12584 10752
rect 12636 10690 12664 11018
rect 12544 10662 12664 10690
rect 12440 10192 12492 10198
rect 12346 10160 12402 10169
rect 12440 10134 12492 10140
rect 12346 10095 12402 10104
rect 12268 9710 12388 9738
rect 12360 9466 12388 9710
rect 12438 9480 12494 9489
rect 12268 9438 12438 9466
rect 11980 9104 12032 9110
rect 11980 9046 12032 9052
rect 11888 8968 11940 8974
rect 11888 8910 11940 8916
rect 12268 8838 12296 9438
rect 12438 9415 12494 9424
rect 12360 9178 12480 9194
rect 12360 9172 12492 9178
rect 12360 9166 12440 9172
rect 12360 8906 12388 9166
rect 12440 9114 12492 9120
rect 12348 8900 12400 8906
rect 12348 8842 12400 8848
rect 12256 8832 12308 8838
rect 12256 8774 12308 8780
rect 12440 8832 12492 8838
rect 12440 8774 12492 8780
rect 11980 8424 12032 8430
rect 11794 8392 11850 8401
rect 11980 8366 12032 8372
rect 12164 8424 12216 8430
rect 12164 8366 12216 8372
rect 11794 8327 11850 8336
rect 11808 8090 11836 8327
rect 11796 8084 11848 8090
rect 11796 8026 11848 8032
rect 11992 7886 12020 8366
rect 11980 7880 12032 7886
rect 11980 7822 12032 7828
rect 12072 7404 12124 7410
rect 12072 7346 12124 7352
rect 11980 7200 12032 7206
rect 11980 7142 12032 7148
rect 11664 6820 11744 6848
rect 11612 6802 11664 6808
rect 11624 6254 11652 6802
rect 11992 6798 12020 7142
rect 11980 6792 12032 6798
rect 11980 6734 12032 6740
rect 11886 6352 11942 6361
rect 11704 6316 11756 6322
rect 11886 6287 11942 6296
rect 11704 6258 11756 6264
rect 11612 6248 11664 6254
rect 11612 6190 11664 6196
rect 11348 5902 11468 5930
rect 11716 5914 11744 6258
rect 11704 5908 11756 5914
rect 11244 5772 11296 5778
rect 11244 5714 11296 5720
rect 11152 5228 11204 5234
rect 11152 5170 11204 5176
rect 10968 5160 11020 5166
rect 10968 5102 11020 5108
rect 10980 4486 11008 5102
rect 10968 4480 11020 4486
rect 10968 4422 11020 4428
rect 11164 4282 11192 5170
rect 11152 4276 11204 4282
rect 11152 4218 11204 4224
rect 11150 3088 11206 3097
rect 11150 3023 11152 3032
rect 11204 3023 11206 3032
rect 11152 2994 11204 3000
rect 11164 2854 11192 2994
rect 11152 2848 11204 2854
rect 11152 2790 11204 2796
rect 10796 2746 10916 2774
rect 10888 2038 10916 2746
rect 10968 2372 11020 2378
rect 10968 2314 11020 2320
rect 10980 2258 11008 2314
rect 10980 2230 11100 2258
rect 10876 2032 10928 2038
rect 10876 1974 10928 1980
rect 11072 800 11100 2230
rect 11348 2106 11376 5902
rect 11704 5850 11756 5856
rect 11900 4690 11928 6287
rect 11992 6118 12020 6734
rect 11980 6112 12032 6118
rect 11980 6054 12032 6060
rect 11992 5574 12020 6054
rect 11980 5568 12032 5574
rect 11980 5510 12032 5516
rect 11888 4684 11940 4690
rect 11888 4626 11940 4632
rect 12084 4010 12112 7346
rect 12176 6186 12204 8366
rect 12348 7812 12400 7818
rect 12348 7754 12400 7760
rect 12360 7546 12388 7754
rect 12348 7540 12400 7546
rect 12348 7482 12400 7488
rect 12256 7336 12308 7342
rect 12256 7278 12308 7284
rect 12348 7336 12400 7342
rect 12348 7278 12400 7284
rect 12268 6322 12296 7278
rect 12256 6316 12308 6322
rect 12256 6258 12308 6264
rect 12164 6180 12216 6186
rect 12164 6122 12216 6128
rect 12360 5658 12388 7278
rect 12452 6866 12480 8774
rect 12440 6860 12492 6866
rect 12440 6802 12492 6808
rect 12268 5630 12388 5658
rect 12268 4078 12296 5630
rect 12348 5568 12400 5574
rect 12348 5510 12400 5516
rect 12256 4072 12308 4078
rect 12256 4014 12308 4020
rect 12072 4004 12124 4010
rect 12072 3946 12124 3952
rect 11612 3936 11664 3942
rect 11612 3878 11664 3884
rect 11624 3058 11652 3878
rect 12360 3534 12388 5510
rect 12348 3528 12400 3534
rect 12348 3470 12400 3476
rect 12544 3058 12572 10662
rect 12728 10266 12756 14214
rect 12820 12238 12848 14214
rect 13452 13932 13504 13938
rect 13452 13874 13504 13880
rect 12950 13628 13258 13637
rect 12950 13626 12956 13628
rect 13012 13626 13036 13628
rect 13092 13626 13116 13628
rect 13172 13626 13196 13628
rect 13252 13626 13258 13628
rect 13012 13574 13014 13626
rect 13194 13574 13196 13626
rect 12950 13572 12956 13574
rect 13012 13572 13036 13574
rect 13092 13572 13116 13574
rect 13172 13572 13196 13574
rect 13252 13572 13258 13574
rect 12950 13563 13258 13572
rect 13464 13274 13492 13874
rect 13544 13864 13596 13870
rect 13544 13806 13596 13812
rect 13556 13394 13584 13806
rect 13544 13388 13596 13394
rect 13544 13330 13596 13336
rect 13464 13246 13584 13274
rect 13452 13184 13504 13190
rect 13452 13126 13504 13132
rect 12992 12844 13044 12850
rect 12992 12786 13044 12792
rect 13360 12844 13412 12850
rect 13360 12786 13412 12792
rect 13004 12646 13032 12786
rect 12992 12640 13044 12646
rect 12992 12582 13044 12588
rect 12950 12540 13258 12549
rect 12950 12538 12956 12540
rect 13012 12538 13036 12540
rect 13092 12538 13116 12540
rect 13172 12538 13196 12540
rect 13252 12538 13258 12540
rect 13012 12486 13014 12538
rect 13194 12486 13196 12538
rect 12950 12484 12956 12486
rect 13012 12484 13036 12486
rect 13092 12484 13116 12486
rect 13172 12484 13196 12486
rect 13252 12484 13258 12486
rect 12950 12475 13258 12484
rect 12808 12232 12860 12238
rect 12808 12174 12860 12180
rect 13372 12102 13400 12786
rect 13360 12096 13412 12102
rect 13360 12038 13412 12044
rect 13268 11892 13320 11898
rect 13268 11834 13320 11840
rect 13280 11558 13308 11834
rect 13358 11792 13414 11801
rect 13358 11727 13414 11736
rect 12808 11552 12860 11558
rect 12808 11494 12860 11500
rect 13268 11552 13320 11558
rect 13268 11494 13320 11500
rect 12716 10260 12768 10266
rect 12716 10202 12768 10208
rect 12624 10056 12676 10062
rect 12624 9998 12676 10004
rect 12636 8430 12664 9998
rect 12820 8650 12848 11494
rect 12950 11452 13258 11461
rect 12950 11450 12956 11452
rect 13012 11450 13036 11452
rect 13092 11450 13116 11452
rect 13172 11450 13196 11452
rect 13252 11450 13258 11452
rect 13012 11398 13014 11450
rect 13194 11398 13196 11450
rect 12950 11396 12956 11398
rect 13012 11396 13036 11398
rect 13092 11396 13116 11398
rect 13172 11396 13196 11398
rect 13252 11396 13258 11398
rect 12950 11387 13258 11396
rect 12992 11348 13044 11354
rect 12992 11290 13044 11296
rect 12900 11280 12952 11286
rect 12900 11222 12952 11228
rect 12912 11082 12940 11222
rect 13004 11082 13032 11290
rect 12900 11076 12952 11082
rect 12900 11018 12952 11024
rect 12992 11076 13044 11082
rect 12992 11018 13044 11024
rect 13372 10606 13400 11727
rect 13464 11336 13492 13126
rect 13556 12073 13584 13246
rect 13648 12442 13676 16458
rect 13740 15162 13768 16612
rect 13924 15978 13952 17190
rect 14004 16788 14056 16794
rect 14004 16730 14056 16736
rect 13912 15972 13964 15978
rect 13912 15914 13964 15920
rect 13728 15156 13780 15162
rect 13728 15098 13780 15104
rect 14016 13682 14044 16730
rect 14096 16652 14148 16658
rect 14096 16594 14148 16600
rect 14108 16454 14136 16594
rect 14096 16448 14148 16454
rect 14096 16390 14148 16396
rect 13832 13654 14044 13682
rect 13728 12640 13780 12646
rect 13726 12608 13728 12617
rect 13780 12608 13782 12617
rect 13726 12543 13782 12552
rect 13636 12436 13688 12442
rect 13636 12378 13688 12384
rect 13636 12096 13688 12102
rect 13542 12064 13598 12073
rect 13636 12038 13688 12044
rect 13542 11999 13598 12008
rect 13464 11308 13584 11336
rect 13452 11212 13504 11218
rect 13452 11154 13504 11160
rect 13360 10600 13412 10606
rect 13360 10542 13412 10548
rect 12950 10364 13258 10373
rect 12950 10362 12956 10364
rect 13012 10362 13036 10364
rect 13092 10362 13116 10364
rect 13172 10362 13196 10364
rect 13252 10362 13258 10364
rect 13012 10310 13014 10362
rect 13194 10310 13196 10362
rect 12950 10308 12956 10310
rect 13012 10308 13036 10310
rect 13092 10308 13116 10310
rect 13172 10308 13196 10310
rect 13252 10308 13258 10310
rect 12950 10299 13258 10308
rect 13372 10130 13400 10542
rect 13360 10124 13412 10130
rect 13360 10066 13412 10072
rect 13268 9648 13320 9654
rect 13268 9590 13320 9596
rect 13280 9382 13308 9590
rect 13360 9512 13412 9518
rect 13360 9454 13412 9460
rect 13268 9376 13320 9382
rect 13268 9318 13320 9324
rect 12950 9276 13258 9285
rect 12950 9274 12956 9276
rect 13012 9274 13036 9276
rect 13092 9274 13116 9276
rect 13172 9274 13196 9276
rect 13252 9274 13258 9276
rect 13012 9222 13014 9274
rect 13194 9222 13196 9274
rect 12950 9220 12956 9222
rect 13012 9220 13036 9222
rect 13092 9220 13116 9222
rect 13172 9220 13196 9222
rect 13252 9220 13258 9222
rect 12950 9211 13258 9220
rect 12728 8622 12848 8650
rect 12624 8424 12676 8430
rect 12624 8366 12676 8372
rect 12636 3466 12664 8366
rect 12728 7546 12756 8622
rect 12808 8492 12860 8498
rect 12808 8434 12860 8440
rect 12820 7954 12848 8434
rect 12950 8188 13258 8197
rect 12950 8186 12956 8188
rect 13012 8186 13036 8188
rect 13092 8186 13116 8188
rect 13172 8186 13196 8188
rect 13252 8186 13258 8188
rect 13012 8134 13014 8186
rect 13194 8134 13196 8186
rect 12950 8132 12956 8134
rect 13012 8132 13036 8134
rect 13092 8132 13116 8134
rect 13172 8132 13196 8134
rect 13252 8132 13258 8134
rect 12950 8123 13258 8132
rect 12808 7948 12860 7954
rect 12808 7890 12860 7896
rect 12716 7540 12768 7546
rect 12716 7482 12768 7488
rect 12728 6934 12756 7482
rect 12820 7002 12848 7890
rect 13372 7886 13400 9454
rect 13464 9042 13492 11154
rect 13556 10996 13584 11308
rect 13648 11150 13676 12038
rect 13726 11928 13782 11937
rect 13832 11898 13860 13654
rect 13912 13524 13964 13530
rect 13912 13466 13964 13472
rect 13726 11863 13782 11872
rect 13820 11892 13872 11898
rect 13636 11144 13688 11150
rect 13636 11086 13688 11092
rect 13556 10968 13676 10996
rect 13544 10464 13596 10470
rect 13544 10406 13596 10412
rect 13556 10062 13584 10406
rect 13544 10056 13596 10062
rect 13544 9998 13596 10004
rect 13556 9722 13584 9998
rect 13544 9716 13596 9722
rect 13544 9658 13596 9664
rect 13544 9444 13596 9450
rect 13544 9386 13596 9392
rect 13452 9036 13504 9042
rect 13452 8978 13504 8984
rect 13452 8832 13504 8838
rect 13452 8774 13504 8780
rect 13464 8634 13492 8774
rect 13452 8628 13504 8634
rect 13452 8570 13504 8576
rect 13556 8294 13584 9386
rect 13648 9110 13676 10968
rect 13740 10810 13768 11863
rect 13820 11834 13872 11840
rect 13820 11280 13872 11286
rect 13820 11222 13872 11228
rect 13728 10804 13780 10810
rect 13728 10746 13780 10752
rect 13832 10742 13860 11222
rect 13820 10736 13872 10742
rect 13820 10678 13872 10684
rect 13728 10668 13780 10674
rect 13728 10610 13780 10616
rect 13740 10266 13768 10610
rect 13728 10260 13780 10266
rect 13728 10202 13780 10208
rect 13820 9920 13872 9926
rect 13820 9862 13872 9868
rect 13726 9752 13782 9761
rect 13832 9722 13860 9862
rect 13726 9687 13782 9696
rect 13820 9716 13872 9722
rect 13636 9104 13688 9110
rect 13636 9046 13688 9052
rect 13740 8922 13768 9687
rect 13820 9658 13872 9664
rect 13820 9580 13872 9586
rect 13820 9522 13872 9528
rect 13648 8894 13768 8922
rect 13544 8288 13596 8294
rect 13544 8230 13596 8236
rect 13360 7880 13412 7886
rect 13360 7822 13412 7828
rect 13648 7342 13676 8894
rect 13728 8832 13780 8838
rect 13728 8774 13780 8780
rect 13636 7336 13688 7342
rect 13636 7278 13688 7284
rect 13360 7268 13412 7274
rect 13360 7210 13412 7216
rect 13452 7268 13504 7274
rect 13452 7210 13504 7216
rect 12950 7100 13258 7109
rect 12950 7098 12956 7100
rect 13012 7098 13036 7100
rect 13092 7098 13116 7100
rect 13172 7098 13196 7100
rect 13252 7098 13258 7100
rect 13012 7046 13014 7098
rect 13194 7046 13196 7098
rect 12950 7044 12956 7046
rect 13012 7044 13036 7046
rect 13092 7044 13116 7046
rect 13172 7044 13196 7046
rect 13252 7044 13258 7046
rect 12950 7035 13258 7044
rect 12808 6996 12860 7002
rect 12808 6938 12860 6944
rect 13372 6934 13400 7210
rect 12716 6928 12768 6934
rect 12716 6870 12768 6876
rect 13360 6928 13412 6934
rect 13360 6870 13412 6876
rect 12992 6656 13044 6662
rect 12992 6598 13044 6604
rect 13360 6656 13412 6662
rect 13360 6598 13412 6604
rect 13004 6458 13032 6598
rect 12992 6452 13044 6458
rect 12992 6394 13044 6400
rect 12950 6012 13258 6021
rect 12950 6010 12956 6012
rect 13012 6010 13036 6012
rect 13092 6010 13116 6012
rect 13172 6010 13196 6012
rect 13252 6010 13258 6012
rect 13012 5958 13014 6010
rect 13194 5958 13196 6010
rect 12950 5956 12956 5958
rect 13012 5956 13036 5958
rect 13092 5956 13116 5958
rect 13172 5956 13196 5958
rect 13252 5956 13258 5958
rect 12950 5947 13258 5956
rect 12716 5704 12768 5710
rect 12716 5646 12768 5652
rect 12728 3942 12756 5646
rect 13268 5296 13320 5302
rect 13268 5238 13320 5244
rect 13280 5098 13308 5238
rect 13268 5092 13320 5098
rect 13268 5034 13320 5040
rect 12808 5024 12860 5030
rect 12808 4966 12860 4972
rect 12820 4826 12848 4966
rect 12950 4924 13258 4933
rect 12950 4922 12956 4924
rect 13012 4922 13036 4924
rect 13092 4922 13116 4924
rect 13172 4922 13196 4924
rect 13252 4922 13258 4924
rect 13012 4870 13014 4922
rect 13194 4870 13196 4922
rect 12950 4868 12956 4870
rect 13012 4868 13036 4870
rect 13092 4868 13116 4870
rect 13172 4868 13196 4870
rect 13252 4868 13258 4870
rect 12950 4859 13258 4868
rect 12808 4820 12860 4826
rect 12808 4762 12860 4768
rect 12992 4140 13044 4146
rect 12992 4082 13044 4088
rect 12808 4072 12860 4078
rect 13004 4049 13032 4082
rect 12808 4014 12860 4020
rect 12990 4040 13046 4049
rect 12716 3936 12768 3942
rect 12716 3878 12768 3884
rect 12624 3460 12676 3466
rect 12624 3402 12676 3408
rect 11612 3052 11664 3058
rect 11612 2994 11664 3000
rect 12532 3052 12584 3058
rect 12532 2994 12584 3000
rect 11624 2774 11652 2994
rect 12164 2984 12216 2990
rect 12164 2926 12216 2932
rect 11796 2848 11848 2854
rect 11796 2790 11848 2796
rect 11440 2746 11652 2774
rect 11336 2100 11388 2106
rect 11336 2042 11388 2048
rect 11440 800 11468 2746
rect 11808 800 11836 2790
rect 12176 800 12204 2926
rect 12348 2440 12400 2446
rect 12400 2400 12572 2428
rect 12348 2382 12400 2388
rect 12544 800 12572 2400
rect 12820 2088 12848 4014
rect 12990 3975 13046 3984
rect 12950 3836 13258 3845
rect 12950 3834 12956 3836
rect 13012 3834 13036 3836
rect 13092 3834 13116 3836
rect 13172 3834 13196 3836
rect 13252 3834 13258 3836
rect 13012 3782 13014 3834
rect 13194 3782 13196 3834
rect 12950 3780 12956 3782
rect 13012 3780 13036 3782
rect 13092 3780 13116 3782
rect 13172 3780 13196 3782
rect 13252 3780 13258 3782
rect 12950 3771 13258 3780
rect 13372 3398 13400 6598
rect 13464 4690 13492 7210
rect 13634 7168 13690 7177
rect 13634 7103 13690 7112
rect 13544 6656 13596 6662
rect 13544 6598 13596 6604
rect 13556 6390 13584 6598
rect 13544 6384 13596 6390
rect 13544 6326 13596 6332
rect 13544 5364 13596 5370
rect 13544 5306 13596 5312
rect 13452 4684 13504 4690
rect 13452 4626 13504 4632
rect 13556 4282 13584 5306
rect 13544 4276 13596 4282
rect 13544 4218 13596 4224
rect 13360 3392 13412 3398
rect 13360 3334 13412 3340
rect 13648 3194 13676 7103
rect 13740 6254 13768 8774
rect 13832 8294 13860 9522
rect 13924 8906 13952 13466
rect 14004 12980 14056 12986
rect 14004 12922 14056 12928
rect 14016 12714 14044 12922
rect 14004 12708 14056 12714
rect 14004 12650 14056 12656
rect 14108 12345 14136 16390
rect 14280 15360 14332 15366
rect 14280 15302 14332 15308
rect 14292 15162 14320 15302
rect 14280 15156 14332 15162
rect 14280 15098 14332 15104
rect 14188 15088 14240 15094
rect 14188 15030 14240 15036
rect 14200 13530 14228 15030
rect 14384 14618 14412 19110
rect 14476 15094 14504 22510
rect 14660 21690 14688 23462
rect 14648 21684 14700 21690
rect 14648 21626 14700 21632
rect 14752 21350 14780 26930
rect 14844 26314 14872 27882
rect 15120 27674 15148 28630
rect 15200 28416 15252 28422
rect 15200 28358 15252 28364
rect 15108 27668 15160 27674
rect 15108 27610 15160 27616
rect 15108 27532 15160 27538
rect 15108 27474 15160 27480
rect 15016 27124 15068 27130
rect 15016 27066 15068 27072
rect 15028 26450 15056 27066
rect 15120 26858 15148 27474
rect 15212 27062 15240 28358
rect 15200 27056 15252 27062
rect 15200 26998 15252 27004
rect 15108 26852 15160 26858
rect 15108 26794 15160 26800
rect 15108 26512 15160 26518
rect 15108 26454 15160 26460
rect 15016 26444 15068 26450
rect 15016 26386 15068 26392
rect 14832 26308 14884 26314
rect 14832 26250 14884 26256
rect 15120 25974 15148 26454
rect 15108 25968 15160 25974
rect 15108 25910 15160 25916
rect 15016 25832 15068 25838
rect 15016 25774 15068 25780
rect 15108 25832 15160 25838
rect 15108 25774 15160 25780
rect 15028 25702 15056 25774
rect 15016 25696 15068 25702
rect 15016 25638 15068 25644
rect 15120 25362 15148 25774
rect 15108 25356 15160 25362
rect 15108 25298 15160 25304
rect 15396 25158 15424 29106
rect 15476 27328 15528 27334
rect 15476 27270 15528 27276
rect 15292 25152 15344 25158
rect 15384 25152 15436 25158
rect 15292 25094 15344 25100
rect 15382 25120 15384 25129
rect 15436 25120 15438 25129
rect 15304 24818 15332 25094
rect 15382 25055 15438 25064
rect 15488 24954 15516 27270
rect 15856 25770 15884 30194
rect 15948 28558 15976 31726
rect 16592 31142 16620 33798
rect 16684 32366 16712 38286
rect 16764 38208 16816 38214
rect 16764 38150 16816 38156
rect 16672 32360 16724 32366
rect 16672 32302 16724 32308
rect 16684 31890 16712 32302
rect 16672 31884 16724 31890
rect 16672 31826 16724 31832
rect 16672 31680 16724 31686
rect 16672 31622 16724 31628
rect 16580 31136 16632 31142
rect 16580 31078 16632 31084
rect 16592 30598 16620 31078
rect 16580 30592 16632 30598
rect 16580 30534 16632 30540
rect 16028 30184 16080 30190
rect 16028 30126 16080 30132
rect 16120 30184 16172 30190
rect 16120 30126 16172 30132
rect 16040 30054 16068 30126
rect 16028 30048 16080 30054
rect 16028 29990 16080 29996
rect 16028 29504 16080 29510
rect 16028 29446 16080 29452
rect 16040 29073 16068 29446
rect 16132 29102 16160 30126
rect 16212 30048 16264 30054
rect 16212 29990 16264 29996
rect 16120 29096 16172 29102
rect 16026 29064 16082 29073
rect 16120 29038 16172 29044
rect 16026 28999 16082 29008
rect 15936 28552 15988 28558
rect 15936 28494 15988 28500
rect 15936 28416 15988 28422
rect 15936 28358 15988 28364
rect 15948 28150 15976 28358
rect 15936 28144 15988 28150
rect 15936 28086 15988 28092
rect 16040 28082 16068 28999
rect 16224 28506 16252 29990
rect 16304 29844 16356 29850
rect 16304 29786 16356 29792
rect 16132 28478 16252 28506
rect 16028 28076 16080 28082
rect 16028 28018 16080 28024
rect 15936 27056 15988 27062
rect 15936 26998 15988 27004
rect 15948 26790 15976 26998
rect 15936 26784 15988 26790
rect 15936 26726 15988 26732
rect 15844 25764 15896 25770
rect 15844 25706 15896 25712
rect 15476 24948 15528 24954
rect 15476 24890 15528 24896
rect 15292 24812 15344 24818
rect 15292 24754 15344 24760
rect 15948 24732 15976 26726
rect 16028 26240 16080 26246
rect 16028 26182 16080 26188
rect 16040 26042 16068 26182
rect 16132 26042 16160 28478
rect 16212 28416 16264 28422
rect 16212 28358 16264 28364
rect 16224 27470 16252 28358
rect 16212 27464 16264 27470
rect 16212 27406 16264 27412
rect 16028 26036 16080 26042
rect 16028 25978 16080 25984
rect 16120 26036 16172 26042
rect 16120 25978 16172 25984
rect 16132 25702 16160 25978
rect 16120 25696 16172 25702
rect 16120 25638 16172 25644
rect 16028 24744 16080 24750
rect 15948 24704 16028 24732
rect 16028 24686 16080 24692
rect 15384 24608 15436 24614
rect 15384 24550 15436 24556
rect 15844 24608 15896 24614
rect 15844 24550 15896 24556
rect 15016 24404 15068 24410
rect 15016 24346 15068 24352
rect 15028 23186 15056 24346
rect 15108 23520 15160 23526
rect 15108 23462 15160 23468
rect 15120 23254 15148 23462
rect 15108 23248 15160 23254
rect 15108 23190 15160 23196
rect 15016 23180 15068 23186
rect 15016 23122 15068 23128
rect 15028 22710 15056 23122
rect 15016 22704 15068 22710
rect 15016 22646 15068 22652
rect 15200 22432 15252 22438
rect 15200 22374 15252 22380
rect 15212 22166 15240 22374
rect 15200 22160 15252 22166
rect 15200 22102 15252 22108
rect 15396 22098 15424 24550
rect 15660 22228 15712 22234
rect 15660 22170 15712 22176
rect 15384 22092 15436 22098
rect 15384 22034 15436 22040
rect 15476 22092 15528 22098
rect 15476 22034 15528 22040
rect 14924 21888 14976 21894
rect 14924 21830 14976 21836
rect 15292 21888 15344 21894
rect 15292 21830 15344 21836
rect 14936 21622 14964 21830
rect 14924 21616 14976 21622
rect 14924 21558 14976 21564
rect 15108 21480 15160 21486
rect 15108 21422 15160 21428
rect 14740 21344 14792 21350
rect 14740 21286 14792 21292
rect 15120 21078 15148 21422
rect 15200 21140 15252 21146
rect 15200 21082 15252 21088
rect 15108 21072 15160 21078
rect 15108 21014 15160 21020
rect 15212 20942 15240 21082
rect 15200 20936 15252 20942
rect 15200 20878 15252 20884
rect 14740 20800 14792 20806
rect 14740 20742 14792 20748
rect 14648 20392 14700 20398
rect 14648 20334 14700 20340
rect 14556 19780 14608 19786
rect 14556 19722 14608 19728
rect 14568 18426 14596 19722
rect 14660 19446 14688 20334
rect 14648 19440 14700 19446
rect 14648 19382 14700 19388
rect 14752 18834 14780 20742
rect 14740 18828 14792 18834
rect 14740 18770 14792 18776
rect 14648 18624 14700 18630
rect 14648 18566 14700 18572
rect 14556 18420 14608 18426
rect 14556 18362 14608 18368
rect 14660 17746 14688 18566
rect 15212 18426 15240 20878
rect 15304 18766 15332 21830
rect 15488 21554 15516 22034
rect 15672 21690 15700 22170
rect 15660 21684 15712 21690
rect 15660 21626 15712 21632
rect 15476 21548 15528 21554
rect 15476 21490 15528 21496
rect 15384 21412 15436 21418
rect 15384 21354 15436 21360
rect 15292 18760 15344 18766
rect 15292 18702 15344 18708
rect 15200 18420 15252 18426
rect 15120 18380 15200 18408
rect 14648 17740 14700 17746
rect 14648 17682 14700 17688
rect 15120 17338 15148 18380
rect 15200 18362 15252 18368
rect 15200 17604 15252 17610
rect 15200 17546 15252 17552
rect 15108 17332 15160 17338
rect 15108 17274 15160 17280
rect 15212 17270 15240 17546
rect 15200 17264 15252 17270
rect 15200 17206 15252 17212
rect 15212 16998 15240 17206
rect 15200 16992 15252 16998
rect 15200 16934 15252 16940
rect 15292 16108 15344 16114
rect 15292 16050 15344 16056
rect 14556 16040 14608 16046
rect 14556 15982 14608 15988
rect 14568 15706 14596 15982
rect 14556 15700 14608 15706
rect 14556 15642 14608 15648
rect 15304 15570 15332 16050
rect 15292 15564 15344 15570
rect 15292 15506 15344 15512
rect 15396 15314 15424 21354
rect 15476 21344 15528 21350
rect 15476 21286 15528 21292
rect 15488 21010 15516 21286
rect 15476 21004 15528 21010
rect 15476 20946 15528 20952
rect 15856 20602 15884 24550
rect 16040 24342 16068 24686
rect 16028 24336 16080 24342
rect 16028 24278 16080 24284
rect 16132 23730 16160 25638
rect 16120 23724 16172 23730
rect 16120 23666 16172 23672
rect 16132 23526 16160 23666
rect 16212 23588 16264 23594
rect 16212 23530 16264 23536
rect 16120 23520 16172 23526
rect 16120 23462 16172 23468
rect 16120 22500 16172 22506
rect 16120 22442 16172 22448
rect 16028 22092 16080 22098
rect 16132 22080 16160 22442
rect 16080 22052 16160 22080
rect 16028 22034 16080 22040
rect 16132 21146 16160 22052
rect 16120 21140 16172 21146
rect 16120 21082 16172 21088
rect 16028 21004 16080 21010
rect 16028 20946 16080 20952
rect 15844 20596 15896 20602
rect 15844 20538 15896 20544
rect 15936 19984 15988 19990
rect 15936 19926 15988 19932
rect 15752 18692 15804 18698
rect 15752 18634 15804 18640
rect 15764 18222 15792 18634
rect 15752 18216 15804 18222
rect 15752 18158 15804 18164
rect 15568 17604 15620 17610
rect 15568 17546 15620 17552
rect 15476 17128 15528 17134
rect 15476 17070 15528 17076
rect 15488 16250 15516 17070
rect 15476 16244 15528 16250
rect 15476 16186 15528 16192
rect 15212 15286 15424 15314
rect 14464 15088 14516 15094
rect 14464 15030 14516 15036
rect 14556 15020 14608 15026
rect 14556 14962 14608 14968
rect 14372 14612 14424 14618
rect 14372 14554 14424 14560
rect 14372 13864 14424 13870
rect 14372 13806 14424 13812
rect 14188 13524 14240 13530
rect 14188 13466 14240 13472
rect 14280 12844 14332 12850
rect 14280 12786 14332 12792
rect 14094 12336 14150 12345
rect 14094 12271 14150 12280
rect 14188 12300 14240 12306
rect 14188 12242 14240 12248
rect 14004 11824 14056 11830
rect 14004 11766 14056 11772
rect 13912 8900 13964 8906
rect 13912 8842 13964 8848
rect 13820 8288 13872 8294
rect 13820 8230 13872 8236
rect 13832 7818 13860 8230
rect 13820 7812 13872 7818
rect 13820 7754 13872 7760
rect 13832 6390 13860 7754
rect 14016 7206 14044 11766
rect 14200 11694 14228 12242
rect 14292 12238 14320 12786
rect 14384 12782 14412 13806
rect 14372 12776 14424 12782
rect 14372 12718 14424 12724
rect 14280 12232 14332 12238
rect 14280 12174 14332 12180
rect 14372 12232 14424 12238
rect 14372 12174 14424 12180
rect 14384 12102 14412 12174
rect 14372 12096 14424 12102
rect 14372 12038 14424 12044
rect 14188 11688 14240 11694
rect 14188 11630 14240 11636
rect 14096 11620 14148 11626
rect 14096 11562 14148 11568
rect 14108 11014 14136 11562
rect 14188 11552 14240 11558
rect 14188 11494 14240 11500
rect 14200 11150 14228 11494
rect 14384 11218 14412 12038
rect 14464 11892 14516 11898
rect 14464 11834 14516 11840
rect 14372 11212 14424 11218
rect 14372 11154 14424 11160
rect 14188 11144 14240 11150
rect 14188 11086 14240 11092
rect 14280 11076 14332 11082
rect 14280 11018 14332 11024
rect 14096 11008 14148 11014
rect 14096 10950 14148 10956
rect 14188 10464 14240 10470
rect 14188 10406 14240 10412
rect 14096 9920 14148 9926
rect 14094 9888 14096 9897
rect 14148 9888 14150 9897
rect 14094 9823 14150 9832
rect 14096 9172 14148 9178
rect 14096 9114 14148 9120
rect 14108 8498 14136 9114
rect 14096 8492 14148 8498
rect 14096 8434 14148 8440
rect 14004 7200 14056 7206
rect 14004 7142 14056 7148
rect 13820 6384 13872 6390
rect 13820 6326 13872 6332
rect 13728 6248 13780 6254
rect 13728 6190 13780 6196
rect 13728 6112 13780 6118
rect 13728 6054 13780 6060
rect 13740 5234 13768 6054
rect 14004 5568 14056 5574
rect 14004 5510 14056 5516
rect 14016 5302 14044 5510
rect 14004 5296 14056 5302
rect 14004 5238 14056 5244
rect 13728 5228 13780 5234
rect 13728 5170 13780 5176
rect 13912 4072 13964 4078
rect 13912 4014 13964 4020
rect 13924 3534 13952 4014
rect 14004 3596 14056 3602
rect 14004 3538 14056 3544
rect 13912 3528 13964 3534
rect 13912 3470 13964 3476
rect 13636 3188 13688 3194
rect 13636 3130 13688 3136
rect 13174 3088 13230 3097
rect 13174 3023 13176 3032
rect 13228 3023 13230 3032
rect 13176 2994 13228 3000
rect 13636 2984 13688 2990
rect 13636 2926 13688 2932
rect 12950 2748 13258 2757
rect 12950 2746 12956 2748
rect 13012 2746 13036 2748
rect 13092 2746 13116 2748
rect 13172 2746 13196 2748
rect 13252 2746 13258 2748
rect 13012 2694 13014 2746
rect 13194 2694 13196 2746
rect 12950 2692 12956 2694
rect 13012 2692 13036 2694
rect 13092 2692 13116 2694
rect 13172 2692 13196 2694
rect 13252 2692 13258 2694
rect 12950 2683 13258 2692
rect 13268 2372 13320 2378
rect 13268 2314 13320 2320
rect 12820 2060 12940 2088
rect 12912 800 12940 2060
rect 13280 800 13308 2314
rect 13648 800 13676 2926
rect 13924 2650 13952 3470
rect 13820 2644 13872 2650
rect 13820 2586 13872 2592
rect 13912 2644 13964 2650
rect 13912 2586 13964 2592
rect 13832 2378 13860 2586
rect 13820 2372 13872 2378
rect 13820 2314 13872 2320
rect 14016 800 14044 3538
rect 14200 2378 14228 10406
rect 14292 9450 14320 11018
rect 14384 10810 14412 11154
rect 14476 11082 14504 11834
rect 14568 11286 14596 14962
rect 14740 14612 14792 14618
rect 14740 14554 14792 14560
rect 14648 14068 14700 14074
rect 14648 14010 14700 14016
rect 14556 11280 14608 11286
rect 14556 11222 14608 11228
rect 14464 11076 14516 11082
rect 14464 11018 14516 11024
rect 14660 10996 14688 14010
rect 14752 12102 14780 14554
rect 15108 14544 15160 14550
rect 15108 14486 15160 14492
rect 14924 13932 14976 13938
rect 14924 13874 14976 13880
rect 14936 13802 14964 13874
rect 14924 13796 14976 13802
rect 14924 13738 14976 13744
rect 14936 13394 14964 13738
rect 15016 13524 15068 13530
rect 15016 13466 15068 13472
rect 14924 13388 14976 13394
rect 14924 13330 14976 13336
rect 15028 12306 15056 13466
rect 15120 12918 15148 14486
rect 15212 14414 15240 15286
rect 15292 15156 15344 15162
rect 15292 15098 15344 15104
rect 15200 14408 15252 14414
rect 15200 14350 15252 14356
rect 15200 13728 15252 13734
rect 15200 13670 15252 13676
rect 15108 12912 15160 12918
rect 15108 12854 15160 12860
rect 15108 12776 15160 12782
rect 15108 12718 15160 12724
rect 15016 12300 15068 12306
rect 15016 12242 15068 12248
rect 14830 12200 14886 12209
rect 14830 12135 14886 12144
rect 14740 12096 14792 12102
rect 14740 12038 14792 12044
rect 14568 10968 14688 10996
rect 14372 10804 14424 10810
rect 14372 10746 14424 10752
rect 14568 10441 14596 10968
rect 14646 10840 14702 10849
rect 14646 10775 14702 10784
rect 14554 10432 14610 10441
rect 14554 10367 14610 10376
rect 14462 10296 14518 10305
rect 14462 10231 14518 10240
rect 14280 9444 14332 9450
rect 14280 9386 14332 9392
rect 14280 8424 14332 8430
rect 14280 8366 14332 8372
rect 14292 3738 14320 8366
rect 14372 6180 14424 6186
rect 14372 6122 14424 6128
rect 14384 5710 14412 6122
rect 14372 5704 14424 5710
rect 14372 5646 14424 5652
rect 14370 4720 14426 4729
rect 14370 4655 14372 4664
rect 14424 4655 14426 4664
rect 14372 4626 14424 4632
rect 14476 4570 14504 10231
rect 14556 8900 14608 8906
rect 14556 8842 14608 8848
rect 14384 4542 14504 4570
rect 14384 4078 14412 4542
rect 14464 4480 14516 4486
rect 14464 4422 14516 4428
rect 14372 4072 14424 4078
rect 14372 4014 14424 4020
rect 14280 3732 14332 3738
rect 14280 3674 14332 3680
rect 14476 2446 14504 4422
rect 14568 3058 14596 8842
rect 14660 4758 14688 10775
rect 14752 10674 14780 12038
rect 14844 11898 14872 12135
rect 14924 12096 14976 12102
rect 14924 12038 14976 12044
rect 14832 11892 14884 11898
rect 14832 11834 14884 11840
rect 14832 11756 14884 11762
rect 14832 11698 14884 11704
rect 14740 10668 14792 10674
rect 14740 10610 14792 10616
rect 14844 10470 14872 11698
rect 14936 11082 14964 12038
rect 15120 11762 15148 12718
rect 15212 11898 15240 13670
rect 15304 13326 15332 15098
rect 15580 14890 15608 17546
rect 15660 17536 15712 17542
rect 15660 17478 15712 17484
rect 15672 16590 15700 17478
rect 15752 16652 15804 16658
rect 15752 16594 15804 16600
rect 15660 16584 15712 16590
rect 15660 16526 15712 16532
rect 15764 16402 15792 16594
rect 15672 16374 15792 16402
rect 15568 14884 15620 14890
rect 15568 14826 15620 14832
rect 15384 14476 15436 14482
rect 15384 14418 15436 14424
rect 15568 14476 15620 14482
rect 15568 14418 15620 14424
rect 15396 13394 15424 14418
rect 15580 13938 15608 14418
rect 15568 13932 15620 13938
rect 15568 13874 15620 13880
rect 15384 13388 15436 13394
rect 15384 13330 15436 13336
rect 15292 13320 15344 13326
rect 15292 13262 15344 13268
rect 15672 13190 15700 16374
rect 15844 16108 15896 16114
rect 15844 16050 15896 16056
rect 15856 13870 15884 16050
rect 15844 13864 15896 13870
rect 15844 13806 15896 13812
rect 15856 13394 15884 13806
rect 15948 13734 15976 19926
rect 16040 19514 16068 20946
rect 16028 19508 16080 19514
rect 16028 19450 16080 19456
rect 16120 18624 16172 18630
rect 16120 18566 16172 18572
rect 16028 15360 16080 15366
rect 16028 15302 16080 15308
rect 16040 14958 16068 15302
rect 16028 14952 16080 14958
rect 16028 14894 16080 14900
rect 16040 14278 16068 14894
rect 16028 14272 16080 14278
rect 16026 14240 16028 14249
rect 16080 14240 16082 14249
rect 16026 14175 16082 14184
rect 15936 13728 15988 13734
rect 15936 13670 15988 13676
rect 15844 13388 15896 13394
rect 15844 13330 15896 13336
rect 15384 13184 15436 13190
rect 15290 13152 15346 13161
rect 15384 13126 15436 13132
rect 15568 13184 15620 13190
rect 15660 13184 15712 13190
rect 15568 13126 15620 13132
rect 15658 13152 15660 13161
rect 15752 13184 15804 13190
rect 15712 13152 15714 13161
rect 15290 13087 15346 13096
rect 15304 12714 15332 13087
rect 15292 12708 15344 12714
rect 15292 12650 15344 12656
rect 15292 12300 15344 12306
rect 15292 12242 15344 12248
rect 15200 11892 15252 11898
rect 15200 11834 15252 11840
rect 15108 11756 15160 11762
rect 15108 11698 15160 11704
rect 15016 11212 15068 11218
rect 15016 11154 15068 11160
rect 14924 11076 14976 11082
rect 14924 11018 14976 11024
rect 14922 10568 14978 10577
rect 14922 10503 14978 10512
rect 14832 10464 14884 10470
rect 14832 10406 14884 10412
rect 14936 10130 14964 10503
rect 14924 10124 14976 10130
rect 14924 10066 14976 10072
rect 15028 7954 15056 11154
rect 15120 9382 15148 11698
rect 15304 11558 15332 12242
rect 15292 11552 15344 11558
rect 15292 11494 15344 11500
rect 15396 11354 15424 13126
rect 15580 12782 15608 13126
rect 15752 13126 15804 13132
rect 15658 13087 15714 13096
rect 15764 12986 15792 13126
rect 15752 12980 15804 12986
rect 15752 12922 15804 12928
rect 15752 12844 15804 12850
rect 15752 12786 15804 12792
rect 15568 12776 15620 12782
rect 15568 12718 15620 12724
rect 15660 12368 15712 12374
rect 15660 12310 15712 12316
rect 15384 11348 15436 11354
rect 15384 11290 15436 11296
rect 15290 11112 15346 11121
rect 15290 11047 15346 11056
rect 15200 9580 15252 9586
rect 15200 9522 15252 9528
rect 15108 9376 15160 9382
rect 15108 9318 15160 9324
rect 15212 9110 15240 9522
rect 15200 9104 15252 9110
rect 15200 9046 15252 9052
rect 15108 8424 15160 8430
rect 15108 8366 15160 8372
rect 15016 7948 15068 7954
rect 15016 7890 15068 7896
rect 15016 7812 15068 7818
rect 15016 7754 15068 7760
rect 15028 7290 15056 7754
rect 15120 7478 15148 8366
rect 15108 7472 15160 7478
rect 15108 7414 15160 7420
rect 15028 7262 15240 7290
rect 15212 7206 15240 7262
rect 15016 7200 15068 7206
rect 15016 7142 15068 7148
rect 15200 7200 15252 7206
rect 15200 7142 15252 7148
rect 15028 6798 15056 7142
rect 15212 7002 15240 7142
rect 15200 6996 15252 7002
rect 15120 6956 15200 6984
rect 15016 6792 15068 6798
rect 15016 6734 15068 6740
rect 15016 6316 15068 6322
rect 15016 6258 15068 6264
rect 14648 4752 14700 4758
rect 14648 4694 14700 4700
rect 15028 3670 15056 6258
rect 15120 5574 15148 6956
rect 15200 6938 15252 6944
rect 15304 6746 15332 11047
rect 15568 10804 15620 10810
rect 15568 10746 15620 10752
rect 15580 10690 15608 10746
rect 15488 10662 15608 10690
rect 15384 10532 15436 10538
rect 15384 10474 15436 10480
rect 15212 6718 15332 6746
rect 15212 6254 15240 6718
rect 15292 6656 15344 6662
rect 15292 6598 15344 6604
rect 15200 6248 15252 6254
rect 15200 6190 15252 6196
rect 15200 5704 15252 5710
rect 15200 5646 15252 5652
rect 15108 5568 15160 5574
rect 15108 5510 15160 5516
rect 15120 5234 15148 5510
rect 15108 5228 15160 5234
rect 15108 5170 15160 5176
rect 15120 4486 15148 5170
rect 15212 5030 15240 5646
rect 15200 5024 15252 5030
rect 15200 4966 15252 4972
rect 15304 4554 15332 6598
rect 15396 5302 15424 10474
rect 15488 9586 15516 10662
rect 15568 10532 15620 10538
rect 15568 10474 15620 10480
rect 15580 10441 15608 10474
rect 15566 10432 15622 10441
rect 15566 10367 15622 10376
rect 15672 10266 15700 12310
rect 15568 10260 15620 10266
rect 15568 10202 15620 10208
rect 15660 10260 15712 10266
rect 15660 10202 15712 10208
rect 15580 10146 15608 10202
rect 15580 10118 15700 10146
rect 15568 10056 15620 10062
rect 15568 9998 15620 10004
rect 15476 9580 15528 9586
rect 15476 9522 15528 9528
rect 15580 9450 15608 9998
rect 15568 9444 15620 9450
rect 15568 9386 15620 9392
rect 15568 8016 15620 8022
rect 15568 7958 15620 7964
rect 15580 7750 15608 7958
rect 15568 7744 15620 7750
rect 15568 7686 15620 7692
rect 15474 7576 15530 7585
rect 15474 7511 15476 7520
rect 15528 7511 15530 7520
rect 15476 7482 15528 7488
rect 15568 7336 15620 7342
rect 15488 7296 15568 7324
rect 15384 5296 15436 5302
rect 15384 5238 15436 5244
rect 15488 5030 15516 7296
rect 15568 7278 15620 7284
rect 15672 6730 15700 10118
rect 15764 9994 15792 12786
rect 15936 12776 15988 12782
rect 15936 12718 15988 12724
rect 15948 12646 15976 12718
rect 15844 12640 15896 12646
rect 15844 12582 15896 12588
rect 15936 12640 15988 12646
rect 15936 12582 15988 12588
rect 15752 9988 15804 9994
rect 15752 9930 15804 9936
rect 15752 9580 15804 9586
rect 15752 9522 15804 9528
rect 15660 6724 15712 6730
rect 15660 6666 15712 6672
rect 15568 6248 15620 6254
rect 15568 6190 15620 6196
rect 15476 5024 15528 5030
rect 15476 4966 15528 4972
rect 15292 4548 15344 4554
rect 15292 4490 15344 4496
rect 15384 4548 15436 4554
rect 15384 4490 15436 4496
rect 15108 4480 15160 4486
rect 15108 4422 15160 4428
rect 15396 4010 15424 4490
rect 15488 4078 15516 4966
rect 15580 4214 15608 6190
rect 15568 4208 15620 4214
rect 15568 4150 15620 4156
rect 15476 4072 15528 4078
rect 15476 4014 15528 4020
rect 15384 4004 15436 4010
rect 15384 3946 15436 3952
rect 15016 3664 15068 3670
rect 14646 3632 14702 3641
rect 15016 3606 15068 3612
rect 14646 3567 14702 3576
rect 15476 3596 15528 3602
rect 14660 3534 14688 3567
rect 15476 3538 15528 3544
rect 14648 3528 14700 3534
rect 14648 3470 14700 3476
rect 14556 3052 14608 3058
rect 14556 2994 14608 3000
rect 14740 2984 14792 2990
rect 14740 2926 14792 2932
rect 14464 2440 14516 2446
rect 14464 2382 14516 2388
rect 14188 2372 14240 2378
rect 14188 2314 14240 2320
rect 14372 2372 14424 2378
rect 14372 2314 14424 2320
rect 14384 800 14412 2314
rect 14752 800 14780 2926
rect 15108 2916 15160 2922
rect 15108 2858 15160 2864
rect 15120 800 15148 2858
rect 15488 800 15516 3538
rect 15764 2854 15792 9522
rect 15856 8634 15884 12582
rect 16132 12434 16160 18566
rect 16224 18358 16252 23530
rect 16316 22710 16344 29786
rect 16580 29504 16632 29510
rect 16500 29452 16580 29458
rect 16500 29446 16632 29452
rect 16500 29430 16620 29446
rect 16500 29306 16528 29430
rect 16488 29300 16540 29306
rect 16488 29242 16540 29248
rect 16580 29300 16632 29306
rect 16580 29242 16632 29248
rect 16396 28552 16448 28558
rect 16396 28494 16448 28500
rect 16408 27878 16436 28494
rect 16488 28416 16540 28422
rect 16488 28358 16540 28364
rect 16396 27872 16448 27878
rect 16396 27814 16448 27820
rect 16408 26994 16436 27814
rect 16500 27470 16528 28358
rect 16488 27464 16540 27470
rect 16488 27406 16540 27412
rect 16488 27328 16540 27334
rect 16488 27270 16540 27276
rect 16396 26988 16448 26994
rect 16396 26930 16448 26936
rect 16500 26790 16528 27270
rect 16488 26784 16540 26790
rect 16488 26726 16540 26732
rect 16592 26314 16620 29242
rect 16684 28082 16712 31622
rect 16776 31278 16804 38150
rect 16868 36530 16896 41414
rect 16960 41386 17080 41414
rect 16868 36502 16988 36530
rect 16856 32428 16908 32434
rect 16856 32370 16908 32376
rect 16868 31890 16896 32370
rect 16856 31884 16908 31890
rect 16856 31826 16908 31832
rect 16868 31482 16896 31826
rect 16856 31476 16908 31482
rect 16856 31418 16908 31424
rect 16764 31272 16816 31278
rect 16764 31214 16816 31220
rect 16960 30122 16988 36502
rect 17052 32570 17080 41386
rect 17144 32586 17172 45526
rect 17512 35290 17540 45834
rect 17500 35284 17552 35290
rect 17500 35226 17552 35232
rect 17408 33992 17460 33998
rect 17408 33934 17460 33940
rect 17144 32570 17264 32586
rect 17040 32564 17092 32570
rect 17040 32506 17092 32512
rect 17132 32564 17264 32570
rect 17184 32558 17264 32564
rect 17132 32506 17184 32512
rect 16948 30116 17000 30122
rect 16948 30058 17000 30064
rect 16856 29504 16908 29510
rect 16856 29446 16908 29452
rect 16672 28076 16724 28082
rect 16672 28018 16724 28024
rect 16580 26308 16632 26314
rect 16580 26250 16632 26256
rect 16672 26240 16724 26246
rect 16672 26182 16724 26188
rect 16488 25696 16540 25702
rect 16488 25638 16540 25644
rect 16396 24948 16448 24954
rect 16396 24890 16448 24896
rect 16408 24410 16436 24890
rect 16396 24404 16448 24410
rect 16396 24346 16448 24352
rect 16304 22704 16356 22710
rect 16304 22646 16356 22652
rect 16500 22080 16528 25638
rect 16316 22052 16528 22080
rect 16316 18834 16344 22052
rect 16580 21548 16632 21554
rect 16580 21490 16632 21496
rect 16488 21140 16540 21146
rect 16488 21082 16540 21088
rect 16396 19508 16448 19514
rect 16396 19450 16448 19456
rect 16304 18828 16356 18834
rect 16304 18770 16356 18776
rect 16212 18352 16264 18358
rect 16212 18294 16264 18300
rect 16224 17066 16252 18294
rect 16304 17128 16356 17134
rect 16304 17070 16356 17076
rect 16212 17060 16264 17066
rect 16212 17002 16264 17008
rect 16224 15094 16252 17002
rect 16212 15088 16264 15094
rect 16212 15030 16264 15036
rect 16316 14906 16344 17070
rect 16408 16454 16436 19450
rect 16500 16658 16528 21082
rect 16592 19922 16620 21490
rect 16580 19916 16632 19922
rect 16580 19858 16632 19864
rect 16592 19310 16620 19858
rect 16684 19334 16712 26182
rect 16868 24750 16896 29446
rect 17052 29306 17080 32506
rect 17132 31748 17184 31754
rect 17132 31690 17184 31696
rect 17144 31482 17172 31690
rect 17132 31476 17184 31482
rect 17132 31418 17184 31424
rect 17040 29300 17092 29306
rect 17040 29242 17092 29248
rect 17052 29102 17080 29242
rect 17236 29170 17264 32558
rect 17420 32434 17448 33934
rect 17408 32428 17460 32434
rect 17408 32370 17460 32376
rect 17316 32360 17368 32366
rect 17316 32302 17368 32308
rect 17328 31686 17356 32302
rect 17604 31754 17632 47942
rect 17950 47900 18258 47909
rect 17950 47898 17956 47900
rect 18012 47898 18036 47900
rect 18092 47898 18116 47900
rect 18172 47898 18196 47900
rect 18252 47898 18258 47900
rect 18012 47846 18014 47898
rect 18194 47846 18196 47898
rect 17950 47844 17956 47846
rect 18012 47844 18036 47846
rect 18092 47844 18116 47846
rect 18172 47844 18196 47846
rect 18252 47844 18258 47846
rect 17950 47835 18258 47844
rect 17950 46812 18258 46821
rect 17950 46810 17956 46812
rect 18012 46810 18036 46812
rect 18092 46810 18116 46812
rect 18172 46810 18196 46812
rect 18252 46810 18258 46812
rect 18012 46758 18014 46810
rect 18194 46758 18196 46810
rect 17950 46756 17956 46758
rect 18012 46756 18036 46758
rect 18092 46756 18116 46758
rect 18172 46756 18196 46758
rect 18252 46756 18258 46758
rect 17950 46747 18258 46756
rect 17950 45724 18258 45733
rect 17950 45722 17956 45724
rect 18012 45722 18036 45724
rect 18092 45722 18116 45724
rect 18172 45722 18196 45724
rect 18252 45722 18258 45724
rect 18012 45670 18014 45722
rect 18194 45670 18196 45722
rect 17950 45668 17956 45670
rect 18012 45668 18036 45670
rect 18092 45668 18116 45670
rect 18172 45668 18196 45670
rect 18252 45668 18258 45670
rect 17950 45659 18258 45668
rect 17950 44636 18258 44645
rect 17950 44634 17956 44636
rect 18012 44634 18036 44636
rect 18092 44634 18116 44636
rect 18172 44634 18196 44636
rect 18252 44634 18258 44636
rect 18012 44582 18014 44634
rect 18194 44582 18196 44634
rect 17950 44580 17956 44582
rect 18012 44580 18036 44582
rect 18092 44580 18116 44582
rect 18172 44580 18196 44582
rect 18252 44580 18258 44582
rect 17950 44571 18258 44580
rect 17950 43548 18258 43557
rect 17950 43546 17956 43548
rect 18012 43546 18036 43548
rect 18092 43546 18116 43548
rect 18172 43546 18196 43548
rect 18252 43546 18258 43548
rect 18012 43494 18014 43546
rect 18194 43494 18196 43546
rect 17950 43492 17956 43494
rect 18012 43492 18036 43494
rect 18092 43492 18116 43494
rect 18172 43492 18196 43494
rect 18252 43492 18258 43494
rect 17950 43483 18258 43492
rect 17950 42460 18258 42469
rect 17950 42458 17956 42460
rect 18012 42458 18036 42460
rect 18092 42458 18116 42460
rect 18172 42458 18196 42460
rect 18252 42458 18258 42460
rect 18012 42406 18014 42458
rect 18194 42406 18196 42458
rect 17950 42404 17956 42406
rect 18012 42404 18036 42406
rect 18092 42404 18116 42406
rect 18172 42404 18196 42406
rect 18252 42404 18258 42406
rect 17950 42395 18258 42404
rect 18800 41414 18828 53994
rect 20364 52494 20392 56200
rect 20720 53984 20772 53990
rect 20720 53926 20772 53932
rect 20352 52488 20404 52494
rect 20352 52430 20404 52436
rect 18972 47252 19024 47258
rect 18972 47194 19024 47200
rect 18708 41386 18828 41414
rect 18984 41414 19012 47194
rect 20732 44946 20760 53926
rect 21364 51264 21416 51270
rect 21364 51206 21416 51212
rect 20904 49768 20956 49774
rect 20904 49710 20956 49716
rect 20720 44940 20772 44946
rect 20720 44882 20772 44888
rect 19432 44872 19484 44878
rect 19432 44814 19484 44820
rect 18984 41386 19104 41414
rect 17950 41372 18258 41381
rect 17950 41370 17956 41372
rect 18012 41370 18036 41372
rect 18092 41370 18116 41372
rect 18172 41370 18196 41372
rect 18252 41370 18258 41372
rect 18012 41318 18014 41370
rect 18194 41318 18196 41370
rect 17950 41316 17956 41318
rect 18012 41316 18036 41318
rect 18092 41316 18116 41318
rect 18172 41316 18196 41318
rect 18252 41316 18258 41318
rect 17950 41307 18258 41316
rect 17950 40284 18258 40293
rect 17950 40282 17956 40284
rect 18012 40282 18036 40284
rect 18092 40282 18116 40284
rect 18172 40282 18196 40284
rect 18252 40282 18258 40284
rect 18012 40230 18014 40282
rect 18194 40230 18196 40282
rect 17950 40228 17956 40230
rect 18012 40228 18036 40230
rect 18092 40228 18116 40230
rect 18172 40228 18196 40230
rect 18252 40228 18258 40230
rect 17950 40219 18258 40228
rect 17950 39196 18258 39205
rect 17950 39194 17956 39196
rect 18012 39194 18036 39196
rect 18092 39194 18116 39196
rect 18172 39194 18196 39196
rect 18252 39194 18258 39196
rect 18012 39142 18014 39194
rect 18194 39142 18196 39194
rect 17950 39140 17956 39142
rect 18012 39140 18036 39142
rect 18092 39140 18116 39142
rect 18172 39140 18196 39142
rect 18252 39140 18258 39142
rect 17950 39131 18258 39140
rect 17950 38108 18258 38117
rect 17950 38106 17956 38108
rect 18012 38106 18036 38108
rect 18092 38106 18116 38108
rect 18172 38106 18196 38108
rect 18252 38106 18258 38108
rect 18012 38054 18014 38106
rect 18194 38054 18196 38106
rect 17950 38052 17956 38054
rect 18012 38052 18036 38054
rect 18092 38052 18116 38054
rect 18172 38052 18196 38054
rect 18252 38052 18258 38054
rect 17950 38043 18258 38052
rect 17950 37020 18258 37029
rect 17950 37018 17956 37020
rect 18012 37018 18036 37020
rect 18092 37018 18116 37020
rect 18172 37018 18196 37020
rect 18252 37018 18258 37020
rect 18012 36966 18014 37018
rect 18194 36966 18196 37018
rect 17950 36964 17956 36966
rect 18012 36964 18036 36966
rect 18092 36964 18116 36966
rect 18172 36964 18196 36966
rect 18252 36964 18258 36966
rect 17950 36955 18258 36964
rect 17950 35932 18258 35941
rect 17950 35930 17956 35932
rect 18012 35930 18036 35932
rect 18092 35930 18116 35932
rect 18172 35930 18196 35932
rect 18252 35930 18258 35932
rect 18012 35878 18014 35930
rect 18194 35878 18196 35930
rect 17950 35876 17956 35878
rect 18012 35876 18036 35878
rect 18092 35876 18116 35878
rect 18172 35876 18196 35878
rect 18252 35876 18258 35878
rect 17950 35867 18258 35876
rect 17950 34844 18258 34853
rect 17950 34842 17956 34844
rect 18012 34842 18036 34844
rect 18092 34842 18116 34844
rect 18172 34842 18196 34844
rect 18252 34842 18258 34844
rect 18012 34790 18014 34842
rect 18194 34790 18196 34842
rect 17950 34788 17956 34790
rect 18012 34788 18036 34790
rect 18092 34788 18116 34790
rect 18172 34788 18196 34790
rect 18252 34788 18258 34790
rect 17950 34779 18258 34788
rect 17950 33756 18258 33765
rect 17950 33754 17956 33756
rect 18012 33754 18036 33756
rect 18092 33754 18116 33756
rect 18172 33754 18196 33756
rect 18252 33754 18258 33756
rect 18012 33702 18014 33754
rect 18194 33702 18196 33754
rect 17950 33700 17956 33702
rect 18012 33700 18036 33702
rect 18092 33700 18116 33702
rect 18172 33700 18196 33702
rect 18252 33700 18258 33702
rect 17950 33691 18258 33700
rect 18604 32904 18656 32910
rect 18604 32846 18656 32852
rect 17684 32768 17736 32774
rect 17684 32710 17736 32716
rect 17696 32502 17724 32710
rect 17950 32668 18258 32677
rect 17950 32666 17956 32668
rect 18012 32666 18036 32668
rect 18092 32666 18116 32668
rect 18172 32666 18196 32668
rect 18252 32666 18258 32668
rect 18012 32614 18014 32666
rect 18194 32614 18196 32666
rect 17950 32612 17956 32614
rect 18012 32612 18036 32614
rect 18092 32612 18116 32614
rect 18172 32612 18196 32614
rect 18252 32612 18258 32614
rect 17950 32603 18258 32612
rect 18420 32564 18472 32570
rect 18420 32506 18472 32512
rect 17684 32496 17736 32502
rect 17684 32438 17736 32444
rect 17868 32224 17920 32230
rect 17868 32166 17920 32172
rect 17880 32026 17908 32166
rect 17868 32020 17920 32026
rect 17868 31962 17920 31968
rect 17880 31754 17908 31962
rect 18432 31754 18460 32506
rect 18616 32026 18644 32846
rect 18604 32020 18656 32026
rect 18604 31962 18656 31968
rect 17512 31726 17632 31754
rect 17696 31726 17908 31754
rect 18420 31748 18472 31754
rect 17316 31680 17368 31686
rect 17316 31622 17368 31628
rect 17316 30592 17368 30598
rect 17316 30534 17368 30540
rect 17224 29164 17276 29170
rect 17224 29106 17276 29112
rect 17040 29096 17092 29102
rect 17040 29038 17092 29044
rect 17052 24834 17080 29038
rect 17132 27532 17184 27538
rect 17132 27474 17184 27480
rect 17144 27334 17172 27474
rect 17132 27328 17184 27334
rect 17132 27270 17184 27276
rect 17144 24886 17172 27270
rect 16960 24806 17080 24834
rect 17132 24880 17184 24886
rect 17132 24822 17184 24828
rect 16856 24744 16908 24750
rect 16856 24686 16908 24692
rect 16960 23662 16988 24806
rect 17040 24676 17092 24682
rect 17040 24618 17092 24624
rect 17052 24206 17080 24618
rect 17040 24200 17092 24206
rect 17040 24142 17092 24148
rect 16948 23656 17000 23662
rect 16948 23598 17000 23604
rect 17132 23656 17184 23662
rect 17132 23598 17184 23604
rect 16948 23520 17000 23526
rect 16948 23462 17000 23468
rect 16764 19712 16816 19718
rect 16764 19654 16816 19660
rect 16776 19514 16804 19654
rect 16960 19514 16988 23462
rect 17144 23322 17172 23598
rect 17132 23316 17184 23322
rect 17132 23258 17184 23264
rect 17040 22976 17092 22982
rect 17040 22918 17092 22924
rect 17052 22098 17080 22918
rect 17144 22778 17172 23258
rect 17132 22772 17184 22778
rect 17132 22714 17184 22720
rect 17040 22092 17092 22098
rect 17040 22034 17092 22040
rect 17052 21146 17080 22034
rect 17040 21140 17092 21146
rect 17040 21082 17092 21088
rect 16764 19508 16816 19514
rect 16764 19450 16816 19456
rect 16948 19508 17000 19514
rect 16948 19450 17000 19456
rect 16580 19304 16632 19310
rect 16684 19306 16804 19334
rect 16580 19246 16632 19252
rect 16672 17740 16724 17746
rect 16672 17682 16724 17688
rect 16580 17060 16632 17066
rect 16580 17002 16632 17008
rect 16488 16652 16540 16658
rect 16488 16594 16540 16600
rect 16396 16448 16448 16454
rect 16396 16390 16448 16396
rect 16592 15434 16620 17002
rect 16684 16998 16712 17682
rect 16776 17678 16804 19306
rect 17236 18834 17264 29106
rect 17328 27878 17356 30534
rect 17408 30048 17460 30054
rect 17408 29990 17460 29996
rect 17420 29714 17448 29990
rect 17408 29708 17460 29714
rect 17408 29650 17460 29656
rect 17512 29152 17540 31726
rect 17696 31142 17724 31726
rect 18420 31690 18472 31696
rect 17950 31580 18258 31589
rect 17950 31578 17956 31580
rect 18012 31578 18036 31580
rect 18092 31578 18116 31580
rect 18172 31578 18196 31580
rect 18252 31578 18258 31580
rect 18012 31526 18014 31578
rect 18194 31526 18196 31578
rect 17950 31524 17956 31526
rect 18012 31524 18036 31526
rect 18092 31524 18116 31526
rect 18172 31524 18196 31526
rect 18252 31524 18258 31526
rect 17950 31515 18258 31524
rect 17684 31136 17736 31142
rect 17684 31078 17736 31084
rect 17512 29124 17632 29152
rect 17408 29096 17460 29102
rect 17460 29073 17540 29084
rect 17460 29064 17554 29073
rect 17460 29056 17498 29064
rect 17408 29038 17460 29044
rect 17498 28999 17554 29008
rect 17408 28484 17460 28490
rect 17408 28426 17460 28432
rect 17420 28218 17448 28426
rect 17408 28212 17460 28218
rect 17408 28154 17460 28160
rect 17512 28014 17540 28999
rect 17408 28008 17460 28014
rect 17408 27950 17460 27956
rect 17500 28008 17552 28014
rect 17500 27950 17552 27956
rect 17316 27872 17368 27878
rect 17316 27814 17368 27820
rect 17328 25294 17356 27814
rect 17420 27334 17448 27950
rect 17500 27464 17552 27470
rect 17500 27406 17552 27412
rect 17408 27328 17460 27334
rect 17408 27270 17460 27276
rect 17316 25288 17368 25294
rect 17316 25230 17368 25236
rect 17132 18828 17184 18834
rect 17132 18770 17184 18776
rect 17224 18828 17276 18834
rect 17224 18770 17276 18776
rect 17144 18630 17172 18770
rect 17040 18624 17092 18630
rect 17040 18566 17092 18572
rect 17132 18624 17184 18630
rect 17132 18566 17184 18572
rect 16856 18284 16908 18290
rect 16856 18226 16908 18232
rect 16764 17672 16816 17678
rect 16764 17614 16816 17620
rect 16764 17536 16816 17542
rect 16764 17478 16816 17484
rect 16672 16992 16724 16998
rect 16670 16960 16672 16969
rect 16724 16960 16726 16969
rect 16670 16895 16726 16904
rect 16672 16788 16724 16794
rect 16672 16730 16724 16736
rect 16684 16697 16712 16730
rect 16670 16688 16726 16697
rect 16670 16623 16726 16632
rect 16580 15428 16632 15434
rect 16580 15370 16632 15376
rect 16224 14878 16344 14906
rect 16224 12918 16252 14878
rect 16304 14272 16356 14278
rect 16304 14214 16356 14220
rect 16580 14272 16632 14278
rect 16580 14214 16632 14220
rect 16316 13977 16344 14214
rect 16488 14068 16540 14074
rect 16488 14010 16540 14016
rect 16302 13968 16358 13977
rect 16302 13903 16358 13912
rect 16304 13728 16356 13734
rect 16304 13670 16356 13676
rect 16212 12912 16264 12918
rect 16212 12854 16264 12860
rect 16040 12406 16160 12434
rect 15934 11792 15990 11801
rect 15934 11727 15990 11736
rect 15948 10810 15976 11727
rect 15936 10804 15988 10810
rect 15936 10746 15988 10752
rect 15934 10432 15990 10441
rect 15934 10367 15990 10376
rect 15844 8628 15896 8634
rect 15844 8570 15896 8576
rect 15948 8401 15976 10367
rect 16040 10198 16068 12406
rect 16316 12238 16344 13670
rect 16396 13320 16448 13326
rect 16396 13262 16448 13268
rect 16304 12232 16356 12238
rect 16304 12174 16356 12180
rect 16120 12096 16172 12102
rect 16120 12038 16172 12044
rect 16212 12096 16264 12102
rect 16212 12038 16264 12044
rect 16132 11830 16160 12038
rect 16120 11824 16172 11830
rect 16120 11766 16172 11772
rect 16120 10804 16172 10810
rect 16120 10746 16172 10752
rect 16132 10577 16160 10746
rect 16118 10568 16174 10577
rect 16118 10503 16174 10512
rect 16028 10192 16080 10198
rect 16028 10134 16080 10140
rect 16118 9888 16174 9897
rect 16118 9823 16174 9832
rect 16132 9586 16160 9823
rect 16120 9580 16172 9586
rect 16120 9522 16172 9528
rect 15934 8392 15990 8401
rect 15934 8327 15990 8336
rect 16028 7744 16080 7750
rect 16028 7686 16080 7692
rect 15844 6928 15896 6934
rect 15844 6870 15896 6876
rect 15856 5166 15884 6870
rect 16040 6866 16068 7686
rect 16120 7200 16172 7206
rect 16120 7142 16172 7148
rect 16028 6860 16080 6866
rect 16028 6802 16080 6808
rect 16028 6724 16080 6730
rect 16028 6666 16080 6672
rect 15844 5160 15896 5166
rect 15844 5102 15896 5108
rect 15844 2984 15896 2990
rect 15844 2926 15896 2932
rect 15752 2848 15804 2854
rect 15752 2790 15804 2796
rect 15856 800 15884 2926
rect 16040 1970 16068 6666
rect 16132 6322 16160 7142
rect 16120 6316 16172 6322
rect 16120 6258 16172 6264
rect 16224 4162 16252 12038
rect 16316 9897 16344 12174
rect 16302 9888 16358 9897
rect 16302 9823 16358 9832
rect 16408 9518 16436 13262
rect 16500 11257 16528 14010
rect 16592 13326 16620 14214
rect 16580 13320 16632 13326
rect 16580 13262 16632 13268
rect 16776 12306 16804 17478
rect 16868 17202 16896 18226
rect 16856 17196 16908 17202
rect 16856 17138 16908 17144
rect 16856 16992 16908 16998
rect 16856 16934 16908 16940
rect 16946 16960 17002 16969
rect 16868 14618 16896 16934
rect 16946 16895 17002 16904
rect 16960 15434 16988 16895
rect 16948 15428 17000 15434
rect 16948 15370 17000 15376
rect 16960 15094 16988 15370
rect 16948 15088 17000 15094
rect 16948 15030 17000 15036
rect 16856 14612 16908 14618
rect 16856 14554 16908 14560
rect 16960 14074 16988 15030
rect 16948 14068 17000 14074
rect 16948 14010 17000 14016
rect 16946 12880 17002 12889
rect 16946 12815 16948 12824
rect 17000 12815 17002 12824
rect 16948 12786 17000 12792
rect 16764 12300 16816 12306
rect 16816 12260 16988 12288
rect 16764 12242 16816 12248
rect 16764 12096 16816 12102
rect 16578 12064 16634 12073
rect 16764 12038 16816 12044
rect 16578 11999 16634 12008
rect 16486 11248 16542 11257
rect 16486 11183 16542 11192
rect 16500 11082 16528 11183
rect 16488 11076 16540 11082
rect 16488 11018 16540 11024
rect 16488 10464 16540 10470
rect 16488 10406 16540 10412
rect 16500 10198 16528 10406
rect 16592 10266 16620 11999
rect 16672 11008 16724 11014
rect 16672 10950 16724 10956
rect 16684 10742 16712 10950
rect 16672 10736 16724 10742
rect 16672 10678 16724 10684
rect 16672 10464 16724 10470
rect 16672 10406 16724 10412
rect 16580 10260 16632 10266
rect 16580 10202 16632 10208
rect 16488 10192 16540 10198
rect 16488 10134 16540 10140
rect 16580 9920 16632 9926
rect 16580 9862 16632 9868
rect 16396 9512 16448 9518
rect 16396 9454 16448 9460
rect 16304 9444 16356 9450
rect 16304 9386 16356 9392
rect 16316 5574 16344 9386
rect 16408 9042 16436 9454
rect 16396 9036 16448 9042
rect 16396 8978 16448 8984
rect 16408 8430 16436 8978
rect 16488 8832 16540 8838
rect 16488 8774 16540 8780
rect 16500 8430 16528 8774
rect 16396 8424 16448 8430
rect 16396 8366 16448 8372
rect 16488 8424 16540 8430
rect 16488 8366 16540 8372
rect 16394 8256 16450 8265
rect 16394 8191 16450 8200
rect 16408 7546 16436 8191
rect 16396 7540 16448 7546
rect 16396 7482 16448 7488
rect 16396 7200 16448 7206
rect 16592 7177 16620 9862
rect 16684 8090 16712 10406
rect 16776 8362 16804 12038
rect 16960 11778 16988 12260
rect 17052 11898 17080 18566
rect 17236 18086 17264 18770
rect 17224 18080 17276 18086
rect 17224 18022 17276 18028
rect 17236 16402 17264 18022
rect 17328 17882 17356 25230
rect 17420 24954 17448 27270
rect 17408 24948 17460 24954
rect 17408 24890 17460 24896
rect 17408 24744 17460 24750
rect 17408 24686 17460 24692
rect 17420 22438 17448 24686
rect 17408 22432 17460 22438
rect 17408 22374 17460 22380
rect 17408 19984 17460 19990
rect 17408 19926 17460 19932
rect 17316 17876 17368 17882
rect 17316 17818 17368 17824
rect 17328 17270 17356 17818
rect 17316 17264 17368 17270
rect 17316 17206 17368 17212
rect 17328 16794 17356 17206
rect 17316 16788 17368 16794
rect 17316 16730 17368 16736
rect 17420 16538 17448 19926
rect 17512 18766 17540 27406
rect 17604 23866 17632 29124
rect 17696 28082 17724 31078
rect 18432 30666 18460 31690
rect 18420 30660 18472 30666
rect 18420 30602 18472 30608
rect 17950 30492 18258 30501
rect 17950 30490 17956 30492
rect 18012 30490 18036 30492
rect 18092 30490 18116 30492
rect 18172 30490 18196 30492
rect 18252 30490 18258 30492
rect 18012 30438 18014 30490
rect 18194 30438 18196 30490
rect 17950 30436 17956 30438
rect 18012 30436 18036 30438
rect 18092 30436 18116 30438
rect 18172 30436 18196 30438
rect 18252 30436 18258 30438
rect 17950 30427 18258 30436
rect 18432 29578 18460 30602
rect 18420 29572 18472 29578
rect 18420 29514 18472 29520
rect 17950 29404 18258 29413
rect 17950 29402 17956 29404
rect 18012 29402 18036 29404
rect 18092 29402 18116 29404
rect 18172 29402 18196 29404
rect 18252 29402 18258 29404
rect 18012 29350 18014 29402
rect 18194 29350 18196 29402
rect 17950 29348 17956 29350
rect 18012 29348 18036 29350
rect 18092 29348 18116 29350
rect 18172 29348 18196 29350
rect 18252 29348 18258 29350
rect 17950 29339 18258 29348
rect 18432 29306 18460 29514
rect 18420 29300 18472 29306
rect 18420 29242 18472 29248
rect 18432 28490 18460 29242
rect 18420 28484 18472 28490
rect 18420 28426 18472 28432
rect 17950 28316 18258 28325
rect 17950 28314 17956 28316
rect 18012 28314 18036 28316
rect 18092 28314 18116 28316
rect 18172 28314 18196 28316
rect 18252 28314 18258 28316
rect 18012 28262 18014 28314
rect 18194 28262 18196 28314
rect 17950 28260 17956 28262
rect 18012 28260 18036 28262
rect 18092 28260 18116 28262
rect 18172 28260 18196 28262
rect 18252 28260 18258 28262
rect 17950 28251 18258 28260
rect 18432 28200 18460 28426
rect 18432 28172 18552 28200
rect 17684 28076 17736 28082
rect 17684 28018 17736 28024
rect 18420 28076 18472 28082
rect 18420 28018 18472 28024
rect 17696 27334 17724 28018
rect 17960 27872 18012 27878
rect 17960 27814 18012 27820
rect 17972 27470 18000 27814
rect 18432 27538 18460 28018
rect 18420 27532 18472 27538
rect 18420 27474 18472 27480
rect 17960 27464 18012 27470
rect 17960 27406 18012 27412
rect 17684 27328 17736 27334
rect 17682 27296 17684 27305
rect 17736 27296 17738 27305
rect 17682 27231 17738 27240
rect 17950 27228 18258 27237
rect 17950 27226 17956 27228
rect 18012 27226 18036 27228
rect 18092 27226 18116 27228
rect 18172 27226 18196 27228
rect 18252 27226 18258 27228
rect 18012 27174 18014 27226
rect 18194 27174 18196 27226
rect 17950 27172 17956 27174
rect 18012 27172 18036 27174
rect 18092 27172 18116 27174
rect 18172 27172 18196 27174
rect 18252 27172 18258 27174
rect 17950 27163 18258 27172
rect 18524 27062 18552 28172
rect 18616 28014 18644 31962
rect 18708 31754 18736 41386
rect 18972 32564 19024 32570
rect 18972 32506 19024 32512
rect 18984 32366 19012 32506
rect 18972 32360 19024 32366
rect 18972 32302 19024 32308
rect 19076 31754 19104 41386
rect 19340 34604 19392 34610
rect 19340 34546 19392 34552
rect 19352 32230 19380 34546
rect 19444 34134 19472 44814
rect 20916 41414 20944 49710
rect 21376 45082 21404 51206
rect 21364 45076 21416 45082
rect 21364 45018 21416 45024
rect 21272 44940 21324 44946
rect 21272 44882 21324 44888
rect 21284 44810 21312 44882
rect 21272 44804 21324 44810
rect 21272 44746 21324 44752
rect 21284 41414 21312 44746
rect 20916 41386 21036 41414
rect 21284 41386 21404 41414
rect 20536 38208 20588 38214
rect 20536 38150 20588 38156
rect 19892 35556 19944 35562
rect 19892 35498 19944 35504
rect 19616 35080 19668 35086
rect 19616 35022 19668 35028
rect 19432 34128 19484 34134
rect 19432 34070 19484 34076
rect 19444 33522 19472 34070
rect 19628 33658 19656 35022
rect 19708 34944 19760 34950
rect 19708 34886 19760 34892
rect 19720 33930 19748 34886
rect 19708 33924 19760 33930
rect 19708 33866 19760 33872
rect 19616 33652 19668 33658
rect 19616 33594 19668 33600
rect 19432 33516 19484 33522
rect 19432 33458 19484 33464
rect 19432 32904 19484 32910
rect 19432 32846 19484 32852
rect 19444 32502 19472 32846
rect 19524 32768 19576 32774
rect 19524 32710 19576 32716
rect 19432 32496 19484 32502
rect 19432 32438 19484 32444
rect 19340 32224 19392 32230
rect 19340 32166 19392 32172
rect 19352 32026 19380 32166
rect 19340 32020 19392 32026
rect 19340 31962 19392 31968
rect 19444 31906 19472 32438
rect 18708 31726 18828 31754
rect 18696 31272 18748 31278
rect 18696 31214 18748 31220
rect 18708 30938 18736 31214
rect 18696 30932 18748 30938
rect 18696 30874 18748 30880
rect 18800 30818 18828 31726
rect 18880 31748 18932 31754
rect 18880 31690 18932 31696
rect 18984 31726 19104 31754
rect 19352 31890 19472 31906
rect 19352 31884 19484 31890
rect 19352 31878 19432 31884
rect 18892 30938 18920 31690
rect 18880 30932 18932 30938
rect 18880 30874 18932 30880
rect 18708 30790 18828 30818
rect 18604 28008 18656 28014
rect 18604 27950 18656 27956
rect 18708 27606 18736 30790
rect 18880 30728 18932 30734
rect 18880 30670 18932 30676
rect 18788 30252 18840 30258
rect 18788 30194 18840 30200
rect 18800 29646 18828 30194
rect 18788 29640 18840 29646
rect 18788 29582 18840 29588
rect 18800 28762 18828 29582
rect 18892 29510 18920 30670
rect 18880 29504 18932 29510
rect 18880 29446 18932 29452
rect 18788 28756 18840 28762
rect 18788 28698 18840 28704
rect 18696 27600 18748 27606
rect 18696 27542 18748 27548
rect 18604 27396 18656 27402
rect 18656 27356 18736 27384
rect 18604 27338 18656 27344
rect 18604 27124 18656 27130
rect 18604 27066 18656 27072
rect 18512 27056 18564 27062
rect 18512 26998 18564 27004
rect 18616 26908 18644 27066
rect 18524 26880 18644 26908
rect 17960 26376 18012 26382
rect 17958 26344 17960 26353
rect 18328 26376 18380 26382
rect 18012 26344 18014 26353
rect 18328 26318 18380 26324
rect 17958 26279 18014 26288
rect 17950 26140 18258 26149
rect 17950 26138 17956 26140
rect 18012 26138 18036 26140
rect 18092 26138 18116 26140
rect 18172 26138 18196 26140
rect 18252 26138 18258 26140
rect 18012 26086 18014 26138
rect 18194 26086 18196 26138
rect 17950 26084 17956 26086
rect 18012 26084 18036 26086
rect 18092 26084 18116 26086
rect 18172 26084 18196 26086
rect 18252 26084 18258 26086
rect 17950 26075 18258 26084
rect 18340 26042 18368 26318
rect 18328 26036 18380 26042
rect 18328 25978 18380 25984
rect 17950 25052 18258 25061
rect 17950 25050 17956 25052
rect 18012 25050 18036 25052
rect 18092 25050 18116 25052
rect 18172 25050 18196 25052
rect 18252 25050 18258 25052
rect 18012 24998 18014 25050
rect 18194 24998 18196 25050
rect 17950 24996 17956 24998
rect 18012 24996 18036 24998
rect 18092 24996 18116 24998
rect 18172 24996 18196 24998
rect 18252 24996 18258 24998
rect 17950 24987 18258 24996
rect 18524 24750 18552 26880
rect 18512 24744 18564 24750
rect 18512 24686 18564 24692
rect 18604 24744 18656 24750
rect 18604 24686 18656 24692
rect 17776 24608 17828 24614
rect 17776 24550 17828 24556
rect 17868 24608 17920 24614
rect 17868 24550 17920 24556
rect 17684 24064 17736 24070
rect 17684 24006 17736 24012
rect 17592 23860 17644 23866
rect 17592 23802 17644 23808
rect 17604 23769 17632 23802
rect 17590 23760 17646 23769
rect 17590 23695 17646 23704
rect 17592 22568 17644 22574
rect 17592 22510 17644 22516
rect 17604 22112 17632 22510
rect 17592 22106 17644 22112
rect 17592 22048 17644 22054
rect 17500 18760 17552 18766
rect 17500 18702 17552 18708
rect 17592 18760 17644 18766
rect 17592 18702 17644 18708
rect 17420 16510 17540 16538
rect 17408 16448 17460 16454
rect 17236 16374 17356 16402
rect 17408 16390 17460 16396
rect 17222 16280 17278 16289
rect 17222 16215 17278 16224
rect 17236 16182 17264 16215
rect 17224 16176 17276 16182
rect 17224 16118 17276 16124
rect 17328 15994 17356 16374
rect 17236 15966 17356 15994
rect 17236 15366 17264 15966
rect 17316 15904 17368 15910
rect 17316 15846 17368 15852
rect 17224 15360 17276 15366
rect 17328 15337 17356 15846
rect 17224 15302 17276 15308
rect 17314 15328 17370 15337
rect 17314 15263 17370 15272
rect 17132 14000 17184 14006
rect 17132 13942 17184 13948
rect 17040 11892 17092 11898
rect 17040 11834 17092 11840
rect 16960 11750 17080 11778
rect 16854 11520 16910 11529
rect 16854 11455 16910 11464
rect 16868 9178 16896 11455
rect 16948 11008 17000 11014
rect 16948 10950 17000 10956
rect 16960 10441 16988 10950
rect 16946 10432 17002 10441
rect 16946 10367 17002 10376
rect 16948 9648 17000 9654
rect 16946 9616 16948 9625
rect 17000 9616 17002 9625
rect 16946 9551 17002 9560
rect 17052 9466 17080 11750
rect 16960 9438 17080 9466
rect 16856 9172 16908 9178
rect 16856 9114 16908 9120
rect 16856 8968 16908 8974
rect 16854 8936 16856 8945
rect 16908 8936 16910 8945
rect 16854 8871 16910 8880
rect 16764 8356 16816 8362
rect 16764 8298 16816 8304
rect 16672 8084 16724 8090
rect 16672 8026 16724 8032
rect 16856 7948 16908 7954
rect 16856 7890 16908 7896
rect 16672 7880 16724 7886
rect 16672 7822 16724 7828
rect 16396 7142 16448 7148
rect 16578 7168 16634 7177
rect 16304 5568 16356 5574
rect 16304 5510 16356 5516
rect 16224 4134 16344 4162
rect 16120 4072 16172 4078
rect 16120 4014 16172 4020
rect 16212 4072 16264 4078
rect 16212 4014 16264 4020
rect 16132 3194 16160 4014
rect 16120 3188 16172 3194
rect 16120 3130 16172 3136
rect 16118 2544 16174 2553
rect 16118 2479 16174 2488
rect 16132 2310 16160 2479
rect 16120 2304 16172 2310
rect 16120 2246 16172 2252
rect 16028 1964 16080 1970
rect 16028 1906 16080 1912
rect 16224 800 16252 4014
rect 16316 3777 16344 4134
rect 16302 3768 16358 3777
rect 16302 3703 16358 3712
rect 16408 2582 16436 7142
rect 16578 7103 16634 7112
rect 16684 4826 16712 7822
rect 16764 6792 16816 6798
rect 16764 6734 16816 6740
rect 16672 4820 16724 4826
rect 16672 4762 16724 4768
rect 16488 4752 16540 4758
rect 16486 4720 16488 4729
rect 16540 4720 16542 4729
rect 16486 4655 16542 4664
rect 16672 4616 16724 4622
rect 16672 4558 16724 4564
rect 16684 3534 16712 4558
rect 16672 3528 16724 3534
rect 16672 3470 16724 3476
rect 16580 3120 16632 3126
rect 16580 3062 16632 3068
rect 16396 2576 16448 2582
rect 16396 2518 16448 2524
rect 16592 800 16620 3062
rect 16776 2446 16804 6734
rect 16868 6322 16896 7890
rect 16960 7342 16988 9438
rect 17040 9376 17092 9382
rect 17040 9318 17092 9324
rect 16948 7336 17000 7342
rect 16948 7278 17000 7284
rect 16948 6860 17000 6866
rect 16948 6802 17000 6808
rect 16856 6316 16908 6322
rect 16856 6258 16908 6264
rect 16868 5234 16896 6258
rect 16856 5228 16908 5234
rect 16856 5170 16908 5176
rect 16868 4690 16896 5170
rect 16960 4826 16988 6802
rect 16948 4820 17000 4826
rect 16948 4762 17000 4768
rect 16856 4684 16908 4690
rect 16856 4626 16908 4632
rect 16856 4004 16908 4010
rect 16856 3946 16908 3952
rect 16764 2440 16816 2446
rect 16764 2382 16816 2388
rect 16868 2106 16896 3946
rect 16960 3534 16988 4762
rect 16948 3528 17000 3534
rect 16948 3470 17000 3476
rect 16948 2848 17000 2854
rect 16948 2790 17000 2796
rect 16856 2100 16908 2106
rect 16856 2042 16908 2048
rect 16960 800 16988 2790
rect 17052 2446 17080 9318
rect 17144 8888 17172 13942
rect 17224 13728 17276 13734
rect 17224 13670 17276 13676
rect 17236 11529 17264 13670
rect 17420 12434 17448 16390
rect 17512 15978 17540 16510
rect 17500 15972 17552 15978
rect 17500 15914 17552 15920
rect 17604 13734 17632 18702
rect 17696 16590 17724 24006
rect 17788 23866 17816 24550
rect 17776 23860 17828 23866
rect 17776 23802 17828 23808
rect 17776 23656 17828 23662
rect 17776 23598 17828 23604
rect 17788 22438 17816 23598
rect 17776 22432 17828 22438
rect 17776 22374 17828 22380
rect 17776 21888 17828 21894
rect 17776 21830 17828 21836
rect 17788 19990 17816 21830
rect 17776 19984 17828 19990
rect 17776 19926 17828 19932
rect 17788 19378 17816 19926
rect 17880 19922 17908 24550
rect 18524 24342 18552 24686
rect 18512 24336 18564 24342
rect 18512 24278 18564 24284
rect 18236 24200 18288 24206
rect 18236 24142 18288 24148
rect 18248 24070 18276 24142
rect 18236 24064 18288 24070
rect 18236 24006 18288 24012
rect 17950 23964 18258 23973
rect 17950 23962 17956 23964
rect 18012 23962 18036 23964
rect 18092 23962 18116 23964
rect 18172 23962 18196 23964
rect 18252 23962 18258 23964
rect 18012 23910 18014 23962
rect 18194 23910 18196 23962
rect 17950 23908 17956 23910
rect 18012 23908 18036 23910
rect 18092 23908 18116 23910
rect 18172 23908 18196 23910
rect 18252 23908 18258 23910
rect 17950 23899 18258 23908
rect 18236 23860 18288 23866
rect 18236 23802 18288 23808
rect 18248 23610 18276 23802
rect 18524 23730 18552 24278
rect 18512 23724 18564 23730
rect 18512 23666 18564 23672
rect 18248 23582 18460 23610
rect 18248 23186 18276 23582
rect 18328 23520 18380 23526
rect 18328 23462 18380 23468
rect 18236 23180 18288 23186
rect 18236 23122 18288 23128
rect 17950 22876 18258 22885
rect 17950 22874 17956 22876
rect 18012 22874 18036 22876
rect 18092 22874 18116 22876
rect 18172 22874 18196 22876
rect 18252 22874 18258 22876
rect 18012 22822 18014 22874
rect 18194 22822 18196 22874
rect 17950 22820 17956 22822
rect 18012 22820 18036 22822
rect 18092 22820 18116 22822
rect 18172 22820 18196 22822
rect 18252 22820 18258 22822
rect 17950 22811 18258 22820
rect 18236 22432 18288 22438
rect 18236 22374 18288 22380
rect 18248 22234 18276 22374
rect 18236 22228 18288 22234
rect 18236 22170 18288 22176
rect 17950 21788 18258 21797
rect 17950 21786 17956 21788
rect 18012 21786 18036 21788
rect 18092 21786 18116 21788
rect 18172 21786 18196 21788
rect 18252 21786 18258 21788
rect 18012 21734 18014 21786
rect 18194 21734 18196 21786
rect 17950 21732 17956 21734
rect 18012 21732 18036 21734
rect 18092 21732 18116 21734
rect 18172 21732 18196 21734
rect 18252 21732 18258 21734
rect 17950 21723 18258 21732
rect 18340 21010 18368 23462
rect 18432 22710 18460 23582
rect 18512 23248 18564 23254
rect 18512 23190 18564 23196
rect 18420 22704 18472 22710
rect 18420 22646 18472 22652
rect 18420 22432 18472 22438
rect 18420 22374 18472 22380
rect 18432 22166 18460 22374
rect 18420 22160 18472 22166
rect 18420 22102 18472 22108
rect 18432 21962 18460 22102
rect 18420 21956 18472 21962
rect 18420 21898 18472 21904
rect 18328 21004 18380 21010
rect 18328 20946 18380 20952
rect 18420 20936 18472 20942
rect 18420 20878 18472 20884
rect 17950 20700 18258 20709
rect 17950 20698 17956 20700
rect 18012 20698 18036 20700
rect 18092 20698 18116 20700
rect 18172 20698 18196 20700
rect 18252 20698 18258 20700
rect 18012 20646 18014 20698
rect 18194 20646 18196 20698
rect 17950 20644 17956 20646
rect 18012 20644 18036 20646
rect 18092 20644 18116 20646
rect 18172 20644 18196 20646
rect 18252 20644 18258 20646
rect 17950 20635 18258 20644
rect 17868 19916 17920 19922
rect 17868 19858 17920 19864
rect 18432 19786 18460 20878
rect 18420 19780 18472 19786
rect 18420 19722 18472 19728
rect 17950 19612 18258 19621
rect 17950 19610 17956 19612
rect 18012 19610 18036 19612
rect 18092 19610 18116 19612
rect 18172 19610 18196 19612
rect 18252 19610 18258 19612
rect 18012 19558 18014 19610
rect 18194 19558 18196 19610
rect 17950 19556 17956 19558
rect 18012 19556 18036 19558
rect 18092 19556 18116 19558
rect 18172 19556 18196 19558
rect 18252 19556 18258 19558
rect 17950 19547 18258 19556
rect 17776 19372 17828 19378
rect 17776 19314 17828 19320
rect 17776 18828 17828 18834
rect 17776 18770 17828 18776
rect 17684 16584 17736 16590
rect 17684 16526 17736 16532
rect 17788 15706 17816 18770
rect 17950 18524 18258 18533
rect 17950 18522 17956 18524
rect 18012 18522 18036 18524
rect 18092 18522 18116 18524
rect 18172 18522 18196 18524
rect 18252 18522 18258 18524
rect 18012 18470 18014 18522
rect 18194 18470 18196 18522
rect 17950 18468 17956 18470
rect 18012 18468 18036 18470
rect 18092 18468 18116 18470
rect 18172 18468 18196 18470
rect 18252 18468 18258 18470
rect 17950 18459 18258 18468
rect 17868 18352 17920 18358
rect 17868 18294 17920 18300
rect 18418 18320 18474 18329
rect 17880 17814 17908 18294
rect 18418 18255 18474 18264
rect 17868 17808 17920 17814
rect 17866 17776 17868 17785
rect 17920 17776 17922 17785
rect 17866 17711 17922 17720
rect 18328 17672 18380 17678
rect 18328 17614 18380 17620
rect 17950 17436 18258 17445
rect 17950 17434 17956 17436
rect 18012 17434 18036 17436
rect 18092 17434 18116 17436
rect 18172 17434 18196 17436
rect 18252 17434 18258 17436
rect 18012 17382 18014 17434
rect 18194 17382 18196 17434
rect 17950 17380 17956 17382
rect 18012 17380 18036 17382
rect 18092 17380 18116 17382
rect 18172 17380 18196 17382
rect 18252 17380 18258 17382
rect 17950 17371 18258 17380
rect 18340 17202 18368 17614
rect 18328 17196 18380 17202
rect 18328 17138 18380 17144
rect 18328 16788 18380 16794
rect 18328 16730 18380 16736
rect 17950 16348 18258 16357
rect 17950 16346 17956 16348
rect 18012 16346 18036 16348
rect 18092 16346 18116 16348
rect 18172 16346 18196 16348
rect 18252 16346 18258 16348
rect 18012 16294 18014 16346
rect 18194 16294 18196 16346
rect 17950 16292 17956 16294
rect 18012 16292 18036 16294
rect 18092 16292 18116 16294
rect 18172 16292 18196 16294
rect 18252 16292 18258 16294
rect 17950 16283 18258 16292
rect 17776 15700 17828 15706
rect 17776 15642 17828 15648
rect 17592 13728 17644 13734
rect 17592 13670 17644 13676
rect 17684 13728 17736 13734
rect 17684 13670 17736 13676
rect 17592 13320 17644 13326
rect 17592 13262 17644 13268
rect 17500 13252 17552 13258
rect 17500 13194 17552 13200
rect 17328 12406 17448 12434
rect 17222 11520 17278 11529
rect 17222 11455 17278 11464
rect 17224 11348 17276 11354
rect 17224 11290 17276 11296
rect 17236 10674 17264 11290
rect 17328 10674 17356 12406
rect 17408 11688 17460 11694
rect 17408 11630 17460 11636
rect 17420 11354 17448 11630
rect 17408 11348 17460 11354
rect 17408 11290 17460 11296
rect 17406 11248 17462 11257
rect 17406 11183 17462 11192
rect 17420 11150 17448 11183
rect 17408 11144 17460 11150
rect 17408 11086 17460 11092
rect 17224 10668 17276 10674
rect 17224 10610 17276 10616
rect 17316 10668 17368 10674
rect 17316 10610 17368 10616
rect 17328 10418 17356 10610
rect 17408 10600 17460 10606
rect 17408 10542 17460 10548
rect 17236 10390 17356 10418
rect 17236 9722 17264 10390
rect 17316 10260 17368 10266
rect 17316 10202 17368 10208
rect 17328 9926 17356 10202
rect 17420 10130 17448 10542
rect 17408 10124 17460 10130
rect 17408 10066 17460 10072
rect 17316 9920 17368 9926
rect 17316 9862 17368 9868
rect 17512 9722 17540 13194
rect 17604 9761 17632 13262
rect 17696 12646 17724 13670
rect 17788 13326 17816 15642
rect 17950 15260 18258 15269
rect 17950 15258 17956 15260
rect 18012 15258 18036 15260
rect 18092 15258 18116 15260
rect 18172 15258 18196 15260
rect 18252 15258 18258 15260
rect 18012 15206 18014 15258
rect 18194 15206 18196 15258
rect 17950 15204 17956 15206
rect 18012 15204 18036 15206
rect 18092 15204 18116 15206
rect 18172 15204 18196 15206
rect 18252 15204 18258 15206
rect 17950 15195 18258 15204
rect 18340 14618 18368 16730
rect 18432 16726 18460 18255
rect 18524 17746 18552 23190
rect 18616 22982 18644 24686
rect 18604 22976 18656 22982
rect 18604 22918 18656 22924
rect 18604 21888 18656 21894
rect 18604 21830 18656 21836
rect 18616 21418 18644 21830
rect 18604 21412 18656 21418
rect 18604 21354 18656 21360
rect 18616 20466 18644 21354
rect 18604 20460 18656 20466
rect 18604 20402 18656 20408
rect 18708 20346 18736 27356
rect 18892 26450 18920 29446
rect 18880 26444 18932 26450
rect 18880 26386 18932 26392
rect 18984 26353 19012 31726
rect 19352 30802 19380 31878
rect 19432 31826 19484 31832
rect 19536 31346 19564 32710
rect 19524 31340 19576 31346
rect 19524 31282 19576 31288
rect 19432 31204 19484 31210
rect 19432 31146 19484 31152
rect 19340 30796 19392 30802
rect 19340 30738 19392 30744
rect 19156 28416 19208 28422
rect 19156 28358 19208 28364
rect 19064 27872 19116 27878
rect 19064 27814 19116 27820
rect 18970 26344 19026 26353
rect 18970 26279 19026 26288
rect 18880 25832 18932 25838
rect 18880 25774 18932 25780
rect 18788 24812 18840 24818
rect 18788 24754 18840 24760
rect 18800 24614 18828 24754
rect 18788 24608 18840 24614
rect 18788 24550 18840 24556
rect 18800 23050 18828 24550
rect 18892 24206 18920 25774
rect 18972 25696 19024 25702
rect 18972 25638 19024 25644
rect 18880 24200 18932 24206
rect 18880 24142 18932 24148
rect 18880 23180 18932 23186
rect 18880 23122 18932 23128
rect 18788 23044 18840 23050
rect 18788 22986 18840 22992
rect 18800 22574 18828 22986
rect 18788 22568 18840 22574
rect 18788 22510 18840 22516
rect 18800 22234 18828 22510
rect 18788 22228 18840 22234
rect 18788 22170 18840 22176
rect 18892 20618 18920 23122
rect 18984 21554 19012 25638
rect 19076 24070 19104 27814
rect 19064 24064 19116 24070
rect 19064 24006 19116 24012
rect 19076 23322 19104 24006
rect 19064 23316 19116 23322
rect 19064 23258 19116 23264
rect 19064 22432 19116 22438
rect 19064 22374 19116 22380
rect 19076 21622 19104 22374
rect 19064 21616 19116 21622
rect 19064 21558 19116 21564
rect 18972 21548 19024 21554
rect 18972 21490 19024 21496
rect 18892 20590 19012 20618
rect 18616 20318 18736 20346
rect 18788 20392 18840 20398
rect 18788 20334 18840 20340
rect 18616 18766 18644 20318
rect 18696 20256 18748 20262
rect 18696 20198 18748 20204
rect 18708 18766 18736 20198
rect 18800 19514 18828 20334
rect 18984 20262 19012 20590
rect 18972 20256 19024 20262
rect 18972 20198 19024 20204
rect 19064 20256 19116 20262
rect 19064 20198 19116 20204
rect 18788 19508 18840 19514
rect 18788 19450 18840 19456
rect 18972 19508 19024 19514
rect 18972 19450 19024 19456
rect 18788 19168 18840 19174
rect 18788 19110 18840 19116
rect 18800 18834 18828 19110
rect 18788 18828 18840 18834
rect 18788 18770 18840 18776
rect 18604 18760 18656 18766
rect 18604 18702 18656 18708
rect 18696 18760 18748 18766
rect 18696 18702 18748 18708
rect 18616 18358 18644 18702
rect 18604 18352 18656 18358
rect 18604 18294 18656 18300
rect 18616 18193 18644 18294
rect 18602 18184 18658 18193
rect 18602 18119 18658 18128
rect 18604 18080 18656 18086
rect 18604 18022 18656 18028
rect 18616 17746 18644 18022
rect 18512 17740 18564 17746
rect 18512 17682 18564 17688
rect 18604 17740 18656 17746
rect 18604 17682 18656 17688
rect 18616 17202 18644 17682
rect 18604 17196 18656 17202
rect 18604 17138 18656 17144
rect 18420 16720 18472 16726
rect 18420 16662 18472 16668
rect 18604 16584 18656 16590
rect 18604 16526 18656 16532
rect 18616 16250 18644 16526
rect 18604 16244 18656 16250
rect 18604 16186 18656 16192
rect 18604 16108 18656 16114
rect 18604 16050 18656 16056
rect 18328 14612 18380 14618
rect 18380 14572 18460 14600
rect 18328 14554 18380 14560
rect 18328 14476 18380 14482
rect 18328 14418 18380 14424
rect 17950 14172 18258 14181
rect 17950 14170 17956 14172
rect 18012 14170 18036 14172
rect 18092 14170 18116 14172
rect 18172 14170 18196 14172
rect 18252 14170 18258 14172
rect 18012 14118 18014 14170
rect 18194 14118 18196 14170
rect 17950 14116 17956 14118
rect 18012 14116 18036 14118
rect 18092 14116 18116 14118
rect 18172 14116 18196 14118
rect 18252 14116 18258 14118
rect 17950 14107 18258 14116
rect 17868 13864 17920 13870
rect 17868 13806 17920 13812
rect 17776 13320 17828 13326
rect 17776 13262 17828 13268
rect 17880 12782 17908 13806
rect 18340 13326 18368 14418
rect 18432 14006 18460 14572
rect 18616 14074 18644 16050
rect 18708 15026 18736 18702
rect 18880 18080 18932 18086
rect 18880 18022 18932 18028
rect 18786 17776 18842 17785
rect 18786 17711 18788 17720
rect 18840 17711 18842 17720
rect 18788 17682 18840 17688
rect 18800 17542 18828 17682
rect 18788 17536 18840 17542
rect 18788 17478 18840 17484
rect 18892 16454 18920 18022
rect 18880 16448 18932 16454
rect 18880 16390 18932 16396
rect 18788 15360 18840 15366
rect 18788 15302 18840 15308
rect 18696 15020 18748 15026
rect 18696 14962 18748 14968
rect 18696 14816 18748 14822
rect 18696 14758 18748 14764
rect 18604 14068 18656 14074
rect 18604 14010 18656 14016
rect 18420 14000 18472 14006
rect 18420 13942 18472 13948
rect 18328 13320 18380 13326
rect 18328 13262 18380 13268
rect 18328 13184 18380 13190
rect 18328 13126 18380 13132
rect 17950 13084 18258 13093
rect 17950 13082 17956 13084
rect 18012 13082 18036 13084
rect 18092 13082 18116 13084
rect 18172 13082 18196 13084
rect 18252 13082 18258 13084
rect 18012 13030 18014 13082
rect 18194 13030 18196 13082
rect 17950 13028 17956 13030
rect 18012 13028 18036 13030
rect 18092 13028 18116 13030
rect 18172 13028 18196 13030
rect 18252 13028 18258 13030
rect 17950 13019 18258 13028
rect 17868 12776 17920 12782
rect 17868 12718 17920 12724
rect 17684 12640 17736 12646
rect 17684 12582 17736 12588
rect 17776 12640 17828 12646
rect 17776 12582 17828 12588
rect 17682 12472 17738 12481
rect 17682 12407 17738 12416
rect 17696 12374 17724 12407
rect 17684 12368 17736 12374
rect 17684 12310 17736 12316
rect 17682 12200 17738 12209
rect 17682 12135 17738 12144
rect 17696 10062 17724 12135
rect 17788 10849 17816 12582
rect 17880 11150 17908 12718
rect 18340 12170 18368 13126
rect 18432 12850 18460 13942
rect 18420 12844 18472 12850
rect 18420 12786 18472 12792
rect 18432 12442 18460 12786
rect 18512 12776 18564 12782
rect 18512 12718 18564 12724
rect 18420 12436 18472 12442
rect 18420 12378 18472 12384
rect 18418 12336 18474 12345
rect 18418 12271 18474 12280
rect 18432 12170 18460 12271
rect 18328 12164 18380 12170
rect 18328 12106 18380 12112
rect 18420 12164 18472 12170
rect 18420 12106 18472 12112
rect 18524 12102 18552 12718
rect 18616 12306 18644 14010
rect 18604 12300 18656 12306
rect 18604 12242 18656 12248
rect 18708 12209 18736 14758
rect 18800 12481 18828 15302
rect 18984 15094 19012 19450
rect 19076 19417 19104 20198
rect 19168 19854 19196 28358
rect 19444 28150 19472 31146
rect 19616 30048 19668 30054
rect 19616 29990 19668 29996
rect 19432 28144 19484 28150
rect 19432 28086 19484 28092
rect 19248 28076 19300 28082
rect 19248 28018 19300 28024
rect 19260 26858 19288 28018
rect 19432 27464 19484 27470
rect 19432 27406 19484 27412
rect 19248 26852 19300 26858
rect 19248 26794 19300 26800
rect 19260 24274 19288 26794
rect 19444 26790 19472 27406
rect 19432 26784 19484 26790
rect 19432 26726 19484 26732
rect 19340 25152 19392 25158
rect 19338 25120 19340 25129
rect 19392 25120 19394 25129
rect 19338 25055 19394 25064
rect 19444 24750 19472 26726
rect 19432 24744 19484 24750
rect 19432 24686 19484 24692
rect 19340 24404 19392 24410
rect 19340 24346 19392 24352
rect 19248 24268 19300 24274
rect 19248 24210 19300 24216
rect 19352 22710 19380 24346
rect 19444 24206 19472 24686
rect 19432 24200 19484 24206
rect 19432 24142 19484 24148
rect 19340 22704 19392 22710
rect 19340 22646 19392 22652
rect 19248 22636 19300 22642
rect 19248 22578 19300 22584
rect 19260 21690 19288 22578
rect 19340 21888 19392 21894
rect 19340 21830 19392 21836
rect 19248 21684 19300 21690
rect 19248 21626 19300 21632
rect 19352 21486 19380 21830
rect 19340 21480 19392 21486
rect 19340 21422 19392 21428
rect 19340 20800 19392 20806
rect 19340 20742 19392 20748
rect 19248 20596 19300 20602
rect 19248 20538 19300 20544
rect 19156 19848 19208 19854
rect 19156 19790 19208 19796
rect 19062 19408 19118 19417
rect 19260 19378 19288 20538
rect 19352 20466 19380 20742
rect 19340 20460 19392 20466
rect 19340 20402 19392 20408
rect 19444 20330 19472 24142
rect 19524 22976 19576 22982
rect 19524 22918 19576 22924
rect 19432 20324 19484 20330
rect 19432 20266 19484 20272
rect 19062 19343 19118 19352
rect 19248 19372 19300 19378
rect 19248 19314 19300 19320
rect 19248 19168 19300 19174
rect 19248 19110 19300 19116
rect 19064 18896 19116 18902
rect 19064 18838 19116 18844
rect 18972 15088 19024 15094
rect 18972 15030 19024 15036
rect 18880 15020 18932 15026
rect 18880 14962 18932 14968
rect 18786 12472 18842 12481
rect 18786 12407 18842 12416
rect 18788 12368 18840 12374
rect 18788 12310 18840 12316
rect 18694 12200 18750 12209
rect 18694 12135 18750 12144
rect 18512 12096 18564 12102
rect 18512 12038 18564 12044
rect 17950 11996 18258 12005
rect 17950 11994 17956 11996
rect 18012 11994 18036 11996
rect 18092 11994 18116 11996
rect 18172 11994 18196 11996
rect 18252 11994 18258 11996
rect 18012 11942 18014 11994
rect 18194 11942 18196 11994
rect 17950 11940 17956 11942
rect 18012 11940 18036 11942
rect 18092 11940 18116 11942
rect 18172 11940 18196 11942
rect 18252 11940 18258 11942
rect 17950 11931 18258 11940
rect 18524 11801 18552 12038
rect 18510 11792 18566 11801
rect 18510 11727 18566 11736
rect 18512 11688 18564 11694
rect 18510 11656 18512 11665
rect 18564 11656 18566 11665
rect 18510 11591 18566 11600
rect 18604 11552 18656 11558
rect 18604 11494 18656 11500
rect 18694 11520 18750 11529
rect 18326 11384 18382 11393
rect 18326 11319 18328 11328
rect 18380 11319 18382 11328
rect 18420 11348 18472 11354
rect 18328 11290 18380 11296
rect 18420 11290 18472 11296
rect 18144 11212 18196 11218
rect 18196 11172 18368 11200
rect 18144 11154 18196 11160
rect 17868 11144 17920 11150
rect 17868 11086 17920 11092
rect 17868 11008 17920 11014
rect 17868 10950 17920 10956
rect 17774 10840 17830 10849
rect 17774 10775 17830 10784
rect 17774 10432 17830 10441
rect 17774 10367 17830 10376
rect 17684 10056 17736 10062
rect 17684 9998 17736 10004
rect 17590 9752 17646 9761
rect 17224 9716 17276 9722
rect 17224 9658 17276 9664
rect 17500 9716 17552 9722
rect 17590 9687 17646 9696
rect 17500 9658 17552 9664
rect 17696 9602 17724 9998
rect 17604 9574 17724 9602
rect 17604 8945 17632 9574
rect 17684 8968 17736 8974
rect 17590 8936 17646 8945
rect 17224 8900 17276 8906
rect 17144 8860 17224 8888
rect 17684 8910 17736 8916
rect 17590 8871 17646 8880
rect 17224 8842 17276 8848
rect 17316 8832 17368 8838
rect 17316 8774 17368 8780
rect 17408 8832 17460 8838
rect 17408 8774 17460 8780
rect 17328 8634 17356 8774
rect 17316 8628 17368 8634
rect 17316 8570 17368 8576
rect 17328 7426 17356 8570
rect 17420 7954 17448 8774
rect 17592 8424 17644 8430
rect 17592 8366 17644 8372
rect 17500 8288 17552 8294
rect 17500 8230 17552 8236
rect 17408 7948 17460 7954
rect 17408 7890 17460 7896
rect 17512 7546 17540 8230
rect 17500 7540 17552 7546
rect 17500 7482 17552 7488
rect 17328 7398 17540 7426
rect 17316 7336 17368 7342
rect 17316 7278 17368 7284
rect 17132 6792 17184 6798
rect 17132 6734 17184 6740
rect 17144 6390 17172 6734
rect 17132 6384 17184 6390
rect 17132 6326 17184 6332
rect 17132 6248 17184 6254
rect 17132 6190 17184 6196
rect 17144 5914 17172 6190
rect 17132 5908 17184 5914
rect 17132 5850 17184 5856
rect 17224 5636 17276 5642
rect 17224 5578 17276 5584
rect 17130 4992 17186 5001
rect 17130 4927 17186 4936
rect 17144 3058 17172 4927
rect 17132 3052 17184 3058
rect 17132 2994 17184 3000
rect 17236 2446 17264 5578
rect 17328 3398 17356 7278
rect 17408 5840 17460 5846
rect 17408 5782 17460 5788
rect 17420 4593 17448 5782
rect 17406 4584 17462 4593
rect 17406 4519 17462 4528
rect 17408 3664 17460 3670
rect 17408 3606 17460 3612
rect 17316 3392 17368 3398
rect 17316 3334 17368 3340
rect 17316 2916 17368 2922
rect 17316 2858 17368 2864
rect 17328 2514 17356 2858
rect 17316 2508 17368 2514
rect 17316 2450 17368 2456
rect 17040 2440 17092 2446
rect 17040 2382 17092 2388
rect 17224 2440 17276 2446
rect 17224 2382 17276 2388
rect 17420 2258 17448 3606
rect 17512 2378 17540 7398
rect 17604 5710 17632 8366
rect 17696 7342 17724 8910
rect 17788 8634 17816 10367
rect 17880 9654 17908 10950
rect 17950 10908 18258 10917
rect 17950 10906 17956 10908
rect 18012 10906 18036 10908
rect 18092 10906 18116 10908
rect 18172 10906 18196 10908
rect 18252 10906 18258 10908
rect 18012 10854 18014 10906
rect 18194 10854 18196 10906
rect 17950 10852 17956 10854
rect 18012 10852 18036 10854
rect 18092 10852 18116 10854
rect 18172 10852 18196 10854
rect 18252 10852 18258 10854
rect 17950 10843 18258 10852
rect 18340 10554 18368 11172
rect 18432 11082 18460 11290
rect 18512 11280 18564 11286
rect 18512 11222 18564 11228
rect 18420 11076 18472 11082
rect 18420 11018 18472 11024
rect 18340 10526 18460 10554
rect 18328 10464 18380 10470
rect 18328 10406 18380 10412
rect 17950 9820 18258 9829
rect 17950 9818 17956 9820
rect 18012 9818 18036 9820
rect 18092 9818 18116 9820
rect 18172 9818 18196 9820
rect 18252 9818 18258 9820
rect 18012 9766 18014 9818
rect 18194 9766 18196 9818
rect 17950 9764 17956 9766
rect 18012 9764 18036 9766
rect 18092 9764 18116 9766
rect 18172 9764 18196 9766
rect 18252 9764 18258 9766
rect 17950 9755 18258 9764
rect 17868 9648 17920 9654
rect 17868 9590 17920 9596
rect 17960 9512 18012 9518
rect 17960 9454 18012 9460
rect 18052 9512 18104 9518
rect 18052 9454 18104 9460
rect 17972 9178 18000 9454
rect 17868 9172 17920 9178
rect 17868 9114 17920 9120
rect 17960 9172 18012 9178
rect 17960 9114 18012 9120
rect 17880 8838 17908 9114
rect 18064 9042 18092 9454
rect 18052 9036 18104 9042
rect 18052 8978 18104 8984
rect 17868 8832 17920 8838
rect 17868 8774 17920 8780
rect 17950 8732 18258 8741
rect 17950 8730 17956 8732
rect 18012 8730 18036 8732
rect 18092 8730 18116 8732
rect 18172 8730 18196 8732
rect 18252 8730 18258 8732
rect 18012 8678 18014 8730
rect 18194 8678 18196 8730
rect 17950 8676 17956 8678
rect 18012 8676 18036 8678
rect 18092 8676 18116 8678
rect 18172 8676 18196 8678
rect 18252 8676 18258 8678
rect 17950 8667 18258 8676
rect 17776 8628 17828 8634
rect 17776 8570 17828 8576
rect 17788 8498 17816 8570
rect 17776 8492 17828 8498
rect 17776 8434 17828 8440
rect 17788 7698 17816 8434
rect 17788 7670 17908 7698
rect 17776 7540 17828 7546
rect 17776 7482 17828 7488
rect 17684 7336 17736 7342
rect 17684 7278 17736 7284
rect 17696 6254 17724 7278
rect 17788 6934 17816 7482
rect 17880 7002 17908 7670
rect 17950 7644 18258 7653
rect 17950 7642 17956 7644
rect 18012 7642 18036 7644
rect 18092 7642 18116 7644
rect 18172 7642 18196 7644
rect 18252 7642 18258 7644
rect 18012 7590 18014 7642
rect 18194 7590 18196 7642
rect 17950 7588 17956 7590
rect 18012 7588 18036 7590
rect 18092 7588 18116 7590
rect 18172 7588 18196 7590
rect 18252 7588 18258 7590
rect 17950 7579 18258 7588
rect 18144 7404 18196 7410
rect 18144 7346 18196 7352
rect 18156 7206 18184 7346
rect 18144 7200 18196 7206
rect 18144 7142 18196 7148
rect 17868 6996 17920 7002
rect 17868 6938 17920 6944
rect 17776 6928 17828 6934
rect 17776 6870 17828 6876
rect 17950 6556 18258 6565
rect 17950 6554 17956 6556
rect 18012 6554 18036 6556
rect 18092 6554 18116 6556
rect 18172 6554 18196 6556
rect 18252 6554 18258 6556
rect 18012 6502 18014 6554
rect 18194 6502 18196 6554
rect 17950 6500 17956 6502
rect 18012 6500 18036 6502
rect 18092 6500 18116 6502
rect 18172 6500 18196 6502
rect 18252 6500 18258 6502
rect 17950 6491 18258 6500
rect 18144 6384 18196 6390
rect 18144 6326 18196 6332
rect 17684 6248 17736 6254
rect 17684 6190 17736 6196
rect 18156 6118 18184 6326
rect 18144 6112 18196 6118
rect 18144 6054 18196 6060
rect 17592 5704 17644 5710
rect 17592 5646 17644 5652
rect 17868 5636 17920 5642
rect 17868 5578 17920 5584
rect 17880 5114 17908 5578
rect 17950 5468 18258 5477
rect 17950 5466 17956 5468
rect 18012 5466 18036 5468
rect 18092 5466 18116 5468
rect 18172 5466 18196 5468
rect 18252 5466 18258 5468
rect 18012 5414 18014 5466
rect 18194 5414 18196 5466
rect 17950 5412 17956 5414
rect 18012 5412 18036 5414
rect 18092 5412 18116 5414
rect 18172 5412 18196 5414
rect 18252 5412 18258 5414
rect 17950 5403 18258 5412
rect 17880 5086 18276 5114
rect 18248 5030 18276 5086
rect 18236 5024 18288 5030
rect 18236 4966 18288 4972
rect 18340 4690 18368 10406
rect 18432 10198 18460 10526
rect 18420 10192 18472 10198
rect 18420 10134 18472 10140
rect 18420 9920 18472 9926
rect 18420 9862 18472 9868
rect 18432 9042 18460 9862
rect 18420 9036 18472 9042
rect 18420 8978 18472 8984
rect 18420 8628 18472 8634
rect 18420 8570 18472 8576
rect 18432 7954 18460 8570
rect 18420 7948 18472 7954
rect 18420 7890 18472 7896
rect 18432 7818 18460 7890
rect 18420 7812 18472 7818
rect 18420 7754 18472 7760
rect 18432 6118 18460 7754
rect 18420 6112 18472 6118
rect 18420 6054 18472 6060
rect 18524 5658 18552 11222
rect 18432 5630 18552 5658
rect 18328 4684 18380 4690
rect 18328 4626 18380 4632
rect 18328 4548 18380 4554
rect 18328 4490 18380 4496
rect 17950 4380 18258 4389
rect 17950 4378 17956 4380
rect 18012 4378 18036 4380
rect 18092 4378 18116 4380
rect 18172 4378 18196 4380
rect 18252 4378 18258 4380
rect 18012 4326 18014 4378
rect 18194 4326 18196 4378
rect 17950 4324 17956 4326
rect 18012 4324 18036 4326
rect 18092 4324 18116 4326
rect 18172 4324 18196 4326
rect 18252 4324 18258 4326
rect 17950 4315 18258 4324
rect 18340 3670 18368 4490
rect 18432 4214 18460 5630
rect 18512 5568 18564 5574
rect 18512 5510 18564 5516
rect 18420 4208 18472 4214
rect 18420 4150 18472 4156
rect 18524 4146 18552 5510
rect 18616 5302 18644 11494
rect 18694 11455 18750 11464
rect 18708 11354 18736 11455
rect 18696 11348 18748 11354
rect 18696 11290 18748 11296
rect 18696 11076 18748 11082
rect 18696 11018 18748 11024
rect 18708 10674 18736 11018
rect 18696 10668 18748 10674
rect 18696 10610 18748 10616
rect 18696 10464 18748 10470
rect 18694 10432 18696 10441
rect 18748 10432 18750 10441
rect 18694 10367 18750 10376
rect 18708 10130 18736 10367
rect 18696 10124 18748 10130
rect 18696 10066 18748 10072
rect 18696 9104 18748 9110
rect 18800 9092 18828 12310
rect 18892 11898 18920 14962
rect 19076 14906 19104 18838
rect 19260 18222 19288 19110
rect 19248 18216 19300 18222
rect 19248 18158 19300 18164
rect 19432 17876 19484 17882
rect 19432 17818 19484 17824
rect 19156 17808 19208 17814
rect 19156 17750 19208 17756
rect 18984 14878 19104 14906
rect 18984 12238 19012 14878
rect 19064 14816 19116 14822
rect 19064 14758 19116 14764
rect 19076 14550 19104 14758
rect 19064 14544 19116 14550
rect 19064 14486 19116 14492
rect 19168 14482 19196 17750
rect 19248 17604 19300 17610
rect 19248 17546 19300 17552
rect 19340 17604 19392 17610
rect 19340 17546 19392 17552
rect 19260 17338 19288 17546
rect 19248 17332 19300 17338
rect 19248 17274 19300 17280
rect 19248 17196 19300 17202
rect 19248 17138 19300 17144
rect 19260 17105 19288 17138
rect 19246 17096 19302 17105
rect 19246 17031 19302 17040
rect 19248 16448 19300 16454
rect 19248 16390 19300 16396
rect 19156 14476 19208 14482
rect 19156 14418 19208 14424
rect 19260 13394 19288 16390
rect 19352 16250 19380 17546
rect 19444 16794 19472 17818
rect 19536 17270 19564 22918
rect 19628 20534 19656 29990
rect 19904 29714 19932 35498
rect 20076 34536 20128 34542
rect 20076 34478 20128 34484
rect 20260 34536 20312 34542
rect 20260 34478 20312 34484
rect 20088 31890 20116 34478
rect 20272 32978 20300 34478
rect 20444 33652 20496 33658
rect 20444 33594 20496 33600
rect 20260 32972 20312 32978
rect 20260 32914 20312 32920
rect 20076 31884 20128 31890
rect 20076 31826 20128 31832
rect 20076 31680 20128 31686
rect 20128 31640 20208 31668
rect 20076 31622 20128 31628
rect 19984 31340 20036 31346
rect 19984 31282 20036 31288
rect 19996 29714 20024 31282
rect 20076 31136 20128 31142
rect 20076 31078 20128 31084
rect 19892 29708 19944 29714
rect 19892 29650 19944 29656
rect 19984 29708 20036 29714
rect 19984 29650 20036 29656
rect 19800 29504 19852 29510
rect 19800 29446 19852 29452
rect 19984 29504 20036 29510
rect 19984 29446 20036 29452
rect 19812 29306 19840 29446
rect 19800 29300 19852 29306
rect 19800 29242 19852 29248
rect 19800 29096 19852 29102
rect 19800 29038 19852 29044
rect 19812 28558 19840 29038
rect 19800 28552 19852 28558
rect 19800 28494 19852 28500
rect 19892 28552 19944 28558
rect 19892 28494 19944 28500
rect 19904 28014 19932 28494
rect 19892 28008 19944 28014
rect 19892 27950 19944 27956
rect 19904 27470 19932 27950
rect 19892 27464 19944 27470
rect 19892 27406 19944 27412
rect 19996 26314 20024 29446
rect 20088 28626 20116 31078
rect 20180 28694 20208 31640
rect 20352 31340 20404 31346
rect 20352 31282 20404 31288
rect 20364 30938 20392 31282
rect 20352 30932 20404 30938
rect 20352 30874 20404 30880
rect 20260 30388 20312 30394
rect 20260 30330 20312 30336
rect 20168 28688 20220 28694
rect 20168 28630 20220 28636
rect 20076 28620 20128 28626
rect 20076 28562 20128 28568
rect 20272 28422 20300 30330
rect 20456 30190 20484 33594
rect 20548 31482 20576 38150
rect 20628 35488 20680 35494
rect 20628 35430 20680 35436
rect 20536 31476 20588 31482
rect 20536 31418 20588 31424
rect 20536 31204 20588 31210
rect 20536 31146 20588 31152
rect 20548 30802 20576 31146
rect 20536 30796 20588 30802
rect 20536 30738 20588 30744
rect 20640 30326 20668 35430
rect 21008 31754 21036 41386
rect 21180 40044 21232 40050
rect 21180 39986 21232 39992
rect 21192 35834 21220 39986
rect 21180 35828 21232 35834
rect 21180 35770 21232 35776
rect 21272 35624 21324 35630
rect 21272 35566 21324 35572
rect 21284 34610 21312 35566
rect 21376 35222 21404 41386
rect 21364 35216 21416 35222
rect 21364 35158 21416 35164
rect 21272 34604 21324 34610
rect 21272 34546 21324 34552
rect 21284 34202 21312 34546
rect 21272 34196 21324 34202
rect 21272 34138 21324 34144
rect 21376 33930 21404 35158
rect 21548 34536 21600 34542
rect 21548 34478 21600 34484
rect 21364 33924 21416 33930
rect 21364 33866 21416 33872
rect 21376 33658 21404 33866
rect 21364 33652 21416 33658
rect 21364 33594 21416 33600
rect 21376 33114 21404 33594
rect 21560 33454 21588 34478
rect 21548 33448 21600 33454
rect 21548 33390 21600 33396
rect 21364 33108 21416 33114
rect 21364 33050 21416 33056
rect 21376 32842 21404 33050
rect 21364 32836 21416 32842
rect 21364 32778 21416 32784
rect 21088 32564 21140 32570
rect 21088 32506 21140 32512
rect 21100 32298 21128 32506
rect 21376 32366 21404 32778
rect 21364 32360 21416 32366
rect 21364 32302 21416 32308
rect 21088 32292 21140 32298
rect 21088 32234 21140 32240
rect 21180 31952 21232 31958
rect 21180 31894 21232 31900
rect 21008 31726 21128 31754
rect 20628 30320 20680 30326
rect 20628 30262 20680 30268
rect 20444 30184 20496 30190
rect 20444 30126 20496 30132
rect 20444 29572 20496 29578
rect 20444 29514 20496 29520
rect 20456 29238 20484 29514
rect 20444 29232 20496 29238
rect 20444 29174 20496 29180
rect 20260 28416 20312 28422
rect 20260 28358 20312 28364
rect 20168 28212 20220 28218
rect 20168 28154 20220 28160
rect 20180 27538 20208 28154
rect 20456 27962 20484 29174
rect 20364 27934 20484 27962
rect 20168 27532 20220 27538
rect 20168 27474 20220 27480
rect 20260 27532 20312 27538
rect 20260 27474 20312 27480
rect 20272 27402 20300 27474
rect 20260 27396 20312 27402
rect 20260 27338 20312 27344
rect 20076 26920 20128 26926
rect 20076 26862 20128 26868
rect 19984 26308 20036 26314
rect 19984 26250 20036 26256
rect 20088 26042 20116 26862
rect 20076 26036 20128 26042
rect 20076 25978 20128 25984
rect 19708 25288 19760 25294
rect 19708 25230 19760 25236
rect 19720 24410 19748 25230
rect 19984 25152 20036 25158
rect 19984 25094 20036 25100
rect 19996 24886 20024 25094
rect 20168 24948 20220 24954
rect 20168 24890 20220 24896
rect 19984 24880 20036 24886
rect 19984 24822 20036 24828
rect 19708 24404 19760 24410
rect 19708 24346 19760 24352
rect 20076 24404 20128 24410
rect 20076 24346 20128 24352
rect 19708 24132 19760 24138
rect 19708 24074 19760 24080
rect 19720 23866 19748 24074
rect 19708 23860 19760 23866
rect 19708 23802 19760 23808
rect 19800 23792 19852 23798
rect 19800 23734 19852 23740
rect 19708 22772 19760 22778
rect 19708 22714 19760 22720
rect 19720 20874 19748 22714
rect 19812 22094 19840 23734
rect 19892 23520 19944 23526
rect 19892 23462 19944 23468
rect 19904 23118 19932 23462
rect 20088 23186 20116 24346
rect 20076 23180 20128 23186
rect 20076 23122 20128 23128
rect 19892 23112 19944 23118
rect 19892 23054 19944 23060
rect 19984 23112 20036 23118
rect 19984 23054 20036 23060
rect 19996 22506 20024 23054
rect 20076 22636 20128 22642
rect 20076 22578 20128 22584
rect 19984 22500 20036 22506
rect 19984 22442 20036 22448
rect 20088 22094 20116 22578
rect 19812 22066 19932 22094
rect 19904 20942 19932 22066
rect 19996 22066 20116 22094
rect 19996 21146 20024 22066
rect 20180 21894 20208 24890
rect 20364 23730 20392 27934
rect 20444 27872 20496 27878
rect 20444 27814 20496 27820
rect 20456 26450 20484 27814
rect 20996 27328 21048 27334
rect 20996 27270 21048 27276
rect 20904 26784 20956 26790
rect 20904 26726 20956 26732
rect 20444 26444 20496 26450
rect 20444 26386 20496 26392
rect 20720 26444 20772 26450
rect 20720 26386 20772 26392
rect 20732 25906 20760 26386
rect 20720 25900 20772 25906
rect 20720 25842 20772 25848
rect 20812 25900 20864 25906
rect 20812 25842 20864 25848
rect 20824 24954 20852 25842
rect 20812 24948 20864 24954
rect 20812 24890 20864 24896
rect 20916 24274 20944 26726
rect 21008 26382 21036 27270
rect 20996 26376 21048 26382
rect 20996 26318 21048 26324
rect 21100 25294 21128 31726
rect 21192 31686 21220 31894
rect 21180 31680 21232 31686
rect 21180 31622 21232 31628
rect 21272 31680 21324 31686
rect 21272 31622 21324 31628
rect 21284 30394 21312 31622
rect 21376 31414 21404 32302
rect 21744 31754 21772 56200
rect 22192 44736 22244 44742
rect 22192 44678 22244 44684
rect 22008 39296 22060 39302
rect 22008 39238 22060 39244
rect 21824 35692 21876 35698
rect 21824 35634 21876 35640
rect 21836 35222 21864 35634
rect 21824 35216 21876 35222
rect 21824 35158 21876 35164
rect 21652 31726 21772 31754
rect 21836 31754 21864 35158
rect 22020 31890 22048 39238
rect 22204 38350 22232 44678
rect 22468 38548 22520 38554
rect 22468 38490 22520 38496
rect 22192 38344 22244 38350
rect 22192 38286 22244 38292
rect 22480 35834 22508 38490
rect 22756 35894 22784 56222
rect 23032 56114 23060 56222
rect 23110 56200 23166 57000
rect 24490 56200 24546 57000
rect 25870 56200 25926 57000
rect 23124 56114 23152 56200
rect 23032 56086 23152 56114
rect 23386 56128 23442 56137
rect 23386 56063 23442 56072
rect 22950 53884 23258 53893
rect 22950 53882 22956 53884
rect 23012 53882 23036 53884
rect 23092 53882 23116 53884
rect 23172 53882 23196 53884
rect 23252 53882 23258 53884
rect 23012 53830 23014 53882
rect 23194 53830 23196 53882
rect 22950 53828 22956 53830
rect 23012 53828 23036 53830
rect 23092 53828 23116 53830
rect 23172 53828 23196 53830
rect 23252 53828 23258 53830
rect 22950 53819 23258 53828
rect 23400 53582 23428 56063
rect 24504 55706 24532 56200
rect 24412 55678 24532 55706
rect 23480 54188 23532 54194
rect 23480 54130 23532 54136
rect 23492 53786 23520 54130
rect 23480 53780 23532 53786
rect 23480 53722 23532 53728
rect 23388 53576 23440 53582
rect 23388 53518 23440 53524
rect 23940 53440 23992 53446
rect 23940 53382 23992 53388
rect 22950 52796 23258 52805
rect 22950 52794 22956 52796
rect 23012 52794 23036 52796
rect 23092 52794 23116 52796
rect 23172 52794 23196 52796
rect 23252 52794 23258 52796
rect 23012 52742 23014 52794
rect 23194 52742 23196 52794
rect 22950 52740 22956 52742
rect 23012 52740 23036 52742
rect 23092 52740 23116 52742
rect 23172 52740 23196 52742
rect 23252 52740 23258 52742
rect 22950 52731 23258 52740
rect 22950 51708 23258 51717
rect 22950 51706 22956 51708
rect 23012 51706 23036 51708
rect 23092 51706 23116 51708
rect 23172 51706 23196 51708
rect 23252 51706 23258 51708
rect 23012 51654 23014 51706
rect 23194 51654 23196 51706
rect 22950 51652 22956 51654
rect 23012 51652 23036 51654
rect 23092 51652 23116 51654
rect 23172 51652 23196 51654
rect 23252 51652 23258 51654
rect 22950 51643 23258 51652
rect 22950 50620 23258 50629
rect 22950 50618 22956 50620
rect 23012 50618 23036 50620
rect 23092 50618 23116 50620
rect 23172 50618 23196 50620
rect 23252 50618 23258 50620
rect 23012 50566 23014 50618
rect 23194 50566 23196 50618
rect 22950 50564 22956 50566
rect 23012 50564 23036 50566
rect 23092 50564 23116 50566
rect 23172 50564 23196 50566
rect 23252 50564 23258 50566
rect 22950 50555 23258 50564
rect 22950 49532 23258 49541
rect 22950 49530 22956 49532
rect 23012 49530 23036 49532
rect 23092 49530 23116 49532
rect 23172 49530 23196 49532
rect 23252 49530 23258 49532
rect 23012 49478 23014 49530
rect 23194 49478 23196 49530
rect 22950 49476 22956 49478
rect 23012 49476 23036 49478
rect 23092 49476 23116 49478
rect 23172 49476 23196 49478
rect 23252 49476 23258 49478
rect 22950 49467 23258 49476
rect 22950 48444 23258 48453
rect 22950 48442 22956 48444
rect 23012 48442 23036 48444
rect 23092 48442 23116 48444
rect 23172 48442 23196 48444
rect 23252 48442 23258 48444
rect 23012 48390 23014 48442
rect 23194 48390 23196 48442
rect 22950 48388 22956 48390
rect 23012 48388 23036 48390
rect 23092 48388 23116 48390
rect 23172 48388 23196 48390
rect 23252 48388 23258 48390
rect 22950 48379 23258 48388
rect 22950 47356 23258 47365
rect 22950 47354 22956 47356
rect 23012 47354 23036 47356
rect 23092 47354 23116 47356
rect 23172 47354 23196 47356
rect 23252 47354 23258 47356
rect 23012 47302 23014 47354
rect 23194 47302 23196 47354
rect 22950 47300 22956 47302
rect 23012 47300 23036 47302
rect 23092 47300 23116 47302
rect 23172 47300 23196 47302
rect 23252 47300 23258 47302
rect 22950 47291 23258 47300
rect 23296 46368 23348 46374
rect 23296 46310 23348 46316
rect 22950 46268 23258 46277
rect 22950 46266 22956 46268
rect 23012 46266 23036 46268
rect 23092 46266 23116 46268
rect 23172 46266 23196 46268
rect 23252 46266 23258 46268
rect 23012 46214 23014 46266
rect 23194 46214 23196 46266
rect 22950 46212 22956 46214
rect 23012 46212 23036 46214
rect 23092 46212 23116 46214
rect 23172 46212 23196 46214
rect 23252 46212 23258 46214
rect 22950 46203 23258 46212
rect 22950 45180 23258 45189
rect 22950 45178 22956 45180
rect 23012 45178 23036 45180
rect 23092 45178 23116 45180
rect 23172 45178 23196 45180
rect 23252 45178 23258 45180
rect 23012 45126 23014 45178
rect 23194 45126 23196 45178
rect 22950 45124 22956 45126
rect 23012 45124 23036 45126
rect 23092 45124 23116 45126
rect 23172 45124 23196 45126
rect 23252 45124 23258 45126
rect 22950 45115 23258 45124
rect 22950 44092 23258 44101
rect 22950 44090 22956 44092
rect 23012 44090 23036 44092
rect 23092 44090 23116 44092
rect 23172 44090 23196 44092
rect 23252 44090 23258 44092
rect 23012 44038 23014 44090
rect 23194 44038 23196 44090
rect 22950 44036 22956 44038
rect 23012 44036 23036 44038
rect 23092 44036 23116 44038
rect 23172 44036 23196 44038
rect 23252 44036 23258 44038
rect 22950 44027 23258 44036
rect 22950 43004 23258 43013
rect 22950 43002 22956 43004
rect 23012 43002 23036 43004
rect 23092 43002 23116 43004
rect 23172 43002 23196 43004
rect 23252 43002 23258 43004
rect 23012 42950 23014 43002
rect 23194 42950 23196 43002
rect 22950 42948 22956 42950
rect 23012 42948 23036 42950
rect 23092 42948 23116 42950
rect 23172 42948 23196 42950
rect 23252 42948 23258 42950
rect 22950 42939 23258 42948
rect 22950 41916 23258 41925
rect 22950 41914 22956 41916
rect 23012 41914 23036 41916
rect 23092 41914 23116 41916
rect 23172 41914 23196 41916
rect 23252 41914 23258 41916
rect 23012 41862 23014 41914
rect 23194 41862 23196 41914
rect 22950 41860 22956 41862
rect 23012 41860 23036 41862
rect 23092 41860 23116 41862
rect 23172 41860 23196 41862
rect 23252 41860 23258 41862
rect 22950 41851 23258 41860
rect 22950 40828 23258 40837
rect 22950 40826 22956 40828
rect 23012 40826 23036 40828
rect 23092 40826 23116 40828
rect 23172 40826 23196 40828
rect 23252 40826 23258 40828
rect 23012 40774 23014 40826
rect 23194 40774 23196 40826
rect 22950 40772 22956 40774
rect 23012 40772 23036 40774
rect 23092 40772 23116 40774
rect 23172 40772 23196 40774
rect 23252 40772 23258 40774
rect 22950 40763 23258 40772
rect 23308 40050 23336 46310
rect 23480 44736 23532 44742
rect 23480 44678 23532 44684
rect 23296 40044 23348 40050
rect 23296 39986 23348 39992
rect 22950 39740 23258 39749
rect 22950 39738 22956 39740
rect 23012 39738 23036 39740
rect 23092 39738 23116 39740
rect 23172 39738 23196 39740
rect 23252 39738 23258 39740
rect 23012 39686 23014 39738
rect 23194 39686 23196 39738
rect 22950 39684 22956 39686
rect 23012 39684 23036 39686
rect 23092 39684 23116 39686
rect 23172 39684 23196 39686
rect 23252 39684 23258 39686
rect 22950 39675 23258 39684
rect 22950 38652 23258 38661
rect 22950 38650 22956 38652
rect 23012 38650 23036 38652
rect 23092 38650 23116 38652
rect 23172 38650 23196 38652
rect 23252 38650 23258 38652
rect 23012 38598 23014 38650
rect 23194 38598 23196 38650
rect 22950 38596 22956 38598
rect 23012 38596 23036 38598
rect 23092 38596 23116 38598
rect 23172 38596 23196 38598
rect 23252 38596 23258 38598
rect 22950 38587 23258 38596
rect 22950 37564 23258 37573
rect 22950 37562 22956 37564
rect 23012 37562 23036 37564
rect 23092 37562 23116 37564
rect 23172 37562 23196 37564
rect 23252 37562 23258 37564
rect 23012 37510 23014 37562
rect 23194 37510 23196 37562
rect 22950 37508 22956 37510
rect 23012 37508 23036 37510
rect 23092 37508 23116 37510
rect 23172 37508 23196 37510
rect 23252 37508 23258 37510
rect 22950 37499 23258 37508
rect 22950 36476 23258 36485
rect 22950 36474 22956 36476
rect 23012 36474 23036 36476
rect 23092 36474 23116 36476
rect 23172 36474 23196 36476
rect 23252 36474 23258 36476
rect 23012 36422 23014 36474
rect 23194 36422 23196 36474
rect 22950 36420 22956 36422
rect 23012 36420 23036 36422
rect 23092 36420 23116 36422
rect 23172 36420 23196 36422
rect 23252 36420 23258 36422
rect 22950 36411 23258 36420
rect 23492 35894 23520 44678
rect 23952 41478 23980 53382
rect 24412 50454 24440 55678
rect 24490 55448 24546 55457
rect 24490 55383 24546 55392
rect 24504 54330 24532 55383
rect 24674 54632 24730 54641
rect 24674 54567 24730 54576
rect 24492 54324 24544 54330
rect 24492 54266 24544 54272
rect 24688 53582 24716 54567
rect 24768 54188 24820 54194
rect 24768 54130 24820 54136
rect 24780 53825 24808 54130
rect 24766 53816 24822 53825
rect 25884 53786 25912 56200
rect 26792 53984 26844 53990
rect 26792 53926 26844 53932
rect 24766 53751 24822 53760
rect 25872 53780 25924 53786
rect 25872 53722 25924 53728
rect 24676 53576 24728 53582
rect 24676 53518 24728 53524
rect 24860 53440 24912 53446
rect 24860 53382 24912 53388
rect 24400 50448 24452 50454
rect 24400 50390 24452 50396
rect 24216 46096 24268 46102
rect 24216 46038 24268 46044
rect 23940 41472 23992 41478
rect 23940 41414 23992 41420
rect 24228 38554 24256 46038
rect 24768 44396 24820 44402
rect 24768 44338 24820 44344
rect 24780 44033 24808 44338
rect 24766 44024 24822 44033
rect 24766 43959 24822 43968
rect 24216 38548 24268 38554
rect 24216 38490 24268 38496
rect 24768 36032 24820 36038
rect 24768 35974 24820 35980
rect 24780 35894 24808 35974
rect 22664 35866 22784 35894
rect 23400 35866 23520 35894
rect 24688 35866 24808 35894
rect 22468 35828 22520 35834
rect 22468 35770 22520 35776
rect 22100 35624 22152 35630
rect 22100 35566 22152 35572
rect 22112 34610 22140 35566
rect 22192 35080 22244 35086
rect 22192 35022 22244 35028
rect 22100 34604 22152 34610
rect 22100 34546 22152 34552
rect 22112 34202 22140 34546
rect 22100 34196 22152 34202
rect 22100 34138 22152 34144
rect 22100 32428 22152 32434
rect 22100 32370 22152 32376
rect 22112 32230 22140 32370
rect 22100 32224 22152 32230
rect 22100 32166 22152 32172
rect 22008 31884 22060 31890
rect 22008 31826 22060 31832
rect 21836 31726 22048 31754
rect 21364 31408 21416 31414
rect 21364 31350 21416 31356
rect 21272 30388 21324 30394
rect 21272 30330 21324 30336
rect 21456 30048 21508 30054
rect 21456 29990 21508 29996
rect 21180 29028 21232 29034
rect 21180 28970 21232 28976
rect 21192 27674 21220 28970
rect 21180 27668 21232 27674
rect 21180 27610 21232 27616
rect 21180 27328 21232 27334
rect 21180 27270 21232 27276
rect 21192 26994 21220 27270
rect 21180 26988 21232 26994
rect 21180 26930 21232 26936
rect 21088 25288 21140 25294
rect 21088 25230 21140 25236
rect 20996 25152 21048 25158
rect 20996 25094 21048 25100
rect 21008 24993 21036 25094
rect 20994 24984 21050 24993
rect 20994 24919 21050 24928
rect 21192 24698 21220 26930
rect 21272 26920 21324 26926
rect 21272 26862 21324 26868
rect 21284 26450 21312 26862
rect 21272 26444 21324 26450
rect 21272 26386 21324 26392
rect 21468 25378 21496 29990
rect 21548 27396 21600 27402
rect 21548 27338 21600 27344
rect 21560 26908 21588 27338
rect 21652 27062 21680 31726
rect 22020 31686 22048 31726
rect 22008 31680 22060 31686
rect 22008 31622 22060 31628
rect 22020 31482 22048 31622
rect 22008 31476 22060 31482
rect 22008 31418 22060 31424
rect 21732 31408 21784 31414
rect 21732 31350 21784 31356
rect 21744 30666 21772 31350
rect 21732 30660 21784 30666
rect 21732 30602 21784 30608
rect 22112 29714 22140 32166
rect 22204 31346 22232 35022
rect 22468 34944 22520 34950
rect 22468 34886 22520 34892
rect 22284 34060 22336 34066
rect 22284 34002 22336 34008
rect 22296 33590 22324 34002
rect 22376 33924 22428 33930
rect 22376 33866 22428 33872
rect 22388 33658 22416 33866
rect 22376 33652 22428 33658
rect 22376 33594 22428 33600
rect 22284 33584 22336 33590
rect 22284 33526 22336 33532
rect 22296 32978 22324 33526
rect 22284 32972 22336 32978
rect 22284 32914 22336 32920
rect 22296 32502 22324 32914
rect 22284 32496 22336 32502
rect 22284 32438 22336 32444
rect 22284 31476 22336 31482
rect 22284 31418 22336 31424
rect 22192 31340 22244 31346
rect 22192 31282 22244 31288
rect 22100 29708 22152 29714
rect 22100 29650 22152 29656
rect 22112 28234 22140 29650
rect 22192 28484 22244 28490
rect 22192 28426 22244 28432
rect 22204 28234 22232 28426
rect 22112 28206 22232 28234
rect 22204 28150 22232 28206
rect 22192 28144 22244 28150
rect 22192 28086 22244 28092
rect 21916 28008 21968 28014
rect 22098 27976 22154 27985
rect 21968 27956 22048 27962
rect 21916 27950 22048 27956
rect 21928 27934 22048 27950
rect 22020 27860 22048 27934
rect 22098 27911 22154 27920
rect 22112 27860 22140 27911
rect 22020 27832 22140 27860
rect 22296 27470 22324 31418
rect 22376 31340 22428 31346
rect 22376 31282 22428 31288
rect 22388 30394 22416 31282
rect 22376 30388 22428 30394
rect 22376 30330 22428 30336
rect 22480 30326 22508 34886
rect 22560 32836 22612 32842
rect 22560 32778 22612 32784
rect 22572 32026 22600 32778
rect 22560 32020 22612 32026
rect 22560 31962 22612 31968
rect 22468 30320 22520 30326
rect 22468 30262 22520 30268
rect 22664 29850 22692 35866
rect 22836 35828 22888 35834
rect 22836 35770 22888 35776
rect 22744 31272 22796 31278
rect 22744 31214 22796 31220
rect 22756 30938 22784 31214
rect 22744 30932 22796 30938
rect 22744 30874 22796 30880
rect 22652 29844 22704 29850
rect 22652 29786 22704 29792
rect 22848 29782 22876 35770
rect 22950 35388 23258 35397
rect 22950 35386 22956 35388
rect 23012 35386 23036 35388
rect 23092 35386 23116 35388
rect 23172 35386 23196 35388
rect 23252 35386 23258 35388
rect 23012 35334 23014 35386
rect 23194 35334 23196 35386
rect 22950 35332 22956 35334
rect 23012 35332 23036 35334
rect 23092 35332 23116 35334
rect 23172 35332 23196 35334
rect 23252 35332 23258 35334
rect 22950 35323 23258 35332
rect 23296 35148 23348 35154
rect 23296 35090 23348 35096
rect 23308 34610 23336 35090
rect 23400 35086 23428 35866
rect 24124 35216 24176 35222
rect 24688 35193 24716 35866
rect 24768 35488 24820 35494
rect 24768 35430 24820 35436
rect 24124 35158 24176 35164
rect 24674 35184 24730 35193
rect 23388 35080 23440 35086
rect 23388 35022 23440 35028
rect 23664 34740 23716 34746
rect 23664 34682 23716 34688
rect 23296 34604 23348 34610
rect 23296 34546 23348 34552
rect 22950 34300 23258 34309
rect 22950 34298 22956 34300
rect 23012 34298 23036 34300
rect 23092 34298 23116 34300
rect 23172 34298 23196 34300
rect 23252 34298 23258 34300
rect 23012 34246 23014 34298
rect 23194 34246 23196 34298
rect 22950 34244 22956 34246
rect 23012 34244 23036 34246
rect 23092 34244 23116 34246
rect 23172 34244 23196 34246
rect 23252 34244 23258 34246
rect 22950 34235 23258 34244
rect 22950 33212 23258 33221
rect 22950 33210 22956 33212
rect 23012 33210 23036 33212
rect 23092 33210 23116 33212
rect 23172 33210 23196 33212
rect 23252 33210 23258 33212
rect 23012 33158 23014 33210
rect 23194 33158 23196 33210
rect 22950 33156 22956 33158
rect 23012 33156 23036 33158
rect 23092 33156 23116 33158
rect 23172 33156 23196 33158
rect 23252 33156 23258 33158
rect 22950 33147 23258 33156
rect 23308 33114 23336 34546
rect 23480 33992 23532 33998
rect 23480 33934 23532 33940
rect 23492 33318 23520 33934
rect 23572 33856 23624 33862
rect 23572 33798 23624 33804
rect 23584 33658 23612 33798
rect 23572 33652 23624 33658
rect 23572 33594 23624 33600
rect 23480 33312 23532 33318
rect 23480 33254 23532 33260
rect 23296 33108 23348 33114
rect 23296 33050 23348 33056
rect 22950 32124 23258 32133
rect 22950 32122 22956 32124
rect 23012 32122 23036 32124
rect 23092 32122 23116 32124
rect 23172 32122 23196 32124
rect 23252 32122 23258 32124
rect 23012 32070 23014 32122
rect 23194 32070 23196 32122
rect 22950 32068 22956 32070
rect 23012 32068 23036 32070
rect 23092 32068 23116 32070
rect 23172 32068 23196 32070
rect 23252 32068 23258 32070
rect 22950 32059 23258 32068
rect 23296 31816 23348 31822
rect 23296 31758 23348 31764
rect 22950 31036 23258 31045
rect 22950 31034 22956 31036
rect 23012 31034 23036 31036
rect 23092 31034 23116 31036
rect 23172 31034 23196 31036
rect 23252 31034 23258 31036
rect 23012 30982 23014 31034
rect 23194 30982 23196 31034
rect 22950 30980 22956 30982
rect 23012 30980 23036 30982
rect 23092 30980 23116 30982
rect 23172 30980 23196 30982
rect 23252 30980 23258 30982
rect 22950 30971 23258 30980
rect 23308 30802 23336 31758
rect 23296 30796 23348 30802
rect 23296 30738 23348 30744
rect 23492 30326 23520 33254
rect 23584 32842 23612 33594
rect 23572 32836 23624 32842
rect 23572 32778 23624 32784
rect 23572 30660 23624 30666
rect 23572 30602 23624 30608
rect 23584 30326 23612 30602
rect 23480 30320 23532 30326
rect 23480 30262 23532 30268
rect 23572 30320 23624 30326
rect 23572 30262 23624 30268
rect 23296 30184 23348 30190
rect 23296 30126 23348 30132
rect 22950 29948 23258 29957
rect 22950 29946 22956 29948
rect 23012 29946 23036 29948
rect 23092 29946 23116 29948
rect 23172 29946 23196 29948
rect 23252 29946 23258 29948
rect 23012 29894 23014 29946
rect 23194 29894 23196 29946
rect 22950 29892 22956 29894
rect 23012 29892 23036 29894
rect 23092 29892 23116 29894
rect 23172 29892 23196 29894
rect 23252 29892 23258 29894
rect 22950 29883 23258 29892
rect 22836 29776 22888 29782
rect 22836 29718 22888 29724
rect 22468 29640 22520 29646
rect 22468 29582 22520 29588
rect 22284 27464 22336 27470
rect 22204 27412 22284 27418
rect 22204 27406 22336 27412
rect 22204 27390 22324 27406
rect 21640 27056 21692 27062
rect 21640 26998 21692 27004
rect 21560 26880 21680 26908
rect 21652 26790 21680 26880
rect 21822 26888 21878 26897
rect 21822 26823 21878 26832
rect 21640 26784 21692 26790
rect 21640 26726 21692 26732
rect 21548 26444 21600 26450
rect 21548 26386 21600 26392
rect 21376 25350 21496 25378
rect 21272 24880 21324 24886
rect 21272 24822 21324 24828
rect 21008 24670 21220 24698
rect 20904 24268 20956 24274
rect 20904 24210 20956 24216
rect 20352 23724 20404 23730
rect 20352 23666 20404 23672
rect 20812 23724 20864 23730
rect 20812 23666 20864 23672
rect 20364 22438 20392 23666
rect 20536 23520 20588 23526
rect 20536 23462 20588 23468
rect 20352 22432 20404 22438
rect 20352 22374 20404 22380
rect 20444 22160 20496 22166
rect 20444 22102 20496 22108
rect 20352 21956 20404 21962
rect 20352 21898 20404 21904
rect 20168 21888 20220 21894
rect 20220 21848 20300 21876
rect 20168 21830 20220 21836
rect 20168 21684 20220 21690
rect 20168 21626 20220 21632
rect 19984 21140 20036 21146
rect 19984 21082 20036 21088
rect 20180 21026 20208 21626
rect 20272 21146 20300 21848
rect 20260 21140 20312 21146
rect 20260 21082 20312 21088
rect 19984 21004 20036 21010
rect 19984 20946 20036 20952
rect 20088 20998 20208 21026
rect 19892 20936 19944 20942
rect 19892 20878 19944 20884
rect 19708 20868 19760 20874
rect 19708 20810 19760 20816
rect 19800 20800 19852 20806
rect 19800 20742 19852 20748
rect 19616 20528 19668 20534
rect 19616 20470 19668 20476
rect 19616 20392 19668 20398
rect 19616 20334 19668 20340
rect 19628 20262 19656 20334
rect 19616 20256 19668 20262
rect 19616 20198 19668 20204
rect 19628 19718 19656 20198
rect 19616 19712 19668 19718
rect 19616 19654 19668 19660
rect 19708 19168 19760 19174
rect 19708 19110 19760 19116
rect 19720 18630 19748 19110
rect 19708 18624 19760 18630
rect 19708 18566 19760 18572
rect 19616 18080 19668 18086
rect 19616 18022 19668 18028
rect 19524 17264 19576 17270
rect 19524 17206 19576 17212
rect 19432 16788 19484 16794
rect 19432 16730 19484 16736
rect 19444 16697 19472 16730
rect 19430 16688 19486 16697
rect 19430 16623 19486 16632
rect 19340 16244 19392 16250
rect 19340 16186 19392 16192
rect 19340 15904 19392 15910
rect 19340 15846 19392 15852
rect 19352 15502 19380 15846
rect 19340 15496 19392 15502
rect 19340 15438 19392 15444
rect 19524 15360 19576 15366
rect 19524 15302 19576 15308
rect 19432 14884 19484 14890
rect 19432 14826 19484 14832
rect 19444 14618 19472 14826
rect 19432 14612 19484 14618
rect 19432 14554 19484 14560
rect 19340 14544 19392 14550
rect 19340 14486 19392 14492
rect 19352 14414 19380 14486
rect 19340 14408 19392 14414
rect 19340 14350 19392 14356
rect 19432 14272 19484 14278
rect 19432 14214 19484 14220
rect 19444 14006 19472 14214
rect 19432 14000 19484 14006
rect 19432 13942 19484 13948
rect 19340 13728 19392 13734
rect 19340 13670 19392 13676
rect 19248 13388 19300 13394
rect 19248 13330 19300 13336
rect 19352 13274 19380 13670
rect 19536 13410 19564 15302
rect 19260 13246 19380 13274
rect 19444 13382 19564 13410
rect 19064 12844 19116 12850
rect 19064 12786 19116 12792
rect 19076 12434 19104 12786
rect 19260 12782 19288 13246
rect 19340 13184 19392 13190
rect 19340 13126 19392 13132
rect 19248 12776 19300 12782
rect 19248 12718 19300 12724
rect 19076 12406 19288 12434
rect 18972 12232 19024 12238
rect 18972 12174 19024 12180
rect 19156 12164 19208 12170
rect 19156 12106 19208 12112
rect 18972 12096 19024 12102
rect 18972 12038 19024 12044
rect 18880 11892 18932 11898
rect 18880 11834 18932 11840
rect 18984 11286 19012 12038
rect 19168 11898 19196 12106
rect 19156 11892 19208 11898
rect 19156 11834 19208 11840
rect 19064 11756 19116 11762
rect 19064 11698 19116 11704
rect 19076 11354 19104 11698
rect 19168 11626 19196 11834
rect 19156 11620 19208 11626
rect 19156 11562 19208 11568
rect 19154 11384 19210 11393
rect 19064 11348 19116 11354
rect 19154 11319 19210 11328
rect 19064 11290 19116 11296
rect 18972 11280 19024 11286
rect 18972 11222 19024 11228
rect 19076 11098 19104 11290
rect 19168 11218 19196 11319
rect 19156 11212 19208 11218
rect 19156 11154 19208 11160
rect 18984 11070 19104 11098
rect 18880 10192 18932 10198
rect 18880 10134 18932 10140
rect 18892 10062 18920 10134
rect 18880 10056 18932 10062
rect 18880 9998 18932 10004
rect 18748 9064 18828 9092
rect 18696 9046 18748 9052
rect 18708 7886 18736 9046
rect 18788 8560 18840 8566
rect 18788 8502 18840 8508
rect 18800 8430 18828 8502
rect 18788 8424 18840 8430
rect 18786 8392 18788 8401
rect 18840 8392 18842 8401
rect 18786 8327 18842 8336
rect 18892 8090 18920 9998
rect 18984 9518 19012 11070
rect 19062 10976 19118 10985
rect 19062 10911 19118 10920
rect 19076 10674 19104 10911
rect 19064 10668 19116 10674
rect 19064 10610 19116 10616
rect 19156 10464 19208 10470
rect 19156 10406 19208 10412
rect 18972 9512 19024 9518
rect 18972 9454 19024 9460
rect 19064 9376 19116 9382
rect 19064 9318 19116 9324
rect 18970 8936 19026 8945
rect 18970 8871 19026 8880
rect 18984 8650 19012 8871
rect 19076 8838 19104 9318
rect 19064 8832 19116 8838
rect 19064 8774 19116 8780
rect 18984 8622 19104 8650
rect 18880 8084 18932 8090
rect 18880 8026 18932 8032
rect 18696 7880 18748 7886
rect 18696 7822 18748 7828
rect 18788 7744 18840 7750
rect 18788 7686 18840 7692
rect 18800 7410 18828 7686
rect 18788 7404 18840 7410
rect 18788 7346 18840 7352
rect 18972 6724 19024 6730
rect 18972 6666 19024 6672
rect 18696 5636 18748 5642
rect 18696 5578 18748 5584
rect 18604 5296 18656 5302
rect 18604 5238 18656 5244
rect 18604 5160 18656 5166
rect 18604 5102 18656 5108
rect 18512 4140 18564 4146
rect 18512 4082 18564 4088
rect 18420 4072 18472 4078
rect 18420 4014 18472 4020
rect 18328 3664 18380 3670
rect 18328 3606 18380 3612
rect 17684 3596 17736 3602
rect 17684 3538 17736 3544
rect 17592 3460 17644 3466
rect 17592 3402 17644 3408
rect 17604 2961 17632 3402
rect 17590 2952 17646 2961
rect 17590 2887 17646 2896
rect 17500 2372 17552 2378
rect 17500 2314 17552 2320
rect 17328 2230 17448 2258
rect 17328 800 17356 2230
rect 17696 800 17724 3538
rect 17950 3292 18258 3301
rect 17950 3290 17956 3292
rect 18012 3290 18036 3292
rect 18092 3290 18116 3292
rect 18172 3290 18196 3292
rect 18252 3290 18258 3292
rect 18012 3238 18014 3290
rect 18194 3238 18196 3290
rect 17950 3236 17956 3238
rect 18012 3236 18036 3238
rect 18092 3236 18116 3238
rect 18172 3236 18196 3238
rect 18252 3236 18258 3238
rect 17950 3227 18258 3236
rect 17950 2204 18258 2213
rect 17950 2202 17956 2204
rect 18012 2202 18036 2204
rect 18092 2202 18116 2204
rect 18172 2202 18196 2204
rect 18252 2202 18258 2204
rect 18012 2150 18014 2202
rect 18194 2150 18196 2202
rect 17950 2148 17956 2150
rect 18012 2148 18036 2150
rect 18092 2148 18116 2150
rect 18172 2148 18196 2150
rect 18252 2148 18258 2150
rect 17950 2139 18258 2148
rect 18432 1170 18460 4014
rect 18616 3738 18644 5102
rect 18604 3732 18656 3738
rect 18604 3674 18656 3680
rect 18708 3670 18736 5578
rect 18788 4684 18840 4690
rect 18788 4626 18840 4632
rect 18696 3664 18748 3670
rect 18696 3606 18748 3612
rect 18512 1828 18564 1834
rect 18512 1770 18564 1776
rect 18340 1142 18460 1170
rect 18064 870 18184 898
rect 18064 800 18092 870
rect 7852 734 8064 762
rect 8114 0 8170 800
rect 8482 0 8538 800
rect 8850 0 8906 800
rect 9218 0 9274 800
rect 9586 0 9642 800
rect 9954 0 10010 800
rect 10322 0 10378 800
rect 10690 0 10746 800
rect 11058 0 11114 800
rect 11426 0 11482 800
rect 11794 0 11850 800
rect 12162 0 12218 800
rect 12530 0 12586 800
rect 12898 0 12954 800
rect 13266 0 13322 800
rect 13634 0 13690 800
rect 14002 0 14058 800
rect 14370 0 14426 800
rect 14738 0 14794 800
rect 15106 0 15162 800
rect 15474 0 15530 800
rect 15842 0 15898 800
rect 16210 0 16266 800
rect 16578 0 16634 800
rect 16946 0 17002 800
rect 17314 0 17370 800
rect 17682 0 17738 800
rect 18050 0 18106 800
rect 18156 762 18184 870
rect 18340 762 18368 1142
rect 18524 1034 18552 1770
rect 18432 1006 18552 1034
rect 18432 800 18460 1006
rect 18800 800 18828 4626
rect 18984 3398 19012 6666
rect 19076 4554 19104 8622
rect 19168 4622 19196 10406
rect 19260 9926 19288 12406
rect 19352 11506 19380 13126
rect 19444 12102 19472 13382
rect 19522 13288 19578 13297
rect 19522 13223 19524 13232
rect 19576 13223 19578 13232
rect 19524 13194 19576 13200
rect 19432 12096 19484 12102
rect 19432 12038 19484 12044
rect 19444 11694 19472 12038
rect 19432 11688 19484 11694
rect 19432 11630 19484 11636
rect 19352 11478 19564 11506
rect 19432 11348 19484 11354
rect 19432 11290 19484 11296
rect 19340 11212 19392 11218
rect 19340 11154 19392 11160
rect 19352 11014 19380 11154
rect 19340 11008 19392 11014
rect 19340 10950 19392 10956
rect 19248 9920 19300 9926
rect 19248 9862 19300 9868
rect 19248 9648 19300 9654
rect 19248 9590 19300 9596
rect 19260 8838 19288 9590
rect 19248 8832 19300 8838
rect 19248 8774 19300 8780
rect 19260 8634 19288 8774
rect 19248 8628 19300 8634
rect 19248 8570 19300 8576
rect 19248 8356 19300 8362
rect 19248 8298 19300 8304
rect 19156 4616 19208 4622
rect 19156 4558 19208 4564
rect 19064 4548 19116 4554
rect 19064 4490 19116 4496
rect 19064 4208 19116 4214
rect 19064 4150 19116 4156
rect 18880 3392 18932 3398
rect 18880 3334 18932 3340
rect 18972 3392 19024 3398
rect 18972 3334 19024 3340
rect 18892 2446 18920 3334
rect 18880 2440 18932 2446
rect 18880 2382 18932 2388
rect 19076 2310 19104 4150
rect 19260 4078 19288 8298
rect 19340 6316 19392 6322
rect 19340 6258 19392 6264
rect 19352 5098 19380 6258
rect 19340 5092 19392 5098
rect 19340 5034 19392 5040
rect 19248 4072 19300 4078
rect 19248 4014 19300 4020
rect 19156 3460 19208 3466
rect 19156 3402 19208 3408
rect 19064 2304 19116 2310
rect 19064 2246 19116 2252
rect 19168 800 19196 3402
rect 19248 3052 19300 3058
rect 19444 3040 19472 11290
rect 19536 5001 19564 11478
rect 19628 10742 19656 18022
rect 19708 16516 19760 16522
rect 19708 16458 19760 16464
rect 19720 16046 19748 16458
rect 19708 16040 19760 16046
rect 19708 15982 19760 15988
rect 19720 15570 19748 15982
rect 19708 15564 19760 15570
rect 19708 15506 19760 15512
rect 19812 15162 19840 20742
rect 19904 20602 19932 20878
rect 19892 20596 19944 20602
rect 19892 20538 19944 20544
rect 19892 20324 19944 20330
rect 19892 20266 19944 20272
rect 19904 19922 19932 20266
rect 19892 19916 19944 19922
rect 19892 19858 19944 19864
rect 19996 16538 20024 20946
rect 20088 18714 20116 20998
rect 20168 19780 20220 19786
rect 20168 19722 20220 19728
rect 20180 18902 20208 19722
rect 20260 19440 20312 19446
rect 20260 19382 20312 19388
rect 20168 18896 20220 18902
rect 20168 18838 20220 18844
rect 20088 18686 20208 18714
rect 20076 18624 20128 18630
rect 20076 18566 20128 18572
rect 20088 18426 20116 18566
rect 20076 18420 20128 18426
rect 20076 18362 20128 18368
rect 20076 18080 20128 18086
rect 20076 18022 20128 18028
rect 19904 16510 20024 16538
rect 19904 15366 19932 16510
rect 19984 16448 20036 16454
rect 19984 16390 20036 16396
rect 19996 16182 20024 16390
rect 19984 16176 20036 16182
rect 19984 16118 20036 16124
rect 19892 15360 19944 15366
rect 19892 15302 19944 15308
rect 19800 15156 19852 15162
rect 19800 15098 19852 15104
rect 19800 14952 19852 14958
rect 19800 14894 19852 14900
rect 19982 14920 20038 14929
rect 19708 14884 19760 14890
rect 19708 14826 19760 14832
rect 19720 11626 19748 14826
rect 19812 14482 19840 14894
rect 19982 14855 20038 14864
rect 19800 14476 19852 14482
rect 19800 14418 19852 14424
rect 19800 14340 19852 14346
rect 19800 14282 19852 14288
rect 19812 14074 19840 14282
rect 19892 14272 19944 14278
rect 19892 14214 19944 14220
rect 19800 14068 19852 14074
rect 19800 14010 19852 14016
rect 19708 11620 19760 11626
rect 19708 11562 19760 11568
rect 19708 11280 19760 11286
rect 19708 11222 19760 11228
rect 19616 10736 19668 10742
rect 19616 10678 19668 10684
rect 19720 10674 19748 11222
rect 19800 11008 19852 11014
rect 19800 10950 19852 10956
rect 19708 10668 19760 10674
rect 19708 10610 19760 10616
rect 19708 10532 19760 10538
rect 19708 10474 19760 10480
rect 19616 10260 19668 10266
rect 19616 10202 19668 10208
rect 19628 9654 19656 10202
rect 19616 9648 19668 9654
rect 19616 9590 19668 9596
rect 19720 8922 19748 10474
rect 19812 10266 19840 10950
rect 19800 10260 19852 10266
rect 19800 10202 19852 10208
rect 19904 10146 19932 14214
rect 19996 11218 20024 14855
rect 20088 14550 20116 18022
rect 20180 15910 20208 18686
rect 20272 18290 20300 19382
rect 20260 18284 20312 18290
rect 20260 18226 20312 18232
rect 20168 15904 20220 15910
rect 20168 15846 20220 15852
rect 20364 15162 20392 21898
rect 20456 21536 20484 22102
rect 20548 21690 20576 23462
rect 20628 22568 20680 22574
rect 20628 22510 20680 22516
rect 20640 21894 20668 22510
rect 20720 22432 20772 22438
rect 20720 22374 20772 22380
rect 20628 21888 20680 21894
rect 20628 21830 20680 21836
rect 20536 21684 20588 21690
rect 20536 21626 20588 21632
rect 20456 21508 20668 21536
rect 20444 21344 20496 21350
rect 20444 21286 20496 21292
rect 20456 19514 20484 21286
rect 20444 19508 20496 19514
rect 20444 19450 20496 19456
rect 20444 18624 20496 18630
rect 20444 18566 20496 18572
rect 20456 18222 20484 18566
rect 20444 18216 20496 18222
rect 20444 18158 20496 18164
rect 20640 16674 20668 21508
rect 20732 19514 20760 22374
rect 20824 22098 20852 23666
rect 21008 23662 21036 24670
rect 21088 24064 21140 24070
rect 21088 24006 21140 24012
rect 21100 23662 21128 24006
rect 20996 23656 21048 23662
rect 20996 23598 21048 23604
rect 21088 23656 21140 23662
rect 21088 23598 21140 23604
rect 20996 23520 21048 23526
rect 20996 23462 21048 23468
rect 21086 23488 21142 23497
rect 20904 22500 20956 22506
rect 20904 22442 20956 22448
rect 20812 22092 20864 22098
rect 20812 22034 20864 22040
rect 20916 21486 20944 22442
rect 20904 21480 20956 21486
rect 20904 21422 20956 21428
rect 20916 20890 20944 21422
rect 20824 20862 20944 20890
rect 20720 19508 20772 19514
rect 20720 19450 20772 19456
rect 20824 19394 20852 20862
rect 20904 20800 20956 20806
rect 20904 20742 20956 20748
rect 20732 19366 20852 19394
rect 20732 18766 20760 19366
rect 20720 18760 20772 18766
rect 20720 18702 20772 18708
rect 20812 18692 20864 18698
rect 20812 18634 20864 18640
rect 20824 17270 20852 18634
rect 20812 17264 20864 17270
rect 20812 17206 20864 17212
rect 20548 16646 20668 16674
rect 20444 16040 20496 16046
rect 20444 15982 20496 15988
rect 20456 15570 20484 15982
rect 20548 15910 20576 16646
rect 20720 16584 20772 16590
rect 20720 16526 20772 16532
rect 20628 16516 20680 16522
rect 20628 16458 20680 16464
rect 20640 16046 20668 16458
rect 20628 16040 20680 16046
rect 20628 15982 20680 15988
rect 20536 15904 20588 15910
rect 20536 15846 20588 15852
rect 20444 15564 20496 15570
rect 20444 15506 20496 15512
rect 20352 15156 20404 15162
rect 20352 15098 20404 15104
rect 20076 14544 20128 14550
rect 20076 14486 20128 14492
rect 20352 14272 20404 14278
rect 20352 14214 20404 14220
rect 20260 13864 20312 13870
rect 20260 13806 20312 13812
rect 20076 13184 20128 13190
rect 20076 13126 20128 13132
rect 20168 13184 20220 13190
rect 20168 13126 20220 13132
rect 20088 12918 20116 13126
rect 20076 12912 20128 12918
rect 20076 12854 20128 12860
rect 20076 12640 20128 12646
rect 20074 12608 20076 12617
rect 20128 12608 20130 12617
rect 20074 12543 20130 12552
rect 20180 11218 20208 13126
rect 20272 12306 20300 13806
rect 20364 12850 20392 14214
rect 20442 14104 20498 14113
rect 20442 14039 20498 14048
rect 20352 12844 20404 12850
rect 20352 12786 20404 12792
rect 20350 12744 20406 12753
rect 20350 12679 20406 12688
rect 20364 12442 20392 12679
rect 20352 12436 20404 12442
rect 20352 12378 20404 12384
rect 20260 12300 20312 12306
rect 20260 12242 20312 12248
rect 19984 11212 20036 11218
rect 19984 11154 20036 11160
rect 20168 11212 20220 11218
rect 20168 11154 20220 11160
rect 19996 10198 20024 11154
rect 20076 10600 20128 10606
rect 20076 10542 20128 10548
rect 20088 10266 20116 10542
rect 20168 10464 20220 10470
rect 20168 10406 20220 10412
rect 20180 10266 20208 10406
rect 20076 10260 20128 10266
rect 20076 10202 20128 10208
rect 20168 10260 20220 10266
rect 20168 10202 20220 10208
rect 19812 10118 19932 10146
rect 19984 10192 20036 10198
rect 19984 10134 20036 10140
rect 19812 9024 19840 10118
rect 20168 9512 20220 9518
rect 20166 9480 20168 9489
rect 20220 9480 20222 9489
rect 20272 9450 20300 12242
rect 20352 12164 20404 12170
rect 20352 12106 20404 12112
rect 20166 9415 20222 9424
rect 20260 9444 20312 9450
rect 19892 9376 19944 9382
rect 19892 9318 19944 9324
rect 19904 9178 19932 9318
rect 19892 9172 19944 9178
rect 19892 9114 19944 9120
rect 19812 8996 19932 9024
rect 19720 8894 19840 8922
rect 19616 8832 19668 8838
rect 19616 8774 19668 8780
rect 19628 8401 19656 8774
rect 19708 8492 19760 8498
rect 19708 8434 19760 8440
rect 19614 8392 19670 8401
rect 19614 8327 19670 8336
rect 19720 6866 19748 8434
rect 19708 6860 19760 6866
rect 19708 6802 19760 6808
rect 19616 6180 19668 6186
rect 19616 6122 19668 6128
rect 19522 4992 19578 5001
rect 19522 4927 19578 4936
rect 19524 3732 19576 3738
rect 19524 3674 19576 3680
rect 19300 3012 19472 3040
rect 19248 2994 19300 3000
rect 19536 800 19564 3674
rect 19628 2446 19656 6122
rect 19720 5234 19748 6802
rect 19812 5574 19840 8894
rect 19904 8634 19932 8996
rect 20180 8634 20208 9415
rect 20260 9386 20312 9392
rect 19892 8628 19944 8634
rect 19892 8570 19944 8576
rect 20168 8628 20220 8634
rect 20168 8570 20220 8576
rect 19800 5568 19852 5574
rect 19800 5510 19852 5516
rect 19708 5228 19760 5234
rect 19708 5170 19760 5176
rect 19904 3194 19932 8570
rect 20272 8566 20300 9386
rect 20260 8560 20312 8566
rect 20260 8502 20312 8508
rect 20168 8084 20220 8090
rect 20168 8026 20220 8032
rect 19984 6724 20036 6730
rect 19984 6666 20036 6672
rect 19996 6118 20024 6666
rect 19984 6112 20036 6118
rect 19984 6054 20036 6060
rect 19996 5778 20024 6054
rect 19984 5772 20036 5778
rect 19984 5714 20036 5720
rect 19996 5556 20024 5714
rect 20076 5568 20128 5574
rect 19996 5528 20076 5556
rect 20076 5510 20128 5516
rect 20088 5302 20116 5510
rect 20076 5296 20128 5302
rect 20076 5238 20128 5244
rect 19984 4004 20036 4010
rect 19984 3946 20036 3952
rect 19892 3188 19944 3194
rect 19892 3130 19944 3136
rect 19892 2848 19944 2854
rect 19892 2790 19944 2796
rect 19904 2514 19932 2790
rect 19892 2508 19944 2514
rect 19892 2450 19944 2456
rect 19616 2440 19668 2446
rect 19616 2382 19668 2388
rect 19996 2088 20024 3946
rect 20180 3126 20208 8026
rect 20364 6186 20392 12106
rect 20456 11762 20484 14039
rect 20548 13734 20576 15846
rect 20732 14414 20760 16526
rect 20812 15088 20864 15094
rect 20812 15030 20864 15036
rect 20720 14408 20772 14414
rect 20720 14350 20772 14356
rect 20536 13728 20588 13734
rect 20536 13670 20588 13676
rect 20628 13728 20680 13734
rect 20628 13670 20680 13676
rect 20536 13524 20588 13530
rect 20536 13466 20588 13472
rect 20548 13190 20576 13466
rect 20536 13184 20588 13190
rect 20536 13126 20588 13132
rect 20548 12918 20576 13126
rect 20536 12912 20588 12918
rect 20536 12854 20588 12860
rect 20640 12434 20668 13670
rect 20720 13252 20772 13258
rect 20720 13194 20772 13200
rect 20548 12406 20668 12434
rect 20444 11756 20496 11762
rect 20444 11698 20496 11704
rect 20456 11014 20484 11698
rect 20444 11008 20496 11014
rect 20444 10950 20496 10956
rect 20548 10792 20576 12406
rect 20628 12164 20680 12170
rect 20628 12106 20680 12112
rect 20640 11898 20668 12106
rect 20628 11892 20680 11898
rect 20628 11834 20680 11840
rect 20732 11830 20760 13194
rect 20720 11824 20772 11830
rect 20720 11766 20772 11772
rect 20824 11694 20852 15030
rect 20916 13326 20944 20742
rect 21008 18358 21036 23462
rect 21086 23423 21142 23432
rect 21100 22778 21128 23423
rect 21088 22772 21140 22778
rect 21088 22714 21140 22720
rect 21100 21418 21128 22714
rect 21180 22228 21232 22234
rect 21180 22170 21232 22176
rect 21088 21412 21140 21418
rect 21088 21354 21140 21360
rect 21192 21026 21220 22170
rect 21284 22030 21312 24822
rect 21376 23526 21404 25350
rect 21560 25294 21588 26386
rect 21652 26246 21680 26726
rect 21640 26240 21692 26246
rect 21640 26182 21692 26188
rect 21652 25702 21680 26182
rect 21640 25696 21692 25702
rect 21640 25638 21692 25644
rect 21456 25288 21508 25294
rect 21456 25230 21508 25236
rect 21548 25288 21600 25294
rect 21548 25230 21600 25236
rect 21468 24410 21496 25230
rect 21560 24750 21588 25230
rect 21652 24818 21680 25638
rect 21640 24812 21692 24818
rect 21640 24754 21692 24760
rect 21548 24744 21600 24750
rect 21548 24686 21600 24692
rect 21652 24682 21680 24754
rect 21640 24676 21692 24682
rect 21640 24618 21692 24624
rect 21456 24404 21508 24410
rect 21456 24346 21508 24352
rect 21652 24138 21680 24618
rect 21836 24614 21864 26823
rect 21916 26308 21968 26314
rect 21916 26250 21968 26256
rect 21928 25770 21956 26250
rect 22204 26246 22232 27390
rect 22284 27328 22336 27334
rect 22284 27270 22336 27276
rect 22192 26240 22244 26246
rect 22192 26182 22244 26188
rect 22192 25900 22244 25906
rect 22192 25842 22244 25848
rect 22204 25809 22232 25842
rect 22190 25800 22246 25809
rect 21916 25764 21968 25770
rect 22190 25735 22246 25744
rect 21916 25706 21968 25712
rect 22008 25696 22060 25702
rect 22008 25638 22060 25644
rect 21824 24608 21876 24614
rect 21824 24550 21876 24556
rect 21640 24132 21692 24138
rect 21640 24074 21692 24080
rect 21652 23526 21680 24074
rect 21364 23520 21416 23526
rect 21364 23462 21416 23468
rect 21640 23520 21692 23526
rect 21640 23462 21692 23468
rect 21364 23044 21416 23050
rect 21364 22986 21416 22992
rect 21272 22024 21324 22030
rect 21272 21966 21324 21972
rect 21100 20998 21220 21026
rect 21100 20942 21128 20998
rect 21088 20936 21140 20942
rect 21088 20878 21140 20884
rect 21088 20800 21140 20806
rect 21088 20742 21140 20748
rect 21100 19242 21128 20742
rect 21192 20466 21220 20998
rect 21376 20806 21404 22986
rect 22020 22982 22048 25638
rect 22192 25152 22244 25158
rect 22192 25094 22244 25100
rect 22100 24608 22152 24614
rect 22100 24550 22152 24556
rect 22008 22976 22060 22982
rect 22008 22918 22060 22924
rect 21824 21956 21876 21962
rect 21824 21898 21876 21904
rect 21732 21344 21784 21350
rect 21732 21286 21784 21292
rect 21364 20800 21416 20806
rect 21364 20742 21416 20748
rect 21180 20460 21232 20466
rect 21180 20402 21232 20408
rect 21456 19508 21508 19514
rect 21456 19450 21508 19456
rect 21088 19236 21140 19242
rect 21088 19178 21140 19184
rect 21272 19168 21324 19174
rect 21272 19110 21324 19116
rect 21180 18760 21232 18766
rect 21180 18702 21232 18708
rect 20996 18352 21048 18358
rect 20996 18294 21048 18300
rect 20996 18216 21048 18222
rect 20996 18158 21048 18164
rect 21008 18086 21036 18158
rect 20996 18080 21048 18086
rect 20996 18022 21048 18028
rect 21008 17610 21036 18022
rect 21192 17882 21220 18702
rect 21180 17876 21232 17882
rect 21180 17818 21232 17824
rect 20996 17604 21048 17610
rect 20996 17546 21048 17552
rect 21178 17368 21234 17377
rect 21178 17303 21180 17312
rect 21232 17303 21234 17312
rect 21180 17274 21232 17280
rect 20996 16584 21048 16590
rect 20996 16526 21048 16532
rect 21008 15366 21036 16526
rect 21284 15858 21312 19110
rect 21364 18080 21416 18086
rect 21362 18048 21364 18057
rect 21416 18048 21418 18057
rect 21362 17983 21418 17992
rect 21364 17604 21416 17610
rect 21364 17546 21416 17552
rect 21376 16182 21404 17546
rect 21364 16176 21416 16182
rect 21364 16118 21416 16124
rect 21192 15830 21312 15858
rect 20996 15360 21048 15366
rect 20996 15302 21048 15308
rect 21008 14958 21036 15302
rect 21088 15020 21140 15026
rect 21088 14962 21140 14968
rect 20996 14952 21048 14958
rect 20996 14894 21048 14900
rect 20904 13320 20956 13326
rect 20904 13262 20956 13268
rect 20996 13184 21048 13190
rect 20996 13126 21048 13132
rect 20902 13016 20958 13025
rect 21008 12986 21036 13126
rect 20902 12951 20904 12960
rect 20956 12951 20958 12960
rect 20996 12980 21048 12986
rect 20904 12922 20956 12928
rect 20996 12922 21048 12928
rect 21100 12714 21128 14962
rect 21088 12708 21140 12714
rect 21088 12650 21140 12656
rect 20812 11688 20864 11694
rect 20812 11630 20864 11636
rect 20720 11552 20772 11558
rect 20720 11494 20772 11500
rect 20628 10804 20680 10810
rect 20548 10764 20628 10792
rect 20548 8090 20576 10764
rect 20628 10746 20680 10752
rect 20628 9920 20680 9926
rect 20626 9888 20628 9897
rect 20680 9888 20682 9897
rect 20626 9823 20682 9832
rect 20732 9738 20760 11494
rect 20812 11280 20864 11286
rect 20812 11222 20864 11228
rect 20824 11121 20852 11222
rect 20996 11144 21048 11150
rect 20810 11112 20866 11121
rect 20996 11086 21048 11092
rect 20810 11047 20866 11056
rect 20904 11008 20956 11014
rect 20904 10950 20956 10956
rect 20916 10810 20944 10950
rect 20904 10804 20956 10810
rect 20904 10746 20956 10752
rect 20812 10192 20864 10198
rect 20812 10134 20864 10140
rect 20640 9710 20760 9738
rect 20536 8084 20588 8090
rect 20536 8026 20588 8032
rect 20352 6180 20404 6186
rect 20352 6122 20404 6128
rect 20260 5772 20312 5778
rect 20640 5760 20668 9710
rect 20824 9466 20852 10134
rect 20916 9994 20944 10746
rect 20904 9988 20956 9994
rect 20904 9930 20956 9936
rect 20732 9438 20852 9466
rect 20732 8537 20760 9438
rect 20812 9376 20864 9382
rect 20812 9318 20864 9324
rect 20718 8528 20774 8537
rect 20718 8463 20774 8472
rect 20260 5714 20312 5720
rect 20548 5732 20668 5760
rect 20168 3120 20220 3126
rect 20168 3062 20220 3068
rect 19904 2060 20024 2088
rect 19904 800 19932 2060
rect 20272 800 20300 5714
rect 20352 5704 20404 5710
rect 20352 5646 20404 5652
rect 20364 3641 20392 5646
rect 20444 5636 20496 5642
rect 20444 5578 20496 5584
rect 20456 5166 20484 5578
rect 20444 5160 20496 5166
rect 20444 5102 20496 5108
rect 20548 4622 20576 5732
rect 20720 5024 20772 5030
rect 20720 4966 20772 4972
rect 20536 4616 20588 4622
rect 20536 4558 20588 4564
rect 20350 3632 20406 3641
rect 20350 3567 20406 3576
rect 20732 2774 20760 4966
rect 20824 3534 20852 9318
rect 20904 5636 20956 5642
rect 20904 5578 20956 5584
rect 20812 3528 20864 3534
rect 20812 3470 20864 3476
rect 20640 2746 20760 2774
rect 20640 800 20668 2746
rect 20916 2650 20944 5578
rect 21008 3534 21036 11086
rect 21192 10985 21220 15830
rect 21468 15484 21496 19450
rect 21640 18352 21692 18358
rect 21640 18294 21692 18300
rect 21652 17882 21680 18294
rect 21640 17876 21692 17882
rect 21640 17818 21692 17824
rect 21548 16448 21600 16454
rect 21548 16390 21600 16396
rect 21560 16250 21588 16390
rect 21548 16244 21600 16250
rect 21548 16186 21600 16192
rect 21640 16244 21692 16250
rect 21640 16186 21692 16192
rect 21652 15706 21680 16186
rect 21640 15700 21692 15706
rect 21640 15642 21692 15648
rect 21284 15456 21496 15484
rect 21284 13818 21312 15456
rect 21640 15360 21692 15366
rect 21640 15302 21692 15308
rect 21456 15088 21508 15094
rect 21456 15030 21508 15036
rect 21364 14272 21416 14278
rect 21364 14214 21416 14220
rect 21376 13938 21404 14214
rect 21364 13932 21416 13938
rect 21364 13874 21416 13880
rect 21284 13790 21404 13818
rect 21272 13728 21324 13734
rect 21272 13670 21324 13676
rect 21178 10976 21234 10985
rect 21178 10911 21234 10920
rect 21088 10056 21140 10062
rect 21088 9998 21140 10004
rect 21180 10056 21232 10062
rect 21180 9998 21232 10004
rect 21100 8090 21128 9998
rect 21088 8084 21140 8090
rect 21088 8026 21140 8032
rect 21192 7392 21220 9998
rect 21284 9654 21312 13670
rect 21376 11150 21404 13790
rect 21468 12918 21496 15030
rect 21456 12912 21508 12918
rect 21456 12854 21508 12860
rect 21548 12844 21600 12850
rect 21548 12786 21600 12792
rect 21456 11756 21508 11762
rect 21456 11698 21508 11704
rect 21364 11144 21416 11150
rect 21364 11086 21416 11092
rect 21364 11008 21416 11014
rect 21364 10950 21416 10956
rect 21272 9648 21324 9654
rect 21272 9590 21324 9596
rect 21100 7364 21220 7392
rect 21100 4758 21128 7364
rect 21376 7290 21404 10950
rect 21468 10810 21496 11698
rect 21560 11354 21588 12786
rect 21548 11348 21600 11354
rect 21548 11290 21600 11296
rect 21456 10804 21508 10810
rect 21456 10746 21508 10752
rect 21468 10130 21496 10746
rect 21456 10124 21508 10130
rect 21456 10066 21508 10072
rect 21456 9988 21508 9994
rect 21456 9930 21508 9936
rect 21468 9722 21496 9930
rect 21456 9716 21508 9722
rect 21456 9658 21508 9664
rect 21456 9036 21508 9042
rect 21456 8978 21508 8984
rect 21468 8294 21496 8978
rect 21456 8288 21508 8294
rect 21456 8230 21508 8236
rect 21548 8084 21600 8090
rect 21548 8026 21600 8032
rect 21192 7262 21404 7290
rect 21088 4752 21140 4758
rect 21088 4694 21140 4700
rect 21192 4282 21220 7262
rect 21272 7200 21324 7206
rect 21272 7142 21324 7148
rect 21180 4276 21232 4282
rect 21180 4218 21232 4224
rect 21088 4208 21140 4214
rect 21088 4150 21140 4156
rect 20996 3528 21048 3534
rect 20996 3470 21048 3476
rect 20904 2644 20956 2650
rect 20904 2586 20956 2592
rect 21100 2088 21128 4150
rect 21284 3194 21312 7142
rect 21560 6934 21588 8026
rect 21548 6928 21600 6934
rect 21548 6870 21600 6876
rect 21548 5568 21600 5574
rect 21362 5536 21418 5545
rect 21548 5510 21600 5516
rect 21362 5471 21418 5480
rect 21376 4622 21404 5471
rect 21456 5024 21508 5030
rect 21456 4966 21508 4972
rect 21468 4622 21496 4966
rect 21364 4616 21416 4622
rect 21364 4558 21416 4564
rect 21456 4616 21508 4622
rect 21456 4558 21508 4564
rect 21364 4276 21416 4282
rect 21364 4218 21416 4224
rect 21272 3188 21324 3194
rect 21272 3130 21324 3136
rect 21376 3058 21404 4218
rect 21468 4078 21496 4558
rect 21560 4146 21588 5510
rect 21548 4140 21600 4146
rect 21548 4082 21600 4088
rect 21456 4072 21508 4078
rect 21456 4014 21508 4020
rect 21560 3942 21588 4082
rect 21548 3936 21600 3942
rect 21548 3878 21600 3884
rect 21364 3052 21416 3058
rect 21364 2994 21416 3000
rect 21364 2848 21416 2854
rect 21364 2790 21416 2796
rect 21272 2644 21324 2650
rect 21272 2586 21324 2592
rect 21008 2060 21128 2088
rect 21008 800 21036 2060
rect 21284 1902 21312 2586
rect 21272 1896 21324 1902
rect 21272 1838 21324 1844
rect 21376 800 21404 2790
rect 21652 2582 21680 15302
rect 21744 14414 21772 21286
rect 21836 20602 21864 21898
rect 22008 21548 22060 21554
rect 22008 21490 22060 21496
rect 22020 21146 22048 21490
rect 22008 21140 22060 21146
rect 22008 21082 22060 21088
rect 22008 20868 22060 20874
rect 22008 20810 22060 20816
rect 21824 20596 21876 20602
rect 21824 20538 21876 20544
rect 22020 20534 22048 20810
rect 22008 20528 22060 20534
rect 22008 20470 22060 20476
rect 22008 19712 22060 19718
rect 22008 19654 22060 19660
rect 22020 19310 22048 19654
rect 22008 19304 22060 19310
rect 22008 19246 22060 19252
rect 21916 18692 21968 18698
rect 21916 18634 21968 18640
rect 21928 18154 21956 18634
rect 22020 18290 22048 19246
rect 22008 18284 22060 18290
rect 22008 18226 22060 18232
rect 21916 18148 21968 18154
rect 21916 18090 21968 18096
rect 21824 17876 21876 17882
rect 21824 17818 21876 17824
rect 21836 14929 21864 17818
rect 21928 17678 21956 18090
rect 21916 17672 21968 17678
rect 22112 17626 22140 24550
rect 22204 24138 22232 25094
rect 22192 24132 22244 24138
rect 22192 24074 22244 24080
rect 22296 23798 22324 27270
rect 22376 26308 22428 26314
rect 22376 26250 22428 26256
rect 22284 23792 22336 23798
rect 22284 23734 22336 23740
rect 22192 23656 22244 23662
rect 22192 23598 22244 23604
rect 22284 23656 22336 23662
rect 22284 23598 22336 23604
rect 22204 21078 22232 23598
rect 22296 23118 22324 23598
rect 22284 23112 22336 23118
rect 22284 23054 22336 23060
rect 22388 22642 22416 26250
rect 22480 26081 22508 29582
rect 22560 29504 22612 29510
rect 22560 29446 22612 29452
rect 22572 29073 22600 29446
rect 23112 29300 23164 29306
rect 23112 29242 23164 29248
rect 23124 29209 23152 29242
rect 23110 29200 23166 29209
rect 22652 29164 22704 29170
rect 23110 29135 23166 29144
rect 22652 29106 22704 29112
rect 22558 29064 22614 29073
rect 22558 28999 22614 29008
rect 22560 28960 22612 28966
rect 22560 28902 22612 28908
rect 22572 28422 22600 28902
rect 22560 28416 22612 28422
rect 22560 28358 22612 28364
rect 22572 26466 22600 28358
rect 22664 27538 22692 29106
rect 22950 28860 23258 28869
rect 22950 28858 22956 28860
rect 23012 28858 23036 28860
rect 23092 28858 23116 28860
rect 23172 28858 23196 28860
rect 23252 28858 23258 28860
rect 23012 28806 23014 28858
rect 23194 28806 23196 28858
rect 22950 28804 22956 28806
rect 23012 28804 23036 28806
rect 23092 28804 23116 28806
rect 23172 28804 23196 28806
rect 23252 28804 23258 28806
rect 22950 28795 23258 28804
rect 22836 28688 22888 28694
rect 22836 28630 22888 28636
rect 22652 27532 22704 27538
rect 22652 27474 22704 27480
rect 22744 27328 22796 27334
rect 22744 27270 22796 27276
rect 22652 26784 22704 26790
rect 22652 26726 22704 26732
rect 22664 26586 22692 26726
rect 22652 26580 22704 26586
rect 22652 26522 22704 26528
rect 22572 26438 22692 26466
rect 22560 26240 22612 26246
rect 22560 26182 22612 26188
rect 22466 26072 22522 26081
rect 22466 26007 22522 26016
rect 22468 25832 22520 25838
rect 22468 25774 22520 25780
rect 22480 23730 22508 25774
rect 22468 23724 22520 23730
rect 22468 23666 22520 23672
rect 22468 23520 22520 23526
rect 22468 23462 22520 23468
rect 22376 22636 22428 22642
rect 22376 22578 22428 22584
rect 22192 21072 22244 21078
rect 22192 21014 22244 21020
rect 22192 20052 22244 20058
rect 22192 19994 22244 20000
rect 22204 18970 22232 19994
rect 22284 19780 22336 19786
rect 22284 19722 22336 19728
rect 22376 19780 22428 19786
rect 22376 19722 22428 19728
rect 22192 18964 22244 18970
rect 22192 18906 22244 18912
rect 22192 18624 22244 18630
rect 22192 18566 22244 18572
rect 22204 18222 22232 18566
rect 22296 18222 22324 19722
rect 22388 18426 22416 19722
rect 22480 19378 22508 23462
rect 22572 21690 22600 26182
rect 22664 23662 22692 26438
rect 22652 23656 22704 23662
rect 22652 23598 22704 23604
rect 22652 23248 22704 23254
rect 22652 23190 22704 23196
rect 22560 21684 22612 21690
rect 22560 21626 22612 21632
rect 22560 21548 22612 21554
rect 22560 21490 22612 21496
rect 22572 19530 22600 21490
rect 22664 20942 22692 23190
rect 22756 21842 22784 27270
rect 22848 24154 22876 28630
rect 23202 28520 23258 28529
rect 23308 28490 23336 30126
rect 23676 29594 23704 34682
rect 23756 34400 23808 34406
rect 23756 34342 23808 34348
rect 23768 33454 23796 34342
rect 23756 33448 23808 33454
rect 23756 33390 23808 33396
rect 23940 32904 23992 32910
rect 23940 32846 23992 32852
rect 23756 32496 23808 32502
rect 23756 32438 23808 32444
rect 23768 31754 23796 32438
rect 23768 31726 23888 31754
rect 23860 31686 23888 31726
rect 23848 31680 23900 31686
rect 23848 31622 23900 31628
rect 23860 31362 23888 31622
rect 23768 31346 23888 31362
rect 23756 31340 23888 31346
rect 23808 31334 23888 31340
rect 23756 31282 23808 31288
rect 23768 30598 23796 31282
rect 23952 31226 23980 32846
rect 24032 32768 24084 32774
rect 24032 32710 24084 32716
rect 23860 31198 23980 31226
rect 23860 30734 23888 31198
rect 23940 31136 23992 31142
rect 23940 31078 23992 31084
rect 23952 30734 23980 31078
rect 23848 30728 23900 30734
rect 23848 30670 23900 30676
rect 23940 30728 23992 30734
rect 23940 30670 23992 30676
rect 23756 30592 23808 30598
rect 23756 30534 23808 30540
rect 23584 29566 23704 29594
rect 23202 28455 23258 28464
rect 23296 28484 23348 28490
rect 23216 28218 23244 28455
rect 23296 28426 23348 28432
rect 23204 28212 23256 28218
rect 23204 28154 23256 28160
rect 23308 27878 23336 28426
rect 23480 27940 23532 27946
rect 23480 27882 23532 27888
rect 23296 27872 23348 27878
rect 23296 27814 23348 27820
rect 23388 27872 23440 27878
rect 23388 27814 23440 27820
rect 22950 27772 23258 27781
rect 22950 27770 22956 27772
rect 23012 27770 23036 27772
rect 23092 27770 23116 27772
rect 23172 27770 23196 27772
rect 23252 27770 23258 27772
rect 23012 27718 23014 27770
rect 23194 27718 23196 27770
rect 22950 27716 22956 27718
rect 23012 27716 23036 27718
rect 23092 27716 23116 27718
rect 23172 27716 23196 27718
rect 23252 27716 23258 27718
rect 22950 27707 23258 27716
rect 23204 26920 23256 26926
rect 23308 26874 23336 27814
rect 23400 27538 23428 27814
rect 23388 27532 23440 27538
rect 23388 27474 23440 27480
rect 23256 26868 23336 26874
rect 23204 26862 23336 26868
rect 23216 26846 23336 26862
rect 22950 26684 23258 26693
rect 22950 26682 22956 26684
rect 23012 26682 23036 26684
rect 23092 26682 23116 26684
rect 23172 26682 23196 26684
rect 23252 26682 23258 26684
rect 23012 26630 23014 26682
rect 23194 26630 23196 26682
rect 22950 26628 22956 26630
rect 23012 26628 23036 26630
rect 23092 26628 23116 26630
rect 23172 26628 23196 26630
rect 23252 26628 23258 26630
rect 22950 26619 23258 26628
rect 23020 26240 23072 26246
rect 23020 26182 23072 26188
rect 23032 25838 23060 26182
rect 23308 25838 23336 26846
rect 23020 25832 23072 25838
rect 23020 25774 23072 25780
rect 23296 25832 23348 25838
rect 23296 25774 23348 25780
rect 22950 25596 23258 25605
rect 22950 25594 22956 25596
rect 23012 25594 23036 25596
rect 23092 25594 23116 25596
rect 23172 25594 23196 25596
rect 23252 25594 23258 25596
rect 23012 25542 23014 25594
rect 23194 25542 23196 25594
rect 22950 25540 22956 25542
rect 23012 25540 23036 25542
rect 23092 25540 23116 25542
rect 23172 25540 23196 25542
rect 23252 25540 23258 25542
rect 22950 25531 23258 25540
rect 23492 24818 23520 27882
rect 23584 27130 23612 29566
rect 23664 29504 23716 29510
rect 23664 29446 23716 29452
rect 23756 29504 23808 29510
rect 23756 29446 23808 29452
rect 23676 27470 23704 29446
rect 23664 27464 23716 27470
rect 23664 27406 23716 27412
rect 23572 27124 23624 27130
rect 23572 27066 23624 27072
rect 23572 26784 23624 26790
rect 23572 26726 23624 26732
rect 23664 26784 23716 26790
rect 23664 26726 23716 26732
rect 23584 26586 23612 26726
rect 23572 26580 23624 26586
rect 23572 26522 23624 26528
rect 23572 25832 23624 25838
rect 23572 25774 23624 25780
rect 23480 24812 23532 24818
rect 23480 24754 23532 24760
rect 23584 24750 23612 25774
rect 23296 24744 23348 24750
rect 23296 24686 23348 24692
rect 23572 24744 23624 24750
rect 23572 24686 23624 24692
rect 22950 24508 23258 24517
rect 22950 24506 22956 24508
rect 23012 24506 23036 24508
rect 23092 24506 23116 24508
rect 23172 24506 23196 24508
rect 23252 24506 23258 24508
rect 23012 24454 23014 24506
rect 23194 24454 23196 24506
rect 22950 24452 22956 24454
rect 23012 24452 23036 24454
rect 23092 24452 23116 24454
rect 23172 24452 23196 24454
rect 23252 24452 23258 24454
rect 22950 24443 23258 24452
rect 23308 24342 23336 24686
rect 23676 24614 23704 26726
rect 23768 26042 23796 29446
rect 23952 27538 23980 30670
rect 23940 27532 23992 27538
rect 23940 27474 23992 27480
rect 24044 27470 24072 32710
rect 24032 27464 24084 27470
rect 24032 27406 24084 27412
rect 24136 27402 24164 35158
rect 24674 35119 24730 35128
rect 24584 35080 24636 35086
rect 24584 35022 24636 35028
rect 24596 34950 24624 35022
rect 24676 35012 24728 35018
rect 24676 34954 24728 34960
rect 24584 34944 24636 34950
rect 24584 34886 24636 34892
rect 24492 34536 24544 34542
rect 24492 34478 24544 34484
rect 24400 33856 24452 33862
rect 24400 33798 24452 33804
rect 24412 33658 24440 33798
rect 24400 33652 24452 33658
rect 24400 33594 24452 33600
rect 24412 29238 24440 33594
rect 24504 31793 24532 34478
rect 24596 32609 24624 34886
rect 24688 34610 24716 34954
rect 24676 34604 24728 34610
rect 24676 34546 24728 34552
rect 24688 33425 24716 34546
rect 24780 34241 24808 35430
rect 24766 34232 24822 34241
rect 24766 34167 24822 34176
rect 24768 33448 24820 33454
rect 24674 33416 24730 33425
rect 24768 33390 24820 33396
rect 24674 33351 24730 33360
rect 24582 32600 24638 32609
rect 24582 32535 24638 32544
rect 24490 31784 24546 31793
rect 24490 31719 24546 31728
rect 24780 31346 24808 33390
rect 24872 32230 24900 53382
rect 25044 53100 25096 53106
rect 25044 53042 25096 53048
rect 25056 53009 25084 53042
rect 25042 53000 25098 53009
rect 25042 52935 25098 52944
rect 26056 52896 26108 52902
rect 26056 52838 26108 52844
rect 24952 52420 25004 52426
rect 24952 52362 25004 52368
rect 24964 52193 24992 52362
rect 24950 52184 25006 52193
rect 24950 52119 25006 52128
rect 25504 51808 25556 51814
rect 25504 51750 25556 51756
rect 25516 51406 25544 51750
rect 25504 51400 25556 51406
rect 25502 51368 25504 51377
rect 25556 51368 25558 51377
rect 25502 51303 25558 51312
rect 24952 50924 25004 50930
rect 24952 50866 25004 50872
rect 24964 50561 24992 50866
rect 25044 50720 25096 50726
rect 25044 50662 25096 50668
rect 24950 50552 25006 50561
rect 25056 50522 25084 50662
rect 24950 50487 25006 50496
rect 25044 50516 25096 50522
rect 25044 50458 25096 50464
rect 25504 50176 25556 50182
rect 25504 50118 25556 50124
rect 25516 49842 25544 50118
rect 25504 49836 25556 49842
rect 25504 49778 25556 49784
rect 25516 49745 25544 49778
rect 25502 49736 25558 49745
rect 25502 49671 25558 49680
rect 25136 49156 25188 49162
rect 25136 49098 25188 49104
rect 25148 48929 25176 49098
rect 25228 49088 25280 49094
rect 25228 49030 25280 49036
rect 25134 48920 25190 48929
rect 25134 48855 25190 48864
rect 25136 48544 25188 48550
rect 25136 48486 25188 48492
rect 25148 48142 25176 48486
rect 25136 48136 25188 48142
rect 25134 48104 25136 48113
rect 25188 48104 25190 48113
rect 25134 48039 25190 48048
rect 25240 47258 25268 49030
rect 25320 47660 25372 47666
rect 25320 47602 25372 47608
rect 25332 47297 25360 47602
rect 25964 47456 26016 47462
rect 25964 47398 26016 47404
rect 25318 47288 25374 47297
rect 25228 47252 25280 47258
rect 25318 47223 25374 47232
rect 25228 47194 25280 47200
rect 25320 46912 25372 46918
rect 25320 46854 25372 46860
rect 25332 46578 25360 46854
rect 25320 46572 25372 46578
rect 25320 46514 25372 46520
rect 25332 46481 25360 46514
rect 25318 46472 25374 46481
rect 25318 46407 25374 46416
rect 25320 45960 25372 45966
rect 25320 45902 25372 45908
rect 25332 45665 25360 45902
rect 25318 45656 25374 45665
rect 25318 45591 25374 45600
rect 25320 45280 25372 45286
rect 25320 45222 25372 45228
rect 25332 44878 25360 45222
rect 25320 44872 25372 44878
rect 25318 44840 25320 44849
rect 25372 44840 25374 44849
rect 25318 44775 25374 44784
rect 25780 44260 25832 44266
rect 25780 44202 25832 44208
rect 25504 43648 25556 43654
rect 25504 43590 25556 43596
rect 25516 43382 25544 43590
rect 25504 43376 25556 43382
rect 25504 43318 25556 43324
rect 25516 43217 25544 43318
rect 25502 43208 25558 43217
rect 25502 43143 25558 43152
rect 25596 43172 25648 43178
rect 25596 43114 25648 43120
rect 25136 42628 25188 42634
rect 25136 42570 25188 42576
rect 25148 42401 25176 42570
rect 25134 42392 25190 42401
rect 25134 42327 25190 42336
rect 25136 42016 25188 42022
rect 25136 41958 25188 41964
rect 25148 41614 25176 41958
rect 25136 41608 25188 41614
rect 25134 41576 25136 41585
rect 25188 41576 25190 41585
rect 25134 41511 25190 41520
rect 25320 41132 25372 41138
rect 25320 41074 25372 41080
rect 25228 40928 25280 40934
rect 25228 40870 25280 40876
rect 25044 40180 25096 40186
rect 25044 40122 25096 40128
rect 24952 35760 25004 35766
rect 24952 35702 25004 35708
rect 24964 35290 24992 35702
rect 24952 35284 25004 35290
rect 24952 35226 25004 35232
rect 24952 33312 25004 33318
rect 24952 33254 25004 33260
rect 24860 32224 24912 32230
rect 24860 32166 24912 32172
rect 24768 31340 24820 31346
rect 24768 31282 24820 31288
rect 24584 30592 24636 30598
rect 24584 30534 24636 30540
rect 24596 30394 24624 30534
rect 24492 30388 24544 30394
rect 24492 30330 24544 30336
rect 24584 30388 24636 30394
rect 24584 30330 24636 30336
rect 24504 30138 24532 30330
rect 24780 30190 24808 31282
rect 24768 30184 24820 30190
rect 24504 30110 24624 30138
rect 24768 30126 24820 30132
rect 24596 29510 24624 30110
rect 24860 29572 24912 29578
rect 24860 29514 24912 29520
rect 24584 29504 24636 29510
rect 24584 29446 24636 29452
rect 24400 29232 24452 29238
rect 24400 29174 24452 29180
rect 24308 28416 24360 28422
rect 24308 28358 24360 28364
rect 24320 28150 24348 28358
rect 24308 28144 24360 28150
rect 24308 28086 24360 28092
rect 24124 27396 24176 27402
rect 24124 27338 24176 27344
rect 24320 27130 24348 28086
rect 24596 28082 24624 29446
rect 24872 29345 24900 29514
rect 24858 29336 24914 29345
rect 24858 29271 24914 29280
rect 24860 29096 24912 29102
rect 24860 29038 24912 29044
rect 24872 28490 24900 29038
rect 24964 28626 24992 33254
rect 25056 32978 25084 40122
rect 25136 37868 25188 37874
rect 25136 37810 25188 37816
rect 25148 37505 25176 37810
rect 25134 37496 25190 37505
rect 25134 37431 25190 37440
rect 25136 36780 25188 36786
rect 25136 36722 25188 36728
rect 25148 36689 25176 36722
rect 25134 36680 25190 36689
rect 25134 36615 25190 36624
rect 25136 34400 25188 34406
rect 25136 34342 25188 34348
rect 25044 32972 25096 32978
rect 25044 32914 25096 32920
rect 25044 29504 25096 29510
rect 25044 29446 25096 29452
rect 24952 28620 25004 28626
rect 24952 28562 25004 28568
rect 24860 28484 24912 28490
rect 24860 28426 24912 28432
rect 24584 28076 24636 28082
rect 24584 28018 24636 28024
rect 24492 27464 24544 27470
rect 24492 27406 24544 27412
rect 24308 27124 24360 27130
rect 24308 27066 24360 27072
rect 23848 26308 23900 26314
rect 23848 26250 23900 26256
rect 23756 26036 23808 26042
rect 23756 25978 23808 25984
rect 23480 24608 23532 24614
rect 23480 24550 23532 24556
rect 23664 24608 23716 24614
rect 23664 24550 23716 24556
rect 23296 24336 23348 24342
rect 23296 24278 23348 24284
rect 22848 24126 22968 24154
rect 22836 24064 22888 24070
rect 22836 24006 22888 24012
rect 22848 22094 22876 24006
rect 22940 23526 22968 24126
rect 23204 23656 23256 23662
rect 23308 23610 23336 24278
rect 23492 24274 23520 24550
rect 23480 24268 23532 24274
rect 23480 24210 23532 24216
rect 23388 23792 23440 23798
rect 23388 23734 23440 23740
rect 23256 23604 23336 23610
rect 23204 23598 23336 23604
rect 23216 23582 23336 23598
rect 22928 23520 22980 23526
rect 22928 23462 22980 23468
rect 22950 23420 23258 23429
rect 22950 23418 22956 23420
rect 23012 23418 23036 23420
rect 23092 23418 23116 23420
rect 23172 23418 23196 23420
rect 23252 23418 23258 23420
rect 23012 23366 23014 23418
rect 23194 23366 23196 23418
rect 22950 23364 22956 23366
rect 23012 23364 23036 23366
rect 23092 23364 23116 23366
rect 23172 23364 23196 23366
rect 23252 23364 23258 23366
rect 22950 23355 23258 23364
rect 22950 22332 23258 22341
rect 22950 22330 22956 22332
rect 23012 22330 23036 22332
rect 23092 22330 23116 22332
rect 23172 22330 23196 22332
rect 23252 22330 23258 22332
rect 23012 22278 23014 22330
rect 23194 22278 23196 22330
rect 22950 22276 22956 22278
rect 23012 22276 23036 22278
rect 23092 22276 23116 22278
rect 23172 22276 23196 22278
rect 23252 22276 23258 22278
rect 22950 22267 23258 22276
rect 23308 22098 23336 23582
rect 23400 22234 23428 23734
rect 23860 23662 23888 26250
rect 24320 25974 24348 27066
rect 24504 26790 24532 27406
rect 24492 26784 24544 26790
rect 24492 26726 24544 26732
rect 24124 25968 24176 25974
rect 24124 25910 24176 25916
rect 24308 25968 24360 25974
rect 24308 25910 24360 25916
rect 23940 25696 23992 25702
rect 23940 25638 23992 25644
rect 23952 24342 23980 25638
rect 24136 24886 24164 25910
rect 24596 25838 24624 28018
rect 24768 28008 24820 28014
rect 24768 27950 24820 27956
rect 24676 26512 24728 26518
rect 24676 26454 24728 26460
rect 24584 25832 24636 25838
rect 24584 25774 24636 25780
rect 24124 24880 24176 24886
rect 24124 24822 24176 24828
rect 23940 24336 23992 24342
rect 23940 24278 23992 24284
rect 24136 24274 24164 24822
rect 24124 24268 24176 24274
rect 24124 24210 24176 24216
rect 24136 24070 24164 24210
rect 24124 24064 24176 24070
rect 24124 24006 24176 24012
rect 23848 23656 23900 23662
rect 23754 23624 23810 23633
rect 23848 23598 23900 23604
rect 23754 23559 23810 23568
rect 23768 23186 23796 23559
rect 24136 23526 24164 24006
rect 24124 23520 24176 23526
rect 24124 23462 24176 23468
rect 23756 23180 23808 23186
rect 23756 23122 23808 23128
rect 23848 23112 23900 23118
rect 23848 23054 23900 23060
rect 23572 22976 23624 22982
rect 23572 22918 23624 22924
rect 23388 22228 23440 22234
rect 23388 22170 23440 22176
rect 22848 22066 22968 22094
rect 22756 21814 22876 21842
rect 22744 21684 22796 21690
rect 22744 21626 22796 21632
rect 22652 20936 22704 20942
rect 22652 20878 22704 20884
rect 22652 20800 22704 20806
rect 22652 20742 22704 20748
rect 22664 19689 22692 20742
rect 22756 20466 22784 21626
rect 22744 20460 22796 20466
rect 22744 20402 22796 20408
rect 22650 19680 22706 19689
rect 22650 19615 22706 19624
rect 22572 19502 22692 19530
rect 22468 19372 22520 19378
rect 22468 19314 22520 19320
rect 22560 19372 22612 19378
rect 22560 19314 22612 19320
rect 22466 19272 22522 19281
rect 22466 19207 22522 19216
rect 22376 18420 22428 18426
rect 22376 18362 22428 18368
rect 22192 18216 22244 18222
rect 22192 18158 22244 18164
rect 22284 18216 22336 18222
rect 22284 18158 22336 18164
rect 21916 17614 21968 17620
rect 22020 17598 22140 17626
rect 22020 16946 22048 17598
rect 22100 17536 22152 17542
rect 22100 17478 22152 17484
rect 22112 17105 22140 17478
rect 22192 17196 22244 17202
rect 22192 17138 22244 17144
rect 22098 17096 22154 17105
rect 22098 17031 22154 17040
rect 22020 16918 22140 16946
rect 21916 16176 21968 16182
rect 21916 16118 21968 16124
rect 21928 15434 21956 16118
rect 21916 15428 21968 15434
rect 21916 15370 21968 15376
rect 21928 15162 21956 15370
rect 21916 15156 21968 15162
rect 21916 15098 21968 15104
rect 21822 14920 21878 14929
rect 21822 14855 21878 14864
rect 21732 14408 21784 14414
rect 21732 14350 21784 14356
rect 22112 14278 22140 16918
rect 22204 14634 22232 17138
rect 22296 16046 22324 18158
rect 22376 16992 22428 16998
rect 22376 16934 22428 16940
rect 22284 16040 22336 16046
rect 22284 15982 22336 15988
rect 22296 15570 22324 15982
rect 22284 15564 22336 15570
rect 22284 15506 22336 15512
rect 22204 14606 22324 14634
rect 22296 14550 22324 14606
rect 22284 14544 22336 14550
rect 22284 14486 22336 14492
rect 22192 14476 22244 14482
rect 22192 14418 22244 14424
rect 22100 14272 22152 14278
rect 22100 14214 22152 14220
rect 21916 13796 21968 13802
rect 21916 13738 21968 13744
rect 21732 13184 21784 13190
rect 21732 13126 21784 13132
rect 21744 12434 21772 13126
rect 21744 12406 21864 12434
rect 21732 12368 21784 12374
rect 21732 12310 21784 12316
rect 21744 11830 21772 12310
rect 21732 11824 21784 11830
rect 21732 11766 21784 11772
rect 21732 11144 21784 11150
rect 21732 11086 21784 11092
rect 21744 8022 21772 11086
rect 21836 10062 21864 12406
rect 21928 12374 21956 13738
rect 21916 12368 21968 12374
rect 21916 12310 21968 12316
rect 22204 12238 22232 14418
rect 22284 14408 22336 14414
rect 22284 14350 22336 14356
rect 22296 12850 22324 14350
rect 22388 12918 22416 16934
rect 22480 15366 22508 19207
rect 22572 18834 22600 19314
rect 22560 18828 22612 18834
rect 22560 18770 22612 18776
rect 22664 17762 22692 19502
rect 22756 19310 22784 20402
rect 22848 19938 22876 21814
rect 22940 21486 22968 22066
rect 23296 22092 23348 22098
rect 23296 22034 23348 22040
rect 23112 22024 23164 22030
rect 23112 21966 23164 21972
rect 23124 21622 23152 21966
rect 23204 21956 23256 21962
rect 23204 21898 23256 21904
rect 23216 21622 23244 21898
rect 23112 21616 23164 21622
rect 23112 21558 23164 21564
rect 23204 21616 23256 21622
rect 23204 21558 23256 21564
rect 23308 21554 23336 22034
rect 23296 21548 23348 21554
rect 23296 21490 23348 21496
rect 22928 21480 22980 21486
rect 22928 21422 22980 21428
rect 23388 21344 23440 21350
rect 23388 21286 23440 21292
rect 22950 21244 23258 21253
rect 22950 21242 22956 21244
rect 23012 21242 23036 21244
rect 23092 21242 23116 21244
rect 23172 21242 23196 21244
rect 23252 21242 23258 21244
rect 23012 21190 23014 21242
rect 23194 21190 23196 21242
rect 22950 21188 22956 21190
rect 23012 21188 23036 21190
rect 23092 21188 23116 21190
rect 23172 21188 23196 21190
rect 23252 21188 23258 21190
rect 22950 21179 23258 21188
rect 23400 21185 23428 21286
rect 23386 21176 23442 21185
rect 23386 21111 23442 21120
rect 23204 20392 23256 20398
rect 23202 20360 23204 20369
rect 23296 20392 23348 20398
rect 23256 20360 23258 20369
rect 23296 20334 23348 20340
rect 23202 20295 23258 20304
rect 22950 20156 23258 20165
rect 22950 20154 22956 20156
rect 23012 20154 23036 20156
rect 23092 20154 23116 20156
rect 23172 20154 23196 20156
rect 23252 20154 23258 20156
rect 23012 20102 23014 20154
rect 23194 20102 23196 20154
rect 22950 20100 22956 20102
rect 23012 20100 23036 20102
rect 23092 20100 23116 20102
rect 23172 20100 23196 20102
rect 23252 20100 23258 20102
rect 22950 20091 23258 20100
rect 22848 19910 22968 19938
rect 22744 19304 22796 19310
rect 22940 19258 22968 19910
rect 23308 19310 23336 20334
rect 23386 19544 23442 19553
rect 23386 19479 23442 19488
rect 22744 19246 22796 19252
rect 22848 19230 22968 19258
rect 23296 19304 23348 19310
rect 23296 19246 23348 19252
rect 22744 19168 22796 19174
rect 22744 19110 22796 19116
rect 22756 18698 22784 19110
rect 22744 18692 22796 18698
rect 22744 18634 22796 18640
rect 22572 17734 22692 17762
rect 22572 16590 22600 17734
rect 22652 17672 22704 17678
rect 22652 17614 22704 17620
rect 22560 16584 22612 16590
rect 22560 16526 22612 16532
rect 22468 15360 22520 15366
rect 22468 15302 22520 15308
rect 22480 15026 22508 15302
rect 22468 15020 22520 15026
rect 22468 14962 22520 14968
rect 22560 14816 22612 14822
rect 22560 14758 22612 14764
rect 22572 14482 22600 14758
rect 22664 14618 22692 17614
rect 22744 16584 22796 16590
rect 22744 16526 22796 16532
rect 22652 14612 22704 14618
rect 22652 14554 22704 14560
rect 22560 14476 22612 14482
rect 22560 14418 22612 14424
rect 22376 12912 22428 12918
rect 22376 12854 22428 12860
rect 22284 12844 22336 12850
rect 22284 12786 22336 12792
rect 22284 12640 22336 12646
rect 22284 12582 22336 12588
rect 22192 12232 22244 12238
rect 22192 12174 22244 12180
rect 22296 12170 22324 12582
rect 21916 12164 21968 12170
rect 21916 12106 21968 12112
rect 22284 12164 22336 12170
rect 22284 12106 22336 12112
rect 21928 10674 21956 12106
rect 22284 11756 22336 11762
rect 22284 11698 22336 11704
rect 21916 10668 21968 10674
rect 21916 10610 21968 10616
rect 21928 10198 21956 10610
rect 22008 10600 22060 10606
rect 22008 10542 22060 10548
rect 21916 10192 21968 10198
rect 22020 10169 22048 10542
rect 21916 10134 21968 10140
rect 22006 10160 22062 10169
rect 21824 10056 21876 10062
rect 21824 9998 21876 10004
rect 21928 9994 21956 10134
rect 22296 10130 22324 11698
rect 22756 10810 22784 16526
rect 22848 13870 22876 19230
rect 22950 19068 23258 19077
rect 22950 19066 22956 19068
rect 23012 19066 23036 19068
rect 23092 19066 23116 19068
rect 23172 19066 23196 19068
rect 23252 19066 23258 19068
rect 23012 19014 23014 19066
rect 23194 19014 23196 19066
rect 22950 19012 22956 19014
rect 23012 19012 23036 19014
rect 23092 19012 23116 19014
rect 23172 19012 23196 19014
rect 23252 19012 23258 19014
rect 22950 19003 23258 19012
rect 23308 18222 23336 19246
rect 23400 18834 23428 19479
rect 23388 18828 23440 18834
rect 23388 18770 23440 18776
rect 23584 18358 23612 22918
rect 23860 22234 23888 23054
rect 23848 22228 23900 22234
rect 23848 22170 23900 22176
rect 24136 21622 24164 23462
rect 24492 22976 24544 22982
rect 24492 22918 24544 22924
rect 24032 21616 24084 21622
rect 24124 21616 24176 21622
rect 24084 21576 24124 21604
rect 24032 21558 24084 21564
rect 24124 21558 24176 21564
rect 24136 21350 24164 21558
rect 24124 21344 24176 21350
rect 24124 21286 24176 21292
rect 23940 20936 23992 20942
rect 23940 20878 23992 20884
rect 23756 20868 23808 20874
rect 23756 20810 23808 20816
rect 23768 19174 23796 20810
rect 23952 19718 23980 20878
rect 24136 20534 24164 21286
rect 24124 20528 24176 20534
rect 24124 20470 24176 20476
rect 24136 19786 24164 20470
rect 24124 19780 24176 19786
rect 24124 19722 24176 19728
rect 23940 19712 23992 19718
rect 23940 19654 23992 19660
rect 23756 19168 23808 19174
rect 23756 19110 23808 19116
rect 23572 18352 23624 18358
rect 23572 18294 23624 18300
rect 23296 18216 23348 18222
rect 23296 18158 23348 18164
rect 23388 18080 23440 18086
rect 23388 18022 23440 18028
rect 22950 17980 23258 17989
rect 22950 17978 22956 17980
rect 23012 17978 23036 17980
rect 23092 17978 23116 17980
rect 23172 17978 23196 17980
rect 23252 17978 23258 17980
rect 23012 17926 23014 17978
rect 23194 17926 23196 17978
rect 22950 17924 22956 17926
rect 23012 17924 23036 17926
rect 23092 17924 23116 17926
rect 23172 17924 23196 17926
rect 23252 17924 23258 17926
rect 22950 17915 23258 17924
rect 23400 17134 23428 18022
rect 23388 17128 23440 17134
rect 23388 17070 23440 17076
rect 22950 16892 23258 16901
rect 22950 16890 22956 16892
rect 23012 16890 23036 16892
rect 23092 16890 23116 16892
rect 23172 16890 23196 16892
rect 23252 16890 23258 16892
rect 23012 16838 23014 16890
rect 23194 16838 23196 16890
rect 22950 16836 22956 16838
rect 23012 16836 23036 16838
rect 23092 16836 23116 16838
rect 23172 16836 23196 16838
rect 23252 16836 23258 16838
rect 22950 16827 23258 16836
rect 23952 16590 23980 19654
rect 24136 19446 24164 19722
rect 24504 19514 24532 22918
rect 24688 22098 24716 26454
rect 24780 26042 24808 27950
rect 25056 26450 25084 29446
rect 25148 28218 25176 34342
rect 25240 33658 25268 40870
rect 25332 40769 25360 41074
rect 25318 40760 25374 40769
rect 25318 40695 25374 40704
rect 25412 40384 25464 40390
rect 25412 40326 25464 40332
rect 25424 40118 25452 40326
rect 25412 40112 25464 40118
rect 25412 40054 25464 40060
rect 25424 39953 25452 40054
rect 25410 39944 25466 39953
rect 25410 39879 25466 39888
rect 25320 39432 25372 39438
rect 25320 39374 25372 39380
rect 25332 39137 25360 39374
rect 25318 39128 25374 39137
rect 25318 39063 25374 39072
rect 25320 38752 25372 38758
rect 25320 38694 25372 38700
rect 25332 38350 25360 38694
rect 25320 38344 25372 38350
rect 25318 38312 25320 38321
rect 25372 38312 25374 38321
rect 25318 38247 25374 38256
rect 25320 37256 25372 37262
rect 25320 37198 25372 37204
rect 25332 35873 25360 37198
rect 25504 36032 25556 36038
rect 25504 35974 25556 35980
rect 25318 35864 25374 35873
rect 25318 35799 25374 35808
rect 25320 35284 25372 35290
rect 25320 35226 25372 35232
rect 25228 33652 25280 33658
rect 25228 33594 25280 33600
rect 25332 32842 25360 35226
rect 25320 32836 25372 32842
rect 25320 32778 25372 32784
rect 25320 32360 25372 32366
rect 25320 32302 25372 32308
rect 25228 32224 25280 32230
rect 25228 32166 25280 32172
rect 25240 31822 25268 32166
rect 25228 31816 25280 31822
rect 25228 31758 25280 31764
rect 25240 28626 25268 31758
rect 25332 31482 25360 32302
rect 25320 31476 25372 31482
rect 25320 31418 25372 31424
rect 25318 30968 25374 30977
rect 25318 30903 25374 30912
rect 25332 29646 25360 30903
rect 25410 30152 25466 30161
rect 25410 30087 25466 30096
rect 25320 29640 25372 29646
rect 25320 29582 25372 29588
rect 25424 29170 25452 30087
rect 25412 29164 25464 29170
rect 25412 29106 25464 29112
rect 25320 29028 25372 29034
rect 25320 28970 25372 28976
rect 25228 28620 25280 28626
rect 25228 28562 25280 28568
rect 25136 28212 25188 28218
rect 25136 28154 25188 28160
rect 25228 27940 25280 27946
rect 25228 27882 25280 27888
rect 25136 27872 25188 27878
rect 25136 27814 25188 27820
rect 25148 27130 25176 27814
rect 25240 27606 25268 27882
rect 25228 27600 25280 27606
rect 25228 27542 25280 27548
rect 25136 27124 25188 27130
rect 25136 27066 25188 27072
rect 25228 26920 25280 26926
rect 25228 26862 25280 26868
rect 25044 26444 25096 26450
rect 25044 26386 25096 26392
rect 25136 26444 25188 26450
rect 25136 26386 25188 26392
rect 25044 26308 25096 26314
rect 25044 26250 25096 26256
rect 24768 26036 24820 26042
rect 24768 25978 24820 25984
rect 24780 25294 24808 25978
rect 24768 25288 24820 25294
rect 24768 25230 24820 25236
rect 24950 25256 25006 25265
rect 24950 25191 24952 25200
rect 25004 25191 25006 25200
rect 24952 25162 25004 25168
rect 24766 24440 24822 24449
rect 24766 24375 24822 24384
rect 24780 22574 24808 24375
rect 24952 24336 25004 24342
rect 24952 24278 25004 24284
rect 24858 22808 24914 22817
rect 24858 22743 24914 22752
rect 24872 22710 24900 22743
rect 24860 22704 24912 22710
rect 24860 22646 24912 22652
rect 24768 22568 24820 22574
rect 24768 22510 24820 22516
rect 24676 22092 24728 22098
rect 24676 22034 24728 22040
rect 24858 21992 24914 22001
rect 24858 21927 24914 21936
rect 24584 21888 24636 21894
rect 24584 21830 24636 21836
rect 24492 19508 24544 19514
rect 24492 19450 24544 19456
rect 24124 19440 24176 19446
rect 24124 19382 24176 19388
rect 24136 19174 24164 19382
rect 24124 19168 24176 19174
rect 24124 19110 24176 19116
rect 24136 18222 24164 19110
rect 24124 18216 24176 18222
rect 24124 18158 24176 18164
rect 24596 18136 24624 21830
rect 24872 21010 24900 21927
rect 24860 21004 24912 21010
rect 24860 20946 24912 20952
rect 24964 20806 24992 24278
rect 25056 23186 25084 26250
rect 25148 23662 25176 26386
rect 25240 25498 25268 26862
rect 25332 26382 25360 28970
rect 25424 28218 25452 29106
rect 25412 28212 25464 28218
rect 25412 28154 25464 28160
rect 25412 27124 25464 27130
rect 25412 27066 25464 27072
rect 25424 26586 25452 27066
rect 25412 26580 25464 26586
rect 25412 26522 25464 26528
rect 25320 26376 25372 26382
rect 25320 26318 25372 26324
rect 25424 26314 25452 26522
rect 25412 26308 25464 26314
rect 25412 26250 25464 26256
rect 25228 25492 25280 25498
rect 25228 25434 25280 25440
rect 25412 24948 25464 24954
rect 25412 24890 25464 24896
rect 25320 24744 25372 24750
rect 25320 24686 25372 24692
rect 25228 24064 25280 24070
rect 25228 24006 25280 24012
rect 25240 23866 25268 24006
rect 25228 23860 25280 23866
rect 25228 23802 25280 23808
rect 25136 23656 25188 23662
rect 25136 23598 25188 23604
rect 25044 23180 25096 23186
rect 25044 23122 25096 23128
rect 25044 23044 25096 23050
rect 25044 22986 25096 22992
rect 24860 20800 24912 20806
rect 24860 20742 24912 20748
rect 24952 20800 25004 20806
rect 24952 20742 25004 20748
rect 24766 18728 24822 18737
rect 24766 18663 24822 18672
rect 24596 18108 24716 18136
rect 24584 17536 24636 17542
rect 24584 17478 24636 17484
rect 24596 17066 24624 17478
rect 24584 17060 24636 17066
rect 24584 17002 24636 17008
rect 23940 16584 23992 16590
rect 23940 16526 23992 16532
rect 23572 15972 23624 15978
rect 23572 15914 23624 15920
rect 22950 15804 23258 15813
rect 22950 15802 22956 15804
rect 23012 15802 23036 15804
rect 23092 15802 23116 15804
rect 23172 15802 23196 15804
rect 23252 15802 23258 15804
rect 23012 15750 23014 15802
rect 23194 15750 23196 15802
rect 22950 15748 22956 15750
rect 23012 15748 23036 15750
rect 23092 15748 23116 15750
rect 23172 15748 23196 15750
rect 23252 15748 23258 15750
rect 22950 15739 23258 15748
rect 23584 15434 23612 15914
rect 23756 15904 23808 15910
rect 23756 15846 23808 15852
rect 23768 15450 23796 15846
rect 23848 15496 23900 15502
rect 23768 15444 23848 15450
rect 23768 15438 23900 15444
rect 23572 15428 23624 15434
rect 23572 15370 23624 15376
rect 23768 15422 23888 15438
rect 23584 15162 23612 15370
rect 23572 15156 23624 15162
rect 23572 15098 23624 15104
rect 23584 14822 23612 15098
rect 23768 14958 23796 15422
rect 23756 14952 23808 14958
rect 23756 14894 23808 14900
rect 23572 14816 23624 14822
rect 23572 14758 23624 14764
rect 23848 14816 23900 14822
rect 23848 14758 23900 14764
rect 22950 14716 23258 14725
rect 22950 14714 22956 14716
rect 23012 14714 23036 14716
rect 23092 14714 23116 14716
rect 23172 14714 23196 14716
rect 23252 14714 23258 14716
rect 23012 14662 23014 14714
rect 23194 14662 23196 14714
rect 22950 14660 22956 14662
rect 23012 14660 23036 14662
rect 23092 14660 23116 14662
rect 23172 14660 23196 14662
rect 23252 14660 23258 14662
rect 22950 14651 23258 14660
rect 23860 14346 23888 14758
rect 24688 14414 24716 18108
rect 24780 17134 24808 18663
rect 24872 18034 24900 20742
rect 25056 20346 25084 22986
rect 24964 20318 25084 20346
rect 24964 20058 24992 20318
rect 25044 20256 25096 20262
rect 25044 20198 25096 20204
rect 24952 20052 25004 20058
rect 24952 19994 25004 20000
rect 24872 18006 24992 18034
rect 24858 17912 24914 17921
rect 24858 17847 24914 17856
rect 24872 17746 24900 17847
rect 24964 17746 24992 18006
rect 24860 17740 24912 17746
rect 24860 17682 24912 17688
rect 24952 17740 25004 17746
rect 24952 17682 25004 17688
rect 24952 17536 25004 17542
rect 24952 17478 25004 17484
rect 24860 17264 24912 17270
rect 24860 17206 24912 17212
rect 24768 17128 24820 17134
rect 24872 17105 24900 17206
rect 24768 17070 24820 17076
rect 24858 17096 24914 17105
rect 24858 17031 24914 17040
rect 24964 16674 24992 17478
rect 24872 16646 24992 16674
rect 24872 16454 24900 16646
rect 24952 16516 25004 16522
rect 24952 16458 25004 16464
rect 24860 16448 24912 16454
rect 24860 16390 24912 16396
rect 24964 16289 24992 16458
rect 24950 16280 25006 16289
rect 25056 16250 25084 20198
rect 25148 19854 25176 23598
rect 25228 23180 25280 23186
rect 25228 23122 25280 23128
rect 25240 20602 25268 23122
rect 25228 20596 25280 20602
rect 25228 20538 25280 20544
rect 25136 19848 25188 19854
rect 25136 19790 25188 19796
rect 25240 19394 25268 20538
rect 25332 20058 25360 24686
rect 25424 22166 25452 24890
rect 25412 22160 25464 22166
rect 25412 22102 25464 22108
rect 25412 21480 25464 21486
rect 25412 21422 25464 21428
rect 25320 20052 25372 20058
rect 25320 19994 25372 20000
rect 25240 19366 25360 19394
rect 25228 19304 25280 19310
rect 25228 19246 25280 19252
rect 25136 19168 25188 19174
rect 25136 19110 25188 19116
rect 25148 17746 25176 19110
rect 25136 17740 25188 17746
rect 25136 17682 25188 17688
rect 24950 16215 25006 16224
rect 25044 16244 25096 16250
rect 25044 16186 25096 16192
rect 25148 16114 25176 17682
rect 25240 16590 25268 19246
rect 25332 18766 25360 19366
rect 25424 18970 25452 21422
rect 25516 20874 25544 35974
rect 25504 20868 25556 20874
rect 25504 20810 25556 20816
rect 25412 18964 25464 18970
rect 25412 18906 25464 18912
rect 25320 18760 25372 18766
rect 25320 18702 25372 18708
rect 25228 16584 25280 16590
rect 25228 16526 25280 16532
rect 25136 16108 25188 16114
rect 25136 16050 25188 16056
rect 24766 15464 24822 15473
rect 24766 15399 24822 15408
rect 24780 14958 24808 15399
rect 24768 14952 24820 14958
rect 24768 14894 24820 14900
rect 25608 14890 25636 43114
rect 25688 37120 25740 37126
rect 25688 37062 25740 37068
rect 25700 18426 25728 37062
rect 25688 18420 25740 18426
rect 25688 18362 25740 18368
rect 25792 16794 25820 44202
rect 25872 41540 25924 41546
rect 25872 41482 25924 41488
rect 25884 22094 25912 41482
rect 25976 29306 26004 47398
rect 26068 32978 26096 52838
rect 26516 52488 26568 52494
rect 26516 52430 26568 52436
rect 26148 42628 26200 42634
rect 26148 42570 26200 42576
rect 26056 32972 26108 32978
rect 26056 32914 26108 32920
rect 26056 32836 26108 32842
rect 26056 32778 26108 32784
rect 25964 29300 26016 29306
rect 25964 29242 26016 29248
rect 26068 27130 26096 32778
rect 26056 27124 26108 27130
rect 26056 27066 26108 27072
rect 26068 23118 26096 27066
rect 26056 23112 26108 23118
rect 26056 23054 26108 23060
rect 25884 22066 26004 22094
rect 25872 20800 25924 20806
rect 25872 20742 25924 20748
rect 25780 16788 25832 16794
rect 25780 16730 25832 16736
rect 25884 16182 25912 20742
rect 25872 16176 25924 16182
rect 25872 16118 25924 16124
rect 25596 14884 25648 14890
rect 25596 14826 25648 14832
rect 25134 14648 25190 14657
rect 25134 14583 25190 14592
rect 24676 14408 24728 14414
rect 24676 14350 24728 14356
rect 23848 14340 23900 14346
rect 23848 14282 23900 14288
rect 24032 14272 24084 14278
rect 24032 14214 24084 14220
rect 24492 14272 24544 14278
rect 24492 14214 24544 14220
rect 25044 14272 25096 14278
rect 25044 14214 25096 14220
rect 22836 13864 22888 13870
rect 22836 13806 22888 13812
rect 22950 13628 23258 13637
rect 22950 13626 22956 13628
rect 23012 13626 23036 13628
rect 23092 13626 23116 13628
rect 23172 13626 23196 13628
rect 23252 13626 23258 13628
rect 23012 13574 23014 13626
rect 23194 13574 23196 13626
rect 22950 13572 22956 13574
rect 23012 13572 23036 13574
rect 23092 13572 23116 13574
rect 23172 13572 23196 13574
rect 23252 13572 23258 13574
rect 22950 13563 23258 13572
rect 24044 13394 24072 14214
rect 24032 13388 24084 13394
rect 24032 13330 24084 13336
rect 23756 13320 23808 13326
rect 23756 13262 23808 13268
rect 23296 13184 23348 13190
rect 23296 13126 23348 13132
rect 23308 12918 23336 13126
rect 23296 12912 23348 12918
rect 23296 12854 23348 12860
rect 22836 12844 22888 12850
rect 22836 12786 22888 12792
rect 22848 11762 22876 12786
rect 22950 12540 23258 12549
rect 22950 12538 22956 12540
rect 23012 12538 23036 12540
rect 23092 12538 23116 12540
rect 23172 12538 23196 12540
rect 23252 12538 23258 12540
rect 23012 12486 23014 12538
rect 23194 12486 23196 12538
rect 22950 12484 22956 12486
rect 23012 12484 23036 12486
rect 23092 12484 23116 12486
rect 23172 12484 23196 12486
rect 23252 12484 23258 12486
rect 22950 12475 23258 12484
rect 23768 12434 23796 13262
rect 24504 12730 24532 14214
rect 24860 14000 24912 14006
rect 24860 13942 24912 13948
rect 24872 13841 24900 13942
rect 24858 13832 24914 13841
rect 24858 13767 24914 13776
rect 24768 13456 24820 13462
rect 24768 13398 24820 13404
rect 24780 12986 24808 13398
rect 24952 13252 25004 13258
rect 24952 13194 25004 13200
rect 24964 13025 24992 13194
rect 24950 13016 25006 13025
rect 24768 12980 24820 12986
rect 24950 12951 25006 12960
rect 24768 12922 24820 12928
rect 24412 12702 24532 12730
rect 23768 12406 23888 12434
rect 23388 12096 23440 12102
rect 23388 12038 23440 12044
rect 23400 11830 23428 12038
rect 23388 11824 23440 11830
rect 23388 11766 23440 11772
rect 22836 11756 22888 11762
rect 22836 11698 22888 11704
rect 22950 11452 23258 11461
rect 22950 11450 22956 11452
rect 23012 11450 23036 11452
rect 23092 11450 23116 11452
rect 23172 11450 23196 11452
rect 23252 11450 23258 11452
rect 23012 11398 23014 11450
rect 23194 11398 23196 11450
rect 22950 11396 22956 11398
rect 23012 11396 23036 11398
rect 23092 11396 23116 11398
rect 23172 11396 23196 11398
rect 23252 11396 23258 11398
rect 22950 11387 23258 11396
rect 23480 11076 23532 11082
rect 23480 11018 23532 11024
rect 22744 10804 22796 10810
rect 22744 10746 22796 10752
rect 23388 10736 23440 10742
rect 23388 10678 23440 10684
rect 22950 10364 23258 10373
rect 22950 10362 22956 10364
rect 23012 10362 23036 10364
rect 23092 10362 23116 10364
rect 23172 10362 23196 10364
rect 23252 10362 23258 10364
rect 23012 10310 23014 10362
rect 23194 10310 23196 10362
rect 22950 10308 22956 10310
rect 23012 10308 23036 10310
rect 23092 10308 23116 10310
rect 23172 10308 23196 10310
rect 23252 10308 23258 10310
rect 22950 10299 23258 10308
rect 22006 10095 22062 10104
rect 22284 10124 22336 10130
rect 22284 10066 22336 10072
rect 21916 9988 21968 9994
rect 21916 9930 21968 9936
rect 21928 9674 21956 9930
rect 21928 9646 22048 9674
rect 21824 8900 21876 8906
rect 21824 8842 21876 8848
rect 21732 8016 21784 8022
rect 21732 7958 21784 7964
rect 21732 4684 21784 4690
rect 21732 4626 21784 4632
rect 21744 3738 21772 4626
rect 21732 3732 21784 3738
rect 21732 3674 21784 3680
rect 21732 2984 21784 2990
rect 21732 2926 21784 2932
rect 21640 2576 21692 2582
rect 21640 2518 21692 2524
rect 21548 2508 21600 2514
rect 21548 2450 21600 2456
rect 21560 1834 21588 2450
rect 21548 1828 21600 1834
rect 21548 1770 21600 1776
rect 21744 800 21772 2926
rect 21836 1601 21864 8842
rect 22020 8566 22048 9646
rect 22100 9580 22152 9586
rect 22100 9522 22152 9528
rect 22008 8560 22060 8566
rect 22008 8502 22060 8508
rect 21916 7540 21968 7546
rect 21916 7482 21968 7488
rect 21928 7426 21956 7482
rect 22112 7426 22140 9522
rect 22296 9450 22324 10066
rect 23018 10024 23074 10033
rect 23018 9959 23074 9968
rect 23032 9586 23060 9959
rect 23294 9752 23350 9761
rect 23294 9687 23350 9696
rect 23308 9654 23336 9687
rect 23296 9648 23348 9654
rect 23296 9590 23348 9596
rect 23020 9580 23072 9586
rect 23020 9522 23072 9528
rect 23400 9466 23428 10678
rect 23492 10674 23520 11018
rect 23480 10668 23532 10674
rect 23480 10610 23532 10616
rect 23664 10600 23716 10606
rect 23664 10542 23716 10548
rect 22284 9444 22336 9450
rect 22284 9386 22336 9392
rect 23308 9438 23428 9466
rect 22950 9276 23258 9285
rect 22950 9274 22956 9276
rect 23012 9274 23036 9276
rect 23092 9274 23116 9276
rect 23172 9274 23196 9276
rect 23252 9274 23258 9276
rect 23012 9222 23014 9274
rect 23194 9222 23196 9274
rect 22950 9220 22956 9222
rect 23012 9220 23036 9222
rect 23092 9220 23116 9222
rect 23172 9220 23196 9222
rect 23252 9220 23258 9222
rect 22950 9211 23258 9220
rect 22376 8968 22428 8974
rect 22376 8910 22428 8916
rect 22192 8424 22244 8430
rect 22192 8366 22244 8372
rect 22284 8424 22336 8430
rect 22284 8366 22336 8372
rect 22204 8294 22232 8366
rect 22192 8288 22244 8294
rect 22192 8230 22244 8236
rect 22192 7880 22244 7886
rect 22192 7822 22244 7828
rect 21928 7398 22140 7426
rect 21916 7336 21968 7342
rect 21916 7278 21968 7284
rect 21928 5137 21956 7278
rect 22008 7268 22060 7274
rect 22008 7210 22060 7216
rect 22020 6882 22048 7210
rect 22100 7200 22152 7206
rect 22100 7142 22152 7148
rect 22112 7002 22140 7142
rect 22100 6996 22152 7002
rect 22100 6938 22152 6944
rect 22020 6854 22140 6882
rect 22112 6458 22140 6854
rect 22100 6452 22152 6458
rect 22100 6394 22152 6400
rect 22100 6180 22152 6186
rect 22100 6122 22152 6128
rect 21914 5128 21970 5137
rect 21914 5063 21970 5072
rect 22112 4264 22140 6122
rect 22020 4236 22140 4264
rect 22020 3890 22048 4236
rect 22100 4140 22152 4146
rect 22100 4082 22152 4088
rect 22112 4049 22140 4082
rect 22098 4040 22154 4049
rect 22098 3975 22154 3984
rect 22020 3862 22140 3890
rect 22112 2496 22140 3862
rect 22204 3194 22232 7822
rect 22296 6866 22324 8366
rect 22284 6860 22336 6866
rect 22284 6802 22336 6808
rect 22284 6452 22336 6458
rect 22284 6394 22336 6400
rect 22296 6066 22324 6394
rect 22388 6225 22416 8910
rect 22652 8832 22704 8838
rect 22652 8774 22704 8780
rect 22664 8566 22692 8774
rect 22652 8560 22704 8566
rect 22652 8502 22704 8508
rect 22744 8424 22796 8430
rect 22744 8366 22796 8372
rect 22560 7948 22612 7954
rect 22560 7890 22612 7896
rect 22468 7404 22520 7410
rect 22468 7346 22520 7352
rect 22480 6361 22508 7346
rect 22466 6352 22522 6361
rect 22466 6287 22522 6296
rect 22468 6248 22520 6254
rect 22374 6216 22430 6225
rect 22468 6190 22520 6196
rect 22374 6151 22430 6160
rect 22296 6038 22416 6066
rect 22284 5704 22336 5710
rect 22284 5646 22336 5652
rect 22296 4282 22324 5646
rect 22388 4321 22416 6038
rect 22374 4312 22430 4321
rect 22284 4276 22336 4282
rect 22374 4247 22430 4256
rect 22284 4218 22336 4224
rect 22192 3188 22244 3194
rect 22192 3130 22244 3136
rect 22480 2990 22508 6190
rect 22468 2984 22520 2990
rect 22468 2926 22520 2932
rect 22112 2468 22324 2496
rect 22008 2440 22060 2446
rect 22008 2382 22060 2388
rect 22098 2408 22154 2417
rect 22020 1970 22048 2382
rect 22098 2343 22100 2352
rect 22152 2343 22154 2352
rect 22100 2314 22152 2320
rect 22008 1964 22060 1970
rect 22008 1906 22060 1912
rect 21822 1592 21878 1601
rect 21822 1527 21878 1536
rect 22296 950 22324 2468
rect 22572 1034 22600 7890
rect 22756 6866 22784 8366
rect 22950 8188 23258 8197
rect 22950 8186 22956 8188
rect 23012 8186 23036 8188
rect 23092 8186 23116 8188
rect 23172 8186 23196 8188
rect 23252 8186 23258 8188
rect 23012 8134 23014 8186
rect 23194 8134 23196 8186
rect 22950 8132 22956 8134
rect 23012 8132 23036 8134
rect 23092 8132 23116 8134
rect 23172 8132 23196 8134
rect 23252 8132 23258 8134
rect 22950 8123 23258 8132
rect 23204 8016 23256 8022
rect 23204 7958 23256 7964
rect 22836 7744 22888 7750
rect 22836 7686 22888 7692
rect 22744 6860 22796 6866
rect 22744 6802 22796 6808
rect 22652 5772 22704 5778
rect 22652 5714 22704 5720
rect 22664 2854 22692 5714
rect 22848 4146 22876 7686
rect 23216 7546 23244 7958
rect 23308 7698 23336 9438
rect 23480 8900 23532 8906
rect 23480 8842 23532 8848
rect 23388 8288 23440 8294
rect 23388 8230 23440 8236
rect 23400 7818 23428 8230
rect 23388 7812 23440 7818
rect 23388 7754 23440 7760
rect 23308 7670 23428 7698
rect 23204 7540 23256 7546
rect 23204 7482 23256 7488
rect 23296 7336 23348 7342
rect 23296 7278 23348 7284
rect 22950 7100 23258 7109
rect 22950 7098 22956 7100
rect 23012 7098 23036 7100
rect 23092 7098 23116 7100
rect 23172 7098 23196 7100
rect 23252 7098 23258 7100
rect 23012 7046 23014 7098
rect 23194 7046 23196 7098
rect 22950 7044 22956 7046
rect 23012 7044 23036 7046
rect 23092 7044 23116 7046
rect 23172 7044 23196 7046
rect 23252 7044 23258 7046
rect 22950 7035 23258 7044
rect 22950 6012 23258 6021
rect 22950 6010 22956 6012
rect 23012 6010 23036 6012
rect 23092 6010 23116 6012
rect 23172 6010 23196 6012
rect 23252 6010 23258 6012
rect 23012 5958 23014 6010
rect 23194 5958 23196 6010
rect 22950 5956 22956 5958
rect 23012 5956 23036 5958
rect 23092 5956 23116 5958
rect 23172 5956 23196 5958
rect 23252 5956 23258 5958
rect 22950 5947 23258 5956
rect 23308 5681 23336 7278
rect 23400 7041 23428 7670
rect 23386 7032 23442 7041
rect 23386 6967 23442 6976
rect 23388 6928 23440 6934
rect 23388 6870 23440 6876
rect 23400 5710 23428 6870
rect 23388 5704 23440 5710
rect 23294 5672 23350 5681
rect 23388 5646 23440 5652
rect 23294 5607 23350 5616
rect 23386 5536 23442 5545
rect 23386 5471 23442 5480
rect 22950 4924 23258 4933
rect 22950 4922 22956 4924
rect 23012 4922 23036 4924
rect 23092 4922 23116 4924
rect 23172 4922 23196 4924
rect 23252 4922 23258 4924
rect 23012 4870 23014 4922
rect 23194 4870 23196 4922
rect 22950 4868 22956 4870
rect 23012 4868 23036 4870
rect 23092 4868 23116 4870
rect 23172 4868 23196 4870
rect 23252 4868 23258 4870
rect 22950 4859 23258 4868
rect 22928 4208 22980 4214
rect 22928 4150 22980 4156
rect 22836 4140 22888 4146
rect 22836 4082 22888 4088
rect 22940 4010 22968 4150
rect 22928 4004 22980 4010
rect 22928 3946 22980 3952
rect 22950 3836 23258 3845
rect 22950 3834 22956 3836
rect 23012 3834 23036 3836
rect 23092 3834 23116 3836
rect 23172 3834 23196 3836
rect 23252 3834 23258 3836
rect 23012 3782 23014 3834
rect 23194 3782 23196 3834
rect 22950 3780 22956 3782
rect 23012 3780 23036 3782
rect 23092 3780 23116 3782
rect 23172 3780 23196 3782
rect 23252 3780 23258 3782
rect 22742 3768 22798 3777
rect 22950 3771 23258 3780
rect 22742 3703 22744 3712
rect 22796 3703 22798 3712
rect 22744 3674 22796 3680
rect 22926 3632 22982 3641
rect 22836 3596 22888 3602
rect 22926 3567 22982 3576
rect 22836 3538 22888 3544
rect 22652 2848 22704 2854
rect 22652 2790 22704 2796
rect 22388 1006 22600 1034
rect 22284 944 22336 950
rect 22112 870 22232 898
rect 22284 886 22336 892
rect 22112 800 22140 870
rect 18156 734 18368 762
rect 18418 0 18474 800
rect 18786 0 18842 800
rect 19154 0 19210 800
rect 19522 0 19578 800
rect 19890 0 19946 800
rect 20258 0 20314 800
rect 20626 0 20682 800
rect 20994 0 21050 800
rect 21362 0 21418 800
rect 21730 0 21786 800
rect 22098 0 22154 800
rect 22204 762 22232 870
rect 22388 762 22416 1006
rect 22468 944 22520 950
rect 22468 886 22520 892
rect 22480 800 22508 886
rect 22848 800 22876 3538
rect 22940 3194 22968 3567
rect 23204 3392 23256 3398
rect 23204 3334 23256 3340
rect 23216 3233 23244 3334
rect 23202 3224 23258 3233
rect 22928 3188 22980 3194
rect 23202 3159 23258 3168
rect 22928 3130 22980 3136
rect 23400 3126 23428 5471
rect 23492 3738 23520 8842
rect 23572 7744 23624 7750
rect 23572 7686 23624 7692
rect 23480 3732 23532 3738
rect 23480 3674 23532 3680
rect 23388 3120 23440 3126
rect 23388 3062 23440 3068
rect 23296 2916 23348 2922
rect 23296 2858 23348 2864
rect 22950 2748 23258 2757
rect 22950 2746 22956 2748
rect 23012 2746 23036 2748
rect 23092 2746 23116 2748
rect 23172 2746 23196 2748
rect 23252 2746 23258 2748
rect 23012 2694 23014 2746
rect 23194 2694 23196 2746
rect 22950 2692 22956 2694
rect 23012 2692 23036 2694
rect 23092 2692 23116 2694
rect 23172 2692 23196 2694
rect 23252 2692 23258 2694
rect 22950 2683 23258 2692
rect 23308 1578 23336 2858
rect 23216 1550 23336 1578
rect 23216 800 23244 1550
rect 23584 800 23612 7686
rect 23676 5234 23704 10542
rect 23756 7200 23808 7206
rect 23756 7142 23808 7148
rect 23664 5228 23716 5234
rect 23664 5170 23716 5176
rect 23768 4826 23796 7142
rect 23756 4820 23808 4826
rect 23756 4762 23808 4768
rect 23860 2650 23888 12406
rect 23938 10704 23994 10713
rect 23938 10639 23940 10648
rect 23992 10639 23994 10648
rect 23940 10610 23992 10616
rect 24412 10266 24440 12702
rect 24780 12238 24808 12922
rect 25056 12900 25084 14214
rect 25148 14006 25176 14583
rect 25136 14000 25188 14006
rect 25136 13942 25188 13948
rect 25136 12912 25188 12918
rect 25056 12872 25136 12900
rect 25136 12854 25188 12860
rect 25148 12646 25176 12854
rect 25976 12753 26004 22066
rect 26160 17882 26188 42570
rect 26240 32972 26292 32978
rect 26240 32914 26292 32920
rect 26252 27538 26280 32914
rect 26528 32570 26556 52430
rect 26608 37732 26660 37738
rect 26608 37674 26660 37680
rect 26516 32564 26568 32570
rect 26516 32506 26568 32512
rect 26240 27532 26292 27538
rect 26240 27474 26292 27480
rect 26148 17876 26200 17882
rect 26148 17818 26200 17824
rect 26620 13802 26648 37674
rect 26700 36644 26752 36650
rect 26700 36586 26752 36592
rect 26712 14113 26740 36586
rect 26804 30054 26832 53926
rect 26792 30048 26844 30054
rect 26792 29990 26844 29996
rect 26698 14104 26754 14113
rect 26698 14039 26754 14048
rect 26608 13796 26660 13802
rect 26608 13738 26660 13744
rect 25962 12744 26018 12753
rect 25962 12679 26018 12688
rect 25136 12640 25188 12646
rect 25136 12582 25188 12588
rect 24768 12232 24820 12238
rect 24768 12174 24820 12180
rect 24950 12200 25006 12209
rect 24950 12135 24952 12144
rect 25004 12135 25006 12144
rect 24952 12106 25004 12112
rect 25148 11830 25176 12582
rect 25136 11824 25188 11830
rect 25136 11766 25188 11772
rect 25148 11558 25176 11766
rect 24584 11552 24636 11558
rect 24584 11494 24636 11500
rect 25136 11552 25188 11558
rect 25136 11494 25188 11500
rect 24596 11150 24624 11494
rect 24766 11384 24822 11393
rect 24766 11319 24822 11328
rect 24584 11144 24636 11150
rect 24584 11086 24636 11092
rect 24780 10606 24808 11319
rect 24768 10600 24820 10606
rect 24674 10568 24730 10577
rect 24768 10542 24820 10548
rect 24674 10503 24730 10512
rect 24400 10260 24452 10266
rect 24400 10202 24452 10208
rect 24124 10192 24176 10198
rect 24124 10134 24176 10140
rect 24032 9920 24084 9926
rect 24032 9862 24084 9868
rect 24044 9518 24072 9862
rect 24032 9512 24084 9518
rect 24032 9454 24084 9460
rect 24044 8974 24072 9454
rect 24032 8968 24084 8974
rect 24032 8910 24084 8916
rect 24032 8560 24084 8566
rect 24136 8548 24164 10134
rect 24084 8520 24164 8548
rect 24032 8502 24084 8508
rect 24044 7750 24072 8502
rect 24032 7744 24084 7750
rect 24032 7686 24084 7692
rect 24044 6662 24072 7686
rect 24032 6656 24084 6662
rect 24032 6598 24084 6604
rect 23940 6316 23992 6322
rect 23940 6258 23992 6264
rect 23952 5914 23980 6258
rect 23940 5908 23992 5914
rect 23940 5850 23992 5856
rect 24044 5574 24072 6598
rect 24032 5568 24084 5574
rect 24032 5510 24084 5516
rect 24216 5568 24268 5574
rect 24216 5510 24268 5516
rect 24044 3942 24072 5510
rect 24228 5370 24256 5510
rect 24216 5364 24268 5370
rect 24216 5306 24268 5312
rect 24032 3936 24084 3942
rect 24032 3878 24084 3884
rect 23938 3496 23994 3505
rect 23938 3431 23994 3440
rect 23848 2644 23900 2650
rect 23848 2586 23900 2592
rect 23952 800 23980 3431
rect 24044 3194 24072 3878
rect 24412 3534 24440 10202
rect 24584 9920 24636 9926
rect 24582 9888 24584 9897
rect 24636 9888 24638 9897
rect 24582 9823 24638 9832
rect 24688 9518 24716 10503
rect 25148 10266 25176 11494
rect 25228 11008 25280 11014
rect 25228 10950 25280 10956
rect 25136 10260 25188 10266
rect 25136 10202 25188 10208
rect 25240 10130 25268 10950
rect 25228 10124 25280 10130
rect 25228 10066 25280 10072
rect 24676 9512 24728 9518
rect 24676 9454 24728 9460
rect 25044 9172 25096 9178
rect 25044 9114 25096 9120
rect 24950 8936 25006 8945
rect 24950 8871 24952 8880
rect 25004 8871 25006 8880
rect 24952 8842 25004 8848
rect 24860 8492 24912 8498
rect 24860 8434 24912 8440
rect 24674 7304 24730 7313
rect 24674 7239 24730 7248
rect 24582 6760 24638 6769
rect 24582 6695 24638 6704
rect 24596 6662 24624 6695
rect 24584 6656 24636 6662
rect 24584 6598 24636 6604
rect 24688 6254 24716 7239
rect 24872 6934 24900 8434
rect 24952 7540 25004 7546
rect 24952 7482 25004 7488
rect 24860 6928 24912 6934
rect 24860 6870 24912 6876
rect 24964 6746 24992 7482
rect 25056 6866 25084 9114
rect 25228 8288 25280 8294
rect 25228 8230 25280 8236
rect 25134 8120 25190 8129
rect 25134 8055 25190 8064
rect 25148 7478 25176 8055
rect 25136 7472 25188 7478
rect 25136 7414 25188 7420
rect 25240 7002 25268 8230
rect 25228 6996 25280 7002
rect 25228 6938 25280 6944
rect 25044 6860 25096 6866
rect 25044 6802 25096 6808
rect 24964 6718 25084 6746
rect 24952 6656 25004 6662
rect 24952 6598 25004 6604
rect 24766 6488 24822 6497
rect 24766 6423 24822 6432
rect 24676 6248 24728 6254
rect 24676 6190 24728 6196
rect 24780 5166 24808 6423
rect 24860 6384 24912 6390
rect 24860 6326 24912 6332
rect 24768 5160 24820 5166
rect 24768 5102 24820 5108
rect 24872 3670 24900 6326
rect 24964 5914 24992 6598
rect 24952 5908 25004 5914
rect 24952 5850 25004 5856
rect 25056 4758 25084 6718
rect 25044 4752 25096 4758
rect 25044 4694 25096 4700
rect 24860 3664 24912 3670
rect 24860 3606 24912 3612
rect 24400 3528 24452 3534
rect 24400 3470 24452 3476
rect 24032 3188 24084 3194
rect 24032 3130 24084 3136
rect 24308 3052 24360 3058
rect 24308 2994 24360 3000
rect 24768 3052 24820 3058
rect 24768 2994 24820 3000
rect 24320 800 24348 2994
rect 24780 2650 24808 2994
rect 24858 2952 24914 2961
rect 24858 2887 24914 2896
rect 24768 2644 24820 2650
rect 24768 2586 24820 2592
rect 24768 2304 24820 2310
rect 24768 2246 24820 2252
rect 24780 2106 24808 2246
rect 24768 2100 24820 2106
rect 24768 2042 24820 2048
rect 22204 734 22416 762
rect 22466 0 22522 800
rect 22834 0 22890 800
rect 23202 0 23258 800
rect 23570 0 23626 800
rect 23938 0 23994 800
rect 24306 0 24362 800
rect 24674 0 24730 800
rect 24872 785 24900 2887
rect 24858 776 24914 785
rect 24858 711 24914 720
rect 25042 0 25098 800
<< via2 >>
rect 2956 53882 3012 53884
rect 3036 53882 3092 53884
rect 3116 53882 3172 53884
rect 3196 53882 3252 53884
rect 2956 53830 3002 53882
rect 3002 53830 3012 53882
rect 3036 53830 3066 53882
rect 3066 53830 3078 53882
rect 3078 53830 3092 53882
rect 3116 53830 3130 53882
rect 3130 53830 3142 53882
rect 3142 53830 3172 53882
rect 3196 53830 3206 53882
rect 3206 53830 3252 53882
rect 2956 53828 3012 53830
rect 3036 53828 3092 53830
rect 3116 53828 3172 53830
rect 3196 53828 3252 53830
rect 2956 52794 3012 52796
rect 3036 52794 3092 52796
rect 3116 52794 3172 52796
rect 3196 52794 3252 52796
rect 2956 52742 3002 52794
rect 3002 52742 3012 52794
rect 3036 52742 3066 52794
rect 3066 52742 3078 52794
rect 3078 52742 3092 52794
rect 3116 52742 3130 52794
rect 3130 52742 3142 52794
rect 3142 52742 3172 52794
rect 3196 52742 3206 52794
rect 3206 52742 3252 52794
rect 2956 52740 3012 52742
rect 3036 52740 3092 52742
rect 3116 52740 3172 52742
rect 3196 52740 3252 52742
rect 2956 51706 3012 51708
rect 3036 51706 3092 51708
rect 3116 51706 3172 51708
rect 3196 51706 3252 51708
rect 2956 51654 3002 51706
rect 3002 51654 3012 51706
rect 3036 51654 3066 51706
rect 3066 51654 3078 51706
rect 3078 51654 3092 51706
rect 3116 51654 3130 51706
rect 3130 51654 3142 51706
rect 3142 51654 3172 51706
rect 3196 51654 3206 51706
rect 3206 51654 3252 51706
rect 2956 51652 3012 51654
rect 3036 51652 3092 51654
rect 3116 51652 3172 51654
rect 3196 51652 3252 51654
rect 7956 54426 8012 54428
rect 8036 54426 8092 54428
rect 8116 54426 8172 54428
rect 8196 54426 8252 54428
rect 7956 54374 8002 54426
rect 8002 54374 8012 54426
rect 8036 54374 8066 54426
rect 8066 54374 8078 54426
rect 8078 54374 8092 54426
rect 8116 54374 8130 54426
rect 8130 54374 8142 54426
rect 8142 54374 8172 54426
rect 8196 54374 8206 54426
rect 8206 54374 8252 54426
rect 7956 54372 8012 54374
rect 8036 54372 8092 54374
rect 8116 54372 8172 54374
rect 8196 54372 8252 54374
rect 7956 53338 8012 53340
rect 8036 53338 8092 53340
rect 8116 53338 8172 53340
rect 8196 53338 8252 53340
rect 7956 53286 8002 53338
rect 8002 53286 8012 53338
rect 8036 53286 8066 53338
rect 8066 53286 8078 53338
rect 8078 53286 8092 53338
rect 8116 53286 8130 53338
rect 8130 53286 8142 53338
rect 8142 53286 8172 53338
rect 8196 53286 8206 53338
rect 8206 53286 8252 53338
rect 7956 53284 8012 53286
rect 8036 53284 8092 53286
rect 8116 53284 8172 53286
rect 8196 53284 8252 53286
rect 7956 52250 8012 52252
rect 8036 52250 8092 52252
rect 8116 52250 8172 52252
rect 8196 52250 8252 52252
rect 7956 52198 8002 52250
rect 8002 52198 8012 52250
rect 8036 52198 8066 52250
rect 8066 52198 8078 52250
rect 8078 52198 8092 52250
rect 8116 52198 8130 52250
rect 8130 52198 8142 52250
rect 8142 52198 8172 52250
rect 8196 52198 8206 52250
rect 8206 52198 8252 52250
rect 7956 52196 8012 52198
rect 8036 52196 8092 52198
rect 8116 52196 8172 52198
rect 8196 52196 8252 52198
rect 2956 50618 3012 50620
rect 3036 50618 3092 50620
rect 3116 50618 3172 50620
rect 3196 50618 3252 50620
rect 2956 50566 3002 50618
rect 3002 50566 3012 50618
rect 3036 50566 3066 50618
rect 3066 50566 3078 50618
rect 3078 50566 3092 50618
rect 3116 50566 3130 50618
rect 3130 50566 3142 50618
rect 3142 50566 3172 50618
rect 3196 50566 3206 50618
rect 3206 50566 3252 50618
rect 2956 50564 3012 50566
rect 3036 50564 3092 50566
rect 3116 50564 3172 50566
rect 3196 50564 3252 50566
rect 2956 49530 3012 49532
rect 3036 49530 3092 49532
rect 3116 49530 3172 49532
rect 3196 49530 3252 49532
rect 2956 49478 3002 49530
rect 3002 49478 3012 49530
rect 3036 49478 3066 49530
rect 3066 49478 3078 49530
rect 3078 49478 3092 49530
rect 3116 49478 3130 49530
rect 3130 49478 3142 49530
rect 3142 49478 3172 49530
rect 3196 49478 3206 49530
rect 3206 49478 3252 49530
rect 2956 49476 3012 49478
rect 3036 49476 3092 49478
rect 3116 49476 3172 49478
rect 3196 49476 3252 49478
rect 7956 51162 8012 51164
rect 8036 51162 8092 51164
rect 8116 51162 8172 51164
rect 8196 51162 8252 51164
rect 7956 51110 8002 51162
rect 8002 51110 8012 51162
rect 8036 51110 8066 51162
rect 8066 51110 8078 51162
rect 8078 51110 8092 51162
rect 8116 51110 8130 51162
rect 8130 51110 8142 51162
rect 8142 51110 8172 51162
rect 8196 51110 8206 51162
rect 8206 51110 8252 51162
rect 7956 51108 8012 51110
rect 8036 51108 8092 51110
rect 8116 51108 8172 51110
rect 8196 51108 8252 51110
rect 7956 50074 8012 50076
rect 8036 50074 8092 50076
rect 8116 50074 8172 50076
rect 8196 50074 8252 50076
rect 7956 50022 8002 50074
rect 8002 50022 8012 50074
rect 8036 50022 8066 50074
rect 8066 50022 8078 50074
rect 8078 50022 8092 50074
rect 8116 50022 8130 50074
rect 8130 50022 8142 50074
rect 8142 50022 8172 50074
rect 8196 50022 8206 50074
rect 8206 50022 8252 50074
rect 7956 50020 8012 50022
rect 8036 50020 8092 50022
rect 8116 50020 8172 50022
rect 8196 50020 8252 50022
rect 7956 48986 8012 48988
rect 8036 48986 8092 48988
rect 8116 48986 8172 48988
rect 8196 48986 8252 48988
rect 7956 48934 8002 48986
rect 8002 48934 8012 48986
rect 8036 48934 8066 48986
rect 8066 48934 8078 48986
rect 8078 48934 8092 48986
rect 8116 48934 8130 48986
rect 8130 48934 8142 48986
rect 8142 48934 8172 48986
rect 8196 48934 8206 48986
rect 8206 48934 8252 48986
rect 7956 48932 8012 48934
rect 8036 48932 8092 48934
rect 8116 48932 8172 48934
rect 8196 48932 8252 48934
rect 2956 48442 3012 48444
rect 3036 48442 3092 48444
rect 3116 48442 3172 48444
rect 3196 48442 3252 48444
rect 2956 48390 3002 48442
rect 3002 48390 3012 48442
rect 3036 48390 3066 48442
rect 3066 48390 3078 48442
rect 3078 48390 3092 48442
rect 3116 48390 3130 48442
rect 3130 48390 3142 48442
rect 3142 48390 3172 48442
rect 3196 48390 3206 48442
rect 3206 48390 3252 48442
rect 2956 48388 3012 48390
rect 3036 48388 3092 48390
rect 3116 48388 3172 48390
rect 3196 48388 3252 48390
rect 2956 47354 3012 47356
rect 3036 47354 3092 47356
rect 3116 47354 3172 47356
rect 3196 47354 3252 47356
rect 2956 47302 3002 47354
rect 3002 47302 3012 47354
rect 3036 47302 3066 47354
rect 3066 47302 3078 47354
rect 3078 47302 3092 47354
rect 3116 47302 3130 47354
rect 3130 47302 3142 47354
rect 3142 47302 3172 47354
rect 3196 47302 3206 47354
rect 3206 47302 3252 47354
rect 2956 47300 3012 47302
rect 3036 47300 3092 47302
rect 3116 47300 3172 47302
rect 3196 47300 3252 47302
rect 2956 46266 3012 46268
rect 3036 46266 3092 46268
rect 3116 46266 3172 46268
rect 3196 46266 3252 46268
rect 2956 46214 3002 46266
rect 3002 46214 3012 46266
rect 3036 46214 3066 46266
rect 3066 46214 3078 46266
rect 3078 46214 3092 46266
rect 3116 46214 3130 46266
rect 3130 46214 3142 46266
rect 3142 46214 3172 46266
rect 3196 46214 3206 46266
rect 3206 46214 3252 46266
rect 2956 46212 3012 46214
rect 3036 46212 3092 46214
rect 3116 46212 3172 46214
rect 3196 46212 3252 46214
rect 2956 45178 3012 45180
rect 3036 45178 3092 45180
rect 3116 45178 3172 45180
rect 3196 45178 3252 45180
rect 2956 45126 3002 45178
rect 3002 45126 3012 45178
rect 3036 45126 3066 45178
rect 3066 45126 3078 45178
rect 3078 45126 3092 45178
rect 3116 45126 3130 45178
rect 3130 45126 3142 45178
rect 3142 45126 3172 45178
rect 3196 45126 3206 45178
rect 3206 45126 3252 45178
rect 2956 45124 3012 45126
rect 3036 45124 3092 45126
rect 3116 45124 3172 45126
rect 3196 45124 3252 45126
rect 2956 44090 3012 44092
rect 3036 44090 3092 44092
rect 3116 44090 3172 44092
rect 3196 44090 3252 44092
rect 2956 44038 3002 44090
rect 3002 44038 3012 44090
rect 3036 44038 3066 44090
rect 3066 44038 3078 44090
rect 3078 44038 3092 44090
rect 3116 44038 3130 44090
rect 3130 44038 3142 44090
rect 3142 44038 3172 44090
rect 3196 44038 3206 44090
rect 3206 44038 3252 44090
rect 2956 44036 3012 44038
rect 3036 44036 3092 44038
rect 3116 44036 3172 44038
rect 3196 44036 3252 44038
rect 2956 43002 3012 43004
rect 3036 43002 3092 43004
rect 3116 43002 3172 43004
rect 3196 43002 3252 43004
rect 2956 42950 3002 43002
rect 3002 42950 3012 43002
rect 3036 42950 3066 43002
rect 3066 42950 3078 43002
rect 3078 42950 3092 43002
rect 3116 42950 3130 43002
rect 3130 42950 3142 43002
rect 3142 42950 3172 43002
rect 3196 42950 3206 43002
rect 3206 42950 3252 43002
rect 2956 42948 3012 42950
rect 3036 42948 3092 42950
rect 3116 42948 3172 42950
rect 3196 42948 3252 42950
rect 2956 41914 3012 41916
rect 3036 41914 3092 41916
rect 3116 41914 3172 41916
rect 3196 41914 3252 41916
rect 2956 41862 3002 41914
rect 3002 41862 3012 41914
rect 3036 41862 3066 41914
rect 3066 41862 3078 41914
rect 3078 41862 3092 41914
rect 3116 41862 3130 41914
rect 3130 41862 3142 41914
rect 3142 41862 3172 41914
rect 3196 41862 3206 41914
rect 3206 41862 3252 41914
rect 2956 41860 3012 41862
rect 3036 41860 3092 41862
rect 3116 41860 3172 41862
rect 3196 41860 3252 41862
rect 2956 40826 3012 40828
rect 3036 40826 3092 40828
rect 3116 40826 3172 40828
rect 3196 40826 3252 40828
rect 2956 40774 3002 40826
rect 3002 40774 3012 40826
rect 3036 40774 3066 40826
rect 3066 40774 3078 40826
rect 3078 40774 3092 40826
rect 3116 40774 3130 40826
rect 3130 40774 3142 40826
rect 3142 40774 3172 40826
rect 3196 40774 3206 40826
rect 3206 40774 3252 40826
rect 2956 40772 3012 40774
rect 3036 40772 3092 40774
rect 3116 40772 3172 40774
rect 3196 40772 3252 40774
rect 2956 39738 3012 39740
rect 3036 39738 3092 39740
rect 3116 39738 3172 39740
rect 3196 39738 3252 39740
rect 2956 39686 3002 39738
rect 3002 39686 3012 39738
rect 3036 39686 3066 39738
rect 3066 39686 3078 39738
rect 3078 39686 3092 39738
rect 3116 39686 3130 39738
rect 3130 39686 3142 39738
rect 3142 39686 3172 39738
rect 3196 39686 3206 39738
rect 3206 39686 3252 39738
rect 2956 39684 3012 39686
rect 3036 39684 3092 39686
rect 3116 39684 3172 39686
rect 3196 39684 3252 39686
rect 7956 47898 8012 47900
rect 8036 47898 8092 47900
rect 8116 47898 8172 47900
rect 8196 47898 8252 47900
rect 7956 47846 8002 47898
rect 8002 47846 8012 47898
rect 8036 47846 8066 47898
rect 8066 47846 8078 47898
rect 8078 47846 8092 47898
rect 8116 47846 8130 47898
rect 8130 47846 8142 47898
rect 8142 47846 8172 47898
rect 8196 47846 8206 47898
rect 8206 47846 8252 47898
rect 7956 47844 8012 47846
rect 8036 47844 8092 47846
rect 8116 47844 8172 47846
rect 8196 47844 8252 47846
rect 7956 46810 8012 46812
rect 8036 46810 8092 46812
rect 8116 46810 8172 46812
rect 8196 46810 8252 46812
rect 7956 46758 8002 46810
rect 8002 46758 8012 46810
rect 8036 46758 8066 46810
rect 8066 46758 8078 46810
rect 8078 46758 8092 46810
rect 8116 46758 8130 46810
rect 8130 46758 8142 46810
rect 8142 46758 8172 46810
rect 8196 46758 8206 46810
rect 8206 46758 8252 46810
rect 7956 46756 8012 46758
rect 8036 46756 8092 46758
rect 8116 46756 8172 46758
rect 8196 46756 8252 46758
rect 7956 45722 8012 45724
rect 8036 45722 8092 45724
rect 8116 45722 8172 45724
rect 8196 45722 8252 45724
rect 7956 45670 8002 45722
rect 8002 45670 8012 45722
rect 8036 45670 8066 45722
rect 8066 45670 8078 45722
rect 8078 45670 8092 45722
rect 8116 45670 8130 45722
rect 8130 45670 8142 45722
rect 8142 45670 8172 45722
rect 8196 45670 8206 45722
rect 8206 45670 8252 45722
rect 7956 45668 8012 45670
rect 8036 45668 8092 45670
rect 8116 45668 8172 45670
rect 8196 45668 8252 45670
rect 7956 44634 8012 44636
rect 8036 44634 8092 44636
rect 8116 44634 8172 44636
rect 8196 44634 8252 44636
rect 7956 44582 8002 44634
rect 8002 44582 8012 44634
rect 8036 44582 8066 44634
rect 8066 44582 8078 44634
rect 8078 44582 8092 44634
rect 8116 44582 8130 44634
rect 8130 44582 8142 44634
rect 8142 44582 8172 44634
rect 8196 44582 8206 44634
rect 8206 44582 8252 44634
rect 7956 44580 8012 44582
rect 8036 44580 8092 44582
rect 8116 44580 8172 44582
rect 8196 44580 8252 44582
rect 7956 43546 8012 43548
rect 8036 43546 8092 43548
rect 8116 43546 8172 43548
rect 8196 43546 8252 43548
rect 7956 43494 8002 43546
rect 8002 43494 8012 43546
rect 8036 43494 8066 43546
rect 8066 43494 8078 43546
rect 8078 43494 8092 43546
rect 8116 43494 8130 43546
rect 8130 43494 8142 43546
rect 8142 43494 8172 43546
rect 8196 43494 8206 43546
rect 8206 43494 8252 43546
rect 7956 43492 8012 43494
rect 8036 43492 8092 43494
rect 8116 43492 8172 43494
rect 8196 43492 8252 43494
rect 7956 42458 8012 42460
rect 8036 42458 8092 42460
rect 8116 42458 8172 42460
rect 8196 42458 8252 42460
rect 7956 42406 8002 42458
rect 8002 42406 8012 42458
rect 8036 42406 8066 42458
rect 8066 42406 8078 42458
rect 8078 42406 8092 42458
rect 8116 42406 8130 42458
rect 8130 42406 8142 42458
rect 8142 42406 8172 42458
rect 8196 42406 8206 42458
rect 8206 42406 8252 42458
rect 7956 42404 8012 42406
rect 8036 42404 8092 42406
rect 8116 42404 8172 42406
rect 8196 42404 8252 42406
rect 7956 41370 8012 41372
rect 8036 41370 8092 41372
rect 8116 41370 8172 41372
rect 8196 41370 8252 41372
rect 7956 41318 8002 41370
rect 8002 41318 8012 41370
rect 8036 41318 8066 41370
rect 8066 41318 8078 41370
rect 8078 41318 8092 41370
rect 8116 41318 8130 41370
rect 8130 41318 8142 41370
rect 8142 41318 8172 41370
rect 8196 41318 8206 41370
rect 8206 41318 8252 41370
rect 7956 41316 8012 41318
rect 8036 41316 8092 41318
rect 8116 41316 8172 41318
rect 8196 41316 8252 41318
rect 7956 40282 8012 40284
rect 8036 40282 8092 40284
rect 8116 40282 8172 40284
rect 8196 40282 8252 40284
rect 7956 40230 8002 40282
rect 8002 40230 8012 40282
rect 8036 40230 8066 40282
rect 8066 40230 8078 40282
rect 8078 40230 8092 40282
rect 8116 40230 8130 40282
rect 8130 40230 8142 40282
rect 8142 40230 8172 40282
rect 8196 40230 8206 40282
rect 8206 40230 8252 40282
rect 7956 40228 8012 40230
rect 8036 40228 8092 40230
rect 8116 40228 8172 40230
rect 8196 40228 8252 40230
rect 7956 39194 8012 39196
rect 8036 39194 8092 39196
rect 8116 39194 8172 39196
rect 8196 39194 8252 39196
rect 7956 39142 8002 39194
rect 8002 39142 8012 39194
rect 8036 39142 8066 39194
rect 8066 39142 8078 39194
rect 8078 39142 8092 39194
rect 8116 39142 8130 39194
rect 8130 39142 8142 39194
rect 8142 39142 8172 39194
rect 8196 39142 8206 39194
rect 8206 39142 8252 39194
rect 7956 39140 8012 39142
rect 8036 39140 8092 39142
rect 8116 39140 8172 39142
rect 8196 39140 8252 39142
rect 2956 38650 3012 38652
rect 3036 38650 3092 38652
rect 3116 38650 3172 38652
rect 3196 38650 3252 38652
rect 2956 38598 3002 38650
rect 3002 38598 3012 38650
rect 3036 38598 3066 38650
rect 3066 38598 3078 38650
rect 3078 38598 3092 38650
rect 3116 38598 3130 38650
rect 3130 38598 3142 38650
rect 3142 38598 3172 38650
rect 3196 38598 3206 38650
rect 3206 38598 3252 38650
rect 2956 38596 3012 38598
rect 3036 38596 3092 38598
rect 3116 38596 3172 38598
rect 3196 38596 3252 38598
rect 7956 38106 8012 38108
rect 8036 38106 8092 38108
rect 8116 38106 8172 38108
rect 8196 38106 8252 38108
rect 7956 38054 8002 38106
rect 8002 38054 8012 38106
rect 8036 38054 8066 38106
rect 8066 38054 8078 38106
rect 8078 38054 8092 38106
rect 8116 38054 8130 38106
rect 8130 38054 8142 38106
rect 8142 38054 8172 38106
rect 8196 38054 8206 38106
rect 8206 38054 8252 38106
rect 7956 38052 8012 38054
rect 8036 38052 8092 38054
rect 8116 38052 8172 38054
rect 8196 38052 8252 38054
rect 2956 37562 3012 37564
rect 3036 37562 3092 37564
rect 3116 37562 3172 37564
rect 3196 37562 3252 37564
rect 2956 37510 3002 37562
rect 3002 37510 3012 37562
rect 3036 37510 3066 37562
rect 3066 37510 3078 37562
rect 3078 37510 3092 37562
rect 3116 37510 3130 37562
rect 3130 37510 3142 37562
rect 3142 37510 3172 37562
rect 3196 37510 3206 37562
rect 3206 37510 3252 37562
rect 2956 37508 3012 37510
rect 3036 37508 3092 37510
rect 3116 37508 3172 37510
rect 3196 37508 3252 37510
rect 7956 37018 8012 37020
rect 8036 37018 8092 37020
rect 8116 37018 8172 37020
rect 8196 37018 8252 37020
rect 7956 36966 8002 37018
rect 8002 36966 8012 37018
rect 8036 36966 8066 37018
rect 8066 36966 8078 37018
rect 8078 36966 8092 37018
rect 8116 36966 8130 37018
rect 8130 36966 8142 37018
rect 8142 36966 8172 37018
rect 8196 36966 8206 37018
rect 8206 36966 8252 37018
rect 7956 36964 8012 36966
rect 8036 36964 8092 36966
rect 8116 36964 8172 36966
rect 8196 36964 8252 36966
rect 2956 36474 3012 36476
rect 3036 36474 3092 36476
rect 3116 36474 3172 36476
rect 3196 36474 3252 36476
rect 2956 36422 3002 36474
rect 3002 36422 3012 36474
rect 3036 36422 3066 36474
rect 3066 36422 3078 36474
rect 3078 36422 3092 36474
rect 3116 36422 3130 36474
rect 3130 36422 3142 36474
rect 3142 36422 3172 36474
rect 3196 36422 3206 36474
rect 3206 36422 3252 36474
rect 2956 36420 3012 36422
rect 3036 36420 3092 36422
rect 3116 36420 3172 36422
rect 3196 36420 3252 36422
rect 7956 35930 8012 35932
rect 8036 35930 8092 35932
rect 8116 35930 8172 35932
rect 8196 35930 8252 35932
rect 7956 35878 8002 35930
rect 8002 35878 8012 35930
rect 8036 35878 8066 35930
rect 8066 35878 8078 35930
rect 8078 35878 8092 35930
rect 8116 35878 8130 35930
rect 8130 35878 8142 35930
rect 8142 35878 8172 35930
rect 8196 35878 8206 35930
rect 8206 35878 8252 35930
rect 7956 35876 8012 35878
rect 8036 35876 8092 35878
rect 8116 35876 8172 35878
rect 8196 35876 8252 35878
rect 2956 35386 3012 35388
rect 3036 35386 3092 35388
rect 3116 35386 3172 35388
rect 3196 35386 3252 35388
rect 2956 35334 3002 35386
rect 3002 35334 3012 35386
rect 3036 35334 3066 35386
rect 3066 35334 3078 35386
rect 3078 35334 3092 35386
rect 3116 35334 3130 35386
rect 3130 35334 3142 35386
rect 3142 35334 3172 35386
rect 3196 35334 3206 35386
rect 3206 35334 3252 35386
rect 2956 35332 3012 35334
rect 3036 35332 3092 35334
rect 3116 35332 3172 35334
rect 3196 35332 3252 35334
rect 7956 34842 8012 34844
rect 8036 34842 8092 34844
rect 8116 34842 8172 34844
rect 8196 34842 8252 34844
rect 7956 34790 8002 34842
rect 8002 34790 8012 34842
rect 8036 34790 8066 34842
rect 8066 34790 8078 34842
rect 8078 34790 8092 34842
rect 8116 34790 8130 34842
rect 8130 34790 8142 34842
rect 8142 34790 8172 34842
rect 8196 34790 8206 34842
rect 8206 34790 8252 34842
rect 7956 34788 8012 34790
rect 8036 34788 8092 34790
rect 8116 34788 8172 34790
rect 8196 34788 8252 34790
rect 2956 34298 3012 34300
rect 3036 34298 3092 34300
rect 3116 34298 3172 34300
rect 3196 34298 3252 34300
rect 2956 34246 3002 34298
rect 3002 34246 3012 34298
rect 3036 34246 3066 34298
rect 3066 34246 3078 34298
rect 3078 34246 3092 34298
rect 3116 34246 3130 34298
rect 3130 34246 3142 34298
rect 3142 34246 3172 34298
rect 3196 34246 3206 34298
rect 3206 34246 3252 34298
rect 2956 34244 3012 34246
rect 3036 34244 3092 34246
rect 3116 34244 3172 34246
rect 3196 34244 3252 34246
rect 7956 33754 8012 33756
rect 8036 33754 8092 33756
rect 8116 33754 8172 33756
rect 8196 33754 8252 33756
rect 7956 33702 8002 33754
rect 8002 33702 8012 33754
rect 8036 33702 8066 33754
rect 8066 33702 8078 33754
rect 8078 33702 8092 33754
rect 8116 33702 8130 33754
rect 8130 33702 8142 33754
rect 8142 33702 8172 33754
rect 8196 33702 8206 33754
rect 8206 33702 8252 33754
rect 7956 33700 8012 33702
rect 8036 33700 8092 33702
rect 8116 33700 8172 33702
rect 8196 33700 8252 33702
rect 2956 33210 3012 33212
rect 3036 33210 3092 33212
rect 3116 33210 3172 33212
rect 3196 33210 3252 33212
rect 2956 33158 3002 33210
rect 3002 33158 3012 33210
rect 3036 33158 3066 33210
rect 3066 33158 3078 33210
rect 3078 33158 3092 33210
rect 3116 33158 3130 33210
rect 3130 33158 3142 33210
rect 3142 33158 3172 33210
rect 3196 33158 3206 33210
rect 3206 33158 3252 33210
rect 2956 33156 3012 33158
rect 3036 33156 3092 33158
rect 3116 33156 3172 33158
rect 3196 33156 3252 33158
rect 7956 32666 8012 32668
rect 8036 32666 8092 32668
rect 8116 32666 8172 32668
rect 8196 32666 8252 32668
rect 7956 32614 8002 32666
rect 8002 32614 8012 32666
rect 8036 32614 8066 32666
rect 8066 32614 8078 32666
rect 8078 32614 8092 32666
rect 8116 32614 8130 32666
rect 8130 32614 8142 32666
rect 8142 32614 8172 32666
rect 8196 32614 8206 32666
rect 8206 32614 8252 32666
rect 7956 32612 8012 32614
rect 8036 32612 8092 32614
rect 8116 32612 8172 32614
rect 8196 32612 8252 32614
rect 2956 32122 3012 32124
rect 3036 32122 3092 32124
rect 3116 32122 3172 32124
rect 3196 32122 3252 32124
rect 2956 32070 3002 32122
rect 3002 32070 3012 32122
rect 3036 32070 3066 32122
rect 3066 32070 3078 32122
rect 3078 32070 3092 32122
rect 3116 32070 3130 32122
rect 3130 32070 3142 32122
rect 3142 32070 3172 32122
rect 3196 32070 3206 32122
rect 3206 32070 3252 32122
rect 2956 32068 3012 32070
rect 3036 32068 3092 32070
rect 3116 32068 3172 32070
rect 3196 32068 3252 32070
rect 7956 31578 8012 31580
rect 8036 31578 8092 31580
rect 8116 31578 8172 31580
rect 8196 31578 8252 31580
rect 7956 31526 8002 31578
rect 8002 31526 8012 31578
rect 8036 31526 8066 31578
rect 8066 31526 8078 31578
rect 8078 31526 8092 31578
rect 8116 31526 8130 31578
rect 8130 31526 8142 31578
rect 8142 31526 8172 31578
rect 8196 31526 8206 31578
rect 8206 31526 8252 31578
rect 7956 31524 8012 31526
rect 8036 31524 8092 31526
rect 8116 31524 8172 31526
rect 8196 31524 8252 31526
rect 2956 31034 3012 31036
rect 3036 31034 3092 31036
rect 3116 31034 3172 31036
rect 3196 31034 3252 31036
rect 2956 30982 3002 31034
rect 3002 30982 3012 31034
rect 3036 30982 3066 31034
rect 3066 30982 3078 31034
rect 3078 30982 3092 31034
rect 3116 30982 3130 31034
rect 3130 30982 3142 31034
rect 3142 30982 3172 31034
rect 3196 30982 3206 31034
rect 3206 30982 3252 31034
rect 2956 30980 3012 30982
rect 3036 30980 3092 30982
rect 3116 30980 3172 30982
rect 3196 30980 3252 30982
rect 7956 30490 8012 30492
rect 8036 30490 8092 30492
rect 8116 30490 8172 30492
rect 8196 30490 8252 30492
rect 7956 30438 8002 30490
rect 8002 30438 8012 30490
rect 8036 30438 8066 30490
rect 8066 30438 8078 30490
rect 8078 30438 8092 30490
rect 8116 30438 8130 30490
rect 8130 30438 8142 30490
rect 8142 30438 8172 30490
rect 8196 30438 8206 30490
rect 8206 30438 8252 30490
rect 7956 30436 8012 30438
rect 8036 30436 8092 30438
rect 8116 30436 8172 30438
rect 8196 30436 8252 30438
rect 2956 29946 3012 29948
rect 3036 29946 3092 29948
rect 3116 29946 3172 29948
rect 3196 29946 3252 29948
rect 2956 29894 3002 29946
rect 3002 29894 3012 29946
rect 3036 29894 3066 29946
rect 3066 29894 3078 29946
rect 3078 29894 3092 29946
rect 3116 29894 3130 29946
rect 3130 29894 3142 29946
rect 3142 29894 3172 29946
rect 3196 29894 3206 29946
rect 3206 29894 3252 29946
rect 2956 29892 3012 29894
rect 3036 29892 3092 29894
rect 3116 29892 3172 29894
rect 3196 29892 3252 29894
rect 7956 29402 8012 29404
rect 8036 29402 8092 29404
rect 8116 29402 8172 29404
rect 8196 29402 8252 29404
rect 7956 29350 8002 29402
rect 8002 29350 8012 29402
rect 8036 29350 8066 29402
rect 8066 29350 8078 29402
rect 8078 29350 8092 29402
rect 8116 29350 8130 29402
rect 8130 29350 8142 29402
rect 8142 29350 8172 29402
rect 8196 29350 8206 29402
rect 8206 29350 8252 29402
rect 7956 29348 8012 29350
rect 8036 29348 8092 29350
rect 8116 29348 8172 29350
rect 8196 29348 8252 29350
rect 2956 28858 3012 28860
rect 3036 28858 3092 28860
rect 3116 28858 3172 28860
rect 3196 28858 3252 28860
rect 2956 28806 3002 28858
rect 3002 28806 3012 28858
rect 3036 28806 3066 28858
rect 3066 28806 3078 28858
rect 3078 28806 3092 28858
rect 3116 28806 3130 28858
rect 3130 28806 3142 28858
rect 3142 28806 3172 28858
rect 3196 28806 3206 28858
rect 3206 28806 3252 28858
rect 2956 28804 3012 28806
rect 3036 28804 3092 28806
rect 3116 28804 3172 28806
rect 3196 28804 3252 28806
rect 7956 28314 8012 28316
rect 8036 28314 8092 28316
rect 8116 28314 8172 28316
rect 8196 28314 8252 28316
rect 7956 28262 8002 28314
rect 8002 28262 8012 28314
rect 8036 28262 8066 28314
rect 8066 28262 8078 28314
rect 8078 28262 8092 28314
rect 8116 28262 8130 28314
rect 8130 28262 8142 28314
rect 8142 28262 8172 28314
rect 8196 28262 8206 28314
rect 8206 28262 8252 28314
rect 7956 28260 8012 28262
rect 8036 28260 8092 28262
rect 8116 28260 8172 28262
rect 8196 28260 8252 28262
rect 2956 27770 3012 27772
rect 3036 27770 3092 27772
rect 3116 27770 3172 27772
rect 3196 27770 3252 27772
rect 2956 27718 3002 27770
rect 3002 27718 3012 27770
rect 3036 27718 3066 27770
rect 3066 27718 3078 27770
rect 3078 27718 3092 27770
rect 3116 27718 3130 27770
rect 3130 27718 3142 27770
rect 3142 27718 3172 27770
rect 3196 27718 3206 27770
rect 3206 27718 3252 27770
rect 2956 27716 3012 27718
rect 3036 27716 3092 27718
rect 3116 27716 3172 27718
rect 3196 27716 3252 27718
rect 7956 27226 8012 27228
rect 8036 27226 8092 27228
rect 8116 27226 8172 27228
rect 8196 27226 8252 27228
rect 7956 27174 8002 27226
rect 8002 27174 8012 27226
rect 8036 27174 8066 27226
rect 8066 27174 8078 27226
rect 8078 27174 8092 27226
rect 8116 27174 8130 27226
rect 8130 27174 8142 27226
rect 8142 27174 8172 27226
rect 8196 27174 8206 27226
rect 8206 27174 8252 27226
rect 7956 27172 8012 27174
rect 8036 27172 8092 27174
rect 8116 27172 8172 27174
rect 8196 27172 8252 27174
rect 2956 26682 3012 26684
rect 3036 26682 3092 26684
rect 3116 26682 3172 26684
rect 3196 26682 3252 26684
rect 2956 26630 3002 26682
rect 3002 26630 3012 26682
rect 3036 26630 3066 26682
rect 3066 26630 3078 26682
rect 3078 26630 3092 26682
rect 3116 26630 3130 26682
rect 3130 26630 3142 26682
rect 3142 26630 3172 26682
rect 3196 26630 3206 26682
rect 3206 26630 3252 26682
rect 2956 26628 3012 26630
rect 3036 26628 3092 26630
rect 3116 26628 3172 26630
rect 3196 26628 3252 26630
rect 7956 26138 8012 26140
rect 8036 26138 8092 26140
rect 8116 26138 8172 26140
rect 8196 26138 8252 26140
rect 7956 26086 8002 26138
rect 8002 26086 8012 26138
rect 8036 26086 8066 26138
rect 8066 26086 8078 26138
rect 8078 26086 8092 26138
rect 8116 26086 8130 26138
rect 8130 26086 8142 26138
rect 8142 26086 8172 26138
rect 8196 26086 8206 26138
rect 8206 26086 8252 26138
rect 7956 26084 8012 26086
rect 8036 26084 8092 26086
rect 8116 26084 8172 26086
rect 8196 26084 8252 26086
rect 2956 25594 3012 25596
rect 3036 25594 3092 25596
rect 3116 25594 3172 25596
rect 3196 25594 3252 25596
rect 2956 25542 3002 25594
rect 3002 25542 3012 25594
rect 3036 25542 3066 25594
rect 3066 25542 3078 25594
rect 3078 25542 3092 25594
rect 3116 25542 3130 25594
rect 3130 25542 3142 25594
rect 3142 25542 3172 25594
rect 3196 25542 3206 25594
rect 3206 25542 3252 25594
rect 2956 25540 3012 25542
rect 3036 25540 3092 25542
rect 3116 25540 3172 25542
rect 3196 25540 3252 25542
rect 7956 25050 8012 25052
rect 8036 25050 8092 25052
rect 8116 25050 8172 25052
rect 8196 25050 8252 25052
rect 7956 24998 8002 25050
rect 8002 24998 8012 25050
rect 8036 24998 8066 25050
rect 8066 24998 8078 25050
rect 8078 24998 8092 25050
rect 8116 24998 8130 25050
rect 8130 24998 8142 25050
rect 8142 24998 8172 25050
rect 8196 24998 8206 25050
rect 8206 24998 8252 25050
rect 7956 24996 8012 24998
rect 8036 24996 8092 24998
rect 8116 24996 8172 24998
rect 8196 24996 8252 24998
rect 2956 24506 3012 24508
rect 3036 24506 3092 24508
rect 3116 24506 3172 24508
rect 3196 24506 3252 24508
rect 2956 24454 3002 24506
rect 3002 24454 3012 24506
rect 3036 24454 3066 24506
rect 3066 24454 3078 24506
rect 3078 24454 3092 24506
rect 3116 24454 3130 24506
rect 3130 24454 3142 24506
rect 3142 24454 3172 24506
rect 3196 24454 3206 24506
rect 3206 24454 3252 24506
rect 2956 24452 3012 24454
rect 3036 24452 3092 24454
rect 3116 24452 3172 24454
rect 3196 24452 3252 24454
rect 7956 23962 8012 23964
rect 8036 23962 8092 23964
rect 8116 23962 8172 23964
rect 8196 23962 8252 23964
rect 7956 23910 8002 23962
rect 8002 23910 8012 23962
rect 8036 23910 8066 23962
rect 8066 23910 8078 23962
rect 8078 23910 8092 23962
rect 8116 23910 8130 23962
rect 8130 23910 8142 23962
rect 8142 23910 8172 23962
rect 8196 23910 8206 23962
rect 8206 23910 8252 23962
rect 7956 23908 8012 23910
rect 8036 23908 8092 23910
rect 8116 23908 8172 23910
rect 8196 23908 8252 23910
rect 2956 23418 3012 23420
rect 3036 23418 3092 23420
rect 3116 23418 3172 23420
rect 3196 23418 3252 23420
rect 2956 23366 3002 23418
rect 3002 23366 3012 23418
rect 3036 23366 3066 23418
rect 3066 23366 3078 23418
rect 3078 23366 3092 23418
rect 3116 23366 3130 23418
rect 3130 23366 3142 23418
rect 3142 23366 3172 23418
rect 3196 23366 3206 23418
rect 3206 23366 3252 23418
rect 2956 23364 3012 23366
rect 3036 23364 3092 23366
rect 3116 23364 3172 23366
rect 3196 23364 3252 23366
rect 7956 22874 8012 22876
rect 8036 22874 8092 22876
rect 8116 22874 8172 22876
rect 8196 22874 8252 22876
rect 7956 22822 8002 22874
rect 8002 22822 8012 22874
rect 8036 22822 8066 22874
rect 8066 22822 8078 22874
rect 8078 22822 8092 22874
rect 8116 22822 8130 22874
rect 8130 22822 8142 22874
rect 8142 22822 8172 22874
rect 8196 22822 8206 22874
rect 8206 22822 8252 22874
rect 7956 22820 8012 22822
rect 8036 22820 8092 22822
rect 8116 22820 8172 22822
rect 8196 22820 8252 22822
rect 2956 22330 3012 22332
rect 3036 22330 3092 22332
rect 3116 22330 3172 22332
rect 3196 22330 3252 22332
rect 2956 22278 3002 22330
rect 3002 22278 3012 22330
rect 3036 22278 3066 22330
rect 3066 22278 3078 22330
rect 3078 22278 3092 22330
rect 3116 22278 3130 22330
rect 3130 22278 3142 22330
rect 3142 22278 3172 22330
rect 3196 22278 3206 22330
rect 3206 22278 3252 22330
rect 2956 22276 3012 22278
rect 3036 22276 3092 22278
rect 3116 22276 3172 22278
rect 3196 22276 3252 22278
rect 2956 21242 3012 21244
rect 3036 21242 3092 21244
rect 3116 21242 3172 21244
rect 3196 21242 3252 21244
rect 2956 21190 3002 21242
rect 3002 21190 3012 21242
rect 3036 21190 3066 21242
rect 3066 21190 3078 21242
rect 3078 21190 3092 21242
rect 3116 21190 3130 21242
rect 3130 21190 3142 21242
rect 3142 21190 3172 21242
rect 3196 21190 3206 21242
rect 3206 21190 3252 21242
rect 2956 21188 3012 21190
rect 3036 21188 3092 21190
rect 3116 21188 3172 21190
rect 3196 21188 3252 21190
rect 2956 20154 3012 20156
rect 3036 20154 3092 20156
rect 3116 20154 3172 20156
rect 3196 20154 3252 20156
rect 2956 20102 3002 20154
rect 3002 20102 3012 20154
rect 3036 20102 3066 20154
rect 3066 20102 3078 20154
rect 3078 20102 3092 20154
rect 3116 20102 3130 20154
rect 3130 20102 3142 20154
rect 3142 20102 3172 20154
rect 3196 20102 3206 20154
rect 3206 20102 3252 20154
rect 2956 20100 3012 20102
rect 3036 20100 3092 20102
rect 3116 20100 3172 20102
rect 3196 20100 3252 20102
rect 2956 19066 3012 19068
rect 3036 19066 3092 19068
rect 3116 19066 3172 19068
rect 3196 19066 3252 19068
rect 2956 19014 3002 19066
rect 3002 19014 3012 19066
rect 3036 19014 3066 19066
rect 3066 19014 3078 19066
rect 3078 19014 3092 19066
rect 3116 19014 3130 19066
rect 3130 19014 3142 19066
rect 3142 19014 3172 19066
rect 3196 19014 3206 19066
rect 3206 19014 3252 19066
rect 2956 19012 3012 19014
rect 3036 19012 3092 19014
rect 3116 19012 3172 19014
rect 3196 19012 3252 19014
rect 2956 17978 3012 17980
rect 3036 17978 3092 17980
rect 3116 17978 3172 17980
rect 3196 17978 3252 17980
rect 2956 17926 3002 17978
rect 3002 17926 3012 17978
rect 3036 17926 3066 17978
rect 3066 17926 3078 17978
rect 3078 17926 3092 17978
rect 3116 17926 3130 17978
rect 3130 17926 3142 17978
rect 3142 17926 3172 17978
rect 3196 17926 3206 17978
rect 3206 17926 3252 17978
rect 2956 17924 3012 17926
rect 3036 17924 3092 17926
rect 3116 17924 3172 17926
rect 3196 17924 3252 17926
rect 2956 16890 3012 16892
rect 3036 16890 3092 16892
rect 3116 16890 3172 16892
rect 3196 16890 3252 16892
rect 2956 16838 3002 16890
rect 3002 16838 3012 16890
rect 3036 16838 3066 16890
rect 3066 16838 3078 16890
rect 3078 16838 3092 16890
rect 3116 16838 3130 16890
rect 3130 16838 3142 16890
rect 3142 16838 3172 16890
rect 3196 16838 3206 16890
rect 3206 16838 3252 16890
rect 2956 16836 3012 16838
rect 3036 16836 3092 16838
rect 3116 16836 3172 16838
rect 3196 16836 3252 16838
rect 2956 15802 3012 15804
rect 3036 15802 3092 15804
rect 3116 15802 3172 15804
rect 3196 15802 3252 15804
rect 2956 15750 3002 15802
rect 3002 15750 3012 15802
rect 3036 15750 3066 15802
rect 3066 15750 3078 15802
rect 3078 15750 3092 15802
rect 3116 15750 3130 15802
rect 3130 15750 3142 15802
rect 3142 15750 3172 15802
rect 3196 15750 3206 15802
rect 3206 15750 3252 15802
rect 2956 15748 3012 15750
rect 3036 15748 3092 15750
rect 3116 15748 3172 15750
rect 3196 15748 3252 15750
rect 2956 14714 3012 14716
rect 3036 14714 3092 14716
rect 3116 14714 3172 14716
rect 3196 14714 3252 14716
rect 2956 14662 3002 14714
rect 3002 14662 3012 14714
rect 3036 14662 3066 14714
rect 3066 14662 3078 14714
rect 3078 14662 3092 14714
rect 3116 14662 3130 14714
rect 3130 14662 3142 14714
rect 3142 14662 3172 14714
rect 3196 14662 3206 14714
rect 3206 14662 3252 14714
rect 2956 14660 3012 14662
rect 3036 14660 3092 14662
rect 3116 14660 3172 14662
rect 3196 14660 3252 14662
rect 2956 13626 3012 13628
rect 3036 13626 3092 13628
rect 3116 13626 3172 13628
rect 3196 13626 3252 13628
rect 2956 13574 3002 13626
rect 3002 13574 3012 13626
rect 3036 13574 3066 13626
rect 3066 13574 3078 13626
rect 3078 13574 3092 13626
rect 3116 13574 3130 13626
rect 3130 13574 3142 13626
rect 3142 13574 3172 13626
rect 3196 13574 3206 13626
rect 3206 13574 3252 13626
rect 2956 13572 3012 13574
rect 3036 13572 3092 13574
rect 3116 13572 3172 13574
rect 3196 13572 3252 13574
rect 2956 12538 3012 12540
rect 3036 12538 3092 12540
rect 3116 12538 3172 12540
rect 3196 12538 3252 12540
rect 2956 12486 3002 12538
rect 3002 12486 3012 12538
rect 3036 12486 3066 12538
rect 3066 12486 3078 12538
rect 3078 12486 3092 12538
rect 3116 12486 3130 12538
rect 3130 12486 3142 12538
rect 3142 12486 3172 12538
rect 3196 12486 3206 12538
rect 3206 12486 3252 12538
rect 2956 12484 3012 12486
rect 3036 12484 3092 12486
rect 3116 12484 3172 12486
rect 3196 12484 3252 12486
rect 2956 11450 3012 11452
rect 3036 11450 3092 11452
rect 3116 11450 3172 11452
rect 3196 11450 3252 11452
rect 2956 11398 3002 11450
rect 3002 11398 3012 11450
rect 3036 11398 3066 11450
rect 3066 11398 3078 11450
rect 3078 11398 3092 11450
rect 3116 11398 3130 11450
rect 3130 11398 3142 11450
rect 3142 11398 3172 11450
rect 3196 11398 3206 11450
rect 3206 11398 3252 11450
rect 2956 11396 3012 11398
rect 3036 11396 3092 11398
rect 3116 11396 3172 11398
rect 3196 11396 3252 11398
rect 2956 10362 3012 10364
rect 3036 10362 3092 10364
rect 3116 10362 3172 10364
rect 3196 10362 3252 10364
rect 2956 10310 3002 10362
rect 3002 10310 3012 10362
rect 3036 10310 3066 10362
rect 3066 10310 3078 10362
rect 3078 10310 3092 10362
rect 3116 10310 3130 10362
rect 3130 10310 3142 10362
rect 3142 10310 3172 10362
rect 3196 10310 3206 10362
rect 3206 10310 3252 10362
rect 2956 10308 3012 10310
rect 3036 10308 3092 10310
rect 3116 10308 3172 10310
rect 3196 10308 3252 10310
rect 2956 9274 3012 9276
rect 3036 9274 3092 9276
rect 3116 9274 3172 9276
rect 3196 9274 3252 9276
rect 2956 9222 3002 9274
rect 3002 9222 3012 9274
rect 3036 9222 3066 9274
rect 3066 9222 3078 9274
rect 3078 9222 3092 9274
rect 3116 9222 3130 9274
rect 3130 9222 3142 9274
rect 3142 9222 3172 9274
rect 3196 9222 3206 9274
rect 3206 9222 3252 9274
rect 2956 9220 3012 9222
rect 3036 9220 3092 9222
rect 3116 9220 3172 9222
rect 3196 9220 3252 9222
rect 3330 8744 3386 8800
rect 2956 8186 3012 8188
rect 3036 8186 3092 8188
rect 3116 8186 3172 8188
rect 3196 8186 3252 8188
rect 2956 8134 3002 8186
rect 3002 8134 3012 8186
rect 3036 8134 3066 8186
rect 3066 8134 3078 8186
rect 3078 8134 3092 8186
rect 3116 8134 3130 8186
rect 3130 8134 3142 8186
rect 3142 8134 3172 8186
rect 3196 8134 3206 8186
rect 3206 8134 3252 8186
rect 2956 8132 3012 8134
rect 3036 8132 3092 8134
rect 3116 8132 3172 8134
rect 3196 8132 3252 8134
rect 2956 7098 3012 7100
rect 3036 7098 3092 7100
rect 3116 7098 3172 7100
rect 3196 7098 3252 7100
rect 2956 7046 3002 7098
rect 3002 7046 3012 7098
rect 3036 7046 3066 7098
rect 3066 7046 3078 7098
rect 3078 7046 3092 7098
rect 3116 7046 3130 7098
rect 3130 7046 3142 7098
rect 3142 7046 3172 7098
rect 3196 7046 3206 7098
rect 3206 7046 3252 7098
rect 2956 7044 3012 7046
rect 3036 7044 3092 7046
rect 3116 7044 3172 7046
rect 3196 7044 3252 7046
rect 2956 6010 3012 6012
rect 3036 6010 3092 6012
rect 3116 6010 3172 6012
rect 3196 6010 3252 6012
rect 2956 5958 3002 6010
rect 3002 5958 3012 6010
rect 3036 5958 3066 6010
rect 3066 5958 3078 6010
rect 3078 5958 3092 6010
rect 3116 5958 3130 6010
rect 3130 5958 3142 6010
rect 3142 5958 3172 6010
rect 3196 5958 3206 6010
rect 3206 5958 3252 6010
rect 2956 5956 3012 5958
rect 3036 5956 3092 5958
rect 3116 5956 3172 5958
rect 3196 5956 3252 5958
rect 2956 4922 3012 4924
rect 3036 4922 3092 4924
rect 3116 4922 3172 4924
rect 3196 4922 3252 4924
rect 2956 4870 3002 4922
rect 3002 4870 3012 4922
rect 3036 4870 3066 4922
rect 3066 4870 3078 4922
rect 3078 4870 3092 4922
rect 3116 4870 3130 4922
rect 3130 4870 3142 4922
rect 3142 4870 3172 4922
rect 3196 4870 3206 4922
rect 3206 4870 3252 4922
rect 2956 4868 3012 4870
rect 3036 4868 3092 4870
rect 3116 4868 3172 4870
rect 3196 4868 3252 4870
rect 2956 3834 3012 3836
rect 3036 3834 3092 3836
rect 3116 3834 3172 3836
rect 3196 3834 3252 3836
rect 2956 3782 3002 3834
rect 3002 3782 3012 3834
rect 3036 3782 3066 3834
rect 3066 3782 3078 3834
rect 3078 3782 3092 3834
rect 3116 3782 3130 3834
rect 3130 3782 3142 3834
rect 3142 3782 3172 3834
rect 3196 3782 3206 3834
rect 3206 3782 3252 3834
rect 2956 3780 3012 3782
rect 3036 3780 3092 3782
rect 3116 3780 3172 3782
rect 3196 3780 3252 3782
rect 2956 2746 3012 2748
rect 3036 2746 3092 2748
rect 3116 2746 3172 2748
rect 3196 2746 3252 2748
rect 2956 2694 3002 2746
rect 3002 2694 3012 2746
rect 3036 2694 3066 2746
rect 3066 2694 3078 2746
rect 3078 2694 3092 2746
rect 3116 2694 3130 2746
rect 3130 2694 3142 2746
rect 3142 2694 3172 2746
rect 3196 2694 3206 2746
rect 3206 2694 3252 2746
rect 2956 2692 3012 2694
rect 3036 2692 3092 2694
rect 3116 2692 3172 2694
rect 3196 2692 3252 2694
rect 3514 6432 3570 6488
rect 3974 4120 4030 4176
rect 3422 1808 3478 1864
rect 7956 21786 8012 21788
rect 8036 21786 8092 21788
rect 8116 21786 8172 21788
rect 8196 21786 8252 21788
rect 7956 21734 8002 21786
rect 8002 21734 8012 21786
rect 8036 21734 8066 21786
rect 8066 21734 8078 21786
rect 8078 21734 8092 21786
rect 8116 21734 8130 21786
rect 8130 21734 8142 21786
rect 8142 21734 8172 21786
rect 8196 21734 8206 21786
rect 8206 21734 8252 21786
rect 7956 21732 8012 21734
rect 8036 21732 8092 21734
rect 8116 21732 8172 21734
rect 8196 21732 8252 21734
rect 7956 20698 8012 20700
rect 8036 20698 8092 20700
rect 8116 20698 8172 20700
rect 8196 20698 8252 20700
rect 7956 20646 8002 20698
rect 8002 20646 8012 20698
rect 8036 20646 8066 20698
rect 8066 20646 8078 20698
rect 8078 20646 8092 20698
rect 8116 20646 8130 20698
rect 8130 20646 8142 20698
rect 8142 20646 8172 20698
rect 8196 20646 8206 20698
rect 8206 20646 8252 20698
rect 7956 20644 8012 20646
rect 8036 20644 8092 20646
rect 8116 20644 8172 20646
rect 8196 20644 8252 20646
rect 7956 19610 8012 19612
rect 8036 19610 8092 19612
rect 8116 19610 8172 19612
rect 8196 19610 8252 19612
rect 7956 19558 8002 19610
rect 8002 19558 8012 19610
rect 8036 19558 8066 19610
rect 8066 19558 8078 19610
rect 8078 19558 8092 19610
rect 8116 19558 8130 19610
rect 8130 19558 8142 19610
rect 8142 19558 8172 19610
rect 8196 19558 8206 19610
rect 8206 19558 8252 19610
rect 7956 19556 8012 19558
rect 8036 19556 8092 19558
rect 8116 19556 8172 19558
rect 8196 19556 8252 19558
rect 7956 18522 8012 18524
rect 8036 18522 8092 18524
rect 8116 18522 8172 18524
rect 8196 18522 8252 18524
rect 7956 18470 8002 18522
rect 8002 18470 8012 18522
rect 8036 18470 8066 18522
rect 8066 18470 8078 18522
rect 8078 18470 8092 18522
rect 8116 18470 8130 18522
rect 8130 18470 8142 18522
rect 8142 18470 8172 18522
rect 8196 18470 8206 18522
rect 8206 18470 8252 18522
rect 7956 18468 8012 18470
rect 8036 18468 8092 18470
rect 8116 18468 8172 18470
rect 8196 18468 8252 18470
rect 7956 17434 8012 17436
rect 8036 17434 8092 17436
rect 8116 17434 8172 17436
rect 8196 17434 8252 17436
rect 7956 17382 8002 17434
rect 8002 17382 8012 17434
rect 8036 17382 8066 17434
rect 8066 17382 8078 17434
rect 8078 17382 8092 17434
rect 8116 17382 8130 17434
rect 8130 17382 8142 17434
rect 8142 17382 8172 17434
rect 8196 17382 8206 17434
rect 8206 17382 8252 17434
rect 7956 17380 8012 17382
rect 8036 17380 8092 17382
rect 8116 17380 8172 17382
rect 8196 17380 8252 17382
rect 7956 16346 8012 16348
rect 8036 16346 8092 16348
rect 8116 16346 8172 16348
rect 8196 16346 8252 16348
rect 7956 16294 8002 16346
rect 8002 16294 8012 16346
rect 8036 16294 8066 16346
rect 8066 16294 8078 16346
rect 8078 16294 8092 16346
rect 8116 16294 8130 16346
rect 8130 16294 8142 16346
rect 8142 16294 8172 16346
rect 8196 16294 8206 16346
rect 8206 16294 8252 16346
rect 7956 16292 8012 16294
rect 8036 16292 8092 16294
rect 8116 16292 8172 16294
rect 8196 16292 8252 16294
rect 7956 15258 8012 15260
rect 8036 15258 8092 15260
rect 8116 15258 8172 15260
rect 8196 15258 8252 15260
rect 7956 15206 8002 15258
rect 8002 15206 8012 15258
rect 8036 15206 8066 15258
rect 8066 15206 8078 15258
rect 8078 15206 8092 15258
rect 8116 15206 8130 15258
rect 8130 15206 8142 15258
rect 8142 15206 8172 15258
rect 8196 15206 8206 15258
rect 8206 15206 8252 15258
rect 7956 15204 8012 15206
rect 8036 15204 8092 15206
rect 8116 15204 8172 15206
rect 8196 15204 8252 15206
rect 7956 14170 8012 14172
rect 8036 14170 8092 14172
rect 8116 14170 8172 14172
rect 8196 14170 8252 14172
rect 7956 14118 8002 14170
rect 8002 14118 8012 14170
rect 8036 14118 8066 14170
rect 8066 14118 8078 14170
rect 8078 14118 8092 14170
rect 8116 14118 8130 14170
rect 8130 14118 8142 14170
rect 8142 14118 8172 14170
rect 8196 14118 8206 14170
rect 8206 14118 8252 14170
rect 7956 14116 8012 14118
rect 8036 14116 8092 14118
rect 8116 14116 8172 14118
rect 8196 14116 8252 14118
rect 7956 13082 8012 13084
rect 8036 13082 8092 13084
rect 8116 13082 8172 13084
rect 8196 13082 8252 13084
rect 7956 13030 8002 13082
rect 8002 13030 8012 13082
rect 8036 13030 8066 13082
rect 8066 13030 8078 13082
rect 8078 13030 8092 13082
rect 8116 13030 8130 13082
rect 8130 13030 8142 13082
rect 8142 13030 8172 13082
rect 8196 13030 8206 13082
rect 8206 13030 8252 13082
rect 7956 13028 8012 13030
rect 8036 13028 8092 13030
rect 8116 13028 8172 13030
rect 8196 13028 8252 13030
rect 7102 2352 7158 2408
rect 17956 54426 18012 54428
rect 18036 54426 18092 54428
rect 18116 54426 18172 54428
rect 18196 54426 18252 54428
rect 17956 54374 18002 54426
rect 18002 54374 18012 54426
rect 18036 54374 18066 54426
rect 18066 54374 18078 54426
rect 18078 54374 18092 54426
rect 18116 54374 18130 54426
rect 18130 54374 18142 54426
rect 18142 54374 18172 54426
rect 18196 54374 18206 54426
rect 18206 54374 18252 54426
rect 17956 54372 18012 54374
rect 18036 54372 18092 54374
rect 18116 54372 18172 54374
rect 18196 54372 18252 54374
rect 12956 53882 13012 53884
rect 13036 53882 13092 53884
rect 13116 53882 13172 53884
rect 13196 53882 13252 53884
rect 12956 53830 13002 53882
rect 13002 53830 13012 53882
rect 13036 53830 13066 53882
rect 13066 53830 13078 53882
rect 13078 53830 13092 53882
rect 13116 53830 13130 53882
rect 13130 53830 13142 53882
rect 13142 53830 13172 53882
rect 13196 53830 13206 53882
rect 13206 53830 13252 53882
rect 12956 53828 13012 53830
rect 13036 53828 13092 53830
rect 13116 53828 13172 53830
rect 13196 53828 13252 53830
rect 12956 52794 13012 52796
rect 13036 52794 13092 52796
rect 13116 52794 13172 52796
rect 13196 52794 13252 52796
rect 12956 52742 13002 52794
rect 13002 52742 13012 52794
rect 13036 52742 13066 52794
rect 13066 52742 13078 52794
rect 13078 52742 13092 52794
rect 13116 52742 13130 52794
rect 13130 52742 13142 52794
rect 13142 52742 13172 52794
rect 13196 52742 13206 52794
rect 13206 52742 13252 52794
rect 12956 52740 13012 52742
rect 13036 52740 13092 52742
rect 13116 52740 13172 52742
rect 13196 52740 13252 52742
rect 12956 51706 13012 51708
rect 13036 51706 13092 51708
rect 13116 51706 13172 51708
rect 13196 51706 13252 51708
rect 12956 51654 13002 51706
rect 13002 51654 13012 51706
rect 13036 51654 13066 51706
rect 13066 51654 13078 51706
rect 13078 51654 13092 51706
rect 13116 51654 13130 51706
rect 13130 51654 13142 51706
rect 13142 51654 13172 51706
rect 13196 51654 13206 51706
rect 13206 51654 13252 51706
rect 12956 51652 13012 51654
rect 13036 51652 13092 51654
rect 13116 51652 13172 51654
rect 13196 51652 13252 51654
rect 12956 50618 13012 50620
rect 13036 50618 13092 50620
rect 13116 50618 13172 50620
rect 13196 50618 13252 50620
rect 12956 50566 13002 50618
rect 13002 50566 13012 50618
rect 13036 50566 13066 50618
rect 13066 50566 13078 50618
rect 13078 50566 13092 50618
rect 13116 50566 13130 50618
rect 13130 50566 13142 50618
rect 13142 50566 13172 50618
rect 13196 50566 13206 50618
rect 13206 50566 13252 50618
rect 12956 50564 13012 50566
rect 13036 50564 13092 50566
rect 13116 50564 13172 50566
rect 13196 50564 13252 50566
rect 12956 49530 13012 49532
rect 13036 49530 13092 49532
rect 13116 49530 13172 49532
rect 13196 49530 13252 49532
rect 12956 49478 13002 49530
rect 13002 49478 13012 49530
rect 13036 49478 13066 49530
rect 13066 49478 13078 49530
rect 13078 49478 13092 49530
rect 13116 49478 13130 49530
rect 13130 49478 13142 49530
rect 13142 49478 13172 49530
rect 13196 49478 13206 49530
rect 13206 49478 13252 49530
rect 12956 49476 13012 49478
rect 13036 49476 13092 49478
rect 13116 49476 13172 49478
rect 13196 49476 13252 49478
rect 12956 48442 13012 48444
rect 13036 48442 13092 48444
rect 13116 48442 13172 48444
rect 13196 48442 13252 48444
rect 12956 48390 13002 48442
rect 13002 48390 13012 48442
rect 13036 48390 13066 48442
rect 13066 48390 13078 48442
rect 13078 48390 13092 48442
rect 13116 48390 13130 48442
rect 13130 48390 13142 48442
rect 13142 48390 13172 48442
rect 13196 48390 13206 48442
rect 13206 48390 13252 48442
rect 12956 48388 13012 48390
rect 13036 48388 13092 48390
rect 13116 48388 13172 48390
rect 13196 48388 13252 48390
rect 12956 47354 13012 47356
rect 13036 47354 13092 47356
rect 13116 47354 13172 47356
rect 13196 47354 13252 47356
rect 12956 47302 13002 47354
rect 13002 47302 13012 47354
rect 13036 47302 13066 47354
rect 13066 47302 13078 47354
rect 13078 47302 13092 47354
rect 13116 47302 13130 47354
rect 13130 47302 13142 47354
rect 13142 47302 13172 47354
rect 13196 47302 13206 47354
rect 13206 47302 13252 47354
rect 12956 47300 13012 47302
rect 13036 47300 13092 47302
rect 13116 47300 13172 47302
rect 13196 47300 13252 47302
rect 12956 46266 13012 46268
rect 13036 46266 13092 46268
rect 13116 46266 13172 46268
rect 13196 46266 13252 46268
rect 12956 46214 13002 46266
rect 13002 46214 13012 46266
rect 13036 46214 13066 46266
rect 13066 46214 13078 46266
rect 13078 46214 13092 46266
rect 13116 46214 13130 46266
rect 13130 46214 13142 46266
rect 13142 46214 13172 46266
rect 13196 46214 13206 46266
rect 13206 46214 13252 46266
rect 12956 46212 13012 46214
rect 13036 46212 13092 46214
rect 13116 46212 13172 46214
rect 13196 46212 13252 46214
rect 12956 45178 13012 45180
rect 13036 45178 13092 45180
rect 13116 45178 13172 45180
rect 13196 45178 13252 45180
rect 12956 45126 13002 45178
rect 13002 45126 13012 45178
rect 13036 45126 13066 45178
rect 13066 45126 13078 45178
rect 13078 45126 13092 45178
rect 13116 45126 13130 45178
rect 13130 45126 13142 45178
rect 13142 45126 13172 45178
rect 13196 45126 13206 45178
rect 13206 45126 13252 45178
rect 12956 45124 13012 45126
rect 13036 45124 13092 45126
rect 13116 45124 13172 45126
rect 13196 45124 13252 45126
rect 12956 44090 13012 44092
rect 13036 44090 13092 44092
rect 13116 44090 13172 44092
rect 13196 44090 13252 44092
rect 12956 44038 13002 44090
rect 13002 44038 13012 44090
rect 13036 44038 13066 44090
rect 13066 44038 13078 44090
rect 13078 44038 13092 44090
rect 13116 44038 13130 44090
rect 13130 44038 13142 44090
rect 13142 44038 13172 44090
rect 13196 44038 13206 44090
rect 13206 44038 13252 44090
rect 12956 44036 13012 44038
rect 13036 44036 13092 44038
rect 13116 44036 13172 44038
rect 13196 44036 13252 44038
rect 12956 43002 13012 43004
rect 13036 43002 13092 43004
rect 13116 43002 13172 43004
rect 13196 43002 13252 43004
rect 12956 42950 13002 43002
rect 13002 42950 13012 43002
rect 13036 42950 13066 43002
rect 13066 42950 13078 43002
rect 13078 42950 13092 43002
rect 13116 42950 13130 43002
rect 13130 42950 13142 43002
rect 13142 42950 13172 43002
rect 13196 42950 13206 43002
rect 13206 42950 13252 43002
rect 12956 42948 13012 42950
rect 13036 42948 13092 42950
rect 13116 42948 13172 42950
rect 13196 42948 13252 42950
rect 12956 41914 13012 41916
rect 13036 41914 13092 41916
rect 13116 41914 13172 41916
rect 13196 41914 13252 41916
rect 12956 41862 13002 41914
rect 13002 41862 13012 41914
rect 13036 41862 13066 41914
rect 13066 41862 13078 41914
rect 13078 41862 13092 41914
rect 13116 41862 13130 41914
rect 13130 41862 13142 41914
rect 13142 41862 13172 41914
rect 13196 41862 13206 41914
rect 13206 41862 13252 41914
rect 12956 41860 13012 41862
rect 13036 41860 13092 41862
rect 13116 41860 13172 41862
rect 13196 41860 13252 41862
rect 12956 40826 13012 40828
rect 13036 40826 13092 40828
rect 13116 40826 13172 40828
rect 13196 40826 13252 40828
rect 12956 40774 13002 40826
rect 13002 40774 13012 40826
rect 13036 40774 13066 40826
rect 13066 40774 13078 40826
rect 13078 40774 13092 40826
rect 13116 40774 13130 40826
rect 13130 40774 13142 40826
rect 13142 40774 13172 40826
rect 13196 40774 13206 40826
rect 13206 40774 13252 40826
rect 12956 40772 13012 40774
rect 13036 40772 13092 40774
rect 13116 40772 13172 40774
rect 13196 40772 13252 40774
rect 12956 39738 13012 39740
rect 13036 39738 13092 39740
rect 13116 39738 13172 39740
rect 13196 39738 13252 39740
rect 12956 39686 13002 39738
rect 13002 39686 13012 39738
rect 13036 39686 13066 39738
rect 13066 39686 13078 39738
rect 13078 39686 13092 39738
rect 13116 39686 13130 39738
rect 13130 39686 13142 39738
rect 13142 39686 13172 39738
rect 13196 39686 13206 39738
rect 13206 39686 13252 39738
rect 12956 39684 13012 39686
rect 13036 39684 13092 39686
rect 13116 39684 13172 39686
rect 13196 39684 13252 39686
rect 12956 38650 13012 38652
rect 13036 38650 13092 38652
rect 13116 38650 13172 38652
rect 13196 38650 13252 38652
rect 12956 38598 13002 38650
rect 13002 38598 13012 38650
rect 13036 38598 13066 38650
rect 13066 38598 13078 38650
rect 13078 38598 13092 38650
rect 13116 38598 13130 38650
rect 13130 38598 13142 38650
rect 13142 38598 13172 38650
rect 13196 38598 13206 38650
rect 13206 38598 13252 38650
rect 12956 38596 13012 38598
rect 13036 38596 13092 38598
rect 13116 38596 13172 38598
rect 13196 38596 13252 38598
rect 12956 37562 13012 37564
rect 13036 37562 13092 37564
rect 13116 37562 13172 37564
rect 13196 37562 13252 37564
rect 12956 37510 13002 37562
rect 13002 37510 13012 37562
rect 13036 37510 13066 37562
rect 13066 37510 13078 37562
rect 13078 37510 13092 37562
rect 13116 37510 13130 37562
rect 13130 37510 13142 37562
rect 13142 37510 13172 37562
rect 13196 37510 13206 37562
rect 13206 37510 13252 37562
rect 12956 37508 13012 37510
rect 13036 37508 13092 37510
rect 13116 37508 13172 37510
rect 13196 37508 13252 37510
rect 12956 36474 13012 36476
rect 13036 36474 13092 36476
rect 13116 36474 13172 36476
rect 13196 36474 13252 36476
rect 12956 36422 13002 36474
rect 13002 36422 13012 36474
rect 13036 36422 13066 36474
rect 13066 36422 13078 36474
rect 13078 36422 13092 36474
rect 13116 36422 13130 36474
rect 13130 36422 13142 36474
rect 13142 36422 13172 36474
rect 13196 36422 13206 36474
rect 13206 36422 13252 36474
rect 12956 36420 13012 36422
rect 13036 36420 13092 36422
rect 13116 36420 13172 36422
rect 13196 36420 13252 36422
rect 12956 35386 13012 35388
rect 13036 35386 13092 35388
rect 13116 35386 13172 35388
rect 13196 35386 13252 35388
rect 12956 35334 13002 35386
rect 13002 35334 13012 35386
rect 13036 35334 13066 35386
rect 13066 35334 13078 35386
rect 13078 35334 13092 35386
rect 13116 35334 13130 35386
rect 13130 35334 13142 35386
rect 13142 35334 13172 35386
rect 13196 35334 13206 35386
rect 13206 35334 13252 35386
rect 12956 35332 13012 35334
rect 13036 35332 13092 35334
rect 13116 35332 13172 35334
rect 13196 35332 13252 35334
rect 12956 34298 13012 34300
rect 13036 34298 13092 34300
rect 13116 34298 13172 34300
rect 13196 34298 13252 34300
rect 12956 34246 13002 34298
rect 13002 34246 13012 34298
rect 13036 34246 13066 34298
rect 13066 34246 13078 34298
rect 13078 34246 13092 34298
rect 13116 34246 13130 34298
rect 13130 34246 13142 34298
rect 13142 34246 13172 34298
rect 13196 34246 13206 34298
rect 13206 34246 13252 34298
rect 12956 34244 13012 34246
rect 13036 34244 13092 34246
rect 13116 34244 13172 34246
rect 13196 34244 13252 34246
rect 12956 33210 13012 33212
rect 13036 33210 13092 33212
rect 13116 33210 13172 33212
rect 13196 33210 13252 33212
rect 12956 33158 13002 33210
rect 13002 33158 13012 33210
rect 13036 33158 13066 33210
rect 13066 33158 13078 33210
rect 13078 33158 13092 33210
rect 13116 33158 13130 33210
rect 13130 33158 13142 33210
rect 13142 33158 13172 33210
rect 13196 33158 13206 33210
rect 13206 33158 13252 33210
rect 12956 33156 13012 33158
rect 13036 33156 13092 33158
rect 13116 33156 13172 33158
rect 13196 33156 13252 33158
rect 12956 32122 13012 32124
rect 13036 32122 13092 32124
rect 13116 32122 13172 32124
rect 13196 32122 13252 32124
rect 12956 32070 13002 32122
rect 13002 32070 13012 32122
rect 13036 32070 13066 32122
rect 13066 32070 13078 32122
rect 13078 32070 13092 32122
rect 13116 32070 13130 32122
rect 13130 32070 13142 32122
rect 13142 32070 13172 32122
rect 13196 32070 13206 32122
rect 13206 32070 13252 32122
rect 12956 32068 13012 32070
rect 13036 32068 13092 32070
rect 13116 32068 13172 32070
rect 13196 32068 13252 32070
rect 12956 31034 13012 31036
rect 13036 31034 13092 31036
rect 13116 31034 13172 31036
rect 13196 31034 13252 31036
rect 12956 30982 13002 31034
rect 13002 30982 13012 31034
rect 13036 30982 13066 31034
rect 13066 30982 13078 31034
rect 13078 30982 13092 31034
rect 13116 30982 13130 31034
rect 13130 30982 13142 31034
rect 13142 30982 13172 31034
rect 13196 30982 13206 31034
rect 13206 30982 13252 31034
rect 12956 30980 13012 30982
rect 13036 30980 13092 30982
rect 13116 30980 13172 30982
rect 13196 30980 13252 30982
rect 12956 29946 13012 29948
rect 13036 29946 13092 29948
rect 13116 29946 13172 29948
rect 13196 29946 13252 29948
rect 12956 29894 13002 29946
rect 13002 29894 13012 29946
rect 13036 29894 13066 29946
rect 13066 29894 13078 29946
rect 13078 29894 13092 29946
rect 13116 29894 13130 29946
rect 13130 29894 13142 29946
rect 13142 29894 13172 29946
rect 13196 29894 13206 29946
rect 13206 29894 13252 29946
rect 12956 29892 13012 29894
rect 13036 29892 13092 29894
rect 13116 29892 13172 29894
rect 13196 29892 13252 29894
rect 7956 11994 8012 11996
rect 8036 11994 8092 11996
rect 8116 11994 8172 11996
rect 8196 11994 8252 11996
rect 7956 11942 8002 11994
rect 8002 11942 8012 11994
rect 8036 11942 8066 11994
rect 8066 11942 8078 11994
rect 8078 11942 8092 11994
rect 8116 11942 8130 11994
rect 8130 11942 8142 11994
rect 8142 11942 8172 11994
rect 8196 11942 8206 11994
rect 8206 11942 8252 11994
rect 7956 11940 8012 11942
rect 8036 11940 8092 11942
rect 8116 11940 8172 11942
rect 8196 11940 8252 11942
rect 7956 10906 8012 10908
rect 8036 10906 8092 10908
rect 8116 10906 8172 10908
rect 8196 10906 8252 10908
rect 7956 10854 8002 10906
rect 8002 10854 8012 10906
rect 8036 10854 8066 10906
rect 8066 10854 8078 10906
rect 8078 10854 8092 10906
rect 8116 10854 8130 10906
rect 8130 10854 8142 10906
rect 8142 10854 8172 10906
rect 8196 10854 8206 10906
rect 8206 10854 8252 10906
rect 7956 10852 8012 10854
rect 8036 10852 8092 10854
rect 8116 10852 8172 10854
rect 8196 10852 8252 10854
rect 8390 9968 8446 10024
rect 7956 9818 8012 9820
rect 8036 9818 8092 9820
rect 8116 9818 8172 9820
rect 8196 9818 8252 9820
rect 7956 9766 8002 9818
rect 8002 9766 8012 9818
rect 8036 9766 8066 9818
rect 8066 9766 8078 9818
rect 8078 9766 8092 9818
rect 8116 9766 8130 9818
rect 8130 9766 8142 9818
rect 8142 9766 8172 9818
rect 8196 9766 8206 9818
rect 8206 9766 8252 9818
rect 7956 9764 8012 9766
rect 8036 9764 8092 9766
rect 8116 9764 8172 9766
rect 8196 9764 8252 9766
rect 7956 8730 8012 8732
rect 8036 8730 8092 8732
rect 8116 8730 8172 8732
rect 8196 8730 8252 8732
rect 7956 8678 8002 8730
rect 8002 8678 8012 8730
rect 8036 8678 8066 8730
rect 8066 8678 8078 8730
rect 8078 8678 8092 8730
rect 8116 8678 8130 8730
rect 8130 8678 8142 8730
rect 8142 8678 8172 8730
rect 8196 8678 8206 8730
rect 8206 8678 8252 8730
rect 7956 8676 8012 8678
rect 8036 8676 8092 8678
rect 8116 8676 8172 8678
rect 8196 8676 8252 8678
rect 8114 8492 8170 8528
rect 8114 8472 8116 8492
rect 8116 8472 8168 8492
rect 8168 8472 8170 8492
rect 7956 7642 8012 7644
rect 8036 7642 8092 7644
rect 8116 7642 8172 7644
rect 8196 7642 8252 7644
rect 7956 7590 8002 7642
rect 8002 7590 8012 7642
rect 8036 7590 8066 7642
rect 8066 7590 8078 7642
rect 8078 7590 8092 7642
rect 8116 7590 8130 7642
rect 8130 7590 8142 7642
rect 8142 7590 8172 7642
rect 8196 7590 8206 7642
rect 8206 7590 8252 7642
rect 7956 7588 8012 7590
rect 8036 7588 8092 7590
rect 8116 7588 8172 7590
rect 8196 7588 8252 7590
rect 7956 6554 8012 6556
rect 8036 6554 8092 6556
rect 8116 6554 8172 6556
rect 8196 6554 8252 6556
rect 7956 6502 8002 6554
rect 8002 6502 8012 6554
rect 8036 6502 8066 6554
rect 8066 6502 8078 6554
rect 8078 6502 8092 6554
rect 8116 6502 8130 6554
rect 8130 6502 8142 6554
rect 8142 6502 8172 6554
rect 8196 6502 8206 6554
rect 8206 6502 8252 6554
rect 7956 6500 8012 6502
rect 8036 6500 8092 6502
rect 8116 6500 8172 6502
rect 8196 6500 8252 6502
rect 7956 5466 8012 5468
rect 8036 5466 8092 5468
rect 8116 5466 8172 5468
rect 8196 5466 8252 5468
rect 7956 5414 8002 5466
rect 8002 5414 8012 5466
rect 8036 5414 8066 5466
rect 8066 5414 8078 5466
rect 8078 5414 8092 5466
rect 8116 5414 8130 5466
rect 8130 5414 8142 5466
rect 8142 5414 8172 5466
rect 8196 5414 8206 5466
rect 8206 5414 8252 5466
rect 7956 5412 8012 5414
rect 8036 5412 8092 5414
rect 8116 5412 8172 5414
rect 8196 5412 8252 5414
rect 7956 4378 8012 4380
rect 8036 4378 8092 4380
rect 8116 4378 8172 4380
rect 8196 4378 8252 4380
rect 7956 4326 8002 4378
rect 8002 4326 8012 4378
rect 8036 4326 8066 4378
rect 8066 4326 8078 4378
rect 8078 4326 8092 4378
rect 8116 4326 8130 4378
rect 8130 4326 8142 4378
rect 8142 4326 8172 4378
rect 8196 4326 8206 4378
rect 8206 4326 8252 4378
rect 7956 4324 8012 4326
rect 8036 4324 8092 4326
rect 8116 4324 8172 4326
rect 8196 4324 8252 4326
rect 7956 3290 8012 3292
rect 8036 3290 8092 3292
rect 8116 3290 8172 3292
rect 8196 3290 8252 3292
rect 7956 3238 8002 3290
rect 8002 3238 8012 3290
rect 8036 3238 8066 3290
rect 8066 3238 8078 3290
rect 8078 3238 8092 3290
rect 8116 3238 8130 3290
rect 8130 3238 8142 3290
rect 8142 3238 8172 3290
rect 8196 3238 8206 3290
rect 8206 3238 8252 3290
rect 7956 3236 8012 3238
rect 8036 3236 8092 3238
rect 8116 3236 8172 3238
rect 8196 3236 8252 3238
rect 8206 2524 8208 2544
rect 8208 2524 8260 2544
rect 8260 2524 8262 2544
rect 8206 2488 8262 2524
rect 7956 2202 8012 2204
rect 8036 2202 8092 2204
rect 8116 2202 8172 2204
rect 8196 2202 8252 2204
rect 7956 2150 8002 2202
rect 8002 2150 8012 2202
rect 8036 2150 8066 2202
rect 8066 2150 8078 2202
rect 8078 2150 8092 2202
rect 8116 2150 8130 2202
rect 8130 2150 8142 2202
rect 8142 2150 8172 2202
rect 8196 2150 8206 2202
rect 8206 2150 8252 2202
rect 7956 2148 8012 2150
rect 8036 2148 8092 2150
rect 8116 2148 8172 2150
rect 8196 2148 8252 2150
rect 10230 15428 10286 15464
rect 10230 15408 10232 15428
rect 10232 15408 10284 15428
rect 10284 15408 10286 15428
rect 9770 4528 9826 4584
rect 9770 3068 9772 3088
rect 9772 3068 9824 3088
rect 9824 3068 9826 3088
rect 9770 3032 9826 3068
rect 12956 28858 13012 28860
rect 13036 28858 13092 28860
rect 13116 28858 13172 28860
rect 13196 28858 13252 28860
rect 12956 28806 13002 28858
rect 13002 28806 13012 28858
rect 13036 28806 13066 28858
rect 13066 28806 13078 28858
rect 13078 28806 13092 28858
rect 13116 28806 13130 28858
rect 13130 28806 13142 28858
rect 13142 28806 13172 28858
rect 13196 28806 13206 28858
rect 13206 28806 13252 28858
rect 12956 28804 13012 28806
rect 13036 28804 13092 28806
rect 13116 28804 13172 28806
rect 13196 28804 13252 28806
rect 11242 10784 11298 10840
rect 10874 10648 10930 10704
rect 12956 27770 13012 27772
rect 13036 27770 13092 27772
rect 13116 27770 13172 27772
rect 13196 27770 13252 27772
rect 12956 27718 13002 27770
rect 13002 27718 13012 27770
rect 13036 27718 13066 27770
rect 13066 27718 13078 27770
rect 13078 27718 13092 27770
rect 13116 27718 13130 27770
rect 13130 27718 13142 27770
rect 13142 27718 13172 27770
rect 13196 27718 13206 27770
rect 13206 27718 13252 27770
rect 12956 27716 13012 27718
rect 13036 27716 13092 27718
rect 13116 27716 13172 27718
rect 13196 27716 13252 27718
rect 12956 26682 13012 26684
rect 13036 26682 13092 26684
rect 13116 26682 13172 26684
rect 13196 26682 13252 26684
rect 12956 26630 13002 26682
rect 13002 26630 13012 26682
rect 13036 26630 13066 26682
rect 13066 26630 13078 26682
rect 13078 26630 13092 26682
rect 13116 26630 13130 26682
rect 13130 26630 13142 26682
rect 13142 26630 13172 26682
rect 13196 26630 13206 26682
rect 13206 26630 13252 26682
rect 12956 26628 13012 26630
rect 13036 26628 13092 26630
rect 13116 26628 13172 26630
rect 13196 26628 13252 26630
rect 17956 53338 18012 53340
rect 18036 53338 18092 53340
rect 18116 53338 18172 53340
rect 18196 53338 18252 53340
rect 17956 53286 18002 53338
rect 18002 53286 18012 53338
rect 18036 53286 18066 53338
rect 18066 53286 18078 53338
rect 18078 53286 18092 53338
rect 18116 53286 18130 53338
rect 18130 53286 18142 53338
rect 18142 53286 18172 53338
rect 18196 53286 18206 53338
rect 18206 53286 18252 53338
rect 17956 53284 18012 53286
rect 18036 53284 18092 53286
rect 18116 53284 18172 53286
rect 18196 53284 18252 53286
rect 17956 52250 18012 52252
rect 18036 52250 18092 52252
rect 18116 52250 18172 52252
rect 18196 52250 18252 52252
rect 17956 52198 18002 52250
rect 18002 52198 18012 52250
rect 18036 52198 18066 52250
rect 18066 52198 18078 52250
rect 18078 52198 18092 52250
rect 18116 52198 18130 52250
rect 18130 52198 18142 52250
rect 18142 52198 18172 52250
rect 18196 52198 18206 52250
rect 18206 52198 18252 52250
rect 17956 52196 18012 52198
rect 18036 52196 18092 52198
rect 18116 52196 18172 52198
rect 18196 52196 18252 52198
rect 17956 51162 18012 51164
rect 18036 51162 18092 51164
rect 18116 51162 18172 51164
rect 18196 51162 18252 51164
rect 17956 51110 18002 51162
rect 18002 51110 18012 51162
rect 18036 51110 18066 51162
rect 18066 51110 18078 51162
rect 18078 51110 18092 51162
rect 18116 51110 18130 51162
rect 18130 51110 18142 51162
rect 18142 51110 18172 51162
rect 18196 51110 18206 51162
rect 18206 51110 18252 51162
rect 17956 51108 18012 51110
rect 18036 51108 18092 51110
rect 18116 51108 18172 51110
rect 18196 51108 18252 51110
rect 17956 50074 18012 50076
rect 18036 50074 18092 50076
rect 18116 50074 18172 50076
rect 18196 50074 18252 50076
rect 17956 50022 18002 50074
rect 18002 50022 18012 50074
rect 18036 50022 18066 50074
rect 18066 50022 18078 50074
rect 18078 50022 18092 50074
rect 18116 50022 18130 50074
rect 18130 50022 18142 50074
rect 18142 50022 18172 50074
rect 18196 50022 18206 50074
rect 18206 50022 18252 50074
rect 17956 50020 18012 50022
rect 18036 50020 18092 50022
rect 18116 50020 18172 50022
rect 18196 50020 18252 50022
rect 17956 48986 18012 48988
rect 18036 48986 18092 48988
rect 18116 48986 18172 48988
rect 18196 48986 18252 48988
rect 17956 48934 18002 48986
rect 18002 48934 18012 48986
rect 18036 48934 18066 48986
rect 18066 48934 18078 48986
rect 18078 48934 18092 48986
rect 18116 48934 18130 48986
rect 18130 48934 18142 48986
rect 18142 48934 18172 48986
rect 18196 48934 18206 48986
rect 18206 48934 18252 48986
rect 17956 48932 18012 48934
rect 18036 48932 18092 48934
rect 18116 48932 18172 48934
rect 18196 48932 18252 48934
rect 12956 25594 13012 25596
rect 13036 25594 13092 25596
rect 13116 25594 13172 25596
rect 13196 25594 13252 25596
rect 12956 25542 13002 25594
rect 13002 25542 13012 25594
rect 13036 25542 13066 25594
rect 13066 25542 13078 25594
rect 13078 25542 13092 25594
rect 13116 25542 13130 25594
rect 13130 25542 13142 25594
rect 13142 25542 13172 25594
rect 13196 25542 13206 25594
rect 13206 25542 13252 25594
rect 12956 25540 13012 25542
rect 13036 25540 13092 25542
rect 13116 25540 13172 25542
rect 13196 25540 13252 25542
rect 12956 24506 13012 24508
rect 13036 24506 13092 24508
rect 13116 24506 13172 24508
rect 13196 24506 13252 24508
rect 12956 24454 13002 24506
rect 13002 24454 13012 24506
rect 13036 24454 13066 24506
rect 13066 24454 13078 24506
rect 13078 24454 13092 24506
rect 13116 24454 13130 24506
rect 13130 24454 13142 24506
rect 13142 24454 13172 24506
rect 13196 24454 13206 24506
rect 13206 24454 13252 24506
rect 12956 24452 13012 24454
rect 13036 24452 13092 24454
rect 13116 24452 13172 24454
rect 13196 24452 13252 24454
rect 12956 23418 13012 23420
rect 13036 23418 13092 23420
rect 13116 23418 13172 23420
rect 13196 23418 13252 23420
rect 12956 23366 13002 23418
rect 13002 23366 13012 23418
rect 13036 23366 13066 23418
rect 13066 23366 13078 23418
rect 13078 23366 13092 23418
rect 13116 23366 13130 23418
rect 13130 23366 13142 23418
rect 13142 23366 13172 23418
rect 13196 23366 13206 23418
rect 13206 23366 13252 23418
rect 12956 23364 13012 23366
rect 13036 23364 13092 23366
rect 13116 23364 13172 23366
rect 13196 23364 13252 23366
rect 12956 22330 13012 22332
rect 13036 22330 13092 22332
rect 13116 22330 13172 22332
rect 13196 22330 13252 22332
rect 12956 22278 13002 22330
rect 13002 22278 13012 22330
rect 13036 22278 13066 22330
rect 13066 22278 13078 22330
rect 13078 22278 13092 22330
rect 13116 22278 13130 22330
rect 13130 22278 13142 22330
rect 13142 22278 13172 22330
rect 13196 22278 13206 22330
rect 13206 22278 13252 22330
rect 12956 22276 13012 22278
rect 13036 22276 13092 22278
rect 13116 22276 13172 22278
rect 13196 22276 13252 22278
rect 12956 21242 13012 21244
rect 13036 21242 13092 21244
rect 13116 21242 13172 21244
rect 13196 21242 13252 21244
rect 12956 21190 13002 21242
rect 13002 21190 13012 21242
rect 13036 21190 13066 21242
rect 13066 21190 13078 21242
rect 13078 21190 13092 21242
rect 13116 21190 13130 21242
rect 13130 21190 13142 21242
rect 13142 21190 13172 21242
rect 13196 21190 13206 21242
rect 13206 21190 13252 21242
rect 12956 21188 13012 21190
rect 13036 21188 13092 21190
rect 13116 21188 13172 21190
rect 13196 21188 13252 21190
rect 12956 20154 13012 20156
rect 13036 20154 13092 20156
rect 13116 20154 13172 20156
rect 13196 20154 13252 20156
rect 12956 20102 13002 20154
rect 13002 20102 13012 20154
rect 13036 20102 13066 20154
rect 13066 20102 13078 20154
rect 13078 20102 13092 20154
rect 13116 20102 13130 20154
rect 13130 20102 13142 20154
rect 13142 20102 13172 20154
rect 13196 20102 13206 20154
rect 13206 20102 13252 20154
rect 12956 20100 13012 20102
rect 13036 20100 13092 20102
rect 13116 20100 13172 20102
rect 13196 20100 13252 20102
rect 11886 12280 11942 12336
rect 10414 6704 10470 6760
rect 10598 6160 10654 6216
rect 10598 3476 10600 3496
rect 10600 3476 10652 3496
rect 10652 3476 10654 3496
rect 10598 3440 10654 3476
rect 11518 7948 11574 7984
rect 11518 7928 11520 7948
rect 11520 7928 11572 7948
rect 11572 7928 11574 7948
rect 12070 12300 12126 12336
rect 12070 12280 12072 12300
rect 12072 12280 12124 12300
rect 12124 12280 12126 12300
rect 12956 19066 13012 19068
rect 13036 19066 13092 19068
rect 13116 19066 13172 19068
rect 13196 19066 13252 19068
rect 12956 19014 13002 19066
rect 13002 19014 13012 19066
rect 13036 19014 13066 19066
rect 13066 19014 13078 19066
rect 13078 19014 13092 19066
rect 13116 19014 13130 19066
rect 13130 19014 13142 19066
rect 13142 19014 13172 19066
rect 13196 19014 13206 19066
rect 13206 19014 13252 19066
rect 12956 19012 13012 19014
rect 13036 19012 13092 19014
rect 13116 19012 13172 19014
rect 13196 19012 13252 19014
rect 12956 17978 13012 17980
rect 13036 17978 13092 17980
rect 13116 17978 13172 17980
rect 13196 17978 13252 17980
rect 12956 17926 13002 17978
rect 13002 17926 13012 17978
rect 13036 17926 13066 17978
rect 13066 17926 13078 17978
rect 13078 17926 13092 17978
rect 13116 17926 13130 17978
rect 13130 17926 13142 17978
rect 13142 17926 13172 17978
rect 13196 17926 13206 17978
rect 13206 17926 13252 17978
rect 12956 17924 13012 17926
rect 13036 17924 13092 17926
rect 13116 17924 13172 17926
rect 13196 17924 13252 17926
rect 12956 16890 13012 16892
rect 13036 16890 13092 16892
rect 13116 16890 13172 16892
rect 13196 16890 13252 16892
rect 12956 16838 13002 16890
rect 13002 16838 13012 16890
rect 13036 16838 13066 16890
rect 13066 16838 13078 16890
rect 13078 16838 13092 16890
rect 13116 16838 13130 16890
rect 13130 16838 13142 16890
rect 13142 16838 13172 16890
rect 13196 16838 13206 16890
rect 13206 16838 13252 16890
rect 12956 16836 13012 16838
rect 13036 16836 13092 16838
rect 13116 16836 13172 16838
rect 13196 16836 13252 16838
rect 13542 16496 13598 16552
rect 12956 15802 13012 15804
rect 13036 15802 13092 15804
rect 13116 15802 13172 15804
rect 13196 15802 13252 15804
rect 12956 15750 13002 15802
rect 13002 15750 13012 15802
rect 13036 15750 13066 15802
rect 13066 15750 13078 15802
rect 13078 15750 13092 15802
rect 13116 15750 13130 15802
rect 13130 15750 13142 15802
rect 13142 15750 13172 15802
rect 13196 15750 13206 15802
rect 13206 15750 13252 15802
rect 12956 15748 13012 15750
rect 13036 15748 13092 15750
rect 13116 15748 13172 15750
rect 13196 15748 13252 15750
rect 12438 11872 12494 11928
rect 13542 14864 13598 14920
rect 12956 14714 13012 14716
rect 13036 14714 13092 14716
rect 13116 14714 13172 14716
rect 13196 14714 13252 14716
rect 12956 14662 13002 14714
rect 13002 14662 13012 14714
rect 13036 14662 13066 14714
rect 13066 14662 13078 14714
rect 13078 14662 13092 14714
rect 13116 14662 13130 14714
rect 13130 14662 13142 14714
rect 13142 14662 13172 14714
rect 13196 14662 13206 14714
rect 13206 14662 13252 14714
rect 12956 14660 13012 14662
rect 13036 14660 13092 14662
rect 13116 14660 13172 14662
rect 13196 14660 13252 14662
rect 12346 10104 12402 10160
rect 12438 9424 12494 9480
rect 11794 8336 11850 8392
rect 11886 6296 11942 6352
rect 11150 3052 11206 3088
rect 11150 3032 11152 3052
rect 11152 3032 11204 3052
rect 11204 3032 11206 3052
rect 12956 13626 13012 13628
rect 13036 13626 13092 13628
rect 13116 13626 13172 13628
rect 13196 13626 13252 13628
rect 12956 13574 13002 13626
rect 13002 13574 13012 13626
rect 13036 13574 13066 13626
rect 13066 13574 13078 13626
rect 13078 13574 13092 13626
rect 13116 13574 13130 13626
rect 13130 13574 13142 13626
rect 13142 13574 13172 13626
rect 13196 13574 13206 13626
rect 13206 13574 13252 13626
rect 12956 13572 13012 13574
rect 13036 13572 13092 13574
rect 13116 13572 13172 13574
rect 13196 13572 13252 13574
rect 12956 12538 13012 12540
rect 13036 12538 13092 12540
rect 13116 12538 13172 12540
rect 13196 12538 13252 12540
rect 12956 12486 13002 12538
rect 13002 12486 13012 12538
rect 13036 12486 13066 12538
rect 13066 12486 13078 12538
rect 13078 12486 13092 12538
rect 13116 12486 13130 12538
rect 13130 12486 13142 12538
rect 13142 12486 13172 12538
rect 13196 12486 13206 12538
rect 13206 12486 13252 12538
rect 12956 12484 13012 12486
rect 13036 12484 13092 12486
rect 13116 12484 13172 12486
rect 13196 12484 13252 12486
rect 13358 11736 13414 11792
rect 12956 11450 13012 11452
rect 13036 11450 13092 11452
rect 13116 11450 13172 11452
rect 13196 11450 13252 11452
rect 12956 11398 13002 11450
rect 13002 11398 13012 11450
rect 13036 11398 13066 11450
rect 13066 11398 13078 11450
rect 13078 11398 13092 11450
rect 13116 11398 13130 11450
rect 13130 11398 13142 11450
rect 13142 11398 13172 11450
rect 13196 11398 13206 11450
rect 13206 11398 13252 11450
rect 12956 11396 13012 11398
rect 13036 11396 13092 11398
rect 13116 11396 13172 11398
rect 13196 11396 13252 11398
rect 13726 12588 13728 12608
rect 13728 12588 13780 12608
rect 13780 12588 13782 12608
rect 13726 12552 13782 12588
rect 13542 12008 13598 12064
rect 12956 10362 13012 10364
rect 13036 10362 13092 10364
rect 13116 10362 13172 10364
rect 13196 10362 13252 10364
rect 12956 10310 13002 10362
rect 13002 10310 13012 10362
rect 13036 10310 13066 10362
rect 13066 10310 13078 10362
rect 13078 10310 13092 10362
rect 13116 10310 13130 10362
rect 13130 10310 13142 10362
rect 13142 10310 13172 10362
rect 13196 10310 13206 10362
rect 13206 10310 13252 10362
rect 12956 10308 13012 10310
rect 13036 10308 13092 10310
rect 13116 10308 13172 10310
rect 13196 10308 13252 10310
rect 12956 9274 13012 9276
rect 13036 9274 13092 9276
rect 13116 9274 13172 9276
rect 13196 9274 13252 9276
rect 12956 9222 13002 9274
rect 13002 9222 13012 9274
rect 13036 9222 13066 9274
rect 13066 9222 13078 9274
rect 13078 9222 13092 9274
rect 13116 9222 13130 9274
rect 13130 9222 13142 9274
rect 13142 9222 13172 9274
rect 13196 9222 13206 9274
rect 13206 9222 13252 9274
rect 12956 9220 13012 9222
rect 13036 9220 13092 9222
rect 13116 9220 13172 9222
rect 13196 9220 13252 9222
rect 12956 8186 13012 8188
rect 13036 8186 13092 8188
rect 13116 8186 13172 8188
rect 13196 8186 13252 8188
rect 12956 8134 13002 8186
rect 13002 8134 13012 8186
rect 13036 8134 13066 8186
rect 13066 8134 13078 8186
rect 13078 8134 13092 8186
rect 13116 8134 13130 8186
rect 13130 8134 13142 8186
rect 13142 8134 13172 8186
rect 13196 8134 13206 8186
rect 13206 8134 13252 8186
rect 12956 8132 13012 8134
rect 13036 8132 13092 8134
rect 13116 8132 13172 8134
rect 13196 8132 13252 8134
rect 13726 11872 13782 11928
rect 13726 9696 13782 9752
rect 12956 7098 13012 7100
rect 13036 7098 13092 7100
rect 13116 7098 13172 7100
rect 13196 7098 13252 7100
rect 12956 7046 13002 7098
rect 13002 7046 13012 7098
rect 13036 7046 13066 7098
rect 13066 7046 13078 7098
rect 13078 7046 13092 7098
rect 13116 7046 13130 7098
rect 13130 7046 13142 7098
rect 13142 7046 13172 7098
rect 13196 7046 13206 7098
rect 13206 7046 13252 7098
rect 12956 7044 13012 7046
rect 13036 7044 13092 7046
rect 13116 7044 13172 7046
rect 13196 7044 13252 7046
rect 12956 6010 13012 6012
rect 13036 6010 13092 6012
rect 13116 6010 13172 6012
rect 13196 6010 13252 6012
rect 12956 5958 13002 6010
rect 13002 5958 13012 6010
rect 13036 5958 13066 6010
rect 13066 5958 13078 6010
rect 13078 5958 13092 6010
rect 13116 5958 13130 6010
rect 13130 5958 13142 6010
rect 13142 5958 13172 6010
rect 13196 5958 13206 6010
rect 13206 5958 13252 6010
rect 12956 5956 13012 5958
rect 13036 5956 13092 5958
rect 13116 5956 13172 5958
rect 13196 5956 13252 5958
rect 12956 4922 13012 4924
rect 13036 4922 13092 4924
rect 13116 4922 13172 4924
rect 13196 4922 13252 4924
rect 12956 4870 13002 4922
rect 13002 4870 13012 4922
rect 13036 4870 13066 4922
rect 13066 4870 13078 4922
rect 13078 4870 13092 4922
rect 13116 4870 13130 4922
rect 13130 4870 13142 4922
rect 13142 4870 13172 4922
rect 13196 4870 13206 4922
rect 13206 4870 13252 4922
rect 12956 4868 13012 4870
rect 13036 4868 13092 4870
rect 13116 4868 13172 4870
rect 13196 4868 13252 4870
rect 12990 3984 13046 4040
rect 12956 3834 13012 3836
rect 13036 3834 13092 3836
rect 13116 3834 13172 3836
rect 13196 3834 13252 3836
rect 12956 3782 13002 3834
rect 13002 3782 13012 3834
rect 13036 3782 13066 3834
rect 13066 3782 13078 3834
rect 13078 3782 13092 3834
rect 13116 3782 13130 3834
rect 13130 3782 13142 3834
rect 13142 3782 13172 3834
rect 13196 3782 13206 3834
rect 13206 3782 13252 3834
rect 12956 3780 13012 3782
rect 13036 3780 13092 3782
rect 13116 3780 13172 3782
rect 13196 3780 13252 3782
rect 13634 7112 13690 7168
rect 15382 25100 15384 25120
rect 15384 25100 15436 25120
rect 15436 25100 15438 25120
rect 15382 25064 15438 25100
rect 16026 29008 16082 29064
rect 14094 12280 14150 12336
rect 14094 9868 14096 9888
rect 14096 9868 14148 9888
rect 14148 9868 14150 9888
rect 14094 9832 14150 9868
rect 13174 3052 13230 3088
rect 13174 3032 13176 3052
rect 13176 3032 13228 3052
rect 13228 3032 13230 3052
rect 12956 2746 13012 2748
rect 13036 2746 13092 2748
rect 13116 2746 13172 2748
rect 13196 2746 13252 2748
rect 12956 2694 13002 2746
rect 13002 2694 13012 2746
rect 13036 2694 13066 2746
rect 13066 2694 13078 2746
rect 13078 2694 13092 2746
rect 13116 2694 13130 2746
rect 13130 2694 13142 2746
rect 13142 2694 13172 2746
rect 13196 2694 13206 2746
rect 13206 2694 13252 2746
rect 12956 2692 13012 2694
rect 13036 2692 13092 2694
rect 13116 2692 13172 2694
rect 13196 2692 13252 2694
rect 14830 12144 14886 12200
rect 14646 10784 14702 10840
rect 14554 10376 14610 10432
rect 14462 10240 14518 10296
rect 14370 4684 14426 4720
rect 14370 4664 14372 4684
rect 14372 4664 14424 4684
rect 14424 4664 14426 4684
rect 16026 14220 16028 14240
rect 16028 14220 16080 14240
rect 16080 14220 16082 14240
rect 16026 14184 16082 14220
rect 15290 13096 15346 13152
rect 15658 13132 15660 13152
rect 15660 13132 15712 13152
rect 15712 13132 15714 13152
rect 14922 10512 14978 10568
rect 15658 13096 15714 13132
rect 15290 11056 15346 11112
rect 15566 10376 15622 10432
rect 15474 7540 15530 7576
rect 15474 7520 15476 7540
rect 15476 7520 15528 7540
rect 15528 7520 15530 7540
rect 14646 3576 14702 3632
rect 17956 47898 18012 47900
rect 18036 47898 18092 47900
rect 18116 47898 18172 47900
rect 18196 47898 18252 47900
rect 17956 47846 18002 47898
rect 18002 47846 18012 47898
rect 18036 47846 18066 47898
rect 18066 47846 18078 47898
rect 18078 47846 18092 47898
rect 18116 47846 18130 47898
rect 18130 47846 18142 47898
rect 18142 47846 18172 47898
rect 18196 47846 18206 47898
rect 18206 47846 18252 47898
rect 17956 47844 18012 47846
rect 18036 47844 18092 47846
rect 18116 47844 18172 47846
rect 18196 47844 18252 47846
rect 17956 46810 18012 46812
rect 18036 46810 18092 46812
rect 18116 46810 18172 46812
rect 18196 46810 18252 46812
rect 17956 46758 18002 46810
rect 18002 46758 18012 46810
rect 18036 46758 18066 46810
rect 18066 46758 18078 46810
rect 18078 46758 18092 46810
rect 18116 46758 18130 46810
rect 18130 46758 18142 46810
rect 18142 46758 18172 46810
rect 18196 46758 18206 46810
rect 18206 46758 18252 46810
rect 17956 46756 18012 46758
rect 18036 46756 18092 46758
rect 18116 46756 18172 46758
rect 18196 46756 18252 46758
rect 17956 45722 18012 45724
rect 18036 45722 18092 45724
rect 18116 45722 18172 45724
rect 18196 45722 18252 45724
rect 17956 45670 18002 45722
rect 18002 45670 18012 45722
rect 18036 45670 18066 45722
rect 18066 45670 18078 45722
rect 18078 45670 18092 45722
rect 18116 45670 18130 45722
rect 18130 45670 18142 45722
rect 18142 45670 18172 45722
rect 18196 45670 18206 45722
rect 18206 45670 18252 45722
rect 17956 45668 18012 45670
rect 18036 45668 18092 45670
rect 18116 45668 18172 45670
rect 18196 45668 18252 45670
rect 17956 44634 18012 44636
rect 18036 44634 18092 44636
rect 18116 44634 18172 44636
rect 18196 44634 18252 44636
rect 17956 44582 18002 44634
rect 18002 44582 18012 44634
rect 18036 44582 18066 44634
rect 18066 44582 18078 44634
rect 18078 44582 18092 44634
rect 18116 44582 18130 44634
rect 18130 44582 18142 44634
rect 18142 44582 18172 44634
rect 18196 44582 18206 44634
rect 18206 44582 18252 44634
rect 17956 44580 18012 44582
rect 18036 44580 18092 44582
rect 18116 44580 18172 44582
rect 18196 44580 18252 44582
rect 17956 43546 18012 43548
rect 18036 43546 18092 43548
rect 18116 43546 18172 43548
rect 18196 43546 18252 43548
rect 17956 43494 18002 43546
rect 18002 43494 18012 43546
rect 18036 43494 18066 43546
rect 18066 43494 18078 43546
rect 18078 43494 18092 43546
rect 18116 43494 18130 43546
rect 18130 43494 18142 43546
rect 18142 43494 18172 43546
rect 18196 43494 18206 43546
rect 18206 43494 18252 43546
rect 17956 43492 18012 43494
rect 18036 43492 18092 43494
rect 18116 43492 18172 43494
rect 18196 43492 18252 43494
rect 17956 42458 18012 42460
rect 18036 42458 18092 42460
rect 18116 42458 18172 42460
rect 18196 42458 18252 42460
rect 17956 42406 18002 42458
rect 18002 42406 18012 42458
rect 18036 42406 18066 42458
rect 18066 42406 18078 42458
rect 18078 42406 18092 42458
rect 18116 42406 18130 42458
rect 18130 42406 18142 42458
rect 18142 42406 18172 42458
rect 18196 42406 18206 42458
rect 18206 42406 18252 42458
rect 17956 42404 18012 42406
rect 18036 42404 18092 42406
rect 18116 42404 18172 42406
rect 18196 42404 18252 42406
rect 17956 41370 18012 41372
rect 18036 41370 18092 41372
rect 18116 41370 18172 41372
rect 18196 41370 18252 41372
rect 17956 41318 18002 41370
rect 18002 41318 18012 41370
rect 18036 41318 18066 41370
rect 18066 41318 18078 41370
rect 18078 41318 18092 41370
rect 18116 41318 18130 41370
rect 18130 41318 18142 41370
rect 18142 41318 18172 41370
rect 18196 41318 18206 41370
rect 18206 41318 18252 41370
rect 17956 41316 18012 41318
rect 18036 41316 18092 41318
rect 18116 41316 18172 41318
rect 18196 41316 18252 41318
rect 17956 40282 18012 40284
rect 18036 40282 18092 40284
rect 18116 40282 18172 40284
rect 18196 40282 18252 40284
rect 17956 40230 18002 40282
rect 18002 40230 18012 40282
rect 18036 40230 18066 40282
rect 18066 40230 18078 40282
rect 18078 40230 18092 40282
rect 18116 40230 18130 40282
rect 18130 40230 18142 40282
rect 18142 40230 18172 40282
rect 18196 40230 18206 40282
rect 18206 40230 18252 40282
rect 17956 40228 18012 40230
rect 18036 40228 18092 40230
rect 18116 40228 18172 40230
rect 18196 40228 18252 40230
rect 17956 39194 18012 39196
rect 18036 39194 18092 39196
rect 18116 39194 18172 39196
rect 18196 39194 18252 39196
rect 17956 39142 18002 39194
rect 18002 39142 18012 39194
rect 18036 39142 18066 39194
rect 18066 39142 18078 39194
rect 18078 39142 18092 39194
rect 18116 39142 18130 39194
rect 18130 39142 18142 39194
rect 18142 39142 18172 39194
rect 18196 39142 18206 39194
rect 18206 39142 18252 39194
rect 17956 39140 18012 39142
rect 18036 39140 18092 39142
rect 18116 39140 18172 39142
rect 18196 39140 18252 39142
rect 17956 38106 18012 38108
rect 18036 38106 18092 38108
rect 18116 38106 18172 38108
rect 18196 38106 18252 38108
rect 17956 38054 18002 38106
rect 18002 38054 18012 38106
rect 18036 38054 18066 38106
rect 18066 38054 18078 38106
rect 18078 38054 18092 38106
rect 18116 38054 18130 38106
rect 18130 38054 18142 38106
rect 18142 38054 18172 38106
rect 18196 38054 18206 38106
rect 18206 38054 18252 38106
rect 17956 38052 18012 38054
rect 18036 38052 18092 38054
rect 18116 38052 18172 38054
rect 18196 38052 18252 38054
rect 17956 37018 18012 37020
rect 18036 37018 18092 37020
rect 18116 37018 18172 37020
rect 18196 37018 18252 37020
rect 17956 36966 18002 37018
rect 18002 36966 18012 37018
rect 18036 36966 18066 37018
rect 18066 36966 18078 37018
rect 18078 36966 18092 37018
rect 18116 36966 18130 37018
rect 18130 36966 18142 37018
rect 18142 36966 18172 37018
rect 18196 36966 18206 37018
rect 18206 36966 18252 37018
rect 17956 36964 18012 36966
rect 18036 36964 18092 36966
rect 18116 36964 18172 36966
rect 18196 36964 18252 36966
rect 17956 35930 18012 35932
rect 18036 35930 18092 35932
rect 18116 35930 18172 35932
rect 18196 35930 18252 35932
rect 17956 35878 18002 35930
rect 18002 35878 18012 35930
rect 18036 35878 18066 35930
rect 18066 35878 18078 35930
rect 18078 35878 18092 35930
rect 18116 35878 18130 35930
rect 18130 35878 18142 35930
rect 18142 35878 18172 35930
rect 18196 35878 18206 35930
rect 18206 35878 18252 35930
rect 17956 35876 18012 35878
rect 18036 35876 18092 35878
rect 18116 35876 18172 35878
rect 18196 35876 18252 35878
rect 17956 34842 18012 34844
rect 18036 34842 18092 34844
rect 18116 34842 18172 34844
rect 18196 34842 18252 34844
rect 17956 34790 18002 34842
rect 18002 34790 18012 34842
rect 18036 34790 18066 34842
rect 18066 34790 18078 34842
rect 18078 34790 18092 34842
rect 18116 34790 18130 34842
rect 18130 34790 18142 34842
rect 18142 34790 18172 34842
rect 18196 34790 18206 34842
rect 18206 34790 18252 34842
rect 17956 34788 18012 34790
rect 18036 34788 18092 34790
rect 18116 34788 18172 34790
rect 18196 34788 18252 34790
rect 17956 33754 18012 33756
rect 18036 33754 18092 33756
rect 18116 33754 18172 33756
rect 18196 33754 18252 33756
rect 17956 33702 18002 33754
rect 18002 33702 18012 33754
rect 18036 33702 18066 33754
rect 18066 33702 18078 33754
rect 18078 33702 18092 33754
rect 18116 33702 18130 33754
rect 18130 33702 18142 33754
rect 18142 33702 18172 33754
rect 18196 33702 18206 33754
rect 18206 33702 18252 33754
rect 17956 33700 18012 33702
rect 18036 33700 18092 33702
rect 18116 33700 18172 33702
rect 18196 33700 18252 33702
rect 17956 32666 18012 32668
rect 18036 32666 18092 32668
rect 18116 32666 18172 32668
rect 18196 32666 18252 32668
rect 17956 32614 18002 32666
rect 18002 32614 18012 32666
rect 18036 32614 18066 32666
rect 18066 32614 18078 32666
rect 18078 32614 18092 32666
rect 18116 32614 18130 32666
rect 18130 32614 18142 32666
rect 18142 32614 18172 32666
rect 18196 32614 18206 32666
rect 18206 32614 18252 32666
rect 17956 32612 18012 32614
rect 18036 32612 18092 32614
rect 18116 32612 18172 32614
rect 18196 32612 18252 32614
rect 17956 31578 18012 31580
rect 18036 31578 18092 31580
rect 18116 31578 18172 31580
rect 18196 31578 18252 31580
rect 17956 31526 18002 31578
rect 18002 31526 18012 31578
rect 18036 31526 18066 31578
rect 18066 31526 18078 31578
rect 18078 31526 18092 31578
rect 18116 31526 18130 31578
rect 18130 31526 18142 31578
rect 18142 31526 18172 31578
rect 18196 31526 18206 31578
rect 18206 31526 18252 31578
rect 17956 31524 18012 31526
rect 18036 31524 18092 31526
rect 18116 31524 18172 31526
rect 18196 31524 18252 31526
rect 17498 29008 17554 29064
rect 16670 16940 16672 16960
rect 16672 16940 16724 16960
rect 16724 16940 16726 16960
rect 16670 16904 16726 16940
rect 16670 16632 16726 16688
rect 16302 13912 16358 13968
rect 15934 11736 15990 11792
rect 15934 10376 15990 10432
rect 16118 10512 16174 10568
rect 16118 9832 16174 9888
rect 15934 8336 15990 8392
rect 16302 9832 16358 9888
rect 16946 16904 17002 16960
rect 16946 12844 17002 12880
rect 16946 12824 16948 12844
rect 16948 12824 17000 12844
rect 17000 12824 17002 12844
rect 16578 12008 16634 12064
rect 16486 11192 16542 11248
rect 16394 8200 16450 8256
rect 17956 30490 18012 30492
rect 18036 30490 18092 30492
rect 18116 30490 18172 30492
rect 18196 30490 18252 30492
rect 17956 30438 18002 30490
rect 18002 30438 18012 30490
rect 18036 30438 18066 30490
rect 18066 30438 18078 30490
rect 18078 30438 18092 30490
rect 18116 30438 18130 30490
rect 18130 30438 18142 30490
rect 18142 30438 18172 30490
rect 18196 30438 18206 30490
rect 18206 30438 18252 30490
rect 17956 30436 18012 30438
rect 18036 30436 18092 30438
rect 18116 30436 18172 30438
rect 18196 30436 18252 30438
rect 17956 29402 18012 29404
rect 18036 29402 18092 29404
rect 18116 29402 18172 29404
rect 18196 29402 18252 29404
rect 17956 29350 18002 29402
rect 18002 29350 18012 29402
rect 18036 29350 18066 29402
rect 18066 29350 18078 29402
rect 18078 29350 18092 29402
rect 18116 29350 18130 29402
rect 18130 29350 18142 29402
rect 18142 29350 18172 29402
rect 18196 29350 18206 29402
rect 18206 29350 18252 29402
rect 17956 29348 18012 29350
rect 18036 29348 18092 29350
rect 18116 29348 18172 29350
rect 18196 29348 18252 29350
rect 17956 28314 18012 28316
rect 18036 28314 18092 28316
rect 18116 28314 18172 28316
rect 18196 28314 18252 28316
rect 17956 28262 18002 28314
rect 18002 28262 18012 28314
rect 18036 28262 18066 28314
rect 18066 28262 18078 28314
rect 18078 28262 18092 28314
rect 18116 28262 18130 28314
rect 18130 28262 18142 28314
rect 18142 28262 18172 28314
rect 18196 28262 18206 28314
rect 18206 28262 18252 28314
rect 17956 28260 18012 28262
rect 18036 28260 18092 28262
rect 18116 28260 18172 28262
rect 18196 28260 18252 28262
rect 17682 27276 17684 27296
rect 17684 27276 17736 27296
rect 17736 27276 17738 27296
rect 17682 27240 17738 27276
rect 17956 27226 18012 27228
rect 18036 27226 18092 27228
rect 18116 27226 18172 27228
rect 18196 27226 18252 27228
rect 17956 27174 18002 27226
rect 18002 27174 18012 27226
rect 18036 27174 18066 27226
rect 18066 27174 18078 27226
rect 18078 27174 18092 27226
rect 18116 27174 18130 27226
rect 18130 27174 18142 27226
rect 18142 27174 18172 27226
rect 18196 27174 18206 27226
rect 18206 27174 18252 27226
rect 17956 27172 18012 27174
rect 18036 27172 18092 27174
rect 18116 27172 18172 27174
rect 18196 27172 18252 27174
rect 17958 26324 17960 26344
rect 17960 26324 18012 26344
rect 18012 26324 18014 26344
rect 17958 26288 18014 26324
rect 17956 26138 18012 26140
rect 18036 26138 18092 26140
rect 18116 26138 18172 26140
rect 18196 26138 18252 26140
rect 17956 26086 18002 26138
rect 18002 26086 18012 26138
rect 18036 26086 18066 26138
rect 18066 26086 18078 26138
rect 18078 26086 18092 26138
rect 18116 26086 18130 26138
rect 18130 26086 18142 26138
rect 18142 26086 18172 26138
rect 18196 26086 18206 26138
rect 18206 26086 18252 26138
rect 17956 26084 18012 26086
rect 18036 26084 18092 26086
rect 18116 26084 18172 26086
rect 18196 26084 18252 26086
rect 17956 25050 18012 25052
rect 18036 25050 18092 25052
rect 18116 25050 18172 25052
rect 18196 25050 18252 25052
rect 17956 24998 18002 25050
rect 18002 24998 18012 25050
rect 18036 24998 18066 25050
rect 18066 24998 18078 25050
rect 18078 24998 18092 25050
rect 18116 24998 18130 25050
rect 18130 24998 18142 25050
rect 18142 24998 18172 25050
rect 18196 24998 18206 25050
rect 18206 24998 18252 25050
rect 17956 24996 18012 24998
rect 18036 24996 18092 24998
rect 18116 24996 18172 24998
rect 18196 24996 18252 24998
rect 17590 23704 17646 23760
rect 17222 16224 17278 16280
rect 17314 15272 17370 15328
rect 16854 11464 16910 11520
rect 16946 10376 17002 10432
rect 16946 9596 16948 9616
rect 16948 9596 17000 9616
rect 17000 9596 17002 9616
rect 16946 9560 17002 9596
rect 16854 8916 16856 8936
rect 16856 8916 16908 8936
rect 16908 8916 16910 8936
rect 16854 8880 16910 8916
rect 16118 2488 16174 2544
rect 16302 3712 16358 3768
rect 16578 7112 16634 7168
rect 16486 4700 16488 4720
rect 16488 4700 16540 4720
rect 16540 4700 16542 4720
rect 16486 4664 16542 4700
rect 17956 23962 18012 23964
rect 18036 23962 18092 23964
rect 18116 23962 18172 23964
rect 18196 23962 18252 23964
rect 17956 23910 18002 23962
rect 18002 23910 18012 23962
rect 18036 23910 18066 23962
rect 18066 23910 18078 23962
rect 18078 23910 18092 23962
rect 18116 23910 18130 23962
rect 18130 23910 18142 23962
rect 18142 23910 18172 23962
rect 18196 23910 18206 23962
rect 18206 23910 18252 23962
rect 17956 23908 18012 23910
rect 18036 23908 18092 23910
rect 18116 23908 18172 23910
rect 18196 23908 18252 23910
rect 17956 22874 18012 22876
rect 18036 22874 18092 22876
rect 18116 22874 18172 22876
rect 18196 22874 18252 22876
rect 17956 22822 18002 22874
rect 18002 22822 18012 22874
rect 18036 22822 18066 22874
rect 18066 22822 18078 22874
rect 18078 22822 18092 22874
rect 18116 22822 18130 22874
rect 18130 22822 18142 22874
rect 18142 22822 18172 22874
rect 18196 22822 18206 22874
rect 18206 22822 18252 22874
rect 17956 22820 18012 22822
rect 18036 22820 18092 22822
rect 18116 22820 18172 22822
rect 18196 22820 18252 22822
rect 17956 21786 18012 21788
rect 18036 21786 18092 21788
rect 18116 21786 18172 21788
rect 18196 21786 18252 21788
rect 17956 21734 18002 21786
rect 18002 21734 18012 21786
rect 18036 21734 18066 21786
rect 18066 21734 18078 21786
rect 18078 21734 18092 21786
rect 18116 21734 18130 21786
rect 18130 21734 18142 21786
rect 18142 21734 18172 21786
rect 18196 21734 18206 21786
rect 18206 21734 18252 21786
rect 17956 21732 18012 21734
rect 18036 21732 18092 21734
rect 18116 21732 18172 21734
rect 18196 21732 18252 21734
rect 17956 20698 18012 20700
rect 18036 20698 18092 20700
rect 18116 20698 18172 20700
rect 18196 20698 18252 20700
rect 17956 20646 18002 20698
rect 18002 20646 18012 20698
rect 18036 20646 18066 20698
rect 18066 20646 18078 20698
rect 18078 20646 18092 20698
rect 18116 20646 18130 20698
rect 18130 20646 18142 20698
rect 18142 20646 18172 20698
rect 18196 20646 18206 20698
rect 18206 20646 18252 20698
rect 17956 20644 18012 20646
rect 18036 20644 18092 20646
rect 18116 20644 18172 20646
rect 18196 20644 18252 20646
rect 17956 19610 18012 19612
rect 18036 19610 18092 19612
rect 18116 19610 18172 19612
rect 18196 19610 18252 19612
rect 17956 19558 18002 19610
rect 18002 19558 18012 19610
rect 18036 19558 18066 19610
rect 18066 19558 18078 19610
rect 18078 19558 18092 19610
rect 18116 19558 18130 19610
rect 18130 19558 18142 19610
rect 18142 19558 18172 19610
rect 18196 19558 18206 19610
rect 18206 19558 18252 19610
rect 17956 19556 18012 19558
rect 18036 19556 18092 19558
rect 18116 19556 18172 19558
rect 18196 19556 18252 19558
rect 17956 18522 18012 18524
rect 18036 18522 18092 18524
rect 18116 18522 18172 18524
rect 18196 18522 18252 18524
rect 17956 18470 18002 18522
rect 18002 18470 18012 18522
rect 18036 18470 18066 18522
rect 18066 18470 18078 18522
rect 18078 18470 18092 18522
rect 18116 18470 18130 18522
rect 18130 18470 18142 18522
rect 18142 18470 18172 18522
rect 18196 18470 18206 18522
rect 18206 18470 18252 18522
rect 17956 18468 18012 18470
rect 18036 18468 18092 18470
rect 18116 18468 18172 18470
rect 18196 18468 18252 18470
rect 18418 18264 18474 18320
rect 17866 17756 17868 17776
rect 17868 17756 17920 17776
rect 17920 17756 17922 17776
rect 17866 17720 17922 17756
rect 17956 17434 18012 17436
rect 18036 17434 18092 17436
rect 18116 17434 18172 17436
rect 18196 17434 18252 17436
rect 17956 17382 18002 17434
rect 18002 17382 18012 17434
rect 18036 17382 18066 17434
rect 18066 17382 18078 17434
rect 18078 17382 18092 17434
rect 18116 17382 18130 17434
rect 18130 17382 18142 17434
rect 18142 17382 18172 17434
rect 18196 17382 18206 17434
rect 18206 17382 18252 17434
rect 17956 17380 18012 17382
rect 18036 17380 18092 17382
rect 18116 17380 18172 17382
rect 18196 17380 18252 17382
rect 17956 16346 18012 16348
rect 18036 16346 18092 16348
rect 18116 16346 18172 16348
rect 18196 16346 18252 16348
rect 17956 16294 18002 16346
rect 18002 16294 18012 16346
rect 18036 16294 18066 16346
rect 18066 16294 18078 16346
rect 18078 16294 18092 16346
rect 18116 16294 18130 16346
rect 18130 16294 18142 16346
rect 18142 16294 18172 16346
rect 18196 16294 18206 16346
rect 18206 16294 18252 16346
rect 17956 16292 18012 16294
rect 18036 16292 18092 16294
rect 18116 16292 18172 16294
rect 18196 16292 18252 16294
rect 17222 11464 17278 11520
rect 17406 11192 17462 11248
rect 17956 15258 18012 15260
rect 18036 15258 18092 15260
rect 18116 15258 18172 15260
rect 18196 15258 18252 15260
rect 17956 15206 18002 15258
rect 18002 15206 18012 15258
rect 18036 15206 18066 15258
rect 18066 15206 18078 15258
rect 18078 15206 18092 15258
rect 18116 15206 18130 15258
rect 18130 15206 18142 15258
rect 18142 15206 18172 15258
rect 18196 15206 18206 15258
rect 18206 15206 18252 15258
rect 17956 15204 18012 15206
rect 18036 15204 18092 15206
rect 18116 15204 18172 15206
rect 18196 15204 18252 15206
rect 18970 26288 19026 26344
rect 18602 18128 18658 18184
rect 17956 14170 18012 14172
rect 18036 14170 18092 14172
rect 18116 14170 18172 14172
rect 18196 14170 18252 14172
rect 17956 14118 18002 14170
rect 18002 14118 18012 14170
rect 18036 14118 18066 14170
rect 18066 14118 18078 14170
rect 18078 14118 18092 14170
rect 18116 14118 18130 14170
rect 18130 14118 18142 14170
rect 18142 14118 18172 14170
rect 18196 14118 18206 14170
rect 18206 14118 18252 14170
rect 17956 14116 18012 14118
rect 18036 14116 18092 14118
rect 18116 14116 18172 14118
rect 18196 14116 18252 14118
rect 18786 17740 18842 17776
rect 18786 17720 18788 17740
rect 18788 17720 18840 17740
rect 18840 17720 18842 17740
rect 17956 13082 18012 13084
rect 18036 13082 18092 13084
rect 18116 13082 18172 13084
rect 18196 13082 18252 13084
rect 17956 13030 18002 13082
rect 18002 13030 18012 13082
rect 18036 13030 18066 13082
rect 18066 13030 18078 13082
rect 18078 13030 18092 13082
rect 18116 13030 18130 13082
rect 18130 13030 18142 13082
rect 18142 13030 18172 13082
rect 18196 13030 18206 13082
rect 18206 13030 18252 13082
rect 17956 13028 18012 13030
rect 18036 13028 18092 13030
rect 18116 13028 18172 13030
rect 18196 13028 18252 13030
rect 17682 12416 17738 12472
rect 17682 12144 17738 12200
rect 18418 12280 18474 12336
rect 19338 25100 19340 25120
rect 19340 25100 19392 25120
rect 19392 25100 19394 25120
rect 19338 25064 19394 25100
rect 19062 19352 19118 19408
rect 18786 12416 18842 12472
rect 18694 12144 18750 12200
rect 17956 11994 18012 11996
rect 18036 11994 18092 11996
rect 18116 11994 18172 11996
rect 18196 11994 18252 11996
rect 17956 11942 18002 11994
rect 18002 11942 18012 11994
rect 18036 11942 18066 11994
rect 18066 11942 18078 11994
rect 18078 11942 18092 11994
rect 18116 11942 18130 11994
rect 18130 11942 18142 11994
rect 18142 11942 18172 11994
rect 18196 11942 18206 11994
rect 18206 11942 18252 11994
rect 17956 11940 18012 11942
rect 18036 11940 18092 11942
rect 18116 11940 18172 11942
rect 18196 11940 18252 11942
rect 18510 11736 18566 11792
rect 18510 11636 18512 11656
rect 18512 11636 18564 11656
rect 18564 11636 18566 11656
rect 18510 11600 18566 11636
rect 18326 11348 18382 11384
rect 18326 11328 18328 11348
rect 18328 11328 18380 11348
rect 18380 11328 18382 11348
rect 17774 10784 17830 10840
rect 17774 10376 17830 10432
rect 17590 9696 17646 9752
rect 17590 8880 17646 8936
rect 17130 4936 17186 4992
rect 17406 4528 17462 4584
rect 17956 10906 18012 10908
rect 18036 10906 18092 10908
rect 18116 10906 18172 10908
rect 18196 10906 18252 10908
rect 17956 10854 18002 10906
rect 18002 10854 18012 10906
rect 18036 10854 18066 10906
rect 18066 10854 18078 10906
rect 18078 10854 18092 10906
rect 18116 10854 18130 10906
rect 18130 10854 18142 10906
rect 18142 10854 18172 10906
rect 18196 10854 18206 10906
rect 18206 10854 18252 10906
rect 17956 10852 18012 10854
rect 18036 10852 18092 10854
rect 18116 10852 18172 10854
rect 18196 10852 18252 10854
rect 17956 9818 18012 9820
rect 18036 9818 18092 9820
rect 18116 9818 18172 9820
rect 18196 9818 18252 9820
rect 17956 9766 18002 9818
rect 18002 9766 18012 9818
rect 18036 9766 18066 9818
rect 18066 9766 18078 9818
rect 18078 9766 18092 9818
rect 18116 9766 18130 9818
rect 18130 9766 18142 9818
rect 18142 9766 18172 9818
rect 18196 9766 18206 9818
rect 18206 9766 18252 9818
rect 17956 9764 18012 9766
rect 18036 9764 18092 9766
rect 18116 9764 18172 9766
rect 18196 9764 18252 9766
rect 17956 8730 18012 8732
rect 18036 8730 18092 8732
rect 18116 8730 18172 8732
rect 18196 8730 18252 8732
rect 17956 8678 18002 8730
rect 18002 8678 18012 8730
rect 18036 8678 18066 8730
rect 18066 8678 18078 8730
rect 18078 8678 18092 8730
rect 18116 8678 18130 8730
rect 18130 8678 18142 8730
rect 18142 8678 18172 8730
rect 18196 8678 18206 8730
rect 18206 8678 18252 8730
rect 17956 8676 18012 8678
rect 18036 8676 18092 8678
rect 18116 8676 18172 8678
rect 18196 8676 18252 8678
rect 17956 7642 18012 7644
rect 18036 7642 18092 7644
rect 18116 7642 18172 7644
rect 18196 7642 18252 7644
rect 17956 7590 18002 7642
rect 18002 7590 18012 7642
rect 18036 7590 18066 7642
rect 18066 7590 18078 7642
rect 18078 7590 18092 7642
rect 18116 7590 18130 7642
rect 18130 7590 18142 7642
rect 18142 7590 18172 7642
rect 18196 7590 18206 7642
rect 18206 7590 18252 7642
rect 17956 7588 18012 7590
rect 18036 7588 18092 7590
rect 18116 7588 18172 7590
rect 18196 7588 18252 7590
rect 17956 6554 18012 6556
rect 18036 6554 18092 6556
rect 18116 6554 18172 6556
rect 18196 6554 18252 6556
rect 17956 6502 18002 6554
rect 18002 6502 18012 6554
rect 18036 6502 18066 6554
rect 18066 6502 18078 6554
rect 18078 6502 18092 6554
rect 18116 6502 18130 6554
rect 18130 6502 18142 6554
rect 18142 6502 18172 6554
rect 18196 6502 18206 6554
rect 18206 6502 18252 6554
rect 17956 6500 18012 6502
rect 18036 6500 18092 6502
rect 18116 6500 18172 6502
rect 18196 6500 18252 6502
rect 17956 5466 18012 5468
rect 18036 5466 18092 5468
rect 18116 5466 18172 5468
rect 18196 5466 18252 5468
rect 17956 5414 18002 5466
rect 18002 5414 18012 5466
rect 18036 5414 18066 5466
rect 18066 5414 18078 5466
rect 18078 5414 18092 5466
rect 18116 5414 18130 5466
rect 18130 5414 18142 5466
rect 18142 5414 18172 5466
rect 18196 5414 18206 5466
rect 18206 5414 18252 5466
rect 17956 5412 18012 5414
rect 18036 5412 18092 5414
rect 18116 5412 18172 5414
rect 18196 5412 18252 5414
rect 17956 4378 18012 4380
rect 18036 4378 18092 4380
rect 18116 4378 18172 4380
rect 18196 4378 18252 4380
rect 17956 4326 18002 4378
rect 18002 4326 18012 4378
rect 18036 4326 18066 4378
rect 18066 4326 18078 4378
rect 18078 4326 18092 4378
rect 18116 4326 18130 4378
rect 18130 4326 18142 4378
rect 18142 4326 18172 4378
rect 18196 4326 18206 4378
rect 18206 4326 18252 4378
rect 17956 4324 18012 4326
rect 18036 4324 18092 4326
rect 18116 4324 18172 4326
rect 18196 4324 18252 4326
rect 18694 11464 18750 11520
rect 18694 10412 18696 10432
rect 18696 10412 18748 10432
rect 18748 10412 18750 10432
rect 18694 10376 18750 10412
rect 19246 17040 19302 17096
rect 23386 56072 23442 56128
rect 22956 53882 23012 53884
rect 23036 53882 23092 53884
rect 23116 53882 23172 53884
rect 23196 53882 23252 53884
rect 22956 53830 23002 53882
rect 23002 53830 23012 53882
rect 23036 53830 23066 53882
rect 23066 53830 23078 53882
rect 23078 53830 23092 53882
rect 23116 53830 23130 53882
rect 23130 53830 23142 53882
rect 23142 53830 23172 53882
rect 23196 53830 23206 53882
rect 23206 53830 23252 53882
rect 22956 53828 23012 53830
rect 23036 53828 23092 53830
rect 23116 53828 23172 53830
rect 23196 53828 23252 53830
rect 22956 52794 23012 52796
rect 23036 52794 23092 52796
rect 23116 52794 23172 52796
rect 23196 52794 23252 52796
rect 22956 52742 23002 52794
rect 23002 52742 23012 52794
rect 23036 52742 23066 52794
rect 23066 52742 23078 52794
rect 23078 52742 23092 52794
rect 23116 52742 23130 52794
rect 23130 52742 23142 52794
rect 23142 52742 23172 52794
rect 23196 52742 23206 52794
rect 23206 52742 23252 52794
rect 22956 52740 23012 52742
rect 23036 52740 23092 52742
rect 23116 52740 23172 52742
rect 23196 52740 23252 52742
rect 22956 51706 23012 51708
rect 23036 51706 23092 51708
rect 23116 51706 23172 51708
rect 23196 51706 23252 51708
rect 22956 51654 23002 51706
rect 23002 51654 23012 51706
rect 23036 51654 23066 51706
rect 23066 51654 23078 51706
rect 23078 51654 23092 51706
rect 23116 51654 23130 51706
rect 23130 51654 23142 51706
rect 23142 51654 23172 51706
rect 23196 51654 23206 51706
rect 23206 51654 23252 51706
rect 22956 51652 23012 51654
rect 23036 51652 23092 51654
rect 23116 51652 23172 51654
rect 23196 51652 23252 51654
rect 22956 50618 23012 50620
rect 23036 50618 23092 50620
rect 23116 50618 23172 50620
rect 23196 50618 23252 50620
rect 22956 50566 23002 50618
rect 23002 50566 23012 50618
rect 23036 50566 23066 50618
rect 23066 50566 23078 50618
rect 23078 50566 23092 50618
rect 23116 50566 23130 50618
rect 23130 50566 23142 50618
rect 23142 50566 23172 50618
rect 23196 50566 23206 50618
rect 23206 50566 23252 50618
rect 22956 50564 23012 50566
rect 23036 50564 23092 50566
rect 23116 50564 23172 50566
rect 23196 50564 23252 50566
rect 22956 49530 23012 49532
rect 23036 49530 23092 49532
rect 23116 49530 23172 49532
rect 23196 49530 23252 49532
rect 22956 49478 23002 49530
rect 23002 49478 23012 49530
rect 23036 49478 23066 49530
rect 23066 49478 23078 49530
rect 23078 49478 23092 49530
rect 23116 49478 23130 49530
rect 23130 49478 23142 49530
rect 23142 49478 23172 49530
rect 23196 49478 23206 49530
rect 23206 49478 23252 49530
rect 22956 49476 23012 49478
rect 23036 49476 23092 49478
rect 23116 49476 23172 49478
rect 23196 49476 23252 49478
rect 22956 48442 23012 48444
rect 23036 48442 23092 48444
rect 23116 48442 23172 48444
rect 23196 48442 23252 48444
rect 22956 48390 23002 48442
rect 23002 48390 23012 48442
rect 23036 48390 23066 48442
rect 23066 48390 23078 48442
rect 23078 48390 23092 48442
rect 23116 48390 23130 48442
rect 23130 48390 23142 48442
rect 23142 48390 23172 48442
rect 23196 48390 23206 48442
rect 23206 48390 23252 48442
rect 22956 48388 23012 48390
rect 23036 48388 23092 48390
rect 23116 48388 23172 48390
rect 23196 48388 23252 48390
rect 22956 47354 23012 47356
rect 23036 47354 23092 47356
rect 23116 47354 23172 47356
rect 23196 47354 23252 47356
rect 22956 47302 23002 47354
rect 23002 47302 23012 47354
rect 23036 47302 23066 47354
rect 23066 47302 23078 47354
rect 23078 47302 23092 47354
rect 23116 47302 23130 47354
rect 23130 47302 23142 47354
rect 23142 47302 23172 47354
rect 23196 47302 23206 47354
rect 23206 47302 23252 47354
rect 22956 47300 23012 47302
rect 23036 47300 23092 47302
rect 23116 47300 23172 47302
rect 23196 47300 23252 47302
rect 22956 46266 23012 46268
rect 23036 46266 23092 46268
rect 23116 46266 23172 46268
rect 23196 46266 23252 46268
rect 22956 46214 23002 46266
rect 23002 46214 23012 46266
rect 23036 46214 23066 46266
rect 23066 46214 23078 46266
rect 23078 46214 23092 46266
rect 23116 46214 23130 46266
rect 23130 46214 23142 46266
rect 23142 46214 23172 46266
rect 23196 46214 23206 46266
rect 23206 46214 23252 46266
rect 22956 46212 23012 46214
rect 23036 46212 23092 46214
rect 23116 46212 23172 46214
rect 23196 46212 23252 46214
rect 22956 45178 23012 45180
rect 23036 45178 23092 45180
rect 23116 45178 23172 45180
rect 23196 45178 23252 45180
rect 22956 45126 23002 45178
rect 23002 45126 23012 45178
rect 23036 45126 23066 45178
rect 23066 45126 23078 45178
rect 23078 45126 23092 45178
rect 23116 45126 23130 45178
rect 23130 45126 23142 45178
rect 23142 45126 23172 45178
rect 23196 45126 23206 45178
rect 23206 45126 23252 45178
rect 22956 45124 23012 45126
rect 23036 45124 23092 45126
rect 23116 45124 23172 45126
rect 23196 45124 23252 45126
rect 22956 44090 23012 44092
rect 23036 44090 23092 44092
rect 23116 44090 23172 44092
rect 23196 44090 23252 44092
rect 22956 44038 23002 44090
rect 23002 44038 23012 44090
rect 23036 44038 23066 44090
rect 23066 44038 23078 44090
rect 23078 44038 23092 44090
rect 23116 44038 23130 44090
rect 23130 44038 23142 44090
rect 23142 44038 23172 44090
rect 23196 44038 23206 44090
rect 23206 44038 23252 44090
rect 22956 44036 23012 44038
rect 23036 44036 23092 44038
rect 23116 44036 23172 44038
rect 23196 44036 23252 44038
rect 22956 43002 23012 43004
rect 23036 43002 23092 43004
rect 23116 43002 23172 43004
rect 23196 43002 23252 43004
rect 22956 42950 23002 43002
rect 23002 42950 23012 43002
rect 23036 42950 23066 43002
rect 23066 42950 23078 43002
rect 23078 42950 23092 43002
rect 23116 42950 23130 43002
rect 23130 42950 23142 43002
rect 23142 42950 23172 43002
rect 23196 42950 23206 43002
rect 23206 42950 23252 43002
rect 22956 42948 23012 42950
rect 23036 42948 23092 42950
rect 23116 42948 23172 42950
rect 23196 42948 23252 42950
rect 22956 41914 23012 41916
rect 23036 41914 23092 41916
rect 23116 41914 23172 41916
rect 23196 41914 23252 41916
rect 22956 41862 23002 41914
rect 23002 41862 23012 41914
rect 23036 41862 23066 41914
rect 23066 41862 23078 41914
rect 23078 41862 23092 41914
rect 23116 41862 23130 41914
rect 23130 41862 23142 41914
rect 23142 41862 23172 41914
rect 23196 41862 23206 41914
rect 23206 41862 23252 41914
rect 22956 41860 23012 41862
rect 23036 41860 23092 41862
rect 23116 41860 23172 41862
rect 23196 41860 23252 41862
rect 22956 40826 23012 40828
rect 23036 40826 23092 40828
rect 23116 40826 23172 40828
rect 23196 40826 23252 40828
rect 22956 40774 23002 40826
rect 23002 40774 23012 40826
rect 23036 40774 23066 40826
rect 23066 40774 23078 40826
rect 23078 40774 23092 40826
rect 23116 40774 23130 40826
rect 23130 40774 23142 40826
rect 23142 40774 23172 40826
rect 23196 40774 23206 40826
rect 23206 40774 23252 40826
rect 22956 40772 23012 40774
rect 23036 40772 23092 40774
rect 23116 40772 23172 40774
rect 23196 40772 23252 40774
rect 22956 39738 23012 39740
rect 23036 39738 23092 39740
rect 23116 39738 23172 39740
rect 23196 39738 23252 39740
rect 22956 39686 23002 39738
rect 23002 39686 23012 39738
rect 23036 39686 23066 39738
rect 23066 39686 23078 39738
rect 23078 39686 23092 39738
rect 23116 39686 23130 39738
rect 23130 39686 23142 39738
rect 23142 39686 23172 39738
rect 23196 39686 23206 39738
rect 23206 39686 23252 39738
rect 22956 39684 23012 39686
rect 23036 39684 23092 39686
rect 23116 39684 23172 39686
rect 23196 39684 23252 39686
rect 22956 38650 23012 38652
rect 23036 38650 23092 38652
rect 23116 38650 23172 38652
rect 23196 38650 23252 38652
rect 22956 38598 23002 38650
rect 23002 38598 23012 38650
rect 23036 38598 23066 38650
rect 23066 38598 23078 38650
rect 23078 38598 23092 38650
rect 23116 38598 23130 38650
rect 23130 38598 23142 38650
rect 23142 38598 23172 38650
rect 23196 38598 23206 38650
rect 23206 38598 23252 38650
rect 22956 38596 23012 38598
rect 23036 38596 23092 38598
rect 23116 38596 23172 38598
rect 23196 38596 23252 38598
rect 22956 37562 23012 37564
rect 23036 37562 23092 37564
rect 23116 37562 23172 37564
rect 23196 37562 23252 37564
rect 22956 37510 23002 37562
rect 23002 37510 23012 37562
rect 23036 37510 23066 37562
rect 23066 37510 23078 37562
rect 23078 37510 23092 37562
rect 23116 37510 23130 37562
rect 23130 37510 23142 37562
rect 23142 37510 23172 37562
rect 23196 37510 23206 37562
rect 23206 37510 23252 37562
rect 22956 37508 23012 37510
rect 23036 37508 23092 37510
rect 23116 37508 23172 37510
rect 23196 37508 23252 37510
rect 22956 36474 23012 36476
rect 23036 36474 23092 36476
rect 23116 36474 23172 36476
rect 23196 36474 23252 36476
rect 22956 36422 23002 36474
rect 23002 36422 23012 36474
rect 23036 36422 23066 36474
rect 23066 36422 23078 36474
rect 23078 36422 23092 36474
rect 23116 36422 23130 36474
rect 23130 36422 23142 36474
rect 23142 36422 23172 36474
rect 23196 36422 23206 36474
rect 23206 36422 23252 36474
rect 22956 36420 23012 36422
rect 23036 36420 23092 36422
rect 23116 36420 23172 36422
rect 23196 36420 23252 36422
rect 24490 55392 24546 55448
rect 24674 54576 24730 54632
rect 24766 53760 24822 53816
rect 24766 43968 24822 44024
rect 20994 24928 21050 24984
rect 22098 27920 22154 27976
rect 22956 35386 23012 35388
rect 23036 35386 23092 35388
rect 23116 35386 23172 35388
rect 23196 35386 23252 35388
rect 22956 35334 23002 35386
rect 23002 35334 23012 35386
rect 23036 35334 23066 35386
rect 23066 35334 23078 35386
rect 23078 35334 23092 35386
rect 23116 35334 23130 35386
rect 23130 35334 23142 35386
rect 23142 35334 23172 35386
rect 23196 35334 23206 35386
rect 23206 35334 23252 35386
rect 22956 35332 23012 35334
rect 23036 35332 23092 35334
rect 23116 35332 23172 35334
rect 23196 35332 23252 35334
rect 22956 34298 23012 34300
rect 23036 34298 23092 34300
rect 23116 34298 23172 34300
rect 23196 34298 23252 34300
rect 22956 34246 23002 34298
rect 23002 34246 23012 34298
rect 23036 34246 23066 34298
rect 23066 34246 23078 34298
rect 23078 34246 23092 34298
rect 23116 34246 23130 34298
rect 23130 34246 23142 34298
rect 23142 34246 23172 34298
rect 23196 34246 23206 34298
rect 23206 34246 23252 34298
rect 22956 34244 23012 34246
rect 23036 34244 23092 34246
rect 23116 34244 23172 34246
rect 23196 34244 23252 34246
rect 22956 33210 23012 33212
rect 23036 33210 23092 33212
rect 23116 33210 23172 33212
rect 23196 33210 23252 33212
rect 22956 33158 23002 33210
rect 23002 33158 23012 33210
rect 23036 33158 23066 33210
rect 23066 33158 23078 33210
rect 23078 33158 23092 33210
rect 23116 33158 23130 33210
rect 23130 33158 23142 33210
rect 23142 33158 23172 33210
rect 23196 33158 23206 33210
rect 23206 33158 23252 33210
rect 22956 33156 23012 33158
rect 23036 33156 23092 33158
rect 23116 33156 23172 33158
rect 23196 33156 23252 33158
rect 22956 32122 23012 32124
rect 23036 32122 23092 32124
rect 23116 32122 23172 32124
rect 23196 32122 23252 32124
rect 22956 32070 23002 32122
rect 23002 32070 23012 32122
rect 23036 32070 23066 32122
rect 23066 32070 23078 32122
rect 23078 32070 23092 32122
rect 23116 32070 23130 32122
rect 23130 32070 23142 32122
rect 23142 32070 23172 32122
rect 23196 32070 23206 32122
rect 23206 32070 23252 32122
rect 22956 32068 23012 32070
rect 23036 32068 23092 32070
rect 23116 32068 23172 32070
rect 23196 32068 23252 32070
rect 22956 31034 23012 31036
rect 23036 31034 23092 31036
rect 23116 31034 23172 31036
rect 23196 31034 23252 31036
rect 22956 30982 23002 31034
rect 23002 30982 23012 31034
rect 23036 30982 23066 31034
rect 23066 30982 23078 31034
rect 23078 30982 23092 31034
rect 23116 30982 23130 31034
rect 23130 30982 23142 31034
rect 23142 30982 23172 31034
rect 23196 30982 23206 31034
rect 23206 30982 23252 31034
rect 22956 30980 23012 30982
rect 23036 30980 23092 30982
rect 23116 30980 23172 30982
rect 23196 30980 23252 30982
rect 22956 29946 23012 29948
rect 23036 29946 23092 29948
rect 23116 29946 23172 29948
rect 23196 29946 23252 29948
rect 22956 29894 23002 29946
rect 23002 29894 23012 29946
rect 23036 29894 23066 29946
rect 23066 29894 23078 29946
rect 23078 29894 23092 29946
rect 23116 29894 23130 29946
rect 23130 29894 23142 29946
rect 23142 29894 23172 29946
rect 23196 29894 23206 29946
rect 23206 29894 23252 29946
rect 22956 29892 23012 29894
rect 23036 29892 23092 29894
rect 23116 29892 23172 29894
rect 23196 29892 23252 29894
rect 21822 26832 21878 26888
rect 19430 16632 19486 16688
rect 19154 11328 19210 11384
rect 18786 8372 18788 8392
rect 18788 8372 18840 8392
rect 18840 8372 18842 8392
rect 18786 8336 18842 8372
rect 19062 10920 19118 10976
rect 18970 8880 19026 8936
rect 17590 2896 17646 2952
rect 17956 3290 18012 3292
rect 18036 3290 18092 3292
rect 18116 3290 18172 3292
rect 18196 3290 18252 3292
rect 17956 3238 18002 3290
rect 18002 3238 18012 3290
rect 18036 3238 18066 3290
rect 18066 3238 18078 3290
rect 18078 3238 18092 3290
rect 18116 3238 18130 3290
rect 18130 3238 18142 3290
rect 18142 3238 18172 3290
rect 18196 3238 18206 3290
rect 18206 3238 18252 3290
rect 17956 3236 18012 3238
rect 18036 3236 18092 3238
rect 18116 3236 18172 3238
rect 18196 3236 18252 3238
rect 17956 2202 18012 2204
rect 18036 2202 18092 2204
rect 18116 2202 18172 2204
rect 18196 2202 18252 2204
rect 17956 2150 18002 2202
rect 18002 2150 18012 2202
rect 18036 2150 18066 2202
rect 18066 2150 18078 2202
rect 18078 2150 18092 2202
rect 18116 2150 18130 2202
rect 18130 2150 18142 2202
rect 18142 2150 18172 2202
rect 18196 2150 18206 2202
rect 18206 2150 18252 2202
rect 17956 2148 18012 2150
rect 18036 2148 18092 2150
rect 18116 2148 18172 2150
rect 18196 2148 18252 2150
rect 19522 13252 19578 13288
rect 19522 13232 19524 13252
rect 19524 13232 19576 13252
rect 19576 13232 19578 13252
rect 19982 14864 20038 14920
rect 20074 12588 20076 12608
rect 20076 12588 20128 12608
rect 20128 12588 20130 12608
rect 20074 12552 20130 12588
rect 20442 14048 20498 14104
rect 20350 12688 20406 12744
rect 20166 9460 20168 9480
rect 20168 9460 20220 9480
rect 20220 9460 20222 9480
rect 20166 9424 20222 9460
rect 19614 8336 19670 8392
rect 19522 4936 19578 4992
rect 21086 23432 21142 23488
rect 22190 25744 22246 25800
rect 21178 17332 21234 17368
rect 21178 17312 21180 17332
rect 21180 17312 21232 17332
rect 21232 17312 21234 17332
rect 21362 18028 21364 18048
rect 21364 18028 21416 18048
rect 21416 18028 21418 18048
rect 21362 17992 21418 18028
rect 20902 12980 20958 13016
rect 20902 12960 20904 12980
rect 20904 12960 20956 12980
rect 20956 12960 20958 12980
rect 20626 9868 20628 9888
rect 20628 9868 20680 9888
rect 20680 9868 20682 9888
rect 20626 9832 20682 9868
rect 20810 11056 20866 11112
rect 20718 8472 20774 8528
rect 20350 3576 20406 3632
rect 21178 10920 21234 10976
rect 21362 5480 21418 5536
rect 23110 29144 23166 29200
rect 22558 29008 22614 29064
rect 22956 28858 23012 28860
rect 23036 28858 23092 28860
rect 23116 28858 23172 28860
rect 23196 28858 23252 28860
rect 22956 28806 23002 28858
rect 23002 28806 23012 28858
rect 23036 28806 23066 28858
rect 23066 28806 23078 28858
rect 23078 28806 23092 28858
rect 23116 28806 23130 28858
rect 23130 28806 23142 28858
rect 23142 28806 23172 28858
rect 23196 28806 23206 28858
rect 23206 28806 23252 28858
rect 22956 28804 23012 28806
rect 23036 28804 23092 28806
rect 23116 28804 23172 28806
rect 23196 28804 23252 28806
rect 22466 26016 22522 26072
rect 23202 28464 23258 28520
rect 22956 27770 23012 27772
rect 23036 27770 23092 27772
rect 23116 27770 23172 27772
rect 23196 27770 23252 27772
rect 22956 27718 23002 27770
rect 23002 27718 23012 27770
rect 23036 27718 23066 27770
rect 23066 27718 23078 27770
rect 23078 27718 23092 27770
rect 23116 27718 23130 27770
rect 23130 27718 23142 27770
rect 23142 27718 23172 27770
rect 23196 27718 23206 27770
rect 23206 27718 23252 27770
rect 22956 27716 23012 27718
rect 23036 27716 23092 27718
rect 23116 27716 23172 27718
rect 23196 27716 23252 27718
rect 22956 26682 23012 26684
rect 23036 26682 23092 26684
rect 23116 26682 23172 26684
rect 23196 26682 23252 26684
rect 22956 26630 23002 26682
rect 23002 26630 23012 26682
rect 23036 26630 23066 26682
rect 23066 26630 23078 26682
rect 23078 26630 23092 26682
rect 23116 26630 23130 26682
rect 23130 26630 23142 26682
rect 23142 26630 23172 26682
rect 23196 26630 23206 26682
rect 23206 26630 23252 26682
rect 22956 26628 23012 26630
rect 23036 26628 23092 26630
rect 23116 26628 23172 26630
rect 23196 26628 23252 26630
rect 22956 25594 23012 25596
rect 23036 25594 23092 25596
rect 23116 25594 23172 25596
rect 23196 25594 23252 25596
rect 22956 25542 23002 25594
rect 23002 25542 23012 25594
rect 23036 25542 23066 25594
rect 23066 25542 23078 25594
rect 23078 25542 23092 25594
rect 23116 25542 23130 25594
rect 23130 25542 23142 25594
rect 23142 25542 23172 25594
rect 23196 25542 23206 25594
rect 23206 25542 23252 25594
rect 22956 25540 23012 25542
rect 23036 25540 23092 25542
rect 23116 25540 23172 25542
rect 23196 25540 23252 25542
rect 22956 24506 23012 24508
rect 23036 24506 23092 24508
rect 23116 24506 23172 24508
rect 23196 24506 23252 24508
rect 22956 24454 23002 24506
rect 23002 24454 23012 24506
rect 23036 24454 23066 24506
rect 23066 24454 23078 24506
rect 23078 24454 23092 24506
rect 23116 24454 23130 24506
rect 23130 24454 23142 24506
rect 23142 24454 23172 24506
rect 23196 24454 23206 24506
rect 23206 24454 23252 24506
rect 22956 24452 23012 24454
rect 23036 24452 23092 24454
rect 23116 24452 23172 24454
rect 23196 24452 23252 24454
rect 24674 35128 24730 35184
rect 24766 34176 24822 34232
rect 24674 33360 24730 33416
rect 24582 32544 24638 32600
rect 24490 31728 24546 31784
rect 25042 52944 25098 53000
rect 24950 52128 25006 52184
rect 25502 51348 25504 51368
rect 25504 51348 25556 51368
rect 25556 51348 25558 51368
rect 25502 51312 25558 51348
rect 24950 50496 25006 50552
rect 25502 49680 25558 49736
rect 25134 48864 25190 48920
rect 25134 48084 25136 48104
rect 25136 48084 25188 48104
rect 25188 48084 25190 48104
rect 25134 48048 25190 48084
rect 25318 47232 25374 47288
rect 25318 46416 25374 46472
rect 25318 45600 25374 45656
rect 25318 44820 25320 44840
rect 25320 44820 25372 44840
rect 25372 44820 25374 44840
rect 25318 44784 25374 44820
rect 25502 43152 25558 43208
rect 25134 42336 25190 42392
rect 25134 41556 25136 41576
rect 25136 41556 25188 41576
rect 25188 41556 25190 41576
rect 25134 41520 25190 41556
rect 24858 29280 24914 29336
rect 25134 37440 25190 37496
rect 25134 36624 25190 36680
rect 22956 23418 23012 23420
rect 23036 23418 23092 23420
rect 23116 23418 23172 23420
rect 23196 23418 23252 23420
rect 22956 23366 23002 23418
rect 23002 23366 23012 23418
rect 23036 23366 23066 23418
rect 23066 23366 23078 23418
rect 23078 23366 23092 23418
rect 23116 23366 23130 23418
rect 23130 23366 23142 23418
rect 23142 23366 23172 23418
rect 23196 23366 23206 23418
rect 23206 23366 23252 23418
rect 22956 23364 23012 23366
rect 23036 23364 23092 23366
rect 23116 23364 23172 23366
rect 23196 23364 23252 23366
rect 22956 22330 23012 22332
rect 23036 22330 23092 22332
rect 23116 22330 23172 22332
rect 23196 22330 23252 22332
rect 22956 22278 23002 22330
rect 23002 22278 23012 22330
rect 23036 22278 23066 22330
rect 23066 22278 23078 22330
rect 23078 22278 23092 22330
rect 23116 22278 23130 22330
rect 23130 22278 23142 22330
rect 23142 22278 23172 22330
rect 23196 22278 23206 22330
rect 23206 22278 23252 22330
rect 22956 22276 23012 22278
rect 23036 22276 23092 22278
rect 23116 22276 23172 22278
rect 23196 22276 23252 22278
rect 23754 23568 23810 23624
rect 22650 19624 22706 19680
rect 22466 19216 22522 19272
rect 22098 17040 22154 17096
rect 21822 14864 21878 14920
rect 22956 21242 23012 21244
rect 23036 21242 23092 21244
rect 23116 21242 23172 21244
rect 23196 21242 23252 21244
rect 22956 21190 23002 21242
rect 23002 21190 23012 21242
rect 23036 21190 23066 21242
rect 23066 21190 23078 21242
rect 23078 21190 23092 21242
rect 23116 21190 23130 21242
rect 23130 21190 23142 21242
rect 23142 21190 23172 21242
rect 23196 21190 23206 21242
rect 23206 21190 23252 21242
rect 22956 21188 23012 21190
rect 23036 21188 23092 21190
rect 23116 21188 23172 21190
rect 23196 21188 23252 21190
rect 23386 21120 23442 21176
rect 23202 20340 23204 20360
rect 23204 20340 23256 20360
rect 23256 20340 23258 20360
rect 23202 20304 23258 20340
rect 22956 20154 23012 20156
rect 23036 20154 23092 20156
rect 23116 20154 23172 20156
rect 23196 20154 23252 20156
rect 22956 20102 23002 20154
rect 23002 20102 23012 20154
rect 23036 20102 23066 20154
rect 23066 20102 23078 20154
rect 23078 20102 23092 20154
rect 23116 20102 23130 20154
rect 23130 20102 23142 20154
rect 23142 20102 23172 20154
rect 23196 20102 23206 20154
rect 23206 20102 23252 20154
rect 22956 20100 23012 20102
rect 23036 20100 23092 20102
rect 23116 20100 23172 20102
rect 23196 20100 23252 20102
rect 23386 19488 23442 19544
rect 22006 10104 22062 10160
rect 22956 19066 23012 19068
rect 23036 19066 23092 19068
rect 23116 19066 23172 19068
rect 23196 19066 23252 19068
rect 22956 19014 23002 19066
rect 23002 19014 23012 19066
rect 23036 19014 23066 19066
rect 23066 19014 23078 19066
rect 23078 19014 23092 19066
rect 23116 19014 23130 19066
rect 23130 19014 23142 19066
rect 23142 19014 23172 19066
rect 23196 19014 23206 19066
rect 23206 19014 23252 19066
rect 22956 19012 23012 19014
rect 23036 19012 23092 19014
rect 23116 19012 23172 19014
rect 23196 19012 23252 19014
rect 22956 17978 23012 17980
rect 23036 17978 23092 17980
rect 23116 17978 23172 17980
rect 23196 17978 23252 17980
rect 22956 17926 23002 17978
rect 23002 17926 23012 17978
rect 23036 17926 23066 17978
rect 23066 17926 23078 17978
rect 23078 17926 23092 17978
rect 23116 17926 23130 17978
rect 23130 17926 23142 17978
rect 23142 17926 23172 17978
rect 23196 17926 23206 17978
rect 23206 17926 23252 17978
rect 22956 17924 23012 17926
rect 23036 17924 23092 17926
rect 23116 17924 23172 17926
rect 23196 17924 23252 17926
rect 22956 16890 23012 16892
rect 23036 16890 23092 16892
rect 23116 16890 23172 16892
rect 23196 16890 23252 16892
rect 22956 16838 23002 16890
rect 23002 16838 23012 16890
rect 23036 16838 23066 16890
rect 23066 16838 23078 16890
rect 23078 16838 23092 16890
rect 23116 16838 23130 16890
rect 23130 16838 23142 16890
rect 23142 16838 23172 16890
rect 23196 16838 23206 16890
rect 23206 16838 23252 16890
rect 22956 16836 23012 16838
rect 23036 16836 23092 16838
rect 23116 16836 23172 16838
rect 23196 16836 23252 16838
rect 25318 40704 25374 40760
rect 25410 39888 25466 39944
rect 25318 39072 25374 39128
rect 25318 38292 25320 38312
rect 25320 38292 25372 38312
rect 25372 38292 25374 38312
rect 25318 38256 25374 38292
rect 25318 35808 25374 35864
rect 25318 30912 25374 30968
rect 25410 30096 25466 30152
rect 24950 25220 25006 25256
rect 24950 25200 24952 25220
rect 24952 25200 25004 25220
rect 25004 25200 25006 25220
rect 24766 24384 24822 24440
rect 24858 22752 24914 22808
rect 24858 21936 24914 21992
rect 24766 18672 24822 18728
rect 22956 15802 23012 15804
rect 23036 15802 23092 15804
rect 23116 15802 23172 15804
rect 23196 15802 23252 15804
rect 22956 15750 23002 15802
rect 23002 15750 23012 15802
rect 23036 15750 23066 15802
rect 23066 15750 23078 15802
rect 23078 15750 23092 15802
rect 23116 15750 23130 15802
rect 23130 15750 23142 15802
rect 23142 15750 23172 15802
rect 23196 15750 23206 15802
rect 23206 15750 23252 15802
rect 22956 15748 23012 15750
rect 23036 15748 23092 15750
rect 23116 15748 23172 15750
rect 23196 15748 23252 15750
rect 22956 14714 23012 14716
rect 23036 14714 23092 14716
rect 23116 14714 23172 14716
rect 23196 14714 23252 14716
rect 22956 14662 23002 14714
rect 23002 14662 23012 14714
rect 23036 14662 23066 14714
rect 23066 14662 23078 14714
rect 23078 14662 23092 14714
rect 23116 14662 23130 14714
rect 23130 14662 23142 14714
rect 23142 14662 23172 14714
rect 23196 14662 23206 14714
rect 23206 14662 23252 14714
rect 22956 14660 23012 14662
rect 23036 14660 23092 14662
rect 23116 14660 23172 14662
rect 23196 14660 23252 14662
rect 24858 17856 24914 17912
rect 24858 17040 24914 17096
rect 24950 16224 25006 16280
rect 24766 15408 24822 15464
rect 25134 14592 25190 14648
rect 22956 13626 23012 13628
rect 23036 13626 23092 13628
rect 23116 13626 23172 13628
rect 23196 13626 23252 13628
rect 22956 13574 23002 13626
rect 23002 13574 23012 13626
rect 23036 13574 23066 13626
rect 23066 13574 23078 13626
rect 23078 13574 23092 13626
rect 23116 13574 23130 13626
rect 23130 13574 23142 13626
rect 23142 13574 23172 13626
rect 23196 13574 23206 13626
rect 23206 13574 23252 13626
rect 22956 13572 23012 13574
rect 23036 13572 23092 13574
rect 23116 13572 23172 13574
rect 23196 13572 23252 13574
rect 22956 12538 23012 12540
rect 23036 12538 23092 12540
rect 23116 12538 23172 12540
rect 23196 12538 23252 12540
rect 22956 12486 23002 12538
rect 23002 12486 23012 12538
rect 23036 12486 23066 12538
rect 23066 12486 23078 12538
rect 23078 12486 23092 12538
rect 23116 12486 23130 12538
rect 23130 12486 23142 12538
rect 23142 12486 23172 12538
rect 23196 12486 23206 12538
rect 23206 12486 23252 12538
rect 22956 12484 23012 12486
rect 23036 12484 23092 12486
rect 23116 12484 23172 12486
rect 23196 12484 23252 12486
rect 24858 13776 24914 13832
rect 24950 12960 25006 13016
rect 22956 11450 23012 11452
rect 23036 11450 23092 11452
rect 23116 11450 23172 11452
rect 23196 11450 23252 11452
rect 22956 11398 23002 11450
rect 23002 11398 23012 11450
rect 23036 11398 23066 11450
rect 23066 11398 23078 11450
rect 23078 11398 23092 11450
rect 23116 11398 23130 11450
rect 23130 11398 23142 11450
rect 23142 11398 23172 11450
rect 23196 11398 23206 11450
rect 23206 11398 23252 11450
rect 22956 11396 23012 11398
rect 23036 11396 23092 11398
rect 23116 11396 23172 11398
rect 23196 11396 23252 11398
rect 22956 10362 23012 10364
rect 23036 10362 23092 10364
rect 23116 10362 23172 10364
rect 23196 10362 23252 10364
rect 22956 10310 23002 10362
rect 23002 10310 23012 10362
rect 23036 10310 23066 10362
rect 23066 10310 23078 10362
rect 23078 10310 23092 10362
rect 23116 10310 23130 10362
rect 23130 10310 23142 10362
rect 23142 10310 23172 10362
rect 23196 10310 23206 10362
rect 23206 10310 23252 10362
rect 22956 10308 23012 10310
rect 23036 10308 23092 10310
rect 23116 10308 23172 10310
rect 23196 10308 23252 10310
rect 23018 9968 23074 10024
rect 23294 9696 23350 9752
rect 22956 9274 23012 9276
rect 23036 9274 23092 9276
rect 23116 9274 23172 9276
rect 23196 9274 23252 9276
rect 22956 9222 23002 9274
rect 23002 9222 23012 9274
rect 23036 9222 23066 9274
rect 23066 9222 23078 9274
rect 23078 9222 23092 9274
rect 23116 9222 23130 9274
rect 23130 9222 23142 9274
rect 23142 9222 23172 9274
rect 23196 9222 23206 9274
rect 23206 9222 23252 9274
rect 22956 9220 23012 9222
rect 23036 9220 23092 9222
rect 23116 9220 23172 9222
rect 23196 9220 23252 9222
rect 21914 5072 21970 5128
rect 22098 3984 22154 4040
rect 22466 6296 22522 6352
rect 22374 6160 22430 6216
rect 22374 4256 22430 4312
rect 22098 2372 22154 2408
rect 22098 2352 22100 2372
rect 22100 2352 22152 2372
rect 22152 2352 22154 2372
rect 21822 1536 21878 1592
rect 22956 8186 23012 8188
rect 23036 8186 23092 8188
rect 23116 8186 23172 8188
rect 23196 8186 23252 8188
rect 22956 8134 23002 8186
rect 23002 8134 23012 8186
rect 23036 8134 23066 8186
rect 23066 8134 23078 8186
rect 23078 8134 23092 8186
rect 23116 8134 23130 8186
rect 23130 8134 23142 8186
rect 23142 8134 23172 8186
rect 23196 8134 23206 8186
rect 23206 8134 23252 8186
rect 22956 8132 23012 8134
rect 23036 8132 23092 8134
rect 23116 8132 23172 8134
rect 23196 8132 23252 8134
rect 22956 7098 23012 7100
rect 23036 7098 23092 7100
rect 23116 7098 23172 7100
rect 23196 7098 23252 7100
rect 22956 7046 23002 7098
rect 23002 7046 23012 7098
rect 23036 7046 23066 7098
rect 23066 7046 23078 7098
rect 23078 7046 23092 7098
rect 23116 7046 23130 7098
rect 23130 7046 23142 7098
rect 23142 7046 23172 7098
rect 23196 7046 23206 7098
rect 23206 7046 23252 7098
rect 22956 7044 23012 7046
rect 23036 7044 23092 7046
rect 23116 7044 23172 7046
rect 23196 7044 23252 7046
rect 22956 6010 23012 6012
rect 23036 6010 23092 6012
rect 23116 6010 23172 6012
rect 23196 6010 23252 6012
rect 22956 5958 23002 6010
rect 23002 5958 23012 6010
rect 23036 5958 23066 6010
rect 23066 5958 23078 6010
rect 23078 5958 23092 6010
rect 23116 5958 23130 6010
rect 23130 5958 23142 6010
rect 23142 5958 23172 6010
rect 23196 5958 23206 6010
rect 23206 5958 23252 6010
rect 22956 5956 23012 5958
rect 23036 5956 23092 5958
rect 23116 5956 23172 5958
rect 23196 5956 23252 5958
rect 23386 6976 23442 7032
rect 23294 5616 23350 5672
rect 23386 5480 23442 5536
rect 22956 4922 23012 4924
rect 23036 4922 23092 4924
rect 23116 4922 23172 4924
rect 23196 4922 23252 4924
rect 22956 4870 23002 4922
rect 23002 4870 23012 4922
rect 23036 4870 23066 4922
rect 23066 4870 23078 4922
rect 23078 4870 23092 4922
rect 23116 4870 23130 4922
rect 23130 4870 23142 4922
rect 23142 4870 23172 4922
rect 23196 4870 23206 4922
rect 23206 4870 23252 4922
rect 22956 4868 23012 4870
rect 23036 4868 23092 4870
rect 23116 4868 23172 4870
rect 23196 4868 23252 4870
rect 22956 3834 23012 3836
rect 23036 3834 23092 3836
rect 23116 3834 23172 3836
rect 23196 3834 23252 3836
rect 22956 3782 23002 3834
rect 23002 3782 23012 3834
rect 23036 3782 23066 3834
rect 23066 3782 23078 3834
rect 23078 3782 23092 3834
rect 23116 3782 23130 3834
rect 23130 3782 23142 3834
rect 23142 3782 23172 3834
rect 23196 3782 23206 3834
rect 23206 3782 23252 3834
rect 22956 3780 23012 3782
rect 23036 3780 23092 3782
rect 23116 3780 23172 3782
rect 23196 3780 23252 3782
rect 22742 3732 22798 3768
rect 22742 3712 22744 3732
rect 22744 3712 22796 3732
rect 22796 3712 22798 3732
rect 22926 3576 22982 3632
rect 23202 3168 23258 3224
rect 22956 2746 23012 2748
rect 23036 2746 23092 2748
rect 23116 2746 23172 2748
rect 23196 2746 23252 2748
rect 22956 2694 23002 2746
rect 23002 2694 23012 2746
rect 23036 2694 23066 2746
rect 23066 2694 23078 2746
rect 23078 2694 23092 2746
rect 23116 2694 23130 2746
rect 23130 2694 23142 2746
rect 23142 2694 23172 2746
rect 23196 2694 23206 2746
rect 23206 2694 23252 2746
rect 22956 2692 23012 2694
rect 23036 2692 23092 2694
rect 23116 2692 23172 2694
rect 23196 2692 23252 2694
rect 23938 10668 23994 10704
rect 23938 10648 23940 10668
rect 23940 10648 23992 10668
rect 23992 10648 23994 10668
rect 26698 14048 26754 14104
rect 25962 12688 26018 12744
rect 24950 12164 25006 12200
rect 24950 12144 24952 12164
rect 24952 12144 25004 12164
rect 25004 12144 25006 12164
rect 24766 11328 24822 11384
rect 24674 10512 24730 10568
rect 23938 3440 23994 3496
rect 24582 9868 24584 9888
rect 24584 9868 24636 9888
rect 24636 9868 24638 9888
rect 24582 9832 24638 9868
rect 24950 8900 25006 8936
rect 24950 8880 24952 8900
rect 24952 8880 25004 8900
rect 25004 8880 25006 8900
rect 24674 7248 24730 7304
rect 24582 6704 24638 6760
rect 25134 8064 25190 8120
rect 24766 6432 24822 6488
rect 24858 2896 24914 2952
rect 24858 720 24914 776
<< metal3 >>
rect 26200 56266 27000 56296
rect 23430 56206 27000 56266
rect 23430 56133 23490 56206
rect 26200 56176 27000 56206
rect 23381 56128 23490 56133
rect 23381 56072 23386 56128
rect 23442 56072 23490 56128
rect 23381 56070 23490 56072
rect 23381 56067 23447 56070
rect 24485 55450 24551 55453
rect 26200 55450 27000 55480
rect 24485 55448 27000 55450
rect 24485 55392 24490 55448
rect 24546 55392 27000 55448
rect 24485 55390 27000 55392
rect 24485 55387 24551 55390
rect 26200 55360 27000 55390
rect 24669 54634 24735 54637
rect 26200 54634 27000 54664
rect 24669 54632 27000 54634
rect 24669 54576 24674 54632
rect 24730 54576 27000 54632
rect 24669 54574 27000 54576
rect 24669 54571 24735 54574
rect 26200 54544 27000 54574
rect 7946 54432 8262 54433
rect 7946 54368 7952 54432
rect 8016 54368 8032 54432
rect 8096 54368 8112 54432
rect 8176 54368 8192 54432
rect 8256 54368 8262 54432
rect 7946 54367 8262 54368
rect 17946 54432 18262 54433
rect 17946 54368 17952 54432
rect 18016 54368 18032 54432
rect 18096 54368 18112 54432
rect 18176 54368 18192 54432
rect 18256 54368 18262 54432
rect 17946 54367 18262 54368
rect 2946 53888 3262 53889
rect 2946 53824 2952 53888
rect 3016 53824 3032 53888
rect 3096 53824 3112 53888
rect 3176 53824 3192 53888
rect 3256 53824 3262 53888
rect 2946 53823 3262 53824
rect 12946 53888 13262 53889
rect 12946 53824 12952 53888
rect 13016 53824 13032 53888
rect 13096 53824 13112 53888
rect 13176 53824 13192 53888
rect 13256 53824 13262 53888
rect 12946 53823 13262 53824
rect 22946 53888 23262 53889
rect 22946 53824 22952 53888
rect 23016 53824 23032 53888
rect 23096 53824 23112 53888
rect 23176 53824 23192 53888
rect 23256 53824 23262 53888
rect 22946 53823 23262 53824
rect 24761 53818 24827 53821
rect 26200 53818 27000 53848
rect 24761 53816 27000 53818
rect 24761 53760 24766 53816
rect 24822 53760 27000 53816
rect 24761 53758 27000 53760
rect 24761 53755 24827 53758
rect 26200 53728 27000 53758
rect 7946 53344 8262 53345
rect 7946 53280 7952 53344
rect 8016 53280 8032 53344
rect 8096 53280 8112 53344
rect 8176 53280 8192 53344
rect 8256 53280 8262 53344
rect 7946 53279 8262 53280
rect 17946 53344 18262 53345
rect 17946 53280 17952 53344
rect 18016 53280 18032 53344
rect 18096 53280 18112 53344
rect 18176 53280 18192 53344
rect 18256 53280 18262 53344
rect 17946 53279 18262 53280
rect 25037 53002 25103 53005
rect 26200 53002 27000 53032
rect 25037 53000 27000 53002
rect 25037 52944 25042 53000
rect 25098 52944 27000 53000
rect 25037 52942 27000 52944
rect 25037 52939 25103 52942
rect 26200 52912 27000 52942
rect 2946 52800 3262 52801
rect 2946 52736 2952 52800
rect 3016 52736 3032 52800
rect 3096 52736 3112 52800
rect 3176 52736 3192 52800
rect 3256 52736 3262 52800
rect 2946 52735 3262 52736
rect 12946 52800 13262 52801
rect 12946 52736 12952 52800
rect 13016 52736 13032 52800
rect 13096 52736 13112 52800
rect 13176 52736 13192 52800
rect 13256 52736 13262 52800
rect 12946 52735 13262 52736
rect 22946 52800 23262 52801
rect 22946 52736 22952 52800
rect 23016 52736 23032 52800
rect 23096 52736 23112 52800
rect 23176 52736 23192 52800
rect 23256 52736 23262 52800
rect 22946 52735 23262 52736
rect 7946 52256 8262 52257
rect 7946 52192 7952 52256
rect 8016 52192 8032 52256
rect 8096 52192 8112 52256
rect 8176 52192 8192 52256
rect 8256 52192 8262 52256
rect 7946 52191 8262 52192
rect 17946 52256 18262 52257
rect 17946 52192 17952 52256
rect 18016 52192 18032 52256
rect 18096 52192 18112 52256
rect 18176 52192 18192 52256
rect 18256 52192 18262 52256
rect 17946 52191 18262 52192
rect 24945 52186 25011 52189
rect 26200 52186 27000 52216
rect 24945 52184 27000 52186
rect 24945 52128 24950 52184
rect 25006 52128 27000 52184
rect 24945 52126 27000 52128
rect 24945 52123 25011 52126
rect 26200 52096 27000 52126
rect 2946 51712 3262 51713
rect 2946 51648 2952 51712
rect 3016 51648 3032 51712
rect 3096 51648 3112 51712
rect 3176 51648 3192 51712
rect 3256 51648 3262 51712
rect 2946 51647 3262 51648
rect 12946 51712 13262 51713
rect 12946 51648 12952 51712
rect 13016 51648 13032 51712
rect 13096 51648 13112 51712
rect 13176 51648 13192 51712
rect 13256 51648 13262 51712
rect 12946 51647 13262 51648
rect 22946 51712 23262 51713
rect 22946 51648 22952 51712
rect 23016 51648 23032 51712
rect 23096 51648 23112 51712
rect 23176 51648 23192 51712
rect 23256 51648 23262 51712
rect 22946 51647 23262 51648
rect 25497 51370 25563 51373
rect 26200 51370 27000 51400
rect 25497 51368 27000 51370
rect 25497 51312 25502 51368
rect 25558 51312 27000 51368
rect 25497 51310 27000 51312
rect 25497 51307 25563 51310
rect 26200 51280 27000 51310
rect 7946 51168 8262 51169
rect 7946 51104 7952 51168
rect 8016 51104 8032 51168
rect 8096 51104 8112 51168
rect 8176 51104 8192 51168
rect 8256 51104 8262 51168
rect 7946 51103 8262 51104
rect 17946 51168 18262 51169
rect 17946 51104 17952 51168
rect 18016 51104 18032 51168
rect 18096 51104 18112 51168
rect 18176 51104 18192 51168
rect 18256 51104 18262 51168
rect 17946 51103 18262 51104
rect 2946 50624 3262 50625
rect 2946 50560 2952 50624
rect 3016 50560 3032 50624
rect 3096 50560 3112 50624
rect 3176 50560 3192 50624
rect 3256 50560 3262 50624
rect 2946 50559 3262 50560
rect 12946 50624 13262 50625
rect 12946 50560 12952 50624
rect 13016 50560 13032 50624
rect 13096 50560 13112 50624
rect 13176 50560 13192 50624
rect 13256 50560 13262 50624
rect 12946 50559 13262 50560
rect 22946 50624 23262 50625
rect 22946 50560 22952 50624
rect 23016 50560 23032 50624
rect 23096 50560 23112 50624
rect 23176 50560 23192 50624
rect 23256 50560 23262 50624
rect 22946 50559 23262 50560
rect 24945 50554 25011 50557
rect 26200 50554 27000 50584
rect 24945 50552 27000 50554
rect 24945 50496 24950 50552
rect 25006 50496 27000 50552
rect 24945 50494 27000 50496
rect 24945 50491 25011 50494
rect 26200 50464 27000 50494
rect 7946 50080 8262 50081
rect 7946 50016 7952 50080
rect 8016 50016 8032 50080
rect 8096 50016 8112 50080
rect 8176 50016 8192 50080
rect 8256 50016 8262 50080
rect 7946 50015 8262 50016
rect 17946 50080 18262 50081
rect 17946 50016 17952 50080
rect 18016 50016 18032 50080
rect 18096 50016 18112 50080
rect 18176 50016 18192 50080
rect 18256 50016 18262 50080
rect 17946 50015 18262 50016
rect 25497 49738 25563 49741
rect 26200 49738 27000 49768
rect 25497 49736 27000 49738
rect 25497 49680 25502 49736
rect 25558 49680 27000 49736
rect 25497 49678 27000 49680
rect 25497 49675 25563 49678
rect 26200 49648 27000 49678
rect 2946 49536 3262 49537
rect 2946 49472 2952 49536
rect 3016 49472 3032 49536
rect 3096 49472 3112 49536
rect 3176 49472 3192 49536
rect 3256 49472 3262 49536
rect 2946 49471 3262 49472
rect 12946 49536 13262 49537
rect 12946 49472 12952 49536
rect 13016 49472 13032 49536
rect 13096 49472 13112 49536
rect 13176 49472 13192 49536
rect 13256 49472 13262 49536
rect 12946 49471 13262 49472
rect 22946 49536 23262 49537
rect 22946 49472 22952 49536
rect 23016 49472 23032 49536
rect 23096 49472 23112 49536
rect 23176 49472 23192 49536
rect 23256 49472 23262 49536
rect 22946 49471 23262 49472
rect 7946 48992 8262 48993
rect 7946 48928 7952 48992
rect 8016 48928 8032 48992
rect 8096 48928 8112 48992
rect 8176 48928 8192 48992
rect 8256 48928 8262 48992
rect 7946 48927 8262 48928
rect 17946 48992 18262 48993
rect 17946 48928 17952 48992
rect 18016 48928 18032 48992
rect 18096 48928 18112 48992
rect 18176 48928 18192 48992
rect 18256 48928 18262 48992
rect 17946 48927 18262 48928
rect 25129 48922 25195 48925
rect 26200 48922 27000 48952
rect 25129 48920 27000 48922
rect 25129 48864 25134 48920
rect 25190 48864 27000 48920
rect 25129 48862 27000 48864
rect 25129 48859 25195 48862
rect 26200 48832 27000 48862
rect 2946 48448 3262 48449
rect 2946 48384 2952 48448
rect 3016 48384 3032 48448
rect 3096 48384 3112 48448
rect 3176 48384 3192 48448
rect 3256 48384 3262 48448
rect 2946 48383 3262 48384
rect 12946 48448 13262 48449
rect 12946 48384 12952 48448
rect 13016 48384 13032 48448
rect 13096 48384 13112 48448
rect 13176 48384 13192 48448
rect 13256 48384 13262 48448
rect 12946 48383 13262 48384
rect 22946 48448 23262 48449
rect 22946 48384 22952 48448
rect 23016 48384 23032 48448
rect 23096 48384 23112 48448
rect 23176 48384 23192 48448
rect 23256 48384 23262 48448
rect 22946 48383 23262 48384
rect 25129 48106 25195 48109
rect 26200 48106 27000 48136
rect 25129 48104 27000 48106
rect 25129 48048 25134 48104
rect 25190 48048 27000 48104
rect 25129 48046 27000 48048
rect 25129 48043 25195 48046
rect 26200 48016 27000 48046
rect 7946 47904 8262 47905
rect 7946 47840 7952 47904
rect 8016 47840 8032 47904
rect 8096 47840 8112 47904
rect 8176 47840 8192 47904
rect 8256 47840 8262 47904
rect 7946 47839 8262 47840
rect 17946 47904 18262 47905
rect 17946 47840 17952 47904
rect 18016 47840 18032 47904
rect 18096 47840 18112 47904
rect 18176 47840 18192 47904
rect 18256 47840 18262 47904
rect 17946 47839 18262 47840
rect 2946 47360 3262 47361
rect 2946 47296 2952 47360
rect 3016 47296 3032 47360
rect 3096 47296 3112 47360
rect 3176 47296 3192 47360
rect 3256 47296 3262 47360
rect 2946 47295 3262 47296
rect 12946 47360 13262 47361
rect 12946 47296 12952 47360
rect 13016 47296 13032 47360
rect 13096 47296 13112 47360
rect 13176 47296 13192 47360
rect 13256 47296 13262 47360
rect 12946 47295 13262 47296
rect 22946 47360 23262 47361
rect 22946 47296 22952 47360
rect 23016 47296 23032 47360
rect 23096 47296 23112 47360
rect 23176 47296 23192 47360
rect 23256 47296 23262 47360
rect 22946 47295 23262 47296
rect 25313 47290 25379 47293
rect 26200 47290 27000 47320
rect 25313 47288 27000 47290
rect 25313 47232 25318 47288
rect 25374 47232 27000 47288
rect 25313 47230 27000 47232
rect 25313 47227 25379 47230
rect 26200 47200 27000 47230
rect 7946 46816 8262 46817
rect 7946 46752 7952 46816
rect 8016 46752 8032 46816
rect 8096 46752 8112 46816
rect 8176 46752 8192 46816
rect 8256 46752 8262 46816
rect 7946 46751 8262 46752
rect 17946 46816 18262 46817
rect 17946 46752 17952 46816
rect 18016 46752 18032 46816
rect 18096 46752 18112 46816
rect 18176 46752 18192 46816
rect 18256 46752 18262 46816
rect 17946 46751 18262 46752
rect 25313 46474 25379 46477
rect 26200 46474 27000 46504
rect 25313 46472 27000 46474
rect 25313 46416 25318 46472
rect 25374 46416 27000 46472
rect 25313 46414 27000 46416
rect 25313 46411 25379 46414
rect 26200 46384 27000 46414
rect 2946 46272 3262 46273
rect 2946 46208 2952 46272
rect 3016 46208 3032 46272
rect 3096 46208 3112 46272
rect 3176 46208 3192 46272
rect 3256 46208 3262 46272
rect 2946 46207 3262 46208
rect 12946 46272 13262 46273
rect 12946 46208 12952 46272
rect 13016 46208 13032 46272
rect 13096 46208 13112 46272
rect 13176 46208 13192 46272
rect 13256 46208 13262 46272
rect 12946 46207 13262 46208
rect 22946 46272 23262 46273
rect 22946 46208 22952 46272
rect 23016 46208 23032 46272
rect 23096 46208 23112 46272
rect 23176 46208 23192 46272
rect 23256 46208 23262 46272
rect 22946 46207 23262 46208
rect 7946 45728 8262 45729
rect 7946 45664 7952 45728
rect 8016 45664 8032 45728
rect 8096 45664 8112 45728
rect 8176 45664 8192 45728
rect 8256 45664 8262 45728
rect 7946 45663 8262 45664
rect 17946 45728 18262 45729
rect 17946 45664 17952 45728
rect 18016 45664 18032 45728
rect 18096 45664 18112 45728
rect 18176 45664 18192 45728
rect 18256 45664 18262 45728
rect 17946 45663 18262 45664
rect 25313 45658 25379 45661
rect 26200 45658 27000 45688
rect 25313 45656 27000 45658
rect 25313 45600 25318 45656
rect 25374 45600 27000 45656
rect 25313 45598 27000 45600
rect 25313 45595 25379 45598
rect 26200 45568 27000 45598
rect 2946 45184 3262 45185
rect 2946 45120 2952 45184
rect 3016 45120 3032 45184
rect 3096 45120 3112 45184
rect 3176 45120 3192 45184
rect 3256 45120 3262 45184
rect 2946 45119 3262 45120
rect 12946 45184 13262 45185
rect 12946 45120 12952 45184
rect 13016 45120 13032 45184
rect 13096 45120 13112 45184
rect 13176 45120 13192 45184
rect 13256 45120 13262 45184
rect 12946 45119 13262 45120
rect 22946 45184 23262 45185
rect 22946 45120 22952 45184
rect 23016 45120 23032 45184
rect 23096 45120 23112 45184
rect 23176 45120 23192 45184
rect 23256 45120 23262 45184
rect 22946 45119 23262 45120
rect 25313 44842 25379 44845
rect 26200 44842 27000 44872
rect 25313 44840 27000 44842
rect 25313 44784 25318 44840
rect 25374 44784 27000 44840
rect 25313 44782 27000 44784
rect 25313 44779 25379 44782
rect 26200 44752 27000 44782
rect 7946 44640 8262 44641
rect 7946 44576 7952 44640
rect 8016 44576 8032 44640
rect 8096 44576 8112 44640
rect 8176 44576 8192 44640
rect 8256 44576 8262 44640
rect 7946 44575 8262 44576
rect 17946 44640 18262 44641
rect 17946 44576 17952 44640
rect 18016 44576 18032 44640
rect 18096 44576 18112 44640
rect 18176 44576 18192 44640
rect 18256 44576 18262 44640
rect 17946 44575 18262 44576
rect 2946 44096 3262 44097
rect 2946 44032 2952 44096
rect 3016 44032 3032 44096
rect 3096 44032 3112 44096
rect 3176 44032 3192 44096
rect 3256 44032 3262 44096
rect 2946 44031 3262 44032
rect 12946 44096 13262 44097
rect 12946 44032 12952 44096
rect 13016 44032 13032 44096
rect 13096 44032 13112 44096
rect 13176 44032 13192 44096
rect 13256 44032 13262 44096
rect 12946 44031 13262 44032
rect 22946 44096 23262 44097
rect 22946 44032 22952 44096
rect 23016 44032 23032 44096
rect 23096 44032 23112 44096
rect 23176 44032 23192 44096
rect 23256 44032 23262 44096
rect 22946 44031 23262 44032
rect 24761 44026 24827 44029
rect 26200 44026 27000 44056
rect 24761 44024 27000 44026
rect 24761 43968 24766 44024
rect 24822 43968 27000 44024
rect 24761 43966 27000 43968
rect 24761 43963 24827 43966
rect 26200 43936 27000 43966
rect 7946 43552 8262 43553
rect 7946 43488 7952 43552
rect 8016 43488 8032 43552
rect 8096 43488 8112 43552
rect 8176 43488 8192 43552
rect 8256 43488 8262 43552
rect 7946 43487 8262 43488
rect 17946 43552 18262 43553
rect 17946 43488 17952 43552
rect 18016 43488 18032 43552
rect 18096 43488 18112 43552
rect 18176 43488 18192 43552
rect 18256 43488 18262 43552
rect 17946 43487 18262 43488
rect 25497 43210 25563 43213
rect 26200 43210 27000 43240
rect 25497 43208 27000 43210
rect 25497 43152 25502 43208
rect 25558 43152 27000 43208
rect 25497 43150 27000 43152
rect 25497 43147 25563 43150
rect 26200 43120 27000 43150
rect 2946 43008 3262 43009
rect 2946 42944 2952 43008
rect 3016 42944 3032 43008
rect 3096 42944 3112 43008
rect 3176 42944 3192 43008
rect 3256 42944 3262 43008
rect 2946 42943 3262 42944
rect 12946 43008 13262 43009
rect 12946 42944 12952 43008
rect 13016 42944 13032 43008
rect 13096 42944 13112 43008
rect 13176 42944 13192 43008
rect 13256 42944 13262 43008
rect 12946 42943 13262 42944
rect 22946 43008 23262 43009
rect 22946 42944 22952 43008
rect 23016 42944 23032 43008
rect 23096 42944 23112 43008
rect 23176 42944 23192 43008
rect 23256 42944 23262 43008
rect 22946 42943 23262 42944
rect 7946 42464 8262 42465
rect 7946 42400 7952 42464
rect 8016 42400 8032 42464
rect 8096 42400 8112 42464
rect 8176 42400 8192 42464
rect 8256 42400 8262 42464
rect 7946 42399 8262 42400
rect 17946 42464 18262 42465
rect 17946 42400 17952 42464
rect 18016 42400 18032 42464
rect 18096 42400 18112 42464
rect 18176 42400 18192 42464
rect 18256 42400 18262 42464
rect 17946 42399 18262 42400
rect 25129 42394 25195 42397
rect 26200 42394 27000 42424
rect 25129 42392 27000 42394
rect 25129 42336 25134 42392
rect 25190 42336 27000 42392
rect 25129 42334 27000 42336
rect 25129 42331 25195 42334
rect 26200 42304 27000 42334
rect 2946 41920 3262 41921
rect 2946 41856 2952 41920
rect 3016 41856 3032 41920
rect 3096 41856 3112 41920
rect 3176 41856 3192 41920
rect 3256 41856 3262 41920
rect 2946 41855 3262 41856
rect 12946 41920 13262 41921
rect 12946 41856 12952 41920
rect 13016 41856 13032 41920
rect 13096 41856 13112 41920
rect 13176 41856 13192 41920
rect 13256 41856 13262 41920
rect 12946 41855 13262 41856
rect 22946 41920 23262 41921
rect 22946 41856 22952 41920
rect 23016 41856 23032 41920
rect 23096 41856 23112 41920
rect 23176 41856 23192 41920
rect 23256 41856 23262 41920
rect 22946 41855 23262 41856
rect 25129 41578 25195 41581
rect 26200 41578 27000 41608
rect 25129 41576 27000 41578
rect 25129 41520 25134 41576
rect 25190 41520 27000 41576
rect 25129 41518 27000 41520
rect 25129 41515 25195 41518
rect 26200 41488 27000 41518
rect 7946 41376 8262 41377
rect 7946 41312 7952 41376
rect 8016 41312 8032 41376
rect 8096 41312 8112 41376
rect 8176 41312 8192 41376
rect 8256 41312 8262 41376
rect 7946 41311 8262 41312
rect 17946 41376 18262 41377
rect 17946 41312 17952 41376
rect 18016 41312 18032 41376
rect 18096 41312 18112 41376
rect 18176 41312 18192 41376
rect 18256 41312 18262 41376
rect 17946 41311 18262 41312
rect 2946 40832 3262 40833
rect 2946 40768 2952 40832
rect 3016 40768 3032 40832
rect 3096 40768 3112 40832
rect 3176 40768 3192 40832
rect 3256 40768 3262 40832
rect 2946 40767 3262 40768
rect 12946 40832 13262 40833
rect 12946 40768 12952 40832
rect 13016 40768 13032 40832
rect 13096 40768 13112 40832
rect 13176 40768 13192 40832
rect 13256 40768 13262 40832
rect 12946 40767 13262 40768
rect 22946 40832 23262 40833
rect 22946 40768 22952 40832
rect 23016 40768 23032 40832
rect 23096 40768 23112 40832
rect 23176 40768 23192 40832
rect 23256 40768 23262 40832
rect 22946 40767 23262 40768
rect 25313 40762 25379 40765
rect 26200 40762 27000 40792
rect 25313 40760 27000 40762
rect 25313 40704 25318 40760
rect 25374 40704 27000 40760
rect 25313 40702 27000 40704
rect 25313 40699 25379 40702
rect 26200 40672 27000 40702
rect 7946 40288 8262 40289
rect 7946 40224 7952 40288
rect 8016 40224 8032 40288
rect 8096 40224 8112 40288
rect 8176 40224 8192 40288
rect 8256 40224 8262 40288
rect 7946 40223 8262 40224
rect 17946 40288 18262 40289
rect 17946 40224 17952 40288
rect 18016 40224 18032 40288
rect 18096 40224 18112 40288
rect 18176 40224 18192 40288
rect 18256 40224 18262 40288
rect 17946 40223 18262 40224
rect 25405 39946 25471 39949
rect 26200 39946 27000 39976
rect 25405 39944 27000 39946
rect 25405 39888 25410 39944
rect 25466 39888 27000 39944
rect 25405 39886 27000 39888
rect 25405 39883 25471 39886
rect 26200 39856 27000 39886
rect 2946 39744 3262 39745
rect 2946 39680 2952 39744
rect 3016 39680 3032 39744
rect 3096 39680 3112 39744
rect 3176 39680 3192 39744
rect 3256 39680 3262 39744
rect 2946 39679 3262 39680
rect 12946 39744 13262 39745
rect 12946 39680 12952 39744
rect 13016 39680 13032 39744
rect 13096 39680 13112 39744
rect 13176 39680 13192 39744
rect 13256 39680 13262 39744
rect 12946 39679 13262 39680
rect 22946 39744 23262 39745
rect 22946 39680 22952 39744
rect 23016 39680 23032 39744
rect 23096 39680 23112 39744
rect 23176 39680 23192 39744
rect 23256 39680 23262 39744
rect 22946 39679 23262 39680
rect 7946 39200 8262 39201
rect 7946 39136 7952 39200
rect 8016 39136 8032 39200
rect 8096 39136 8112 39200
rect 8176 39136 8192 39200
rect 8256 39136 8262 39200
rect 7946 39135 8262 39136
rect 17946 39200 18262 39201
rect 17946 39136 17952 39200
rect 18016 39136 18032 39200
rect 18096 39136 18112 39200
rect 18176 39136 18192 39200
rect 18256 39136 18262 39200
rect 17946 39135 18262 39136
rect 25313 39130 25379 39133
rect 26200 39130 27000 39160
rect 25313 39128 27000 39130
rect 25313 39072 25318 39128
rect 25374 39072 27000 39128
rect 25313 39070 27000 39072
rect 25313 39067 25379 39070
rect 26200 39040 27000 39070
rect 2946 38656 3262 38657
rect 2946 38592 2952 38656
rect 3016 38592 3032 38656
rect 3096 38592 3112 38656
rect 3176 38592 3192 38656
rect 3256 38592 3262 38656
rect 2946 38591 3262 38592
rect 12946 38656 13262 38657
rect 12946 38592 12952 38656
rect 13016 38592 13032 38656
rect 13096 38592 13112 38656
rect 13176 38592 13192 38656
rect 13256 38592 13262 38656
rect 12946 38591 13262 38592
rect 22946 38656 23262 38657
rect 22946 38592 22952 38656
rect 23016 38592 23032 38656
rect 23096 38592 23112 38656
rect 23176 38592 23192 38656
rect 23256 38592 23262 38656
rect 22946 38591 23262 38592
rect 25313 38314 25379 38317
rect 26200 38314 27000 38344
rect 25313 38312 27000 38314
rect 25313 38256 25318 38312
rect 25374 38256 27000 38312
rect 25313 38254 27000 38256
rect 25313 38251 25379 38254
rect 26200 38224 27000 38254
rect 7946 38112 8262 38113
rect 7946 38048 7952 38112
rect 8016 38048 8032 38112
rect 8096 38048 8112 38112
rect 8176 38048 8192 38112
rect 8256 38048 8262 38112
rect 7946 38047 8262 38048
rect 17946 38112 18262 38113
rect 17946 38048 17952 38112
rect 18016 38048 18032 38112
rect 18096 38048 18112 38112
rect 18176 38048 18192 38112
rect 18256 38048 18262 38112
rect 17946 38047 18262 38048
rect 2946 37568 3262 37569
rect 2946 37504 2952 37568
rect 3016 37504 3032 37568
rect 3096 37504 3112 37568
rect 3176 37504 3192 37568
rect 3256 37504 3262 37568
rect 2946 37503 3262 37504
rect 12946 37568 13262 37569
rect 12946 37504 12952 37568
rect 13016 37504 13032 37568
rect 13096 37504 13112 37568
rect 13176 37504 13192 37568
rect 13256 37504 13262 37568
rect 12946 37503 13262 37504
rect 22946 37568 23262 37569
rect 22946 37504 22952 37568
rect 23016 37504 23032 37568
rect 23096 37504 23112 37568
rect 23176 37504 23192 37568
rect 23256 37504 23262 37568
rect 22946 37503 23262 37504
rect 25129 37498 25195 37501
rect 26200 37498 27000 37528
rect 25129 37496 27000 37498
rect 25129 37440 25134 37496
rect 25190 37440 27000 37496
rect 25129 37438 27000 37440
rect 25129 37435 25195 37438
rect 26200 37408 27000 37438
rect 7946 37024 8262 37025
rect 7946 36960 7952 37024
rect 8016 36960 8032 37024
rect 8096 36960 8112 37024
rect 8176 36960 8192 37024
rect 8256 36960 8262 37024
rect 7946 36959 8262 36960
rect 17946 37024 18262 37025
rect 17946 36960 17952 37024
rect 18016 36960 18032 37024
rect 18096 36960 18112 37024
rect 18176 36960 18192 37024
rect 18256 36960 18262 37024
rect 17946 36959 18262 36960
rect 25129 36682 25195 36685
rect 26200 36682 27000 36712
rect 25129 36680 27000 36682
rect 25129 36624 25134 36680
rect 25190 36624 27000 36680
rect 25129 36622 27000 36624
rect 25129 36619 25195 36622
rect 26200 36592 27000 36622
rect 2946 36480 3262 36481
rect 2946 36416 2952 36480
rect 3016 36416 3032 36480
rect 3096 36416 3112 36480
rect 3176 36416 3192 36480
rect 3256 36416 3262 36480
rect 2946 36415 3262 36416
rect 12946 36480 13262 36481
rect 12946 36416 12952 36480
rect 13016 36416 13032 36480
rect 13096 36416 13112 36480
rect 13176 36416 13192 36480
rect 13256 36416 13262 36480
rect 12946 36415 13262 36416
rect 22946 36480 23262 36481
rect 22946 36416 22952 36480
rect 23016 36416 23032 36480
rect 23096 36416 23112 36480
rect 23176 36416 23192 36480
rect 23256 36416 23262 36480
rect 22946 36415 23262 36416
rect 7946 35936 8262 35937
rect 7946 35872 7952 35936
rect 8016 35872 8032 35936
rect 8096 35872 8112 35936
rect 8176 35872 8192 35936
rect 8256 35872 8262 35936
rect 7946 35871 8262 35872
rect 17946 35936 18262 35937
rect 17946 35872 17952 35936
rect 18016 35872 18032 35936
rect 18096 35872 18112 35936
rect 18176 35872 18192 35936
rect 18256 35872 18262 35936
rect 17946 35871 18262 35872
rect 25313 35866 25379 35869
rect 26200 35866 27000 35896
rect 25313 35864 27000 35866
rect 25313 35808 25318 35864
rect 25374 35808 27000 35864
rect 25313 35806 27000 35808
rect 25313 35803 25379 35806
rect 26200 35776 27000 35806
rect 2946 35392 3262 35393
rect 2946 35328 2952 35392
rect 3016 35328 3032 35392
rect 3096 35328 3112 35392
rect 3176 35328 3192 35392
rect 3256 35328 3262 35392
rect 2946 35327 3262 35328
rect 12946 35392 13262 35393
rect 12946 35328 12952 35392
rect 13016 35328 13032 35392
rect 13096 35328 13112 35392
rect 13176 35328 13192 35392
rect 13256 35328 13262 35392
rect 12946 35327 13262 35328
rect 22946 35392 23262 35393
rect 22946 35328 22952 35392
rect 23016 35328 23032 35392
rect 23096 35328 23112 35392
rect 23176 35328 23192 35392
rect 23256 35328 23262 35392
rect 22946 35327 23262 35328
rect 24669 35186 24735 35189
rect 24669 35184 24778 35186
rect 24669 35128 24674 35184
rect 24730 35128 24778 35184
rect 24669 35123 24778 35128
rect 24718 35050 24778 35123
rect 26200 35050 27000 35080
rect 24718 34990 27000 35050
rect 26200 34960 27000 34990
rect 7946 34848 8262 34849
rect 7946 34784 7952 34848
rect 8016 34784 8032 34848
rect 8096 34784 8112 34848
rect 8176 34784 8192 34848
rect 8256 34784 8262 34848
rect 7946 34783 8262 34784
rect 17946 34848 18262 34849
rect 17946 34784 17952 34848
rect 18016 34784 18032 34848
rect 18096 34784 18112 34848
rect 18176 34784 18192 34848
rect 18256 34784 18262 34848
rect 17946 34783 18262 34784
rect 2946 34304 3262 34305
rect 2946 34240 2952 34304
rect 3016 34240 3032 34304
rect 3096 34240 3112 34304
rect 3176 34240 3192 34304
rect 3256 34240 3262 34304
rect 2946 34239 3262 34240
rect 12946 34304 13262 34305
rect 12946 34240 12952 34304
rect 13016 34240 13032 34304
rect 13096 34240 13112 34304
rect 13176 34240 13192 34304
rect 13256 34240 13262 34304
rect 12946 34239 13262 34240
rect 22946 34304 23262 34305
rect 22946 34240 22952 34304
rect 23016 34240 23032 34304
rect 23096 34240 23112 34304
rect 23176 34240 23192 34304
rect 23256 34240 23262 34304
rect 22946 34239 23262 34240
rect 24761 34234 24827 34237
rect 26200 34234 27000 34264
rect 24761 34232 27000 34234
rect 24761 34176 24766 34232
rect 24822 34176 27000 34232
rect 24761 34174 27000 34176
rect 24761 34171 24827 34174
rect 26200 34144 27000 34174
rect 7946 33760 8262 33761
rect 7946 33696 7952 33760
rect 8016 33696 8032 33760
rect 8096 33696 8112 33760
rect 8176 33696 8192 33760
rect 8256 33696 8262 33760
rect 7946 33695 8262 33696
rect 17946 33760 18262 33761
rect 17946 33696 17952 33760
rect 18016 33696 18032 33760
rect 18096 33696 18112 33760
rect 18176 33696 18192 33760
rect 18256 33696 18262 33760
rect 17946 33695 18262 33696
rect 24669 33418 24735 33421
rect 26200 33418 27000 33448
rect 24669 33416 27000 33418
rect 24669 33360 24674 33416
rect 24730 33360 27000 33416
rect 24669 33358 27000 33360
rect 24669 33355 24735 33358
rect 26200 33328 27000 33358
rect 2946 33216 3262 33217
rect 2946 33152 2952 33216
rect 3016 33152 3032 33216
rect 3096 33152 3112 33216
rect 3176 33152 3192 33216
rect 3256 33152 3262 33216
rect 2946 33151 3262 33152
rect 12946 33216 13262 33217
rect 12946 33152 12952 33216
rect 13016 33152 13032 33216
rect 13096 33152 13112 33216
rect 13176 33152 13192 33216
rect 13256 33152 13262 33216
rect 12946 33151 13262 33152
rect 22946 33216 23262 33217
rect 22946 33152 22952 33216
rect 23016 33152 23032 33216
rect 23096 33152 23112 33216
rect 23176 33152 23192 33216
rect 23256 33152 23262 33216
rect 22946 33151 23262 33152
rect 7946 32672 8262 32673
rect 7946 32608 7952 32672
rect 8016 32608 8032 32672
rect 8096 32608 8112 32672
rect 8176 32608 8192 32672
rect 8256 32608 8262 32672
rect 7946 32607 8262 32608
rect 17946 32672 18262 32673
rect 17946 32608 17952 32672
rect 18016 32608 18032 32672
rect 18096 32608 18112 32672
rect 18176 32608 18192 32672
rect 18256 32608 18262 32672
rect 17946 32607 18262 32608
rect 24577 32602 24643 32605
rect 26200 32602 27000 32632
rect 24577 32600 27000 32602
rect 24577 32544 24582 32600
rect 24638 32544 27000 32600
rect 24577 32542 27000 32544
rect 24577 32539 24643 32542
rect 26200 32512 27000 32542
rect 2946 32128 3262 32129
rect 2946 32064 2952 32128
rect 3016 32064 3032 32128
rect 3096 32064 3112 32128
rect 3176 32064 3192 32128
rect 3256 32064 3262 32128
rect 2946 32063 3262 32064
rect 12946 32128 13262 32129
rect 12946 32064 12952 32128
rect 13016 32064 13032 32128
rect 13096 32064 13112 32128
rect 13176 32064 13192 32128
rect 13256 32064 13262 32128
rect 12946 32063 13262 32064
rect 22946 32128 23262 32129
rect 22946 32064 22952 32128
rect 23016 32064 23032 32128
rect 23096 32064 23112 32128
rect 23176 32064 23192 32128
rect 23256 32064 23262 32128
rect 22946 32063 23262 32064
rect 24485 31786 24551 31789
rect 26200 31786 27000 31816
rect 24485 31784 27000 31786
rect 24485 31728 24490 31784
rect 24546 31728 27000 31784
rect 24485 31726 27000 31728
rect 24485 31723 24551 31726
rect 26200 31696 27000 31726
rect 7946 31584 8262 31585
rect 7946 31520 7952 31584
rect 8016 31520 8032 31584
rect 8096 31520 8112 31584
rect 8176 31520 8192 31584
rect 8256 31520 8262 31584
rect 7946 31519 8262 31520
rect 17946 31584 18262 31585
rect 17946 31520 17952 31584
rect 18016 31520 18032 31584
rect 18096 31520 18112 31584
rect 18176 31520 18192 31584
rect 18256 31520 18262 31584
rect 17946 31519 18262 31520
rect 2946 31040 3262 31041
rect 2946 30976 2952 31040
rect 3016 30976 3032 31040
rect 3096 30976 3112 31040
rect 3176 30976 3192 31040
rect 3256 30976 3262 31040
rect 2946 30975 3262 30976
rect 12946 31040 13262 31041
rect 12946 30976 12952 31040
rect 13016 30976 13032 31040
rect 13096 30976 13112 31040
rect 13176 30976 13192 31040
rect 13256 30976 13262 31040
rect 12946 30975 13262 30976
rect 22946 31040 23262 31041
rect 22946 30976 22952 31040
rect 23016 30976 23032 31040
rect 23096 30976 23112 31040
rect 23176 30976 23192 31040
rect 23256 30976 23262 31040
rect 22946 30975 23262 30976
rect 25313 30970 25379 30973
rect 26200 30970 27000 31000
rect 25313 30968 27000 30970
rect 25313 30912 25318 30968
rect 25374 30912 27000 30968
rect 25313 30910 27000 30912
rect 25313 30907 25379 30910
rect 26200 30880 27000 30910
rect 7946 30496 8262 30497
rect 7946 30432 7952 30496
rect 8016 30432 8032 30496
rect 8096 30432 8112 30496
rect 8176 30432 8192 30496
rect 8256 30432 8262 30496
rect 7946 30431 8262 30432
rect 17946 30496 18262 30497
rect 17946 30432 17952 30496
rect 18016 30432 18032 30496
rect 18096 30432 18112 30496
rect 18176 30432 18192 30496
rect 18256 30432 18262 30496
rect 17946 30431 18262 30432
rect 25405 30154 25471 30157
rect 26200 30154 27000 30184
rect 25405 30152 27000 30154
rect 25405 30096 25410 30152
rect 25466 30096 27000 30152
rect 25405 30094 27000 30096
rect 25405 30091 25471 30094
rect 26200 30064 27000 30094
rect 2946 29952 3262 29953
rect 2946 29888 2952 29952
rect 3016 29888 3032 29952
rect 3096 29888 3112 29952
rect 3176 29888 3192 29952
rect 3256 29888 3262 29952
rect 2946 29887 3262 29888
rect 12946 29952 13262 29953
rect 12946 29888 12952 29952
rect 13016 29888 13032 29952
rect 13096 29888 13112 29952
rect 13176 29888 13192 29952
rect 13256 29888 13262 29952
rect 12946 29887 13262 29888
rect 22946 29952 23262 29953
rect 22946 29888 22952 29952
rect 23016 29888 23032 29952
rect 23096 29888 23112 29952
rect 23176 29888 23192 29952
rect 23256 29888 23262 29952
rect 22946 29887 23262 29888
rect 7946 29408 8262 29409
rect 7946 29344 7952 29408
rect 8016 29344 8032 29408
rect 8096 29344 8112 29408
rect 8176 29344 8192 29408
rect 8256 29344 8262 29408
rect 7946 29343 8262 29344
rect 17946 29408 18262 29409
rect 17946 29344 17952 29408
rect 18016 29344 18032 29408
rect 18096 29344 18112 29408
rect 18176 29344 18192 29408
rect 18256 29344 18262 29408
rect 17946 29343 18262 29344
rect 24853 29338 24919 29341
rect 26200 29338 27000 29368
rect 24853 29336 27000 29338
rect 24853 29280 24858 29336
rect 24914 29280 27000 29336
rect 24853 29278 27000 29280
rect 24853 29275 24919 29278
rect 26200 29248 27000 29278
rect 21214 29140 21220 29204
rect 21284 29202 21290 29204
rect 23105 29202 23171 29205
rect 21284 29200 23171 29202
rect 21284 29144 23110 29200
rect 23166 29144 23171 29200
rect 21284 29142 23171 29144
rect 21284 29140 21290 29142
rect 23105 29139 23171 29142
rect 16021 29066 16087 29069
rect 17493 29066 17559 29069
rect 16021 29064 17559 29066
rect 16021 29008 16026 29064
rect 16082 29008 17498 29064
rect 17554 29008 17559 29064
rect 16021 29006 17559 29008
rect 16021 29003 16087 29006
rect 17493 29003 17559 29006
rect 22553 29066 22619 29069
rect 22686 29066 22692 29068
rect 22553 29064 22692 29066
rect 22553 29008 22558 29064
rect 22614 29008 22692 29064
rect 22553 29006 22692 29008
rect 22553 29003 22619 29006
rect 22686 29004 22692 29006
rect 22756 29004 22762 29068
rect 2946 28864 3262 28865
rect 2946 28800 2952 28864
rect 3016 28800 3032 28864
rect 3096 28800 3112 28864
rect 3176 28800 3192 28864
rect 3256 28800 3262 28864
rect 2946 28799 3262 28800
rect 12946 28864 13262 28865
rect 12946 28800 12952 28864
rect 13016 28800 13032 28864
rect 13096 28800 13112 28864
rect 13176 28800 13192 28864
rect 13256 28800 13262 28864
rect 12946 28799 13262 28800
rect 22946 28864 23262 28865
rect 22946 28800 22952 28864
rect 23016 28800 23032 28864
rect 23096 28800 23112 28864
rect 23176 28800 23192 28864
rect 23256 28800 23262 28864
rect 22946 28799 23262 28800
rect 23197 28522 23263 28525
rect 26200 28522 27000 28552
rect 23197 28520 27000 28522
rect 23197 28464 23202 28520
rect 23258 28464 27000 28520
rect 23197 28462 27000 28464
rect 23197 28459 23263 28462
rect 26200 28432 27000 28462
rect 7946 28320 8262 28321
rect 7946 28256 7952 28320
rect 8016 28256 8032 28320
rect 8096 28256 8112 28320
rect 8176 28256 8192 28320
rect 8256 28256 8262 28320
rect 7946 28255 8262 28256
rect 17946 28320 18262 28321
rect 17946 28256 17952 28320
rect 18016 28256 18032 28320
rect 18096 28256 18112 28320
rect 18176 28256 18192 28320
rect 18256 28256 18262 28320
rect 17946 28255 18262 28256
rect 22093 27978 22159 27981
rect 22093 27976 23490 27978
rect 22093 27920 22098 27976
rect 22154 27920 23490 27976
rect 22093 27918 23490 27920
rect 22093 27915 22159 27918
rect 2946 27776 3262 27777
rect 2946 27712 2952 27776
rect 3016 27712 3032 27776
rect 3096 27712 3112 27776
rect 3176 27712 3192 27776
rect 3256 27712 3262 27776
rect 2946 27711 3262 27712
rect 12946 27776 13262 27777
rect 12946 27712 12952 27776
rect 13016 27712 13032 27776
rect 13096 27712 13112 27776
rect 13176 27712 13192 27776
rect 13256 27712 13262 27776
rect 12946 27711 13262 27712
rect 22946 27776 23262 27777
rect 22946 27712 22952 27776
rect 23016 27712 23032 27776
rect 23096 27712 23112 27776
rect 23176 27712 23192 27776
rect 23256 27712 23262 27776
rect 22946 27711 23262 27712
rect 23430 27706 23490 27918
rect 26200 27706 27000 27736
rect 23430 27646 27000 27706
rect 26200 27616 27000 27646
rect 17677 27300 17743 27301
rect 17677 27298 17724 27300
rect 17632 27296 17724 27298
rect 17632 27240 17682 27296
rect 17632 27238 17724 27240
rect 17677 27236 17724 27238
rect 17788 27236 17794 27300
rect 17677 27235 17743 27236
rect 7946 27232 8262 27233
rect 7946 27168 7952 27232
rect 8016 27168 8032 27232
rect 8096 27168 8112 27232
rect 8176 27168 8192 27232
rect 8256 27168 8262 27232
rect 7946 27167 8262 27168
rect 17946 27232 18262 27233
rect 17946 27168 17952 27232
rect 18016 27168 18032 27232
rect 18096 27168 18112 27232
rect 18176 27168 18192 27232
rect 18256 27168 18262 27232
rect 17946 27167 18262 27168
rect 21817 26890 21883 26893
rect 26200 26890 27000 26920
rect 21817 26888 27000 26890
rect 21817 26832 21822 26888
rect 21878 26832 27000 26888
rect 21817 26830 27000 26832
rect 21817 26827 21883 26830
rect 26200 26800 27000 26830
rect 2946 26688 3262 26689
rect 2946 26624 2952 26688
rect 3016 26624 3032 26688
rect 3096 26624 3112 26688
rect 3176 26624 3192 26688
rect 3256 26624 3262 26688
rect 2946 26623 3262 26624
rect 12946 26688 13262 26689
rect 12946 26624 12952 26688
rect 13016 26624 13032 26688
rect 13096 26624 13112 26688
rect 13176 26624 13192 26688
rect 13256 26624 13262 26688
rect 12946 26623 13262 26624
rect 22946 26688 23262 26689
rect 22946 26624 22952 26688
rect 23016 26624 23032 26688
rect 23096 26624 23112 26688
rect 23176 26624 23192 26688
rect 23256 26624 23262 26688
rect 22946 26623 23262 26624
rect 17953 26346 18019 26349
rect 18638 26346 18644 26348
rect 17953 26344 18644 26346
rect 17953 26288 17958 26344
rect 18014 26288 18644 26344
rect 17953 26286 18644 26288
rect 17953 26283 18019 26286
rect 18638 26284 18644 26286
rect 18708 26346 18714 26348
rect 18965 26346 19031 26349
rect 18708 26344 19031 26346
rect 18708 26288 18970 26344
rect 19026 26288 19031 26344
rect 18708 26286 19031 26288
rect 18708 26284 18714 26286
rect 18965 26283 19031 26286
rect 7946 26144 8262 26145
rect 7946 26080 7952 26144
rect 8016 26080 8032 26144
rect 8096 26080 8112 26144
rect 8176 26080 8192 26144
rect 8256 26080 8262 26144
rect 7946 26079 8262 26080
rect 17946 26144 18262 26145
rect 17946 26080 17952 26144
rect 18016 26080 18032 26144
rect 18096 26080 18112 26144
rect 18176 26080 18192 26144
rect 18256 26080 18262 26144
rect 17946 26079 18262 26080
rect 22461 26074 22527 26077
rect 26200 26074 27000 26104
rect 22461 26072 27000 26074
rect 22461 26016 22466 26072
rect 22522 26016 27000 26072
rect 22461 26014 27000 26016
rect 22461 26011 22527 26014
rect 26200 25984 27000 26014
rect 22185 25804 22251 25805
rect 22134 25740 22140 25804
rect 22204 25802 22251 25804
rect 22204 25800 22296 25802
rect 22246 25744 22296 25800
rect 22204 25742 22296 25744
rect 22204 25740 22251 25742
rect 22185 25739 22251 25740
rect 2946 25600 3262 25601
rect 2946 25536 2952 25600
rect 3016 25536 3032 25600
rect 3096 25536 3112 25600
rect 3176 25536 3192 25600
rect 3256 25536 3262 25600
rect 2946 25535 3262 25536
rect 12946 25600 13262 25601
rect 12946 25536 12952 25600
rect 13016 25536 13032 25600
rect 13096 25536 13112 25600
rect 13176 25536 13192 25600
rect 13256 25536 13262 25600
rect 12946 25535 13262 25536
rect 22946 25600 23262 25601
rect 22946 25536 22952 25600
rect 23016 25536 23032 25600
rect 23096 25536 23112 25600
rect 23176 25536 23192 25600
rect 23256 25536 23262 25600
rect 22946 25535 23262 25536
rect 24945 25258 25011 25261
rect 26200 25258 27000 25288
rect 24945 25256 27000 25258
rect 24945 25200 24950 25256
rect 25006 25200 27000 25256
rect 24945 25198 27000 25200
rect 24945 25195 25011 25198
rect 26200 25168 27000 25198
rect 15377 25124 15443 25125
rect 15326 25060 15332 25124
rect 15396 25122 15443 25124
rect 19333 25124 19399 25125
rect 19333 25122 19380 25124
rect 15396 25120 15488 25122
rect 15438 25064 15488 25120
rect 15396 25062 15488 25064
rect 19288 25120 19380 25122
rect 19288 25064 19338 25120
rect 19288 25062 19380 25064
rect 15396 25060 15443 25062
rect 15377 25059 15443 25060
rect 19333 25060 19380 25062
rect 19444 25060 19450 25124
rect 19333 25059 19399 25060
rect 7946 25056 8262 25057
rect 7946 24992 7952 25056
rect 8016 24992 8032 25056
rect 8096 24992 8112 25056
rect 8176 24992 8192 25056
rect 8256 24992 8262 25056
rect 7946 24991 8262 24992
rect 17946 25056 18262 25057
rect 17946 24992 17952 25056
rect 18016 24992 18032 25056
rect 18096 24992 18112 25056
rect 18176 24992 18192 25056
rect 18256 24992 18262 25056
rect 17946 24991 18262 24992
rect 20989 24988 21055 24989
rect 20989 24984 21036 24988
rect 21100 24986 21106 24988
rect 20989 24928 20994 24984
rect 20989 24924 21036 24928
rect 21100 24926 21146 24986
rect 21100 24924 21106 24926
rect 20989 24923 21055 24924
rect 2946 24512 3262 24513
rect 2946 24448 2952 24512
rect 3016 24448 3032 24512
rect 3096 24448 3112 24512
rect 3176 24448 3192 24512
rect 3256 24448 3262 24512
rect 2946 24447 3262 24448
rect 12946 24512 13262 24513
rect 12946 24448 12952 24512
rect 13016 24448 13032 24512
rect 13096 24448 13112 24512
rect 13176 24448 13192 24512
rect 13256 24448 13262 24512
rect 12946 24447 13262 24448
rect 22946 24512 23262 24513
rect 22946 24448 22952 24512
rect 23016 24448 23032 24512
rect 23096 24448 23112 24512
rect 23176 24448 23192 24512
rect 23256 24448 23262 24512
rect 22946 24447 23262 24448
rect 24761 24442 24827 24445
rect 26200 24442 27000 24472
rect 24761 24440 27000 24442
rect 24761 24384 24766 24440
rect 24822 24384 27000 24440
rect 24761 24382 27000 24384
rect 24761 24379 24827 24382
rect 26200 24352 27000 24382
rect 7946 23968 8262 23969
rect 7946 23904 7952 23968
rect 8016 23904 8032 23968
rect 8096 23904 8112 23968
rect 8176 23904 8192 23968
rect 8256 23904 8262 23968
rect 7946 23903 8262 23904
rect 17946 23968 18262 23969
rect 17946 23904 17952 23968
rect 18016 23904 18032 23968
rect 18096 23904 18112 23968
rect 18176 23904 18192 23968
rect 18256 23904 18262 23968
rect 17946 23903 18262 23904
rect 17166 23700 17172 23764
rect 17236 23762 17242 23764
rect 17585 23762 17651 23765
rect 17236 23760 17651 23762
rect 17236 23704 17590 23760
rect 17646 23704 17651 23760
rect 17236 23702 17651 23704
rect 17236 23700 17242 23702
rect 17585 23699 17651 23702
rect 23749 23626 23815 23629
rect 26200 23626 27000 23656
rect 23749 23624 27000 23626
rect 23749 23568 23754 23624
rect 23810 23568 27000 23624
rect 23749 23566 27000 23568
rect 23749 23563 23815 23566
rect 26200 23536 27000 23566
rect 21081 23490 21147 23493
rect 22134 23490 22140 23492
rect 21081 23488 22140 23490
rect 21081 23432 21086 23488
rect 21142 23432 22140 23488
rect 21081 23430 22140 23432
rect 21081 23427 21147 23430
rect 22134 23428 22140 23430
rect 22204 23428 22210 23492
rect 2946 23424 3262 23425
rect 2946 23360 2952 23424
rect 3016 23360 3032 23424
rect 3096 23360 3112 23424
rect 3176 23360 3192 23424
rect 3256 23360 3262 23424
rect 2946 23359 3262 23360
rect 12946 23424 13262 23425
rect 12946 23360 12952 23424
rect 13016 23360 13032 23424
rect 13096 23360 13112 23424
rect 13176 23360 13192 23424
rect 13256 23360 13262 23424
rect 12946 23359 13262 23360
rect 22946 23424 23262 23425
rect 22946 23360 22952 23424
rect 23016 23360 23032 23424
rect 23096 23360 23112 23424
rect 23176 23360 23192 23424
rect 23256 23360 23262 23424
rect 22946 23359 23262 23360
rect 7946 22880 8262 22881
rect 7946 22816 7952 22880
rect 8016 22816 8032 22880
rect 8096 22816 8112 22880
rect 8176 22816 8192 22880
rect 8256 22816 8262 22880
rect 7946 22815 8262 22816
rect 17946 22880 18262 22881
rect 17946 22816 17952 22880
rect 18016 22816 18032 22880
rect 18096 22816 18112 22880
rect 18176 22816 18192 22880
rect 18256 22816 18262 22880
rect 17946 22815 18262 22816
rect 24853 22810 24919 22813
rect 26200 22810 27000 22840
rect 24853 22808 27000 22810
rect 24853 22752 24858 22808
rect 24914 22752 27000 22808
rect 24853 22750 27000 22752
rect 24853 22747 24919 22750
rect 26200 22720 27000 22750
rect 2946 22336 3262 22337
rect 2946 22272 2952 22336
rect 3016 22272 3032 22336
rect 3096 22272 3112 22336
rect 3176 22272 3192 22336
rect 3256 22272 3262 22336
rect 2946 22271 3262 22272
rect 12946 22336 13262 22337
rect 12946 22272 12952 22336
rect 13016 22272 13032 22336
rect 13096 22272 13112 22336
rect 13176 22272 13192 22336
rect 13256 22272 13262 22336
rect 12946 22271 13262 22272
rect 22946 22336 23262 22337
rect 22946 22272 22952 22336
rect 23016 22272 23032 22336
rect 23096 22272 23112 22336
rect 23176 22272 23192 22336
rect 23256 22272 23262 22336
rect 22946 22271 23262 22272
rect 24853 21994 24919 21997
rect 26200 21994 27000 22024
rect 24853 21992 27000 21994
rect 24853 21936 24858 21992
rect 24914 21936 27000 21992
rect 24853 21934 27000 21936
rect 24853 21931 24919 21934
rect 26200 21904 27000 21934
rect 7946 21792 8262 21793
rect 7946 21728 7952 21792
rect 8016 21728 8032 21792
rect 8096 21728 8112 21792
rect 8176 21728 8192 21792
rect 8256 21728 8262 21792
rect 7946 21727 8262 21728
rect 17946 21792 18262 21793
rect 17946 21728 17952 21792
rect 18016 21728 18032 21792
rect 18096 21728 18112 21792
rect 18176 21728 18192 21792
rect 18256 21728 18262 21792
rect 17946 21727 18262 21728
rect 2946 21248 3262 21249
rect 2946 21184 2952 21248
rect 3016 21184 3032 21248
rect 3096 21184 3112 21248
rect 3176 21184 3192 21248
rect 3256 21184 3262 21248
rect 2946 21183 3262 21184
rect 12946 21248 13262 21249
rect 12946 21184 12952 21248
rect 13016 21184 13032 21248
rect 13096 21184 13112 21248
rect 13176 21184 13192 21248
rect 13256 21184 13262 21248
rect 12946 21183 13262 21184
rect 22946 21248 23262 21249
rect 22946 21184 22952 21248
rect 23016 21184 23032 21248
rect 23096 21184 23112 21248
rect 23176 21184 23192 21248
rect 23256 21184 23262 21248
rect 22946 21183 23262 21184
rect 23381 21178 23447 21181
rect 26200 21178 27000 21208
rect 23381 21176 27000 21178
rect 23381 21120 23386 21176
rect 23442 21120 27000 21176
rect 23381 21118 27000 21120
rect 23381 21115 23447 21118
rect 26200 21088 27000 21118
rect 7946 20704 8262 20705
rect 7946 20640 7952 20704
rect 8016 20640 8032 20704
rect 8096 20640 8112 20704
rect 8176 20640 8192 20704
rect 8256 20640 8262 20704
rect 7946 20639 8262 20640
rect 17946 20704 18262 20705
rect 17946 20640 17952 20704
rect 18016 20640 18032 20704
rect 18096 20640 18112 20704
rect 18176 20640 18192 20704
rect 18256 20640 18262 20704
rect 17946 20639 18262 20640
rect 23197 20362 23263 20365
rect 26200 20362 27000 20392
rect 23197 20360 27000 20362
rect 23197 20304 23202 20360
rect 23258 20304 27000 20360
rect 23197 20302 27000 20304
rect 23197 20299 23263 20302
rect 26200 20272 27000 20302
rect 2946 20160 3262 20161
rect 2946 20096 2952 20160
rect 3016 20096 3032 20160
rect 3096 20096 3112 20160
rect 3176 20096 3192 20160
rect 3256 20096 3262 20160
rect 2946 20095 3262 20096
rect 12946 20160 13262 20161
rect 12946 20096 12952 20160
rect 13016 20096 13032 20160
rect 13096 20096 13112 20160
rect 13176 20096 13192 20160
rect 13256 20096 13262 20160
rect 12946 20095 13262 20096
rect 22946 20160 23262 20161
rect 22946 20096 22952 20160
rect 23016 20096 23032 20160
rect 23096 20096 23112 20160
rect 23176 20096 23192 20160
rect 23256 20096 23262 20160
rect 22946 20095 23262 20096
rect 22645 19682 22711 19685
rect 22510 19680 22711 19682
rect 22510 19624 22650 19680
rect 22706 19624 22711 19680
rect 22510 19622 22711 19624
rect 7946 19616 8262 19617
rect 7946 19552 7952 19616
rect 8016 19552 8032 19616
rect 8096 19552 8112 19616
rect 8176 19552 8192 19616
rect 8256 19552 8262 19616
rect 7946 19551 8262 19552
rect 17946 19616 18262 19617
rect 17946 19552 17952 19616
rect 18016 19552 18032 19616
rect 18096 19552 18112 19616
rect 18176 19552 18192 19616
rect 18256 19552 18262 19616
rect 17946 19551 18262 19552
rect 19057 19410 19123 19413
rect 19190 19410 19196 19412
rect 19057 19408 19196 19410
rect 19057 19352 19062 19408
rect 19118 19352 19196 19408
rect 19057 19350 19196 19352
rect 19057 19347 19123 19350
rect 19190 19348 19196 19350
rect 19260 19348 19266 19412
rect 22510 19277 22570 19622
rect 22645 19619 22711 19622
rect 23381 19546 23447 19549
rect 26200 19546 27000 19576
rect 23381 19544 27000 19546
rect 23381 19488 23386 19544
rect 23442 19488 27000 19544
rect 23381 19486 27000 19488
rect 23381 19483 23447 19486
rect 26200 19456 27000 19486
rect 22461 19272 22570 19277
rect 22461 19216 22466 19272
rect 22522 19216 22570 19272
rect 22461 19214 22570 19216
rect 22461 19211 22527 19214
rect 2946 19072 3262 19073
rect 2946 19008 2952 19072
rect 3016 19008 3032 19072
rect 3096 19008 3112 19072
rect 3176 19008 3192 19072
rect 3256 19008 3262 19072
rect 2946 19007 3262 19008
rect 12946 19072 13262 19073
rect 12946 19008 12952 19072
rect 13016 19008 13032 19072
rect 13096 19008 13112 19072
rect 13176 19008 13192 19072
rect 13256 19008 13262 19072
rect 12946 19007 13262 19008
rect 22946 19072 23262 19073
rect 22946 19008 22952 19072
rect 23016 19008 23032 19072
rect 23096 19008 23112 19072
rect 23176 19008 23192 19072
rect 23256 19008 23262 19072
rect 22946 19007 23262 19008
rect 24761 18730 24827 18733
rect 26200 18730 27000 18760
rect 24761 18728 27000 18730
rect 24761 18672 24766 18728
rect 24822 18672 27000 18728
rect 24761 18670 27000 18672
rect 24761 18667 24827 18670
rect 26200 18640 27000 18670
rect 7946 18528 8262 18529
rect 7946 18464 7952 18528
rect 8016 18464 8032 18528
rect 8096 18464 8112 18528
rect 8176 18464 8192 18528
rect 8256 18464 8262 18528
rect 7946 18463 8262 18464
rect 17946 18528 18262 18529
rect 17946 18464 17952 18528
rect 18016 18464 18032 18528
rect 18096 18464 18112 18528
rect 18176 18464 18192 18528
rect 18256 18464 18262 18528
rect 17946 18463 18262 18464
rect 18413 18322 18479 18325
rect 18638 18322 18644 18324
rect 18413 18320 18644 18322
rect 18413 18264 18418 18320
rect 18474 18264 18644 18320
rect 18413 18262 18644 18264
rect 18413 18259 18479 18262
rect 18638 18260 18644 18262
rect 18708 18260 18714 18324
rect 18597 18188 18663 18189
rect 18597 18184 18644 18188
rect 18708 18186 18714 18188
rect 18597 18128 18602 18184
rect 18597 18124 18644 18128
rect 18708 18126 18754 18186
rect 18708 18124 18714 18126
rect 18597 18123 18663 18124
rect 21357 18052 21423 18053
rect 21357 18048 21404 18052
rect 21468 18050 21474 18052
rect 21357 17992 21362 18048
rect 21357 17988 21404 17992
rect 21468 17990 21514 18050
rect 21468 17988 21474 17990
rect 21357 17987 21423 17988
rect 2946 17984 3262 17985
rect 2946 17920 2952 17984
rect 3016 17920 3032 17984
rect 3096 17920 3112 17984
rect 3176 17920 3192 17984
rect 3256 17920 3262 17984
rect 2946 17919 3262 17920
rect 12946 17984 13262 17985
rect 12946 17920 12952 17984
rect 13016 17920 13032 17984
rect 13096 17920 13112 17984
rect 13176 17920 13192 17984
rect 13256 17920 13262 17984
rect 12946 17919 13262 17920
rect 22946 17984 23262 17985
rect 22946 17920 22952 17984
rect 23016 17920 23032 17984
rect 23096 17920 23112 17984
rect 23176 17920 23192 17984
rect 23256 17920 23262 17984
rect 22946 17919 23262 17920
rect 24853 17914 24919 17917
rect 26200 17914 27000 17944
rect 24853 17912 27000 17914
rect 24853 17856 24858 17912
rect 24914 17856 27000 17912
rect 24853 17854 27000 17856
rect 24853 17851 24919 17854
rect 26200 17824 27000 17854
rect 17861 17778 17927 17781
rect 18781 17778 18847 17781
rect 17861 17776 18847 17778
rect 17861 17720 17866 17776
rect 17922 17720 18786 17776
rect 18842 17720 18847 17776
rect 17861 17718 18847 17720
rect 17861 17715 17927 17718
rect 18781 17715 18847 17718
rect 7946 17440 8262 17441
rect 7946 17376 7952 17440
rect 8016 17376 8032 17440
rect 8096 17376 8112 17440
rect 8176 17376 8192 17440
rect 8256 17376 8262 17440
rect 7946 17375 8262 17376
rect 17946 17440 18262 17441
rect 17946 17376 17952 17440
rect 18016 17376 18032 17440
rect 18096 17376 18112 17440
rect 18176 17376 18192 17440
rect 18256 17376 18262 17440
rect 17946 17375 18262 17376
rect 21173 17372 21239 17373
rect 21173 17370 21220 17372
rect 21128 17368 21220 17370
rect 21128 17312 21178 17368
rect 21128 17310 21220 17312
rect 21173 17308 21220 17310
rect 21284 17308 21290 17372
rect 21173 17307 21239 17308
rect 16798 17036 16804 17100
rect 16868 17098 16874 17100
rect 19241 17098 19307 17101
rect 16868 17096 19307 17098
rect 16868 17040 19246 17096
rect 19302 17040 19307 17096
rect 16868 17038 19307 17040
rect 16868 17036 16874 17038
rect 19241 17035 19307 17038
rect 22093 17100 22159 17101
rect 22093 17096 22140 17100
rect 22204 17098 22210 17100
rect 24853 17098 24919 17101
rect 26200 17098 27000 17128
rect 22093 17040 22098 17096
rect 22093 17036 22140 17040
rect 22204 17038 22250 17098
rect 24853 17096 27000 17098
rect 24853 17040 24858 17096
rect 24914 17040 27000 17096
rect 24853 17038 27000 17040
rect 22204 17036 22210 17038
rect 22093 17035 22159 17036
rect 24853 17035 24919 17038
rect 26200 17008 27000 17038
rect 16665 16962 16731 16965
rect 16941 16962 17007 16965
rect 16665 16960 17007 16962
rect 16665 16904 16670 16960
rect 16726 16904 16946 16960
rect 17002 16904 17007 16960
rect 16665 16902 17007 16904
rect 16665 16899 16731 16902
rect 16941 16899 17007 16902
rect 2946 16896 3262 16897
rect 2946 16832 2952 16896
rect 3016 16832 3032 16896
rect 3096 16832 3112 16896
rect 3176 16832 3192 16896
rect 3256 16832 3262 16896
rect 2946 16831 3262 16832
rect 12946 16896 13262 16897
rect 12946 16832 12952 16896
rect 13016 16832 13032 16896
rect 13096 16832 13112 16896
rect 13176 16832 13192 16896
rect 13256 16832 13262 16896
rect 12946 16831 13262 16832
rect 22946 16896 23262 16897
rect 22946 16832 22952 16896
rect 23016 16832 23032 16896
rect 23096 16832 23112 16896
rect 23176 16832 23192 16896
rect 23256 16832 23262 16896
rect 22946 16831 23262 16832
rect 13486 16628 13492 16692
rect 13556 16690 13562 16692
rect 16665 16690 16731 16693
rect 13556 16688 16731 16690
rect 13556 16632 16670 16688
rect 16726 16632 16731 16688
rect 13556 16630 16731 16632
rect 13556 16628 13562 16630
rect 16665 16627 16731 16630
rect 19425 16690 19491 16693
rect 19558 16690 19564 16692
rect 19425 16688 19564 16690
rect 19425 16632 19430 16688
rect 19486 16632 19564 16688
rect 19425 16630 19564 16632
rect 19425 16627 19491 16630
rect 19558 16628 19564 16630
rect 19628 16628 19634 16692
rect 13537 16554 13603 16557
rect 13670 16554 13676 16556
rect 13537 16552 13676 16554
rect 13537 16496 13542 16552
rect 13598 16496 13676 16552
rect 13537 16494 13676 16496
rect 13537 16491 13603 16494
rect 13670 16492 13676 16494
rect 13740 16492 13746 16556
rect 7946 16352 8262 16353
rect 7946 16288 7952 16352
rect 8016 16288 8032 16352
rect 8096 16288 8112 16352
rect 8176 16288 8192 16352
rect 8256 16288 8262 16352
rect 7946 16287 8262 16288
rect 17946 16352 18262 16353
rect 17946 16288 17952 16352
rect 18016 16288 18032 16352
rect 18096 16288 18112 16352
rect 18176 16288 18192 16352
rect 18256 16288 18262 16352
rect 17946 16287 18262 16288
rect 17217 16284 17283 16285
rect 17166 16220 17172 16284
rect 17236 16282 17283 16284
rect 24945 16282 25011 16285
rect 26200 16282 27000 16312
rect 17236 16280 17328 16282
rect 17278 16224 17328 16280
rect 17236 16222 17328 16224
rect 24945 16280 27000 16282
rect 24945 16224 24950 16280
rect 25006 16224 27000 16280
rect 24945 16222 27000 16224
rect 17236 16220 17283 16222
rect 17217 16219 17283 16220
rect 24945 16219 25011 16222
rect 26200 16192 27000 16222
rect 2946 15808 3262 15809
rect 2946 15744 2952 15808
rect 3016 15744 3032 15808
rect 3096 15744 3112 15808
rect 3176 15744 3192 15808
rect 3256 15744 3262 15808
rect 2946 15743 3262 15744
rect 12946 15808 13262 15809
rect 12946 15744 12952 15808
rect 13016 15744 13032 15808
rect 13096 15744 13112 15808
rect 13176 15744 13192 15808
rect 13256 15744 13262 15808
rect 12946 15743 13262 15744
rect 22946 15808 23262 15809
rect 22946 15744 22952 15808
rect 23016 15744 23032 15808
rect 23096 15744 23112 15808
rect 23176 15744 23192 15808
rect 23256 15744 23262 15808
rect 22946 15743 23262 15744
rect 10225 15466 10291 15469
rect 13670 15466 13676 15468
rect 10225 15464 13676 15466
rect 10225 15408 10230 15464
rect 10286 15408 13676 15464
rect 10225 15406 13676 15408
rect 10225 15403 10291 15406
rect 13670 15404 13676 15406
rect 13740 15404 13746 15468
rect 24761 15466 24827 15469
rect 26200 15466 27000 15496
rect 24761 15464 27000 15466
rect 24761 15408 24766 15464
rect 24822 15408 27000 15464
rect 24761 15406 27000 15408
rect 24761 15403 24827 15406
rect 26200 15376 27000 15406
rect 17309 15332 17375 15333
rect 17309 15328 17356 15332
rect 17420 15330 17426 15332
rect 17309 15272 17314 15328
rect 17309 15268 17356 15272
rect 17420 15270 17466 15330
rect 17420 15268 17426 15270
rect 17309 15267 17375 15268
rect 7946 15264 8262 15265
rect 7946 15200 7952 15264
rect 8016 15200 8032 15264
rect 8096 15200 8112 15264
rect 8176 15200 8192 15264
rect 8256 15200 8262 15264
rect 7946 15199 8262 15200
rect 17946 15264 18262 15265
rect 17946 15200 17952 15264
rect 18016 15200 18032 15264
rect 18096 15200 18112 15264
rect 18176 15200 18192 15264
rect 18256 15200 18262 15264
rect 17946 15199 18262 15200
rect 13537 14922 13603 14925
rect 19977 14922 20043 14925
rect 21817 14922 21883 14925
rect 13537 14920 21883 14922
rect 13537 14864 13542 14920
rect 13598 14864 19982 14920
rect 20038 14864 21822 14920
rect 21878 14864 21883 14920
rect 13537 14862 21883 14864
rect 13537 14859 13603 14862
rect 19977 14859 20043 14862
rect 21817 14859 21883 14862
rect 2946 14720 3262 14721
rect 2946 14656 2952 14720
rect 3016 14656 3032 14720
rect 3096 14656 3112 14720
rect 3176 14656 3192 14720
rect 3256 14656 3262 14720
rect 2946 14655 3262 14656
rect 12946 14720 13262 14721
rect 12946 14656 12952 14720
rect 13016 14656 13032 14720
rect 13096 14656 13112 14720
rect 13176 14656 13192 14720
rect 13256 14656 13262 14720
rect 12946 14655 13262 14656
rect 22946 14720 23262 14721
rect 22946 14656 22952 14720
rect 23016 14656 23032 14720
rect 23096 14656 23112 14720
rect 23176 14656 23192 14720
rect 23256 14656 23262 14720
rect 22946 14655 23262 14656
rect 25129 14650 25195 14653
rect 26200 14650 27000 14680
rect 25129 14648 27000 14650
rect 25129 14592 25134 14648
rect 25190 14592 27000 14648
rect 25129 14590 27000 14592
rect 25129 14587 25195 14590
rect 26200 14560 27000 14590
rect 16021 14244 16087 14245
rect 16021 14242 16068 14244
rect 15976 14240 16068 14242
rect 15976 14184 16026 14240
rect 15976 14182 16068 14184
rect 16021 14180 16068 14182
rect 16132 14180 16138 14244
rect 16021 14179 16087 14180
rect 7946 14176 8262 14177
rect 7946 14112 7952 14176
rect 8016 14112 8032 14176
rect 8096 14112 8112 14176
rect 8176 14112 8192 14176
rect 8256 14112 8262 14176
rect 7946 14111 8262 14112
rect 17946 14176 18262 14177
rect 17946 14112 17952 14176
rect 18016 14112 18032 14176
rect 18096 14112 18112 14176
rect 18176 14112 18192 14176
rect 18256 14112 18262 14176
rect 17946 14111 18262 14112
rect 20437 14106 20503 14109
rect 26693 14106 26759 14109
rect 19290 14104 26759 14106
rect 19290 14048 20442 14104
rect 20498 14048 26698 14104
rect 26754 14048 26759 14104
rect 19290 14046 26759 14048
rect 16297 13970 16363 13973
rect 19290 13970 19350 14046
rect 20437 14043 20503 14046
rect 26693 14043 26759 14046
rect 16297 13968 19350 13970
rect 16297 13912 16302 13968
rect 16358 13912 19350 13968
rect 16297 13910 19350 13912
rect 16297 13907 16363 13910
rect 24853 13834 24919 13837
rect 26200 13834 27000 13864
rect 24853 13832 27000 13834
rect 24853 13776 24858 13832
rect 24914 13776 27000 13832
rect 24853 13774 27000 13776
rect 24853 13771 24919 13774
rect 26200 13744 27000 13774
rect 2946 13632 3262 13633
rect 2946 13568 2952 13632
rect 3016 13568 3032 13632
rect 3096 13568 3112 13632
rect 3176 13568 3192 13632
rect 3256 13568 3262 13632
rect 2946 13567 3262 13568
rect 12946 13632 13262 13633
rect 12946 13568 12952 13632
rect 13016 13568 13032 13632
rect 13096 13568 13112 13632
rect 13176 13568 13192 13632
rect 13256 13568 13262 13632
rect 12946 13567 13262 13568
rect 22946 13632 23262 13633
rect 22946 13568 22952 13632
rect 23016 13568 23032 13632
rect 23096 13568 23112 13632
rect 23176 13568 23192 13632
rect 23256 13568 23262 13632
rect 22946 13567 23262 13568
rect 19517 13292 19583 13293
rect 19517 13290 19564 13292
rect 19472 13288 19564 13290
rect 19472 13232 19522 13288
rect 19472 13230 19564 13232
rect 19517 13228 19564 13230
rect 19628 13228 19634 13292
rect 19517 13227 19583 13228
rect 15285 13154 15351 13157
rect 15653 13154 15719 13157
rect 15285 13152 15719 13154
rect 15285 13096 15290 13152
rect 15346 13096 15658 13152
rect 15714 13096 15719 13152
rect 15285 13094 15719 13096
rect 15285 13091 15351 13094
rect 15653 13091 15719 13094
rect 7946 13088 8262 13089
rect 7946 13024 7952 13088
rect 8016 13024 8032 13088
rect 8096 13024 8112 13088
rect 8176 13024 8192 13088
rect 8256 13024 8262 13088
rect 7946 13023 8262 13024
rect 17946 13088 18262 13089
rect 17946 13024 17952 13088
rect 18016 13024 18032 13088
rect 18096 13024 18112 13088
rect 18176 13024 18192 13088
rect 18256 13024 18262 13088
rect 17946 13023 18262 13024
rect 20897 13018 20963 13021
rect 22686 13018 22692 13020
rect 20897 13016 22692 13018
rect 20897 12960 20902 13016
rect 20958 12960 22692 13016
rect 20897 12958 22692 12960
rect 20897 12955 20963 12958
rect 22686 12956 22692 12958
rect 22756 12956 22762 13020
rect 24945 13018 25011 13021
rect 26200 13018 27000 13048
rect 24945 13016 27000 13018
rect 24945 12960 24950 13016
rect 25006 12960 27000 13016
rect 24945 12958 27000 12960
rect 24945 12955 25011 12958
rect 26200 12928 27000 12958
rect 16941 12882 17007 12885
rect 18638 12882 18644 12884
rect 16941 12880 18644 12882
rect 16941 12824 16946 12880
rect 17002 12824 18644 12880
rect 16941 12822 18644 12824
rect 16941 12819 17007 12822
rect 18638 12820 18644 12822
rect 18708 12820 18714 12884
rect 20345 12746 20411 12749
rect 25957 12746 26023 12749
rect 13862 12744 26023 12746
rect 13862 12688 20350 12744
rect 20406 12688 25962 12744
rect 26018 12688 26023 12744
rect 13862 12686 26023 12688
rect 13721 12610 13787 12613
rect 13862 12610 13922 12686
rect 20345 12683 20411 12686
rect 25957 12683 26023 12686
rect 13721 12608 13922 12610
rect 13721 12552 13726 12608
rect 13782 12552 13922 12608
rect 13721 12550 13922 12552
rect 20069 12612 20135 12613
rect 20069 12608 20116 12612
rect 20180 12610 20186 12612
rect 20069 12552 20074 12608
rect 13721 12547 13787 12550
rect 20069 12548 20116 12552
rect 20180 12550 20226 12610
rect 20180 12548 20186 12550
rect 20069 12547 20135 12548
rect 2946 12544 3262 12545
rect 2946 12480 2952 12544
rect 3016 12480 3032 12544
rect 3096 12480 3112 12544
rect 3176 12480 3192 12544
rect 3256 12480 3262 12544
rect 2946 12479 3262 12480
rect 12946 12544 13262 12545
rect 12946 12480 12952 12544
rect 13016 12480 13032 12544
rect 13096 12480 13112 12544
rect 13176 12480 13192 12544
rect 13256 12480 13262 12544
rect 12946 12479 13262 12480
rect 22946 12544 23262 12545
rect 22946 12480 22952 12544
rect 23016 12480 23032 12544
rect 23096 12480 23112 12544
rect 23176 12480 23192 12544
rect 23256 12480 23262 12544
rect 22946 12479 23262 12480
rect 17677 12474 17743 12477
rect 18781 12474 18847 12477
rect 17677 12472 18847 12474
rect 17677 12416 17682 12472
rect 17738 12416 18786 12472
rect 18842 12416 18847 12472
rect 17677 12414 18847 12416
rect 17677 12411 17743 12414
rect 18781 12411 18847 12414
rect 11881 12338 11947 12341
rect 12065 12338 12131 12341
rect 11881 12336 12131 12338
rect 11881 12280 11886 12336
rect 11942 12280 12070 12336
rect 12126 12280 12131 12336
rect 11881 12278 12131 12280
rect 11881 12275 11947 12278
rect 12065 12275 12131 12278
rect 14089 12338 14155 12341
rect 18413 12338 18479 12341
rect 14089 12336 18479 12338
rect 14089 12280 14094 12336
rect 14150 12280 18418 12336
rect 18474 12280 18479 12336
rect 14089 12278 18479 12280
rect 14089 12275 14155 12278
rect 18413 12275 18479 12278
rect 14825 12202 14891 12205
rect 17677 12202 17743 12205
rect 18689 12202 18755 12205
rect 14825 12200 18755 12202
rect 14825 12144 14830 12200
rect 14886 12144 17682 12200
rect 17738 12144 18694 12200
rect 18750 12144 18755 12200
rect 14825 12142 18755 12144
rect 14825 12139 14891 12142
rect 17677 12139 17743 12142
rect 18689 12139 18755 12142
rect 24945 12202 25011 12205
rect 26200 12202 27000 12232
rect 24945 12200 27000 12202
rect 24945 12144 24950 12200
rect 25006 12144 27000 12200
rect 24945 12142 27000 12144
rect 24945 12139 25011 12142
rect 26200 12112 27000 12142
rect 13537 12066 13603 12069
rect 16573 12066 16639 12069
rect 13537 12064 16639 12066
rect 13537 12008 13542 12064
rect 13598 12008 16578 12064
rect 16634 12008 16639 12064
rect 13537 12006 16639 12008
rect 13537 12003 13603 12006
rect 16573 12003 16639 12006
rect 7946 12000 8262 12001
rect 7946 11936 7952 12000
rect 8016 11936 8032 12000
rect 8096 11936 8112 12000
rect 8176 11936 8192 12000
rect 8256 11936 8262 12000
rect 7946 11935 8262 11936
rect 17946 12000 18262 12001
rect 17946 11936 17952 12000
rect 18016 11936 18032 12000
rect 18096 11936 18112 12000
rect 18176 11936 18192 12000
rect 18256 11936 18262 12000
rect 17946 11935 18262 11936
rect 12433 11930 12499 11933
rect 13721 11930 13787 11933
rect 12433 11928 13787 11930
rect 12433 11872 12438 11928
rect 12494 11872 13726 11928
rect 13782 11872 13787 11928
rect 12433 11870 13787 11872
rect 12433 11867 12499 11870
rect 13721 11867 13787 11870
rect 13353 11794 13419 11797
rect 13670 11794 13676 11796
rect 13353 11792 13676 11794
rect 13353 11736 13358 11792
rect 13414 11736 13676 11792
rect 13353 11734 13676 11736
rect 13353 11731 13419 11734
rect 13670 11732 13676 11734
rect 13740 11732 13746 11796
rect 15929 11794 15995 11797
rect 18505 11794 18571 11797
rect 15929 11792 18571 11794
rect 15929 11736 15934 11792
rect 15990 11736 18510 11792
rect 18566 11736 18571 11792
rect 15929 11734 18571 11736
rect 15929 11731 15995 11734
rect 18505 11731 18571 11734
rect 14958 11596 14964 11660
rect 15028 11658 15034 11660
rect 18505 11658 18571 11661
rect 15028 11656 18571 11658
rect 15028 11600 18510 11656
rect 18566 11600 18571 11656
rect 15028 11598 18571 11600
rect 15028 11596 15034 11598
rect 18505 11595 18571 11598
rect 16849 11522 16915 11525
rect 17217 11522 17283 11525
rect 18689 11524 18755 11525
rect 16849 11520 17283 11522
rect 16849 11464 16854 11520
rect 16910 11464 17222 11520
rect 17278 11464 17283 11520
rect 16849 11462 17283 11464
rect 16849 11459 16915 11462
rect 17217 11459 17283 11462
rect 18638 11460 18644 11524
rect 18708 11522 18755 11524
rect 18708 11520 18800 11522
rect 18750 11464 18800 11520
rect 18708 11462 18800 11464
rect 18708 11460 18755 11462
rect 18689 11459 18755 11460
rect 2946 11456 3262 11457
rect 2946 11392 2952 11456
rect 3016 11392 3032 11456
rect 3096 11392 3112 11456
rect 3176 11392 3192 11456
rect 3256 11392 3262 11456
rect 2946 11391 3262 11392
rect 12946 11456 13262 11457
rect 12946 11392 12952 11456
rect 13016 11392 13032 11456
rect 13096 11392 13112 11456
rect 13176 11392 13192 11456
rect 13256 11392 13262 11456
rect 12946 11391 13262 11392
rect 22946 11456 23262 11457
rect 22946 11392 22952 11456
rect 23016 11392 23032 11456
rect 23096 11392 23112 11456
rect 23176 11392 23192 11456
rect 23256 11392 23262 11456
rect 22946 11391 23262 11392
rect 18321 11386 18387 11389
rect 19149 11386 19215 11389
rect 18321 11384 19215 11386
rect 18321 11328 18326 11384
rect 18382 11328 19154 11384
rect 19210 11328 19215 11384
rect 18321 11326 19215 11328
rect 18321 11323 18387 11326
rect 19149 11323 19215 11326
rect 24761 11386 24827 11389
rect 26200 11386 27000 11416
rect 24761 11384 27000 11386
rect 24761 11328 24766 11384
rect 24822 11328 27000 11384
rect 24761 11326 27000 11328
rect 24761 11323 24827 11326
rect 26200 11296 27000 11326
rect 16481 11250 16547 11253
rect 17401 11250 17467 11253
rect 16481 11248 17467 11250
rect 16481 11192 16486 11248
rect 16542 11192 17406 11248
rect 17462 11192 17467 11248
rect 16481 11190 17467 11192
rect 16481 11187 16547 11190
rect 17401 11187 17467 11190
rect 15285 11114 15351 11117
rect 20805 11114 20871 11117
rect 15285 11112 20871 11114
rect 15285 11056 15290 11112
rect 15346 11056 20810 11112
rect 20866 11056 20871 11112
rect 15285 11054 20871 11056
rect 15285 11051 15351 11054
rect 20805 11051 20871 11054
rect 19057 10978 19123 10981
rect 21173 10978 21239 10981
rect 19057 10976 21239 10978
rect 19057 10920 19062 10976
rect 19118 10920 21178 10976
rect 21234 10920 21239 10976
rect 19057 10918 21239 10920
rect 19057 10915 19123 10918
rect 21173 10915 21239 10918
rect 7946 10912 8262 10913
rect 7946 10848 7952 10912
rect 8016 10848 8032 10912
rect 8096 10848 8112 10912
rect 8176 10848 8192 10912
rect 8256 10848 8262 10912
rect 7946 10847 8262 10848
rect 17946 10912 18262 10913
rect 17946 10848 17952 10912
rect 18016 10848 18032 10912
rect 18096 10848 18112 10912
rect 18176 10848 18192 10912
rect 18256 10848 18262 10912
rect 17946 10847 18262 10848
rect 11237 10842 11303 10845
rect 14641 10842 14707 10845
rect 17769 10842 17835 10845
rect 11237 10840 17835 10842
rect 11237 10784 11242 10840
rect 11298 10784 14646 10840
rect 14702 10784 17774 10840
rect 17830 10784 17835 10840
rect 11237 10782 17835 10784
rect 11237 10779 11303 10782
rect 14641 10779 14707 10782
rect 17769 10779 17835 10782
rect 10869 10706 10935 10709
rect 23933 10706 23999 10709
rect 10869 10704 23999 10706
rect 10869 10648 10874 10704
rect 10930 10648 23938 10704
rect 23994 10648 23999 10704
rect 10869 10646 23999 10648
rect 10869 10643 10935 10646
rect 23933 10643 23999 10646
rect 14917 10570 14983 10573
rect 16113 10570 16179 10573
rect 14917 10568 16179 10570
rect 14917 10512 14922 10568
rect 14978 10512 16118 10568
rect 16174 10512 16179 10568
rect 14917 10510 16179 10512
rect 14917 10507 14983 10510
rect 16113 10507 16179 10510
rect 24669 10570 24735 10573
rect 26200 10570 27000 10600
rect 24669 10568 27000 10570
rect 24669 10512 24674 10568
rect 24730 10512 27000 10568
rect 24669 10510 27000 10512
rect 24669 10507 24735 10510
rect 26200 10480 27000 10510
rect 14549 10434 14615 10437
rect 15561 10434 15627 10437
rect 14549 10432 15627 10434
rect 14549 10376 14554 10432
rect 14610 10376 15566 10432
rect 15622 10376 15627 10432
rect 14549 10374 15627 10376
rect 14549 10371 14615 10374
rect 15561 10371 15627 10374
rect 15929 10434 15995 10437
rect 16941 10434 17007 10437
rect 17769 10436 17835 10437
rect 17718 10434 17724 10436
rect 15929 10432 17007 10434
rect 15929 10376 15934 10432
rect 15990 10376 16946 10432
rect 17002 10376 17007 10432
rect 15929 10374 17007 10376
rect 17678 10374 17724 10434
rect 17788 10434 17835 10436
rect 18689 10434 18755 10437
rect 17788 10432 18755 10434
rect 17830 10376 18694 10432
rect 18750 10376 18755 10432
rect 15929 10371 15995 10374
rect 16941 10371 17007 10374
rect 17718 10372 17724 10374
rect 17788 10374 18755 10376
rect 17788 10372 17835 10374
rect 17769 10371 17835 10372
rect 18689 10371 18755 10374
rect 2946 10368 3262 10369
rect 2946 10304 2952 10368
rect 3016 10304 3032 10368
rect 3096 10304 3112 10368
rect 3176 10304 3192 10368
rect 3256 10304 3262 10368
rect 2946 10303 3262 10304
rect 12946 10368 13262 10369
rect 12946 10304 12952 10368
rect 13016 10304 13032 10368
rect 13096 10304 13112 10368
rect 13176 10304 13192 10368
rect 13256 10304 13262 10368
rect 12946 10303 13262 10304
rect 22946 10368 23262 10369
rect 22946 10304 22952 10368
rect 23016 10304 23032 10368
rect 23096 10304 23112 10368
rect 23176 10304 23192 10368
rect 23256 10304 23262 10368
rect 22946 10303 23262 10304
rect 14457 10298 14523 10301
rect 16798 10298 16804 10300
rect 14457 10296 16804 10298
rect 14457 10240 14462 10296
rect 14518 10240 16804 10296
rect 14457 10238 16804 10240
rect 14457 10235 14523 10238
rect 16798 10236 16804 10238
rect 16868 10236 16874 10300
rect 12341 10162 12407 10165
rect 22001 10162 22067 10165
rect 12341 10160 22067 10162
rect 12341 10104 12346 10160
rect 12402 10104 22006 10160
rect 22062 10104 22067 10160
rect 12341 10102 22067 10104
rect 12341 10099 12407 10102
rect 22001 10099 22067 10102
rect 8385 10026 8451 10029
rect 23013 10026 23079 10029
rect 8385 10024 23079 10026
rect 8385 9968 8390 10024
rect 8446 9968 23018 10024
rect 23074 9968 23079 10024
rect 8385 9966 23079 9968
rect 8385 9963 8451 9966
rect 23013 9963 23079 9966
rect 14089 9890 14155 9893
rect 14958 9890 14964 9892
rect 14089 9888 14964 9890
rect 14089 9832 14094 9888
rect 14150 9832 14964 9888
rect 14089 9830 14964 9832
rect 14089 9827 14155 9830
rect 14958 9828 14964 9830
rect 15028 9828 15034 9892
rect 16113 9890 16179 9893
rect 16297 9890 16363 9893
rect 16113 9888 16363 9890
rect 16113 9832 16118 9888
rect 16174 9832 16302 9888
rect 16358 9832 16363 9888
rect 16113 9830 16363 9832
rect 16113 9827 16179 9830
rect 16297 9827 16363 9830
rect 20621 9890 20687 9893
rect 24577 9890 24643 9893
rect 20621 9888 24643 9890
rect 20621 9832 20626 9888
rect 20682 9832 24582 9888
rect 24638 9832 24643 9888
rect 20621 9830 24643 9832
rect 20621 9827 20687 9830
rect 24577 9827 24643 9830
rect 7946 9824 8262 9825
rect 7946 9760 7952 9824
rect 8016 9760 8032 9824
rect 8096 9760 8112 9824
rect 8176 9760 8192 9824
rect 8256 9760 8262 9824
rect 7946 9759 8262 9760
rect 17946 9824 18262 9825
rect 17946 9760 17952 9824
rect 18016 9760 18032 9824
rect 18096 9760 18112 9824
rect 18176 9760 18192 9824
rect 18256 9760 18262 9824
rect 17946 9759 18262 9760
rect 13721 9754 13787 9757
rect 17585 9754 17651 9757
rect 13721 9752 17651 9754
rect 13721 9696 13726 9752
rect 13782 9696 17590 9752
rect 17646 9696 17651 9752
rect 13721 9694 17651 9696
rect 13721 9691 13787 9694
rect 17585 9691 17651 9694
rect 23289 9754 23355 9757
rect 26200 9754 27000 9784
rect 23289 9752 27000 9754
rect 23289 9696 23294 9752
rect 23350 9696 27000 9752
rect 23289 9694 27000 9696
rect 23289 9691 23355 9694
rect 26200 9664 27000 9694
rect 16941 9618 17007 9621
rect 19190 9618 19196 9620
rect 16941 9616 19196 9618
rect 16941 9560 16946 9616
rect 17002 9560 19196 9616
rect 16941 9558 19196 9560
rect 16941 9555 17007 9558
rect 19190 9556 19196 9558
rect 19260 9556 19266 9620
rect 12433 9482 12499 9485
rect 20161 9482 20227 9485
rect 12433 9480 20227 9482
rect 12433 9424 12438 9480
rect 12494 9424 20166 9480
rect 20222 9424 20227 9480
rect 12433 9422 20227 9424
rect 12433 9419 12499 9422
rect 20161 9419 20227 9422
rect 2946 9280 3262 9281
rect 2946 9216 2952 9280
rect 3016 9216 3032 9280
rect 3096 9216 3112 9280
rect 3176 9216 3192 9280
rect 3256 9216 3262 9280
rect 2946 9215 3262 9216
rect 12946 9280 13262 9281
rect 12946 9216 12952 9280
rect 13016 9216 13032 9280
rect 13096 9216 13112 9280
rect 13176 9216 13192 9280
rect 13256 9216 13262 9280
rect 12946 9215 13262 9216
rect 22946 9280 23262 9281
rect 22946 9216 22952 9280
rect 23016 9216 23032 9280
rect 23096 9216 23112 9280
rect 23176 9216 23192 9280
rect 23256 9216 23262 9280
rect 22946 9215 23262 9216
rect 16849 8938 16915 8941
rect 17585 8938 17651 8941
rect 18965 8938 19031 8941
rect 16849 8936 19031 8938
rect 16849 8880 16854 8936
rect 16910 8880 17590 8936
rect 17646 8880 18970 8936
rect 19026 8880 19031 8936
rect 16849 8878 19031 8880
rect 16849 8875 16915 8878
rect 17585 8875 17651 8878
rect 18965 8875 19031 8878
rect 24945 8938 25011 8941
rect 26200 8938 27000 8968
rect 24945 8936 27000 8938
rect 24945 8880 24950 8936
rect 25006 8880 27000 8936
rect 24945 8878 27000 8880
rect 24945 8875 25011 8878
rect 26200 8848 27000 8878
rect 0 8802 800 8832
rect 3325 8802 3391 8805
rect 0 8800 3391 8802
rect 0 8744 3330 8800
rect 3386 8744 3391 8800
rect 0 8742 3391 8744
rect 0 8712 800 8742
rect 3325 8739 3391 8742
rect 7946 8736 8262 8737
rect 7946 8672 7952 8736
rect 8016 8672 8032 8736
rect 8096 8672 8112 8736
rect 8176 8672 8192 8736
rect 8256 8672 8262 8736
rect 7946 8671 8262 8672
rect 17946 8736 18262 8737
rect 17946 8672 17952 8736
rect 18016 8672 18032 8736
rect 18096 8672 18112 8736
rect 18176 8672 18192 8736
rect 18256 8672 18262 8736
rect 17946 8671 18262 8672
rect 8109 8530 8175 8533
rect 20713 8530 20779 8533
rect 8109 8528 20779 8530
rect 8109 8472 8114 8528
rect 8170 8472 20718 8528
rect 20774 8472 20779 8528
rect 8109 8470 20779 8472
rect 8109 8467 8175 8470
rect 20713 8467 20779 8470
rect 11789 8394 11855 8397
rect 15929 8394 15995 8397
rect 18781 8394 18847 8397
rect 19609 8396 19675 8397
rect 19558 8394 19564 8396
rect 11789 8392 15995 8394
rect 11789 8336 11794 8392
rect 11850 8336 15934 8392
rect 15990 8336 15995 8392
rect 11789 8334 15995 8336
rect 11789 8331 11855 8334
rect 15929 8331 15995 8334
rect 16438 8392 18847 8394
rect 16438 8336 18786 8392
rect 18842 8336 18847 8392
rect 16438 8334 18847 8336
rect 19518 8334 19564 8394
rect 19628 8392 19675 8396
rect 19670 8336 19675 8392
rect 16438 8261 16498 8334
rect 18781 8331 18847 8334
rect 19558 8332 19564 8334
rect 19628 8332 19675 8336
rect 19609 8331 19675 8332
rect 16389 8256 16498 8261
rect 16389 8200 16394 8256
rect 16450 8200 16498 8256
rect 16389 8198 16498 8200
rect 16389 8195 16455 8198
rect 2946 8192 3262 8193
rect 2946 8128 2952 8192
rect 3016 8128 3032 8192
rect 3096 8128 3112 8192
rect 3176 8128 3192 8192
rect 3256 8128 3262 8192
rect 2946 8127 3262 8128
rect 12946 8192 13262 8193
rect 12946 8128 12952 8192
rect 13016 8128 13032 8192
rect 13096 8128 13112 8192
rect 13176 8128 13192 8192
rect 13256 8128 13262 8192
rect 12946 8127 13262 8128
rect 22946 8192 23262 8193
rect 22946 8128 22952 8192
rect 23016 8128 23032 8192
rect 23096 8128 23112 8192
rect 23176 8128 23192 8192
rect 23256 8128 23262 8192
rect 22946 8127 23262 8128
rect 25129 8122 25195 8125
rect 26200 8122 27000 8152
rect 25129 8120 27000 8122
rect 25129 8064 25134 8120
rect 25190 8064 27000 8120
rect 25129 8062 27000 8064
rect 25129 8059 25195 8062
rect 26200 8032 27000 8062
rect 11513 7986 11579 7989
rect 15326 7986 15332 7988
rect 11513 7984 15332 7986
rect 11513 7928 11518 7984
rect 11574 7928 15332 7984
rect 11513 7926 15332 7928
rect 11513 7923 11579 7926
rect 15326 7924 15332 7926
rect 15396 7924 15402 7988
rect 7946 7648 8262 7649
rect 7946 7584 7952 7648
rect 8016 7584 8032 7648
rect 8096 7584 8112 7648
rect 8176 7584 8192 7648
rect 8256 7584 8262 7648
rect 7946 7583 8262 7584
rect 17946 7648 18262 7649
rect 17946 7584 17952 7648
rect 18016 7584 18032 7648
rect 18096 7584 18112 7648
rect 18176 7584 18192 7648
rect 18256 7584 18262 7648
rect 17946 7583 18262 7584
rect 15326 7516 15332 7580
rect 15396 7578 15402 7580
rect 15469 7578 15535 7581
rect 15396 7576 15535 7578
rect 15396 7520 15474 7576
rect 15530 7520 15535 7576
rect 15396 7518 15535 7520
rect 15396 7516 15402 7518
rect 15469 7515 15535 7518
rect 24669 7306 24735 7309
rect 26200 7306 27000 7336
rect 24669 7304 27000 7306
rect 24669 7248 24674 7304
rect 24730 7248 27000 7304
rect 24669 7246 27000 7248
rect 24669 7243 24735 7246
rect 26200 7216 27000 7246
rect 13629 7170 13695 7173
rect 16573 7170 16639 7173
rect 13629 7168 16639 7170
rect 13629 7112 13634 7168
rect 13690 7112 16578 7168
rect 16634 7112 16639 7168
rect 13629 7110 16639 7112
rect 13629 7107 13695 7110
rect 16573 7107 16639 7110
rect 2946 7104 3262 7105
rect 2946 7040 2952 7104
rect 3016 7040 3032 7104
rect 3096 7040 3112 7104
rect 3176 7040 3192 7104
rect 3256 7040 3262 7104
rect 2946 7039 3262 7040
rect 12946 7104 13262 7105
rect 12946 7040 12952 7104
rect 13016 7040 13032 7104
rect 13096 7040 13112 7104
rect 13176 7040 13192 7104
rect 13256 7040 13262 7104
rect 12946 7039 13262 7040
rect 22946 7104 23262 7105
rect 22946 7040 22952 7104
rect 23016 7040 23032 7104
rect 23096 7040 23112 7104
rect 23176 7040 23192 7104
rect 23256 7040 23262 7104
rect 22946 7039 23262 7040
rect 23381 7036 23447 7037
rect 23381 7032 23428 7036
rect 23492 7034 23498 7036
rect 23381 6976 23386 7032
rect 23381 6972 23428 6976
rect 23492 6974 23538 7034
rect 23492 6972 23498 6974
rect 23381 6971 23447 6972
rect 10409 6762 10475 6765
rect 24577 6762 24643 6765
rect 10409 6760 24643 6762
rect 10409 6704 10414 6760
rect 10470 6704 24582 6760
rect 24638 6704 24643 6760
rect 10409 6702 24643 6704
rect 10409 6699 10475 6702
rect 24577 6699 24643 6702
rect 7946 6560 8262 6561
rect 0 6490 800 6520
rect 7946 6496 7952 6560
rect 8016 6496 8032 6560
rect 8096 6496 8112 6560
rect 8176 6496 8192 6560
rect 8256 6496 8262 6560
rect 7946 6495 8262 6496
rect 17946 6560 18262 6561
rect 17946 6496 17952 6560
rect 18016 6496 18032 6560
rect 18096 6496 18112 6560
rect 18176 6496 18192 6560
rect 18256 6496 18262 6560
rect 17946 6495 18262 6496
rect 3509 6490 3575 6493
rect 0 6488 3575 6490
rect 0 6432 3514 6488
rect 3570 6432 3575 6488
rect 0 6430 3575 6432
rect 0 6400 800 6430
rect 3509 6427 3575 6430
rect 24761 6490 24827 6493
rect 26200 6490 27000 6520
rect 24761 6488 27000 6490
rect 24761 6432 24766 6488
rect 24822 6432 27000 6488
rect 24761 6430 27000 6432
rect 24761 6427 24827 6430
rect 26200 6400 27000 6430
rect 11881 6354 11947 6357
rect 22461 6354 22527 6357
rect 11881 6352 22527 6354
rect 11881 6296 11886 6352
rect 11942 6296 22466 6352
rect 22522 6296 22527 6352
rect 11881 6294 22527 6296
rect 11881 6291 11947 6294
rect 22461 6291 22527 6294
rect 10593 6218 10659 6221
rect 22369 6218 22435 6221
rect 10593 6216 22435 6218
rect 10593 6160 10598 6216
rect 10654 6160 22374 6216
rect 22430 6160 22435 6216
rect 10593 6158 22435 6160
rect 10593 6155 10659 6158
rect 22369 6155 22435 6158
rect 2946 6016 3262 6017
rect 2946 5952 2952 6016
rect 3016 5952 3032 6016
rect 3096 5952 3112 6016
rect 3176 5952 3192 6016
rect 3256 5952 3262 6016
rect 2946 5951 3262 5952
rect 12946 6016 13262 6017
rect 12946 5952 12952 6016
rect 13016 5952 13032 6016
rect 13096 5952 13112 6016
rect 13176 5952 13192 6016
rect 13256 5952 13262 6016
rect 12946 5951 13262 5952
rect 22946 6016 23262 6017
rect 22946 5952 22952 6016
rect 23016 5952 23032 6016
rect 23096 5952 23112 6016
rect 23176 5952 23192 6016
rect 23256 5952 23262 6016
rect 22946 5951 23262 5952
rect 23289 5674 23355 5677
rect 26200 5674 27000 5704
rect 23289 5672 27000 5674
rect 23289 5616 23294 5672
rect 23350 5616 27000 5672
rect 23289 5614 27000 5616
rect 23289 5611 23355 5614
rect 26200 5584 27000 5614
rect 21357 5540 21423 5541
rect 23381 5540 23447 5541
rect 21357 5536 21404 5540
rect 21468 5538 21474 5540
rect 21357 5480 21362 5536
rect 21357 5476 21404 5480
rect 21468 5478 21514 5538
rect 23381 5536 23428 5540
rect 23492 5538 23498 5540
rect 23381 5480 23386 5536
rect 21468 5476 21474 5478
rect 23381 5476 23428 5480
rect 23492 5478 23538 5538
rect 23492 5476 23498 5478
rect 21357 5475 21423 5476
rect 23381 5475 23447 5476
rect 7946 5472 8262 5473
rect 7946 5408 7952 5472
rect 8016 5408 8032 5472
rect 8096 5408 8112 5472
rect 8176 5408 8192 5472
rect 8256 5408 8262 5472
rect 7946 5407 8262 5408
rect 17946 5472 18262 5473
rect 17946 5408 17952 5472
rect 18016 5408 18032 5472
rect 18096 5408 18112 5472
rect 18176 5408 18192 5472
rect 18256 5408 18262 5472
rect 17946 5407 18262 5408
rect 21909 5130 21975 5133
rect 21909 5128 24226 5130
rect 21909 5072 21914 5128
rect 21970 5072 24226 5128
rect 21909 5070 24226 5072
rect 21909 5067 21975 5070
rect 17125 4994 17191 4997
rect 19517 4994 19583 4997
rect 17125 4992 19583 4994
rect 17125 4936 17130 4992
rect 17186 4936 19522 4992
rect 19578 4936 19583 4992
rect 17125 4934 19583 4936
rect 17125 4931 17191 4934
rect 19517 4931 19583 4934
rect 2946 4928 3262 4929
rect 2946 4864 2952 4928
rect 3016 4864 3032 4928
rect 3096 4864 3112 4928
rect 3176 4864 3192 4928
rect 3256 4864 3262 4928
rect 2946 4863 3262 4864
rect 12946 4928 13262 4929
rect 12946 4864 12952 4928
rect 13016 4864 13032 4928
rect 13096 4864 13112 4928
rect 13176 4864 13192 4928
rect 13256 4864 13262 4928
rect 12946 4863 13262 4864
rect 22946 4928 23262 4929
rect 22946 4864 22952 4928
rect 23016 4864 23032 4928
rect 23096 4864 23112 4928
rect 23176 4864 23192 4928
rect 23256 4864 23262 4928
rect 22946 4863 23262 4864
rect 24166 4858 24226 5070
rect 26200 4858 27000 4888
rect 24166 4798 27000 4858
rect 26200 4768 27000 4798
rect 14365 4722 14431 4725
rect 16481 4722 16547 4725
rect 14365 4720 16547 4722
rect 14365 4664 14370 4720
rect 14426 4664 16486 4720
rect 16542 4664 16547 4720
rect 14365 4662 16547 4664
rect 14365 4659 14431 4662
rect 16481 4659 16547 4662
rect 9765 4586 9831 4589
rect 17401 4586 17467 4589
rect 9765 4584 17467 4586
rect 9765 4528 9770 4584
rect 9826 4528 17406 4584
rect 17462 4528 17467 4584
rect 9765 4526 17467 4528
rect 9765 4523 9831 4526
rect 17401 4523 17467 4526
rect 7946 4384 8262 4385
rect 7946 4320 7952 4384
rect 8016 4320 8032 4384
rect 8096 4320 8112 4384
rect 8176 4320 8192 4384
rect 8256 4320 8262 4384
rect 7946 4319 8262 4320
rect 17946 4384 18262 4385
rect 17946 4320 17952 4384
rect 18016 4320 18032 4384
rect 18096 4320 18112 4384
rect 18176 4320 18192 4384
rect 18256 4320 18262 4384
rect 17946 4319 18262 4320
rect 22369 4314 22435 4317
rect 22326 4312 22435 4314
rect 22326 4256 22374 4312
rect 22430 4256 22435 4312
rect 22326 4251 22435 4256
rect 0 4178 800 4208
rect 3969 4178 4035 4181
rect 0 4176 4035 4178
rect 0 4120 3974 4176
rect 4030 4120 4035 4176
rect 0 4118 4035 4120
rect 0 4088 800 4118
rect 3969 4115 4035 4118
rect 12985 4042 13051 4045
rect 22093 4044 22159 4045
rect 20110 4042 20116 4044
rect 12985 4040 20116 4042
rect 12985 3984 12990 4040
rect 13046 3984 20116 4040
rect 12985 3982 20116 3984
rect 12985 3979 13051 3982
rect 20110 3980 20116 3982
rect 20180 3980 20186 4044
rect 22093 4040 22140 4044
rect 22204 4042 22210 4044
rect 22326 4042 22386 4251
rect 26200 4042 27000 4072
rect 22093 3984 22098 4040
rect 22093 3980 22140 3984
rect 22204 3982 22250 4042
rect 22326 3982 27000 4042
rect 22204 3980 22210 3982
rect 22093 3979 22159 3980
rect 26200 3952 27000 3982
rect 2946 3840 3262 3841
rect 2946 3776 2952 3840
rect 3016 3776 3032 3840
rect 3096 3776 3112 3840
rect 3176 3776 3192 3840
rect 3256 3776 3262 3840
rect 2946 3775 3262 3776
rect 12946 3840 13262 3841
rect 12946 3776 12952 3840
rect 13016 3776 13032 3840
rect 13096 3776 13112 3840
rect 13176 3776 13192 3840
rect 13256 3776 13262 3840
rect 12946 3775 13262 3776
rect 22946 3840 23262 3841
rect 22946 3776 22952 3840
rect 23016 3776 23032 3840
rect 23096 3776 23112 3840
rect 23176 3776 23192 3840
rect 23256 3776 23262 3840
rect 22946 3775 23262 3776
rect 16297 3770 16363 3773
rect 22737 3770 22803 3773
rect 16297 3768 22803 3770
rect 16297 3712 16302 3768
rect 16358 3712 22742 3768
rect 22798 3712 22803 3768
rect 16297 3710 22803 3712
rect 16297 3707 16363 3710
rect 22737 3707 22803 3710
rect 14641 3634 14707 3637
rect 17350 3634 17356 3636
rect 14641 3632 17356 3634
rect 14641 3576 14646 3632
rect 14702 3576 17356 3632
rect 14641 3574 17356 3576
rect 14641 3571 14707 3574
rect 17350 3572 17356 3574
rect 17420 3572 17426 3636
rect 19558 3634 19564 3636
rect 17542 3574 19564 3634
rect 10593 3498 10659 3501
rect 17542 3498 17602 3574
rect 19558 3572 19564 3574
rect 19628 3572 19634 3636
rect 20345 3634 20411 3637
rect 22921 3634 22987 3637
rect 20345 3632 22987 3634
rect 20345 3576 20350 3632
rect 20406 3576 22926 3632
rect 22982 3576 22987 3632
rect 20345 3574 22987 3576
rect 20345 3571 20411 3574
rect 22921 3571 22987 3574
rect 10593 3496 17602 3498
rect 10593 3440 10598 3496
rect 10654 3440 17602 3496
rect 10593 3438 17602 3440
rect 10593 3435 10659 3438
rect 19374 3436 19380 3500
rect 19444 3498 19450 3500
rect 23933 3498 23999 3501
rect 19444 3496 23999 3498
rect 19444 3440 23938 3496
rect 23994 3440 23999 3496
rect 19444 3438 23999 3440
rect 19444 3436 19450 3438
rect 23933 3435 23999 3438
rect 7946 3296 8262 3297
rect 7946 3232 7952 3296
rect 8016 3232 8032 3296
rect 8096 3232 8112 3296
rect 8176 3232 8192 3296
rect 8256 3232 8262 3296
rect 7946 3231 8262 3232
rect 17946 3296 18262 3297
rect 17946 3232 17952 3296
rect 18016 3232 18032 3296
rect 18096 3232 18112 3296
rect 18176 3232 18192 3296
rect 18256 3232 18262 3296
rect 17946 3231 18262 3232
rect 23197 3226 23263 3229
rect 26200 3226 27000 3256
rect 23197 3224 27000 3226
rect 23197 3168 23202 3224
rect 23258 3168 27000 3224
rect 23197 3166 27000 3168
rect 23197 3163 23263 3166
rect 26200 3136 27000 3166
rect 9765 3090 9831 3093
rect 11145 3090 11211 3093
rect 9765 3088 11211 3090
rect 9765 3032 9770 3088
rect 9826 3032 11150 3088
rect 11206 3032 11211 3088
rect 9765 3030 11211 3032
rect 9765 3027 9831 3030
rect 11145 3027 11211 3030
rect 13169 3090 13235 3093
rect 13486 3090 13492 3092
rect 13169 3088 13492 3090
rect 13169 3032 13174 3088
rect 13230 3032 13492 3088
rect 13169 3030 13492 3032
rect 13169 3027 13235 3030
rect 13486 3028 13492 3030
rect 13556 3028 13562 3092
rect 17585 2954 17651 2957
rect 24853 2954 24919 2957
rect 17585 2952 24919 2954
rect 17585 2896 17590 2952
rect 17646 2896 24858 2952
rect 24914 2896 24919 2952
rect 17585 2894 24919 2896
rect 17585 2891 17651 2894
rect 24853 2891 24919 2894
rect 2946 2752 3262 2753
rect 2946 2688 2952 2752
rect 3016 2688 3032 2752
rect 3096 2688 3112 2752
rect 3176 2688 3192 2752
rect 3256 2688 3262 2752
rect 2946 2687 3262 2688
rect 12946 2752 13262 2753
rect 12946 2688 12952 2752
rect 13016 2688 13032 2752
rect 13096 2688 13112 2752
rect 13176 2688 13192 2752
rect 13256 2688 13262 2752
rect 12946 2687 13262 2688
rect 22946 2752 23262 2753
rect 22946 2688 22952 2752
rect 23016 2688 23032 2752
rect 23096 2688 23112 2752
rect 23176 2688 23192 2752
rect 23256 2688 23262 2752
rect 22946 2687 23262 2688
rect 8201 2546 8267 2549
rect 14958 2546 14964 2548
rect 8201 2544 14964 2546
rect 8201 2488 8206 2544
rect 8262 2488 14964 2544
rect 8201 2486 14964 2488
rect 8201 2483 8267 2486
rect 14958 2484 14964 2486
rect 15028 2484 15034 2548
rect 16113 2546 16179 2549
rect 21030 2546 21036 2548
rect 16113 2544 21036 2546
rect 16113 2488 16118 2544
rect 16174 2488 21036 2544
rect 16113 2486 21036 2488
rect 16113 2483 16179 2486
rect 21030 2484 21036 2486
rect 21100 2484 21106 2548
rect 7097 2410 7163 2413
rect 16062 2410 16068 2412
rect 7097 2408 16068 2410
rect 7097 2352 7102 2408
rect 7158 2352 16068 2408
rect 7097 2350 16068 2352
rect 7097 2347 7163 2350
rect 16062 2348 16068 2350
rect 16132 2348 16138 2412
rect 22093 2410 22159 2413
rect 26200 2410 27000 2440
rect 22093 2408 27000 2410
rect 22093 2352 22098 2408
rect 22154 2352 27000 2408
rect 22093 2350 27000 2352
rect 22093 2347 22159 2350
rect 26200 2320 27000 2350
rect 7946 2208 8262 2209
rect 7946 2144 7952 2208
rect 8016 2144 8032 2208
rect 8096 2144 8112 2208
rect 8176 2144 8192 2208
rect 8256 2144 8262 2208
rect 7946 2143 8262 2144
rect 17946 2208 18262 2209
rect 17946 2144 17952 2208
rect 18016 2144 18032 2208
rect 18096 2144 18112 2208
rect 18176 2144 18192 2208
rect 18256 2144 18262 2208
rect 17946 2143 18262 2144
rect 0 1866 800 1896
rect 3417 1866 3483 1869
rect 0 1864 3483 1866
rect 0 1808 3422 1864
rect 3478 1808 3483 1864
rect 0 1806 3483 1808
rect 0 1776 800 1806
rect 3417 1803 3483 1806
rect 21817 1594 21883 1597
rect 26200 1594 27000 1624
rect 21817 1592 27000 1594
rect 21817 1536 21822 1592
rect 21878 1536 27000 1592
rect 21817 1534 27000 1536
rect 21817 1531 21883 1534
rect 26200 1504 27000 1534
rect 24853 778 24919 781
rect 26200 778 27000 808
rect 24853 776 27000 778
rect 24853 720 24858 776
rect 24914 720 27000 776
rect 24853 718 27000 720
rect 24853 715 24919 718
rect 26200 688 27000 718
<< via3 >>
rect 7952 54428 8016 54432
rect 7952 54372 7956 54428
rect 7956 54372 8012 54428
rect 8012 54372 8016 54428
rect 7952 54368 8016 54372
rect 8032 54428 8096 54432
rect 8032 54372 8036 54428
rect 8036 54372 8092 54428
rect 8092 54372 8096 54428
rect 8032 54368 8096 54372
rect 8112 54428 8176 54432
rect 8112 54372 8116 54428
rect 8116 54372 8172 54428
rect 8172 54372 8176 54428
rect 8112 54368 8176 54372
rect 8192 54428 8256 54432
rect 8192 54372 8196 54428
rect 8196 54372 8252 54428
rect 8252 54372 8256 54428
rect 8192 54368 8256 54372
rect 17952 54428 18016 54432
rect 17952 54372 17956 54428
rect 17956 54372 18012 54428
rect 18012 54372 18016 54428
rect 17952 54368 18016 54372
rect 18032 54428 18096 54432
rect 18032 54372 18036 54428
rect 18036 54372 18092 54428
rect 18092 54372 18096 54428
rect 18032 54368 18096 54372
rect 18112 54428 18176 54432
rect 18112 54372 18116 54428
rect 18116 54372 18172 54428
rect 18172 54372 18176 54428
rect 18112 54368 18176 54372
rect 18192 54428 18256 54432
rect 18192 54372 18196 54428
rect 18196 54372 18252 54428
rect 18252 54372 18256 54428
rect 18192 54368 18256 54372
rect 2952 53884 3016 53888
rect 2952 53828 2956 53884
rect 2956 53828 3012 53884
rect 3012 53828 3016 53884
rect 2952 53824 3016 53828
rect 3032 53884 3096 53888
rect 3032 53828 3036 53884
rect 3036 53828 3092 53884
rect 3092 53828 3096 53884
rect 3032 53824 3096 53828
rect 3112 53884 3176 53888
rect 3112 53828 3116 53884
rect 3116 53828 3172 53884
rect 3172 53828 3176 53884
rect 3112 53824 3176 53828
rect 3192 53884 3256 53888
rect 3192 53828 3196 53884
rect 3196 53828 3252 53884
rect 3252 53828 3256 53884
rect 3192 53824 3256 53828
rect 12952 53884 13016 53888
rect 12952 53828 12956 53884
rect 12956 53828 13012 53884
rect 13012 53828 13016 53884
rect 12952 53824 13016 53828
rect 13032 53884 13096 53888
rect 13032 53828 13036 53884
rect 13036 53828 13092 53884
rect 13092 53828 13096 53884
rect 13032 53824 13096 53828
rect 13112 53884 13176 53888
rect 13112 53828 13116 53884
rect 13116 53828 13172 53884
rect 13172 53828 13176 53884
rect 13112 53824 13176 53828
rect 13192 53884 13256 53888
rect 13192 53828 13196 53884
rect 13196 53828 13252 53884
rect 13252 53828 13256 53884
rect 13192 53824 13256 53828
rect 22952 53884 23016 53888
rect 22952 53828 22956 53884
rect 22956 53828 23012 53884
rect 23012 53828 23016 53884
rect 22952 53824 23016 53828
rect 23032 53884 23096 53888
rect 23032 53828 23036 53884
rect 23036 53828 23092 53884
rect 23092 53828 23096 53884
rect 23032 53824 23096 53828
rect 23112 53884 23176 53888
rect 23112 53828 23116 53884
rect 23116 53828 23172 53884
rect 23172 53828 23176 53884
rect 23112 53824 23176 53828
rect 23192 53884 23256 53888
rect 23192 53828 23196 53884
rect 23196 53828 23252 53884
rect 23252 53828 23256 53884
rect 23192 53824 23256 53828
rect 7952 53340 8016 53344
rect 7952 53284 7956 53340
rect 7956 53284 8012 53340
rect 8012 53284 8016 53340
rect 7952 53280 8016 53284
rect 8032 53340 8096 53344
rect 8032 53284 8036 53340
rect 8036 53284 8092 53340
rect 8092 53284 8096 53340
rect 8032 53280 8096 53284
rect 8112 53340 8176 53344
rect 8112 53284 8116 53340
rect 8116 53284 8172 53340
rect 8172 53284 8176 53340
rect 8112 53280 8176 53284
rect 8192 53340 8256 53344
rect 8192 53284 8196 53340
rect 8196 53284 8252 53340
rect 8252 53284 8256 53340
rect 8192 53280 8256 53284
rect 17952 53340 18016 53344
rect 17952 53284 17956 53340
rect 17956 53284 18012 53340
rect 18012 53284 18016 53340
rect 17952 53280 18016 53284
rect 18032 53340 18096 53344
rect 18032 53284 18036 53340
rect 18036 53284 18092 53340
rect 18092 53284 18096 53340
rect 18032 53280 18096 53284
rect 18112 53340 18176 53344
rect 18112 53284 18116 53340
rect 18116 53284 18172 53340
rect 18172 53284 18176 53340
rect 18112 53280 18176 53284
rect 18192 53340 18256 53344
rect 18192 53284 18196 53340
rect 18196 53284 18252 53340
rect 18252 53284 18256 53340
rect 18192 53280 18256 53284
rect 2952 52796 3016 52800
rect 2952 52740 2956 52796
rect 2956 52740 3012 52796
rect 3012 52740 3016 52796
rect 2952 52736 3016 52740
rect 3032 52796 3096 52800
rect 3032 52740 3036 52796
rect 3036 52740 3092 52796
rect 3092 52740 3096 52796
rect 3032 52736 3096 52740
rect 3112 52796 3176 52800
rect 3112 52740 3116 52796
rect 3116 52740 3172 52796
rect 3172 52740 3176 52796
rect 3112 52736 3176 52740
rect 3192 52796 3256 52800
rect 3192 52740 3196 52796
rect 3196 52740 3252 52796
rect 3252 52740 3256 52796
rect 3192 52736 3256 52740
rect 12952 52796 13016 52800
rect 12952 52740 12956 52796
rect 12956 52740 13012 52796
rect 13012 52740 13016 52796
rect 12952 52736 13016 52740
rect 13032 52796 13096 52800
rect 13032 52740 13036 52796
rect 13036 52740 13092 52796
rect 13092 52740 13096 52796
rect 13032 52736 13096 52740
rect 13112 52796 13176 52800
rect 13112 52740 13116 52796
rect 13116 52740 13172 52796
rect 13172 52740 13176 52796
rect 13112 52736 13176 52740
rect 13192 52796 13256 52800
rect 13192 52740 13196 52796
rect 13196 52740 13252 52796
rect 13252 52740 13256 52796
rect 13192 52736 13256 52740
rect 22952 52796 23016 52800
rect 22952 52740 22956 52796
rect 22956 52740 23012 52796
rect 23012 52740 23016 52796
rect 22952 52736 23016 52740
rect 23032 52796 23096 52800
rect 23032 52740 23036 52796
rect 23036 52740 23092 52796
rect 23092 52740 23096 52796
rect 23032 52736 23096 52740
rect 23112 52796 23176 52800
rect 23112 52740 23116 52796
rect 23116 52740 23172 52796
rect 23172 52740 23176 52796
rect 23112 52736 23176 52740
rect 23192 52796 23256 52800
rect 23192 52740 23196 52796
rect 23196 52740 23252 52796
rect 23252 52740 23256 52796
rect 23192 52736 23256 52740
rect 7952 52252 8016 52256
rect 7952 52196 7956 52252
rect 7956 52196 8012 52252
rect 8012 52196 8016 52252
rect 7952 52192 8016 52196
rect 8032 52252 8096 52256
rect 8032 52196 8036 52252
rect 8036 52196 8092 52252
rect 8092 52196 8096 52252
rect 8032 52192 8096 52196
rect 8112 52252 8176 52256
rect 8112 52196 8116 52252
rect 8116 52196 8172 52252
rect 8172 52196 8176 52252
rect 8112 52192 8176 52196
rect 8192 52252 8256 52256
rect 8192 52196 8196 52252
rect 8196 52196 8252 52252
rect 8252 52196 8256 52252
rect 8192 52192 8256 52196
rect 17952 52252 18016 52256
rect 17952 52196 17956 52252
rect 17956 52196 18012 52252
rect 18012 52196 18016 52252
rect 17952 52192 18016 52196
rect 18032 52252 18096 52256
rect 18032 52196 18036 52252
rect 18036 52196 18092 52252
rect 18092 52196 18096 52252
rect 18032 52192 18096 52196
rect 18112 52252 18176 52256
rect 18112 52196 18116 52252
rect 18116 52196 18172 52252
rect 18172 52196 18176 52252
rect 18112 52192 18176 52196
rect 18192 52252 18256 52256
rect 18192 52196 18196 52252
rect 18196 52196 18252 52252
rect 18252 52196 18256 52252
rect 18192 52192 18256 52196
rect 2952 51708 3016 51712
rect 2952 51652 2956 51708
rect 2956 51652 3012 51708
rect 3012 51652 3016 51708
rect 2952 51648 3016 51652
rect 3032 51708 3096 51712
rect 3032 51652 3036 51708
rect 3036 51652 3092 51708
rect 3092 51652 3096 51708
rect 3032 51648 3096 51652
rect 3112 51708 3176 51712
rect 3112 51652 3116 51708
rect 3116 51652 3172 51708
rect 3172 51652 3176 51708
rect 3112 51648 3176 51652
rect 3192 51708 3256 51712
rect 3192 51652 3196 51708
rect 3196 51652 3252 51708
rect 3252 51652 3256 51708
rect 3192 51648 3256 51652
rect 12952 51708 13016 51712
rect 12952 51652 12956 51708
rect 12956 51652 13012 51708
rect 13012 51652 13016 51708
rect 12952 51648 13016 51652
rect 13032 51708 13096 51712
rect 13032 51652 13036 51708
rect 13036 51652 13092 51708
rect 13092 51652 13096 51708
rect 13032 51648 13096 51652
rect 13112 51708 13176 51712
rect 13112 51652 13116 51708
rect 13116 51652 13172 51708
rect 13172 51652 13176 51708
rect 13112 51648 13176 51652
rect 13192 51708 13256 51712
rect 13192 51652 13196 51708
rect 13196 51652 13252 51708
rect 13252 51652 13256 51708
rect 13192 51648 13256 51652
rect 22952 51708 23016 51712
rect 22952 51652 22956 51708
rect 22956 51652 23012 51708
rect 23012 51652 23016 51708
rect 22952 51648 23016 51652
rect 23032 51708 23096 51712
rect 23032 51652 23036 51708
rect 23036 51652 23092 51708
rect 23092 51652 23096 51708
rect 23032 51648 23096 51652
rect 23112 51708 23176 51712
rect 23112 51652 23116 51708
rect 23116 51652 23172 51708
rect 23172 51652 23176 51708
rect 23112 51648 23176 51652
rect 23192 51708 23256 51712
rect 23192 51652 23196 51708
rect 23196 51652 23252 51708
rect 23252 51652 23256 51708
rect 23192 51648 23256 51652
rect 7952 51164 8016 51168
rect 7952 51108 7956 51164
rect 7956 51108 8012 51164
rect 8012 51108 8016 51164
rect 7952 51104 8016 51108
rect 8032 51164 8096 51168
rect 8032 51108 8036 51164
rect 8036 51108 8092 51164
rect 8092 51108 8096 51164
rect 8032 51104 8096 51108
rect 8112 51164 8176 51168
rect 8112 51108 8116 51164
rect 8116 51108 8172 51164
rect 8172 51108 8176 51164
rect 8112 51104 8176 51108
rect 8192 51164 8256 51168
rect 8192 51108 8196 51164
rect 8196 51108 8252 51164
rect 8252 51108 8256 51164
rect 8192 51104 8256 51108
rect 17952 51164 18016 51168
rect 17952 51108 17956 51164
rect 17956 51108 18012 51164
rect 18012 51108 18016 51164
rect 17952 51104 18016 51108
rect 18032 51164 18096 51168
rect 18032 51108 18036 51164
rect 18036 51108 18092 51164
rect 18092 51108 18096 51164
rect 18032 51104 18096 51108
rect 18112 51164 18176 51168
rect 18112 51108 18116 51164
rect 18116 51108 18172 51164
rect 18172 51108 18176 51164
rect 18112 51104 18176 51108
rect 18192 51164 18256 51168
rect 18192 51108 18196 51164
rect 18196 51108 18252 51164
rect 18252 51108 18256 51164
rect 18192 51104 18256 51108
rect 2952 50620 3016 50624
rect 2952 50564 2956 50620
rect 2956 50564 3012 50620
rect 3012 50564 3016 50620
rect 2952 50560 3016 50564
rect 3032 50620 3096 50624
rect 3032 50564 3036 50620
rect 3036 50564 3092 50620
rect 3092 50564 3096 50620
rect 3032 50560 3096 50564
rect 3112 50620 3176 50624
rect 3112 50564 3116 50620
rect 3116 50564 3172 50620
rect 3172 50564 3176 50620
rect 3112 50560 3176 50564
rect 3192 50620 3256 50624
rect 3192 50564 3196 50620
rect 3196 50564 3252 50620
rect 3252 50564 3256 50620
rect 3192 50560 3256 50564
rect 12952 50620 13016 50624
rect 12952 50564 12956 50620
rect 12956 50564 13012 50620
rect 13012 50564 13016 50620
rect 12952 50560 13016 50564
rect 13032 50620 13096 50624
rect 13032 50564 13036 50620
rect 13036 50564 13092 50620
rect 13092 50564 13096 50620
rect 13032 50560 13096 50564
rect 13112 50620 13176 50624
rect 13112 50564 13116 50620
rect 13116 50564 13172 50620
rect 13172 50564 13176 50620
rect 13112 50560 13176 50564
rect 13192 50620 13256 50624
rect 13192 50564 13196 50620
rect 13196 50564 13252 50620
rect 13252 50564 13256 50620
rect 13192 50560 13256 50564
rect 22952 50620 23016 50624
rect 22952 50564 22956 50620
rect 22956 50564 23012 50620
rect 23012 50564 23016 50620
rect 22952 50560 23016 50564
rect 23032 50620 23096 50624
rect 23032 50564 23036 50620
rect 23036 50564 23092 50620
rect 23092 50564 23096 50620
rect 23032 50560 23096 50564
rect 23112 50620 23176 50624
rect 23112 50564 23116 50620
rect 23116 50564 23172 50620
rect 23172 50564 23176 50620
rect 23112 50560 23176 50564
rect 23192 50620 23256 50624
rect 23192 50564 23196 50620
rect 23196 50564 23252 50620
rect 23252 50564 23256 50620
rect 23192 50560 23256 50564
rect 7952 50076 8016 50080
rect 7952 50020 7956 50076
rect 7956 50020 8012 50076
rect 8012 50020 8016 50076
rect 7952 50016 8016 50020
rect 8032 50076 8096 50080
rect 8032 50020 8036 50076
rect 8036 50020 8092 50076
rect 8092 50020 8096 50076
rect 8032 50016 8096 50020
rect 8112 50076 8176 50080
rect 8112 50020 8116 50076
rect 8116 50020 8172 50076
rect 8172 50020 8176 50076
rect 8112 50016 8176 50020
rect 8192 50076 8256 50080
rect 8192 50020 8196 50076
rect 8196 50020 8252 50076
rect 8252 50020 8256 50076
rect 8192 50016 8256 50020
rect 17952 50076 18016 50080
rect 17952 50020 17956 50076
rect 17956 50020 18012 50076
rect 18012 50020 18016 50076
rect 17952 50016 18016 50020
rect 18032 50076 18096 50080
rect 18032 50020 18036 50076
rect 18036 50020 18092 50076
rect 18092 50020 18096 50076
rect 18032 50016 18096 50020
rect 18112 50076 18176 50080
rect 18112 50020 18116 50076
rect 18116 50020 18172 50076
rect 18172 50020 18176 50076
rect 18112 50016 18176 50020
rect 18192 50076 18256 50080
rect 18192 50020 18196 50076
rect 18196 50020 18252 50076
rect 18252 50020 18256 50076
rect 18192 50016 18256 50020
rect 2952 49532 3016 49536
rect 2952 49476 2956 49532
rect 2956 49476 3012 49532
rect 3012 49476 3016 49532
rect 2952 49472 3016 49476
rect 3032 49532 3096 49536
rect 3032 49476 3036 49532
rect 3036 49476 3092 49532
rect 3092 49476 3096 49532
rect 3032 49472 3096 49476
rect 3112 49532 3176 49536
rect 3112 49476 3116 49532
rect 3116 49476 3172 49532
rect 3172 49476 3176 49532
rect 3112 49472 3176 49476
rect 3192 49532 3256 49536
rect 3192 49476 3196 49532
rect 3196 49476 3252 49532
rect 3252 49476 3256 49532
rect 3192 49472 3256 49476
rect 12952 49532 13016 49536
rect 12952 49476 12956 49532
rect 12956 49476 13012 49532
rect 13012 49476 13016 49532
rect 12952 49472 13016 49476
rect 13032 49532 13096 49536
rect 13032 49476 13036 49532
rect 13036 49476 13092 49532
rect 13092 49476 13096 49532
rect 13032 49472 13096 49476
rect 13112 49532 13176 49536
rect 13112 49476 13116 49532
rect 13116 49476 13172 49532
rect 13172 49476 13176 49532
rect 13112 49472 13176 49476
rect 13192 49532 13256 49536
rect 13192 49476 13196 49532
rect 13196 49476 13252 49532
rect 13252 49476 13256 49532
rect 13192 49472 13256 49476
rect 22952 49532 23016 49536
rect 22952 49476 22956 49532
rect 22956 49476 23012 49532
rect 23012 49476 23016 49532
rect 22952 49472 23016 49476
rect 23032 49532 23096 49536
rect 23032 49476 23036 49532
rect 23036 49476 23092 49532
rect 23092 49476 23096 49532
rect 23032 49472 23096 49476
rect 23112 49532 23176 49536
rect 23112 49476 23116 49532
rect 23116 49476 23172 49532
rect 23172 49476 23176 49532
rect 23112 49472 23176 49476
rect 23192 49532 23256 49536
rect 23192 49476 23196 49532
rect 23196 49476 23252 49532
rect 23252 49476 23256 49532
rect 23192 49472 23256 49476
rect 7952 48988 8016 48992
rect 7952 48932 7956 48988
rect 7956 48932 8012 48988
rect 8012 48932 8016 48988
rect 7952 48928 8016 48932
rect 8032 48988 8096 48992
rect 8032 48932 8036 48988
rect 8036 48932 8092 48988
rect 8092 48932 8096 48988
rect 8032 48928 8096 48932
rect 8112 48988 8176 48992
rect 8112 48932 8116 48988
rect 8116 48932 8172 48988
rect 8172 48932 8176 48988
rect 8112 48928 8176 48932
rect 8192 48988 8256 48992
rect 8192 48932 8196 48988
rect 8196 48932 8252 48988
rect 8252 48932 8256 48988
rect 8192 48928 8256 48932
rect 17952 48988 18016 48992
rect 17952 48932 17956 48988
rect 17956 48932 18012 48988
rect 18012 48932 18016 48988
rect 17952 48928 18016 48932
rect 18032 48988 18096 48992
rect 18032 48932 18036 48988
rect 18036 48932 18092 48988
rect 18092 48932 18096 48988
rect 18032 48928 18096 48932
rect 18112 48988 18176 48992
rect 18112 48932 18116 48988
rect 18116 48932 18172 48988
rect 18172 48932 18176 48988
rect 18112 48928 18176 48932
rect 18192 48988 18256 48992
rect 18192 48932 18196 48988
rect 18196 48932 18252 48988
rect 18252 48932 18256 48988
rect 18192 48928 18256 48932
rect 2952 48444 3016 48448
rect 2952 48388 2956 48444
rect 2956 48388 3012 48444
rect 3012 48388 3016 48444
rect 2952 48384 3016 48388
rect 3032 48444 3096 48448
rect 3032 48388 3036 48444
rect 3036 48388 3092 48444
rect 3092 48388 3096 48444
rect 3032 48384 3096 48388
rect 3112 48444 3176 48448
rect 3112 48388 3116 48444
rect 3116 48388 3172 48444
rect 3172 48388 3176 48444
rect 3112 48384 3176 48388
rect 3192 48444 3256 48448
rect 3192 48388 3196 48444
rect 3196 48388 3252 48444
rect 3252 48388 3256 48444
rect 3192 48384 3256 48388
rect 12952 48444 13016 48448
rect 12952 48388 12956 48444
rect 12956 48388 13012 48444
rect 13012 48388 13016 48444
rect 12952 48384 13016 48388
rect 13032 48444 13096 48448
rect 13032 48388 13036 48444
rect 13036 48388 13092 48444
rect 13092 48388 13096 48444
rect 13032 48384 13096 48388
rect 13112 48444 13176 48448
rect 13112 48388 13116 48444
rect 13116 48388 13172 48444
rect 13172 48388 13176 48444
rect 13112 48384 13176 48388
rect 13192 48444 13256 48448
rect 13192 48388 13196 48444
rect 13196 48388 13252 48444
rect 13252 48388 13256 48444
rect 13192 48384 13256 48388
rect 22952 48444 23016 48448
rect 22952 48388 22956 48444
rect 22956 48388 23012 48444
rect 23012 48388 23016 48444
rect 22952 48384 23016 48388
rect 23032 48444 23096 48448
rect 23032 48388 23036 48444
rect 23036 48388 23092 48444
rect 23092 48388 23096 48444
rect 23032 48384 23096 48388
rect 23112 48444 23176 48448
rect 23112 48388 23116 48444
rect 23116 48388 23172 48444
rect 23172 48388 23176 48444
rect 23112 48384 23176 48388
rect 23192 48444 23256 48448
rect 23192 48388 23196 48444
rect 23196 48388 23252 48444
rect 23252 48388 23256 48444
rect 23192 48384 23256 48388
rect 7952 47900 8016 47904
rect 7952 47844 7956 47900
rect 7956 47844 8012 47900
rect 8012 47844 8016 47900
rect 7952 47840 8016 47844
rect 8032 47900 8096 47904
rect 8032 47844 8036 47900
rect 8036 47844 8092 47900
rect 8092 47844 8096 47900
rect 8032 47840 8096 47844
rect 8112 47900 8176 47904
rect 8112 47844 8116 47900
rect 8116 47844 8172 47900
rect 8172 47844 8176 47900
rect 8112 47840 8176 47844
rect 8192 47900 8256 47904
rect 8192 47844 8196 47900
rect 8196 47844 8252 47900
rect 8252 47844 8256 47900
rect 8192 47840 8256 47844
rect 17952 47900 18016 47904
rect 17952 47844 17956 47900
rect 17956 47844 18012 47900
rect 18012 47844 18016 47900
rect 17952 47840 18016 47844
rect 18032 47900 18096 47904
rect 18032 47844 18036 47900
rect 18036 47844 18092 47900
rect 18092 47844 18096 47900
rect 18032 47840 18096 47844
rect 18112 47900 18176 47904
rect 18112 47844 18116 47900
rect 18116 47844 18172 47900
rect 18172 47844 18176 47900
rect 18112 47840 18176 47844
rect 18192 47900 18256 47904
rect 18192 47844 18196 47900
rect 18196 47844 18252 47900
rect 18252 47844 18256 47900
rect 18192 47840 18256 47844
rect 2952 47356 3016 47360
rect 2952 47300 2956 47356
rect 2956 47300 3012 47356
rect 3012 47300 3016 47356
rect 2952 47296 3016 47300
rect 3032 47356 3096 47360
rect 3032 47300 3036 47356
rect 3036 47300 3092 47356
rect 3092 47300 3096 47356
rect 3032 47296 3096 47300
rect 3112 47356 3176 47360
rect 3112 47300 3116 47356
rect 3116 47300 3172 47356
rect 3172 47300 3176 47356
rect 3112 47296 3176 47300
rect 3192 47356 3256 47360
rect 3192 47300 3196 47356
rect 3196 47300 3252 47356
rect 3252 47300 3256 47356
rect 3192 47296 3256 47300
rect 12952 47356 13016 47360
rect 12952 47300 12956 47356
rect 12956 47300 13012 47356
rect 13012 47300 13016 47356
rect 12952 47296 13016 47300
rect 13032 47356 13096 47360
rect 13032 47300 13036 47356
rect 13036 47300 13092 47356
rect 13092 47300 13096 47356
rect 13032 47296 13096 47300
rect 13112 47356 13176 47360
rect 13112 47300 13116 47356
rect 13116 47300 13172 47356
rect 13172 47300 13176 47356
rect 13112 47296 13176 47300
rect 13192 47356 13256 47360
rect 13192 47300 13196 47356
rect 13196 47300 13252 47356
rect 13252 47300 13256 47356
rect 13192 47296 13256 47300
rect 22952 47356 23016 47360
rect 22952 47300 22956 47356
rect 22956 47300 23012 47356
rect 23012 47300 23016 47356
rect 22952 47296 23016 47300
rect 23032 47356 23096 47360
rect 23032 47300 23036 47356
rect 23036 47300 23092 47356
rect 23092 47300 23096 47356
rect 23032 47296 23096 47300
rect 23112 47356 23176 47360
rect 23112 47300 23116 47356
rect 23116 47300 23172 47356
rect 23172 47300 23176 47356
rect 23112 47296 23176 47300
rect 23192 47356 23256 47360
rect 23192 47300 23196 47356
rect 23196 47300 23252 47356
rect 23252 47300 23256 47356
rect 23192 47296 23256 47300
rect 7952 46812 8016 46816
rect 7952 46756 7956 46812
rect 7956 46756 8012 46812
rect 8012 46756 8016 46812
rect 7952 46752 8016 46756
rect 8032 46812 8096 46816
rect 8032 46756 8036 46812
rect 8036 46756 8092 46812
rect 8092 46756 8096 46812
rect 8032 46752 8096 46756
rect 8112 46812 8176 46816
rect 8112 46756 8116 46812
rect 8116 46756 8172 46812
rect 8172 46756 8176 46812
rect 8112 46752 8176 46756
rect 8192 46812 8256 46816
rect 8192 46756 8196 46812
rect 8196 46756 8252 46812
rect 8252 46756 8256 46812
rect 8192 46752 8256 46756
rect 17952 46812 18016 46816
rect 17952 46756 17956 46812
rect 17956 46756 18012 46812
rect 18012 46756 18016 46812
rect 17952 46752 18016 46756
rect 18032 46812 18096 46816
rect 18032 46756 18036 46812
rect 18036 46756 18092 46812
rect 18092 46756 18096 46812
rect 18032 46752 18096 46756
rect 18112 46812 18176 46816
rect 18112 46756 18116 46812
rect 18116 46756 18172 46812
rect 18172 46756 18176 46812
rect 18112 46752 18176 46756
rect 18192 46812 18256 46816
rect 18192 46756 18196 46812
rect 18196 46756 18252 46812
rect 18252 46756 18256 46812
rect 18192 46752 18256 46756
rect 2952 46268 3016 46272
rect 2952 46212 2956 46268
rect 2956 46212 3012 46268
rect 3012 46212 3016 46268
rect 2952 46208 3016 46212
rect 3032 46268 3096 46272
rect 3032 46212 3036 46268
rect 3036 46212 3092 46268
rect 3092 46212 3096 46268
rect 3032 46208 3096 46212
rect 3112 46268 3176 46272
rect 3112 46212 3116 46268
rect 3116 46212 3172 46268
rect 3172 46212 3176 46268
rect 3112 46208 3176 46212
rect 3192 46268 3256 46272
rect 3192 46212 3196 46268
rect 3196 46212 3252 46268
rect 3252 46212 3256 46268
rect 3192 46208 3256 46212
rect 12952 46268 13016 46272
rect 12952 46212 12956 46268
rect 12956 46212 13012 46268
rect 13012 46212 13016 46268
rect 12952 46208 13016 46212
rect 13032 46268 13096 46272
rect 13032 46212 13036 46268
rect 13036 46212 13092 46268
rect 13092 46212 13096 46268
rect 13032 46208 13096 46212
rect 13112 46268 13176 46272
rect 13112 46212 13116 46268
rect 13116 46212 13172 46268
rect 13172 46212 13176 46268
rect 13112 46208 13176 46212
rect 13192 46268 13256 46272
rect 13192 46212 13196 46268
rect 13196 46212 13252 46268
rect 13252 46212 13256 46268
rect 13192 46208 13256 46212
rect 22952 46268 23016 46272
rect 22952 46212 22956 46268
rect 22956 46212 23012 46268
rect 23012 46212 23016 46268
rect 22952 46208 23016 46212
rect 23032 46268 23096 46272
rect 23032 46212 23036 46268
rect 23036 46212 23092 46268
rect 23092 46212 23096 46268
rect 23032 46208 23096 46212
rect 23112 46268 23176 46272
rect 23112 46212 23116 46268
rect 23116 46212 23172 46268
rect 23172 46212 23176 46268
rect 23112 46208 23176 46212
rect 23192 46268 23256 46272
rect 23192 46212 23196 46268
rect 23196 46212 23252 46268
rect 23252 46212 23256 46268
rect 23192 46208 23256 46212
rect 7952 45724 8016 45728
rect 7952 45668 7956 45724
rect 7956 45668 8012 45724
rect 8012 45668 8016 45724
rect 7952 45664 8016 45668
rect 8032 45724 8096 45728
rect 8032 45668 8036 45724
rect 8036 45668 8092 45724
rect 8092 45668 8096 45724
rect 8032 45664 8096 45668
rect 8112 45724 8176 45728
rect 8112 45668 8116 45724
rect 8116 45668 8172 45724
rect 8172 45668 8176 45724
rect 8112 45664 8176 45668
rect 8192 45724 8256 45728
rect 8192 45668 8196 45724
rect 8196 45668 8252 45724
rect 8252 45668 8256 45724
rect 8192 45664 8256 45668
rect 17952 45724 18016 45728
rect 17952 45668 17956 45724
rect 17956 45668 18012 45724
rect 18012 45668 18016 45724
rect 17952 45664 18016 45668
rect 18032 45724 18096 45728
rect 18032 45668 18036 45724
rect 18036 45668 18092 45724
rect 18092 45668 18096 45724
rect 18032 45664 18096 45668
rect 18112 45724 18176 45728
rect 18112 45668 18116 45724
rect 18116 45668 18172 45724
rect 18172 45668 18176 45724
rect 18112 45664 18176 45668
rect 18192 45724 18256 45728
rect 18192 45668 18196 45724
rect 18196 45668 18252 45724
rect 18252 45668 18256 45724
rect 18192 45664 18256 45668
rect 2952 45180 3016 45184
rect 2952 45124 2956 45180
rect 2956 45124 3012 45180
rect 3012 45124 3016 45180
rect 2952 45120 3016 45124
rect 3032 45180 3096 45184
rect 3032 45124 3036 45180
rect 3036 45124 3092 45180
rect 3092 45124 3096 45180
rect 3032 45120 3096 45124
rect 3112 45180 3176 45184
rect 3112 45124 3116 45180
rect 3116 45124 3172 45180
rect 3172 45124 3176 45180
rect 3112 45120 3176 45124
rect 3192 45180 3256 45184
rect 3192 45124 3196 45180
rect 3196 45124 3252 45180
rect 3252 45124 3256 45180
rect 3192 45120 3256 45124
rect 12952 45180 13016 45184
rect 12952 45124 12956 45180
rect 12956 45124 13012 45180
rect 13012 45124 13016 45180
rect 12952 45120 13016 45124
rect 13032 45180 13096 45184
rect 13032 45124 13036 45180
rect 13036 45124 13092 45180
rect 13092 45124 13096 45180
rect 13032 45120 13096 45124
rect 13112 45180 13176 45184
rect 13112 45124 13116 45180
rect 13116 45124 13172 45180
rect 13172 45124 13176 45180
rect 13112 45120 13176 45124
rect 13192 45180 13256 45184
rect 13192 45124 13196 45180
rect 13196 45124 13252 45180
rect 13252 45124 13256 45180
rect 13192 45120 13256 45124
rect 22952 45180 23016 45184
rect 22952 45124 22956 45180
rect 22956 45124 23012 45180
rect 23012 45124 23016 45180
rect 22952 45120 23016 45124
rect 23032 45180 23096 45184
rect 23032 45124 23036 45180
rect 23036 45124 23092 45180
rect 23092 45124 23096 45180
rect 23032 45120 23096 45124
rect 23112 45180 23176 45184
rect 23112 45124 23116 45180
rect 23116 45124 23172 45180
rect 23172 45124 23176 45180
rect 23112 45120 23176 45124
rect 23192 45180 23256 45184
rect 23192 45124 23196 45180
rect 23196 45124 23252 45180
rect 23252 45124 23256 45180
rect 23192 45120 23256 45124
rect 7952 44636 8016 44640
rect 7952 44580 7956 44636
rect 7956 44580 8012 44636
rect 8012 44580 8016 44636
rect 7952 44576 8016 44580
rect 8032 44636 8096 44640
rect 8032 44580 8036 44636
rect 8036 44580 8092 44636
rect 8092 44580 8096 44636
rect 8032 44576 8096 44580
rect 8112 44636 8176 44640
rect 8112 44580 8116 44636
rect 8116 44580 8172 44636
rect 8172 44580 8176 44636
rect 8112 44576 8176 44580
rect 8192 44636 8256 44640
rect 8192 44580 8196 44636
rect 8196 44580 8252 44636
rect 8252 44580 8256 44636
rect 8192 44576 8256 44580
rect 17952 44636 18016 44640
rect 17952 44580 17956 44636
rect 17956 44580 18012 44636
rect 18012 44580 18016 44636
rect 17952 44576 18016 44580
rect 18032 44636 18096 44640
rect 18032 44580 18036 44636
rect 18036 44580 18092 44636
rect 18092 44580 18096 44636
rect 18032 44576 18096 44580
rect 18112 44636 18176 44640
rect 18112 44580 18116 44636
rect 18116 44580 18172 44636
rect 18172 44580 18176 44636
rect 18112 44576 18176 44580
rect 18192 44636 18256 44640
rect 18192 44580 18196 44636
rect 18196 44580 18252 44636
rect 18252 44580 18256 44636
rect 18192 44576 18256 44580
rect 2952 44092 3016 44096
rect 2952 44036 2956 44092
rect 2956 44036 3012 44092
rect 3012 44036 3016 44092
rect 2952 44032 3016 44036
rect 3032 44092 3096 44096
rect 3032 44036 3036 44092
rect 3036 44036 3092 44092
rect 3092 44036 3096 44092
rect 3032 44032 3096 44036
rect 3112 44092 3176 44096
rect 3112 44036 3116 44092
rect 3116 44036 3172 44092
rect 3172 44036 3176 44092
rect 3112 44032 3176 44036
rect 3192 44092 3256 44096
rect 3192 44036 3196 44092
rect 3196 44036 3252 44092
rect 3252 44036 3256 44092
rect 3192 44032 3256 44036
rect 12952 44092 13016 44096
rect 12952 44036 12956 44092
rect 12956 44036 13012 44092
rect 13012 44036 13016 44092
rect 12952 44032 13016 44036
rect 13032 44092 13096 44096
rect 13032 44036 13036 44092
rect 13036 44036 13092 44092
rect 13092 44036 13096 44092
rect 13032 44032 13096 44036
rect 13112 44092 13176 44096
rect 13112 44036 13116 44092
rect 13116 44036 13172 44092
rect 13172 44036 13176 44092
rect 13112 44032 13176 44036
rect 13192 44092 13256 44096
rect 13192 44036 13196 44092
rect 13196 44036 13252 44092
rect 13252 44036 13256 44092
rect 13192 44032 13256 44036
rect 22952 44092 23016 44096
rect 22952 44036 22956 44092
rect 22956 44036 23012 44092
rect 23012 44036 23016 44092
rect 22952 44032 23016 44036
rect 23032 44092 23096 44096
rect 23032 44036 23036 44092
rect 23036 44036 23092 44092
rect 23092 44036 23096 44092
rect 23032 44032 23096 44036
rect 23112 44092 23176 44096
rect 23112 44036 23116 44092
rect 23116 44036 23172 44092
rect 23172 44036 23176 44092
rect 23112 44032 23176 44036
rect 23192 44092 23256 44096
rect 23192 44036 23196 44092
rect 23196 44036 23252 44092
rect 23252 44036 23256 44092
rect 23192 44032 23256 44036
rect 7952 43548 8016 43552
rect 7952 43492 7956 43548
rect 7956 43492 8012 43548
rect 8012 43492 8016 43548
rect 7952 43488 8016 43492
rect 8032 43548 8096 43552
rect 8032 43492 8036 43548
rect 8036 43492 8092 43548
rect 8092 43492 8096 43548
rect 8032 43488 8096 43492
rect 8112 43548 8176 43552
rect 8112 43492 8116 43548
rect 8116 43492 8172 43548
rect 8172 43492 8176 43548
rect 8112 43488 8176 43492
rect 8192 43548 8256 43552
rect 8192 43492 8196 43548
rect 8196 43492 8252 43548
rect 8252 43492 8256 43548
rect 8192 43488 8256 43492
rect 17952 43548 18016 43552
rect 17952 43492 17956 43548
rect 17956 43492 18012 43548
rect 18012 43492 18016 43548
rect 17952 43488 18016 43492
rect 18032 43548 18096 43552
rect 18032 43492 18036 43548
rect 18036 43492 18092 43548
rect 18092 43492 18096 43548
rect 18032 43488 18096 43492
rect 18112 43548 18176 43552
rect 18112 43492 18116 43548
rect 18116 43492 18172 43548
rect 18172 43492 18176 43548
rect 18112 43488 18176 43492
rect 18192 43548 18256 43552
rect 18192 43492 18196 43548
rect 18196 43492 18252 43548
rect 18252 43492 18256 43548
rect 18192 43488 18256 43492
rect 2952 43004 3016 43008
rect 2952 42948 2956 43004
rect 2956 42948 3012 43004
rect 3012 42948 3016 43004
rect 2952 42944 3016 42948
rect 3032 43004 3096 43008
rect 3032 42948 3036 43004
rect 3036 42948 3092 43004
rect 3092 42948 3096 43004
rect 3032 42944 3096 42948
rect 3112 43004 3176 43008
rect 3112 42948 3116 43004
rect 3116 42948 3172 43004
rect 3172 42948 3176 43004
rect 3112 42944 3176 42948
rect 3192 43004 3256 43008
rect 3192 42948 3196 43004
rect 3196 42948 3252 43004
rect 3252 42948 3256 43004
rect 3192 42944 3256 42948
rect 12952 43004 13016 43008
rect 12952 42948 12956 43004
rect 12956 42948 13012 43004
rect 13012 42948 13016 43004
rect 12952 42944 13016 42948
rect 13032 43004 13096 43008
rect 13032 42948 13036 43004
rect 13036 42948 13092 43004
rect 13092 42948 13096 43004
rect 13032 42944 13096 42948
rect 13112 43004 13176 43008
rect 13112 42948 13116 43004
rect 13116 42948 13172 43004
rect 13172 42948 13176 43004
rect 13112 42944 13176 42948
rect 13192 43004 13256 43008
rect 13192 42948 13196 43004
rect 13196 42948 13252 43004
rect 13252 42948 13256 43004
rect 13192 42944 13256 42948
rect 22952 43004 23016 43008
rect 22952 42948 22956 43004
rect 22956 42948 23012 43004
rect 23012 42948 23016 43004
rect 22952 42944 23016 42948
rect 23032 43004 23096 43008
rect 23032 42948 23036 43004
rect 23036 42948 23092 43004
rect 23092 42948 23096 43004
rect 23032 42944 23096 42948
rect 23112 43004 23176 43008
rect 23112 42948 23116 43004
rect 23116 42948 23172 43004
rect 23172 42948 23176 43004
rect 23112 42944 23176 42948
rect 23192 43004 23256 43008
rect 23192 42948 23196 43004
rect 23196 42948 23252 43004
rect 23252 42948 23256 43004
rect 23192 42944 23256 42948
rect 7952 42460 8016 42464
rect 7952 42404 7956 42460
rect 7956 42404 8012 42460
rect 8012 42404 8016 42460
rect 7952 42400 8016 42404
rect 8032 42460 8096 42464
rect 8032 42404 8036 42460
rect 8036 42404 8092 42460
rect 8092 42404 8096 42460
rect 8032 42400 8096 42404
rect 8112 42460 8176 42464
rect 8112 42404 8116 42460
rect 8116 42404 8172 42460
rect 8172 42404 8176 42460
rect 8112 42400 8176 42404
rect 8192 42460 8256 42464
rect 8192 42404 8196 42460
rect 8196 42404 8252 42460
rect 8252 42404 8256 42460
rect 8192 42400 8256 42404
rect 17952 42460 18016 42464
rect 17952 42404 17956 42460
rect 17956 42404 18012 42460
rect 18012 42404 18016 42460
rect 17952 42400 18016 42404
rect 18032 42460 18096 42464
rect 18032 42404 18036 42460
rect 18036 42404 18092 42460
rect 18092 42404 18096 42460
rect 18032 42400 18096 42404
rect 18112 42460 18176 42464
rect 18112 42404 18116 42460
rect 18116 42404 18172 42460
rect 18172 42404 18176 42460
rect 18112 42400 18176 42404
rect 18192 42460 18256 42464
rect 18192 42404 18196 42460
rect 18196 42404 18252 42460
rect 18252 42404 18256 42460
rect 18192 42400 18256 42404
rect 2952 41916 3016 41920
rect 2952 41860 2956 41916
rect 2956 41860 3012 41916
rect 3012 41860 3016 41916
rect 2952 41856 3016 41860
rect 3032 41916 3096 41920
rect 3032 41860 3036 41916
rect 3036 41860 3092 41916
rect 3092 41860 3096 41916
rect 3032 41856 3096 41860
rect 3112 41916 3176 41920
rect 3112 41860 3116 41916
rect 3116 41860 3172 41916
rect 3172 41860 3176 41916
rect 3112 41856 3176 41860
rect 3192 41916 3256 41920
rect 3192 41860 3196 41916
rect 3196 41860 3252 41916
rect 3252 41860 3256 41916
rect 3192 41856 3256 41860
rect 12952 41916 13016 41920
rect 12952 41860 12956 41916
rect 12956 41860 13012 41916
rect 13012 41860 13016 41916
rect 12952 41856 13016 41860
rect 13032 41916 13096 41920
rect 13032 41860 13036 41916
rect 13036 41860 13092 41916
rect 13092 41860 13096 41916
rect 13032 41856 13096 41860
rect 13112 41916 13176 41920
rect 13112 41860 13116 41916
rect 13116 41860 13172 41916
rect 13172 41860 13176 41916
rect 13112 41856 13176 41860
rect 13192 41916 13256 41920
rect 13192 41860 13196 41916
rect 13196 41860 13252 41916
rect 13252 41860 13256 41916
rect 13192 41856 13256 41860
rect 22952 41916 23016 41920
rect 22952 41860 22956 41916
rect 22956 41860 23012 41916
rect 23012 41860 23016 41916
rect 22952 41856 23016 41860
rect 23032 41916 23096 41920
rect 23032 41860 23036 41916
rect 23036 41860 23092 41916
rect 23092 41860 23096 41916
rect 23032 41856 23096 41860
rect 23112 41916 23176 41920
rect 23112 41860 23116 41916
rect 23116 41860 23172 41916
rect 23172 41860 23176 41916
rect 23112 41856 23176 41860
rect 23192 41916 23256 41920
rect 23192 41860 23196 41916
rect 23196 41860 23252 41916
rect 23252 41860 23256 41916
rect 23192 41856 23256 41860
rect 7952 41372 8016 41376
rect 7952 41316 7956 41372
rect 7956 41316 8012 41372
rect 8012 41316 8016 41372
rect 7952 41312 8016 41316
rect 8032 41372 8096 41376
rect 8032 41316 8036 41372
rect 8036 41316 8092 41372
rect 8092 41316 8096 41372
rect 8032 41312 8096 41316
rect 8112 41372 8176 41376
rect 8112 41316 8116 41372
rect 8116 41316 8172 41372
rect 8172 41316 8176 41372
rect 8112 41312 8176 41316
rect 8192 41372 8256 41376
rect 8192 41316 8196 41372
rect 8196 41316 8252 41372
rect 8252 41316 8256 41372
rect 8192 41312 8256 41316
rect 17952 41372 18016 41376
rect 17952 41316 17956 41372
rect 17956 41316 18012 41372
rect 18012 41316 18016 41372
rect 17952 41312 18016 41316
rect 18032 41372 18096 41376
rect 18032 41316 18036 41372
rect 18036 41316 18092 41372
rect 18092 41316 18096 41372
rect 18032 41312 18096 41316
rect 18112 41372 18176 41376
rect 18112 41316 18116 41372
rect 18116 41316 18172 41372
rect 18172 41316 18176 41372
rect 18112 41312 18176 41316
rect 18192 41372 18256 41376
rect 18192 41316 18196 41372
rect 18196 41316 18252 41372
rect 18252 41316 18256 41372
rect 18192 41312 18256 41316
rect 2952 40828 3016 40832
rect 2952 40772 2956 40828
rect 2956 40772 3012 40828
rect 3012 40772 3016 40828
rect 2952 40768 3016 40772
rect 3032 40828 3096 40832
rect 3032 40772 3036 40828
rect 3036 40772 3092 40828
rect 3092 40772 3096 40828
rect 3032 40768 3096 40772
rect 3112 40828 3176 40832
rect 3112 40772 3116 40828
rect 3116 40772 3172 40828
rect 3172 40772 3176 40828
rect 3112 40768 3176 40772
rect 3192 40828 3256 40832
rect 3192 40772 3196 40828
rect 3196 40772 3252 40828
rect 3252 40772 3256 40828
rect 3192 40768 3256 40772
rect 12952 40828 13016 40832
rect 12952 40772 12956 40828
rect 12956 40772 13012 40828
rect 13012 40772 13016 40828
rect 12952 40768 13016 40772
rect 13032 40828 13096 40832
rect 13032 40772 13036 40828
rect 13036 40772 13092 40828
rect 13092 40772 13096 40828
rect 13032 40768 13096 40772
rect 13112 40828 13176 40832
rect 13112 40772 13116 40828
rect 13116 40772 13172 40828
rect 13172 40772 13176 40828
rect 13112 40768 13176 40772
rect 13192 40828 13256 40832
rect 13192 40772 13196 40828
rect 13196 40772 13252 40828
rect 13252 40772 13256 40828
rect 13192 40768 13256 40772
rect 22952 40828 23016 40832
rect 22952 40772 22956 40828
rect 22956 40772 23012 40828
rect 23012 40772 23016 40828
rect 22952 40768 23016 40772
rect 23032 40828 23096 40832
rect 23032 40772 23036 40828
rect 23036 40772 23092 40828
rect 23092 40772 23096 40828
rect 23032 40768 23096 40772
rect 23112 40828 23176 40832
rect 23112 40772 23116 40828
rect 23116 40772 23172 40828
rect 23172 40772 23176 40828
rect 23112 40768 23176 40772
rect 23192 40828 23256 40832
rect 23192 40772 23196 40828
rect 23196 40772 23252 40828
rect 23252 40772 23256 40828
rect 23192 40768 23256 40772
rect 7952 40284 8016 40288
rect 7952 40228 7956 40284
rect 7956 40228 8012 40284
rect 8012 40228 8016 40284
rect 7952 40224 8016 40228
rect 8032 40284 8096 40288
rect 8032 40228 8036 40284
rect 8036 40228 8092 40284
rect 8092 40228 8096 40284
rect 8032 40224 8096 40228
rect 8112 40284 8176 40288
rect 8112 40228 8116 40284
rect 8116 40228 8172 40284
rect 8172 40228 8176 40284
rect 8112 40224 8176 40228
rect 8192 40284 8256 40288
rect 8192 40228 8196 40284
rect 8196 40228 8252 40284
rect 8252 40228 8256 40284
rect 8192 40224 8256 40228
rect 17952 40284 18016 40288
rect 17952 40228 17956 40284
rect 17956 40228 18012 40284
rect 18012 40228 18016 40284
rect 17952 40224 18016 40228
rect 18032 40284 18096 40288
rect 18032 40228 18036 40284
rect 18036 40228 18092 40284
rect 18092 40228 18096 40284
rect 18032 40224 18096 40228
rect 18112 40284 18176 40288
rect 18112 40228 18116 40284
rect 18116 40228 18172 40284
rect 18172 40228 18176 40284
rect 18112 40224 18176 40228
rect 18192 40284 18256 40288
rect 18192 40228 18196 40284
rect 18196 40228 18252 40284
rect 18252 40228 18256 40284
rect 18192 40224 18256 40228
rect 2952 39740 3016 39744
rect 2952 39684 2956 39740
rect 2956 39684 3012 39740
rect 3012 39684 3016 39740
rect 2952 39680 3016 39684
rect 3032 39740 3096 39744
rect 3032 39684 3036 39740
rect 3036 39684 3092 39740
rect 3092 39684 3096 39740
rect 3032 39680 3096 39684
rect 3112 39740 3176 39744
rect 3112 39684 3116 39740
rect 3116 39684 3172 39740
rect 3172 39684 3176 39740
rect 3112 39680 3176 39684
rect 3192 39740 3256 39744
rect 3192 39684 3196 39740
rect 3196 39684 3252 39740
rect 3252 39684 3256 39740
rect 3192 39680 3256 39684
rect 12952 39740 13016 39744
rect 12952 39684 12956 39740
rect 12956 39684 13012 39740
rect 13012 39684 13016 39740
rect 12952 39680 13016 39684
rect 13032 39740 13096 39744
rect 13032 39684 13036 39740
rect 13036 39684 13092 39740
rect 13092 39684 13096 39740
rect 13032 39680 13096 39684
rect 13112 39740 13176 39744
rect 13112 39684 13116 39740
rect 13116 39684 13172 39740
rect 13172 39684 13176 39740
rect 13112 39680 13176 39684
rect 13192 39740 13256 39744
rect 13192 39684 13196 39740
rect 13196 39684 13252 39740
rect 13252 39684 13256 39740
rect 13192 39680 13256 39684
rect 22952 39740 23016 39744
rect 22952 39684 22956 39740
rect 22956 39684 23012 39740
rect 23012 39684 23016 39740
rect 22952 39680 23016 39684
rect 23032 39740 23096 39744
rect 23032 39684 23036 39740
rect 23036 39684 23092 39740
rect 23092 39684 23096 39740
rect 23032 39680 23096 39684
rect 23112 39740 23176 39744
rect 23112 39684 23116 39740
rect 23116 39684 23172 39740
rect 23172 39684 23176 39740
rect 23112 39680 23176 39684
rect 23192 39740 23256 39744
rect 23192 39684 23196 39740
rect 23196 39684 23252 39740
rect 23252 39684 23256 39740
rect 23192 39680 23256 39684
rect 7952 39196 8016 39200
rect 7952 39140 7956 39196
rect 7956 39140 8012 39196
rect 8012 39140 8016 39196
rect 7952 39136 8016 39140
rect 8032 39196 8096 39200
rect 8032 39140 8036 39196
rect 8036 39140 8092 39196
rect 8092 39140 8096 39196
rect 8032 39136 8096 39140
rect 8112 39196 8176 39200
rect 8112 39140 8116 39196
rect 8116 39140 8172 39196
rect 8172 39140 8176 39196
rect 8112 39136 8176 39140
rect 8192 39196 8256 39200
rect 8192 39140 8196 39196
rect 8196 39140 8252 39196
rect 8252 39140 8256 39196
rect 8192 39136 8256 39140
rect 17952 39196 18016 39200
rect 17952 39140 17956 39196
rect 17956 39140 18012 39196
rect 18012 39140 18016 39196
rect 17952 39136 18016 39140
rect 18032 39196 18096 39200
rect 18032 39140 18036 39196
rect 18036 39140 18092 39196
rect 18092 39140 18096 39196
rect 18032 39136 18096 39140
rect 18112 39196 18176 39200
rect 18112 39140 18116 39196
rect 18116 39140 18172 39196
rect 18172 39140 18176 39196
rect 18112 39136 18176 39140
rect 18192 39196 18256 39200
rect 18192 39140 18196 39196
rect 18196 39140 18252 39196
rect 18252 39140 18256 39196
rect 18192 39136 18256 39140
rect 2952 38652 3016 38656
rect 2952 38596 2956 38652
rect 2956 38596 3012 38652
rect 3012 38596 3016 38652
rect 2952 38592 3016 38596
rect 3032 38652 3096 38656
rect 3032 38596 3036 38652
rect 3036 38596 3092 38652
rect 3092 38596 3096 38652
rect 3032 38592 3096 38596
rect 3112 38652 3176 38656
rect 3112 38596 3116 38652
rect 3116 38596 3172 38652
rect 3172 38596 3176 38652
rect 3112 38592 3176 38596
rect 3192 38652 3256 38656
rect 3192 38596 3196 38652
rect 3196 38596 3252 38652
rect 3252 38596 3256 38652
rect 3192 38592 3256 38596
rect 12952 38652 13016 38656
rect 12952 38596 12956 38652
rect 12956 38596 13012 38652
rect 13012 38596 13016 38652
rect 12952 38592 13016 38596
rect 13032 38652 13096 38656
rect 13032 38596 13036 38652
rect 13036 38596 13092 38652
rect 13092 38596 13096 38652
rect 13032 38592 13096 38596
rect 13112 38652 13176 38656
rect 13112 38596 13116 38652
rect 13116 38596 13172 38652
rect 13172 38596 13176 38652
rect 13112 38592 13176 38596
rect 13192 38652 13256 38656
rect 13192 38596 13196 38652
rect 13196 38596 13252 38652
rect 13252 38596 13256 38652
rect 13192 38592 13256 38596
rect 22952 38652 23016 38656
rect 22952 38596 22956 38652
rect 22956 38596 23012 38652
rect 23012 38596 23016 38652
rect 22952 38592 23016 38596
rect 23032 38652 23096 38656
rect 23032 38596 23036 38652
rect 23036 38596 23092 38652
rect 23092 38596 23096 38652
rect 23032 38592 23096 38596
rect 23112 38652 23176 38656
rect 23112 38596 23116 38652
rect 23116 38596 23172 38652
rect 23172 38596 23176 38652
rect 23112 38592 23176 38596
rect 23192 38652 23256 38656
rect 23192 38596 23196 38652
rect 23196 38596 23252 38652
rect 23252 38596 23256 38652
rect 23192 38592 23256 38596
rect 7952 38108 8016 38112
rect 7952 38052 7956 38108
rect 7956 38052 8012 38108
rect 8012 38052 8016 38108
rect 7952 38048 8016 38052
rect 8032 38108 8096 38112
rect 8032 38052 8036 38108
rect 8036 38052 8092 38108
rect 8092 38052 8096 38108
rect 8032 38048 8096 38052
rect 8112 38108 8176 38112
rect 8112 38052 8116 38108
rect 8116 38052 8172 38108
rect 8172 38052 8176 38108
rect 8112 38048 8176 38052
rect 8192 38108 8256 38112
rect 8192 38052 8196 38108
rect 8196 38052 8252 38108
rect 8252 38052 8256 38108
rect 8192 38048 8256 38052
rect 17952 38108 18016 38112
rect 17952 38052 17956 38108
rect 17956 38052 18012 38108
rect 18012 38052 18016 38108
rect 17952 38048 18016 38052
rect 18032 38108 18096 38112
rect 18032 38052 18036 38108
rect 18036 38052 18092 38108
rect 18092 38052 18096 38108
rect 18032 38048 18096 38052
rect 18112 38108 18176 38112
rect 18112 38052 18116 38108
rect 18116 38052 18172 38108
rect 18172 38052 18176 38108
rect 18112 38048 18176 38052
rect 18192 38108 18256 38112
rect 18192 38052 18196 38108
rect 18196 38052 18252 38108
rect 18252 38052 18256 38108
rect 18192 38048 18256 38052
rect 2952 37564 3016 37568
rect 2952 37508 2956 37564
rect 2956 37508 3012 37564
rect 3012 37508 3016 37564
rect 2952 37504 3016 37508
rect 3032 37564 3096 37568
rect 3032 37508 3036 37564
rect 3036 37508 3092 37564
rect 3092 37508 3096 37564
rect 3032 37504 3096 37508
rect 3112 37564 3176 37568
rect 3112 37508 3116 37564
rect 3116 37508 3172 37564
rect 3172 37508 3176 37564
rect 3112 37504 3176 37508
rect 3192 37564 3256 37568
rect 3192 37508 3196 37564
rect 3196 37508 3252 37564
rect 3252 37508 3256 37564
rect 3192 37504 3256 37508
rect 12952 37564 13016 37568
rect 12952 37508 12956 37564
rect 12956 37508 13012 37564
rect 13012 37508 13016 37564
rect 12952 37504 13016 37508
rect 13032 37564 13096 37568
rect 13032 37508 13036 37564
rect 13036 37508 13092 37564
rect 13092 37508 13096 37564
rect 13032 37504 13096 37508
rect 13112 37564 13176 37568
rect 13112 37508 13116 37564
rect 13116 37508 13172 37564
rect 13172 37508 13176 37564
rect 13112 37504 13176 37508
rect 13192 37564 13256 37568
rect 13192 37508 13196 37564
rect 13196 37508 13252 37564
rect 13252 37508 13256 37564
rect 13192 37504 13256 37508
rect 22952 37564 23016 37568
rect 22952 37508 22956 37564
rect 22956 37508 23012 37564
rect 23012 37508 23016 37564
rect 22952 37504 23016 37508
rect 23032 37564 23096 37568
rect 23032 37508 23036 37564
rect 23036 37508 23092 37564
rect 23092 37508 23096 37564
rect 23032 37504 23096 37508
rect 23112 37564 23176 37568
rect 23112 37508 23116 37564
rect 23116 37508 23172 37564
rect 23172 37508 23176 37564
rect 23112 37504 23176 37508
rect 23192 37564 23256 37568
rect 23192 37508 23196 37564
rect 23196 37508 23252 37564
rect 23252 37508 23256 37564
rect 23192 37504 23256 37508
rect 7952 37020 8016 37024
rect 7952 36964 7956 37020
rect 7956 36964 8012 37020
rect 8012 36964 8016 37020
rect 7952 36960 8016 36964
rect 8032 37020 8096 37024
rect 8032 36964 8036 37020
rect 8036 36964 8092 37020
rect 8092 36964 8096 37020
rect 8032 36960 8096 36964
rect 8112 37020 8176 37024
rect 8112 36964 8116 37020
rect 8116 36964 8172 37020
rect 8172 36964 8176 37020
rect 8112 36960 8176 36964
rect 8192 37020 8256 37024
rect 8192 36964 8196 37020
rect 8196 36964 8252 37020
rect 8252 36964 8256 37020
rect 8192 36960 8256 36964
rect 17952 37020 18016 37024
rect 17952 36964 17956 37020
rect 17956 36964 18012 37020
rect 18012 36964 18016 37020
rect 17952 36960 18016 36964
rect 18032 37020 18096 37024
rect 18032 36964 18036 37020
rect 18036 36964 18092 37020
rect 18092 36964 18096 37020
rect 18032 36960 18096 36964
rect 18112 37020 18176 37024
rect 18112 36964 18116 37020
rect 18116 36964 18172 37020
rect 18172 36964 18176 37020
rect 18112 36960 18176 36964
rect 18192 37020 18256 37024
rect 18192 36964 18196 37020
rect 18196 36964 18252 37020
rect 18252 36964 18256 37020
rect 18192 36960 18256 36964
rect 2952 36476 3016 36480
rect 2952 36420 2956 36476
rect 2956 36420 3012 36476
rect 3012 36420 3016 36476
rect 2952 36416 3016 36420
rect 3032 36476 3096 36480
rect 3032 36420 3036 36476
rect 3036 36420 3092 36476
rect 3092 36420 3096 36476
rect 3032 36416 3096 36420
rect 3112 36476 3176 36480
rect 3112 36420 3116 36476
rect 3116 36420 3172 36476
rect 3172 36420 3176 36476
rect 3112 36416 3176 36420
rect 3192 36476 3256 36480
rect 3192 36420 3196 36476
rect 3196 36420 3252 36476
rect 3252 36420 3256 36476
rect 3192 36416 3256 36420
rect 12952 36476 13016 36480
rect 12952 36420 12956 36476
rect 12956 36420 13012 36476
rect 13012 36420 13016 36476
rect 12952 36416 13016 36420
rect 13032 36476 13096 36480
rect 13032 36420 13036 36476
rect 13036 36420 13092 36476
rect 13092 36420 13096 36476
rect 13032 36416 13096 36420
rect 13112 36476 13176 36480
rect 13112 36420 13116 36476
rect 13116 36420 13172 36476
rect 13172 36420 13176 36476
rect 13112 36416 13176 36420
rect 13192 36476 13256 36480
rect 13192 36420 13196 36476
rect 13196 36420 13252 36476
rect 13252 36420 13256 36476
rect 13192 36416 13256 36420
rect 22952 36476 23016 36480
rect 22952 36420 22956 36476
rect 22956 36420 23012 36476
rect 23012 36420 23016 36476
rect 22952 36416 23016 36420
rect 23032 36476 23096 36480
rect 23032 36420 23036 36476
rect 23036 36420 23092 36476
rect 23092 36420 23096 36476
rect 23032 36416 23096 36420
rect 23112 36476 23176 36480
rect 23112 36420 23116 36476
rect 23116 36420 23172 36476
rect 23172 36420 23176 36476
rect 23112 36416 23176 36420
rect 23192 36476 23256 36480
rect 23192 36420 23196 36476
rect 23196 36420 23252 36476
rect 23252 36420 23256 36476
rect 23192 36416 23256 36420
rect 7952 35932 8016 35936
rect 7952 35876 7956 35932
rect 7956 35876 8012 35932
rect 8012 35876 8016 35932
rect 7952 35872 8016 35876
rect 8032 35932 8096 35936
rect 8032 35876 8036 35932
rect 8036 35876 8092 35932
rect 8092 35876 8096 35932
rect 8032 35872 8096 35876
rect 8112 35932 8176 35936
rect 8112 35876 8116 35932
rect 8116 35876 8172 35932
rect 8172 35876 8176 35932
rect 8112 35872 8176 35876
rect 8192 35932 8256 35936
rect 8192 35876 8196 35932
rect 8196 35876 8252 35932
rect 8252 35876 8256 35932
rect 8192 35872 8256 35876
rect 17952 35932 18016 35936
rect 17952 35876 17956 35932
rect 17956 35876 18012 35932
rect 18012 35876 18016 35932
rect 17952 35872 18016 35876
rect 18032 35932 18096 35936
rect 18032 35876 18036 35932
rect 18036 35876 18092 35932
rect 18092 35876 18096 35932
rect 18032 35872 18096 35876
rect 18112 35932 18176 35936
rect 18112 35876 18116 35932
rect 18116 35876 18172 35932
rect 18172 35876 18176 35932
rect 18112 35872 18176 35876
rect 18192 35932 18256 35936
rect 18192 35876 18196 35932
rect 18196 35876 18252 35932
rect 18252 35876 18256 35932
rect 18192 35872 18256 35876
rect 2952 35388 3016 35392
rect 2952 35332 2956 35388
rect 2956 35332 3012 35388
rect 3012 35332 3016 35388
rect 2952 35328 3016 35332
rect 3032 35388 3096 35392
rect 3032 35332 3036 35388
rect 3036 35332 3092 35388
rect 3092 35332 3096 35388
rect 3032 35328 3096 35332
rect 3112 35388 3176 35392
rect 3112 35332 3116 35388
rect 3116 35332 3172 35388
rect 3172 35332 3176 35388
rect 3112 35328 3176 35332
rect 3192 35388 3256 35392
rect 3192 35332 3196 35388
rect 3196 35332 3252 35388
rect 3252 35332 3256 35388
rect 3192 35328 3256 35332
rect 12952 35388 13016 35392
rect 12952 35332 12956 35388
rect 12956 35332 13012 35388
rect 13012 35332 13016 35388
rect 12952 35328 13016 35332
rect 13032 35388 13096 35392
rect 13032 35332 13036 35388
rect 13036 35332 13092 35388
rect 13092 35332 13096 35388
rect 13032 35328 13096 35332
rect 13112 35388 13176 35392
rect 13112 35332 13116 35388
rect 13116 35332 13172 35388
rect 13172 35332 13176 35388
rect 13112 35328 13176 35332
rect 13192 35388 13256 35392
rect 13192 35332 13196 35388
rect 13196 35332 13252 35388
rect 13252 35332 13256 35388
rect 13192 35328 13256 35332
rect 22952 35388 23016 35392
rect 22952 35332 22956 35388
rect 22956 35332 23012 35388
rect 23012 35332 23016 35388
rect 22952 35328 23016 35332
rect 23032 35388 23096 35392
rect 23032 35332 23036 35388
rect 23036 35332 23092 35388
rect 23092 35332 23096 35388
rect 23032 35328 23096 35332
rect 23112 35388 23176 35392
rect 23112 35332 23116 35388
rect 23116 35332 23172 35388
rect 23172 35332 23176 35388
rect 23112 35328 23176 35332
rect 23192 35388 23256 35392
rect 23192 35332 23196 35388
rect 23196 35332 23252 35388
rect 23252 35332 23256 35388
rect 23192 35328 23256 35332
rect 7952 34844 8016 34848
rect 7952 34788 7956 34844
rect 7956 34788 8012 34844
rect 8012 34788 8016 34844
rect 7952 34784 8016 34788
rect 8032 34844 8096 34848
rect 8032 34788 8036 34844
rect 8036 34788 8092 34844
rect 8092 34788 8096 34844
rect 8032 34784 8096 34788
rect 8112 34844 8176 34848
rect 8112 34788 8116 34844
rect 8116 34788 8172 34844
rect 8172 34788 8176 34844
rect 8112 34784 8176 34788
rect 8192 34844 8256 34848
rect 8192 34788 8196 34844
rect 8196 34788 8252 34844
rect 8252 34788 8256 34844
rect 8192 34784 8256 34788
rect 17952 34844 18016 34848
rect 17952 34788 17956 34844
rect 17956 34788 18012 34844
rect 18012 34788 18016 34844
rect 17952 34784 18016 34788
rect 18032 34844 18096 34848
rect 18032 34788 18036 34844
rect 18036 34788 18092 34844
rect 18092 34788 18096 34844
rect 18032 34784 18096 34788
rect 18112 34844 18176 34848
rect 18112 34788 18116 34844
rect 18116 34788 18172 34844
rect 18172 34788 18176 34844
rect 18112 34784 18176 34788
rect 18192 34844 18256 34848
rect 18192 34788 18196 34844
rect 18196 34788 18252 34844
rect 18252 34788 18256 34844
rect 18192 34784 18256 34788
rect 2952 34300 3016 34304
rect 2952 34244 2956 34300
rect 2956 34244 3012 34300
rect 3012 34244 3016 34300
rect 2952 34240 3016 34244
rect 3032 34300 3096 34304
rect 3032 34244 3036 34300
rect 3036 34244 3092 34300
rect 3092 34244 3096 34300
rect 3032 34240 3096 34244
rect 3112 34300 3176 34304
rect 3112 34244 3116 34300
rect 3116 34244 3172 34300
rect 3172 34244 3176 34300
rect 3112 34240 3176 34244
rect 3192 34300 3256 34304
rect 3192 34244 3196 34300
rect 3196 34244 3252 34300
rect 3252 34244 3256 34300
rect 3192 34240 3256 34244
rect 12952 34300 13016 34304
rect 12952 34244 12956 34300
rect 12956 34244 13012 34300
rect 13012 34244 13016 34300
rect 12952 34240 13016 34244
rect 13032 34300 13096 34304
rect 13032 34244 13036 34300
rect 13036 34244 13092 34300
rect 13092 34244 13096 34300
rect 13032 34240 13096 34244
rect 13112 34300 13176 34304
rect 13112 34244 13116 34300
rect 13116 34244 13172 34300
rect 13172 34244 13176 34300
rect 13112 34240 13176 34244
rect 13192 34300 13256 34304
rect 13192 34244 13196 34300
rect 13196 34244 13252 34300
rect 13252 34244 13256 34300
rect 13192 34240 13256 34244
rect 22952 34300 23016 34304
rect 22952 34244 22956 34300
rect 22956 34244 23012 34300
rect 23012 34244 23016 34300
rect 22952 34240 23016 34244
rect 23032 34300 23096 34304
rect 23032 34244 23036 34300
rect 23036 34244 23092 34300
rect 23092 34244 23096 34300
rect 23032 34240 23096 34244
rect 23112 34300 23176 34304
rect 23112 34244 23116 34300
rect 23116 34244 23172 34300
rect 23172 34244 23176 34300
rect 23112 34240 23176 34244
rect 23192 34300 23256 34304
rect 23192 34244 23196 34300
rect 23196 34244 23252 34300
rect 23252 34244 23256 34300
rect 23192 34240 23256 34244
rect 7952 33756 8016 33760
rect 7952 33700 7956 33756
rect 7956 33700 8012 33756
rect 8012 33700 8016 33756
rect 7952 33696 8016 33700
rect 8032 33756 8096 33760
rect 8032 33700 8036 33756
rect 8036 33700 8092 33756
rect 8092 33700 8096 33756
rect 8032 33696 8096 33700
rect 8112 33756 8176 33760
rect 8112 33700 8116 33756
rect 8116 33700 8172 33756
rect 8172 33700 8176 33756
rect 8112 33696 8176 33700
rect 8192 33756 8256 33760
rect 8192 33700 8196 33756
rect 8196 33700 8252 33756
rect 8252 33700 8256 33756
rect 8192 33696 8256 33700
rect 17952 33756 18016 33760
rect 17952 33700 17956 33756
rect 17956 33700 18012 33756
rect 18012 33700 18016 33756
rect 17952 33696 18016 33700
rect 18032 33756 18096 33760
rect 18032 33700 18036 33756
rect 18036 33700 18092 33756
rect 18092 33700 18096 33756
rect 18032 33696 18096 33700
rect 18112 33756 18176 33760
rect 18112 33700 18116 33756
rect 18116 33700 18172 33756
rect 18172 33700 18176 33756
rect 18112 33696 18176 33700
rect 18192 33756 18256 33760
rect 18192 33700 18196 33756
rect 18196 33700 18252 33756
rect 18252 33700 18256 33756
rect 18192 33696 18256 33700
rect 2952 33212 3016 33216
rect 2952 33156 2956 33212
rect 2956 33156 3012 33212
rect 3012 33156 3016 33212
rect 2952 33152 3016 33156
rect 3032 33212 3096 33216
rect 3032 33156 3036 33212
rect 3036 33156 3092 33212
rect 3092 33156 3096 33212
rect 3032 33152 3096 33156
rect 3112 33212 3176 33216
rect 3112 33156 3116 33212
rect 3116 33156 3172 33212
rect 3172 33156 3176 33212
rect 3112 33152 3176 33156
rect 3192 33212 3256 33216
rect 3192 33156 3196 33212
rect 3196 33156 3252 33212
rect 3252 33156 3256 33212
rect 3192 33152 3256 33156
rect 12952 33212 13016 33216
rect 12952 33156 12956 33212
rect 12956 33156 13012 33212
rect 13012 33156 13016 33212
rect 12952 33152 13016 33156
rect 13032 33212 13096 33216
rect 13032 33156 13036 33212
rect 13036 33156 13092 33212
rect 13092 33156 13096 33212
rect 13032 33152 13096 33156
rect 13112 33212 13176 33216
rect 13112 33156 13116 33212
rect 13116 33156 13172 33212
rect 13172 33156 13176 33212
rect 13112 33152 13176 33156
rect 13192 33212 13256 33216
rect 13192 33156 13196 33212
rect 13196 33156 13252 33212
rect 13252 33156 13256 33212
rect 13192 33152 13256 33156
rect 22952 33212 23016 33216
rect 22952 33156 22956 33212
rect 22956 33156 23012 33212
rect 23012 33156 23016 33212
rect 22952 33152 23016 33156
rect 23032 33212 23096 33216
rect 23032 33156 23036 33212
rect 23036 33156 23092 33212
rect 23092 33156 23096 33212
rect 23032 33152 23096 33156
rect 23112 33212 23176 33216
rect 23112 33156 23116 33212
rect 23116 33156 23172 33212
rect 23172 33156 23176 33212
rect 23112 33152 23176 33156
rect 23192 33212 23256 33216
rect 23192 33156 23196 33212
rect 23196 33156 23252 33212
rect 23252 33156 23256 33212
rect 23192 33152 23256 33156
rect 7952 32668 8016 32672
rect 7952 32612 7956 32668
rect 7956 32612 8012 32668
rect 8012 32612 8016 32668
rect 7952 32608 8016 32612
rect 8032 32668 8096 32672
rect 8032 32612 8036 32668
rect 8036 32612 8092 32668
rect 8092 32612 8096 32668
rect 8032 32608 8096 32612
rect 8112 32668 8176 32672
rect 8112 32612 8116 32668
rect 8116 32612 8172 32668
rect 8172 32612 8176 32668
rect 8112 32608 8176 32612
rect 8192 32668 8256 32672
rect 8192 32612 8196 32668
rect 8196 32612 8252 32668
rect 8252 32612 8256 32668
rect 8192 32608 8256 32612
rect 17952 32668 18016 32672
rect 17952 32612 17956 32668
rect 17956 32612 18012 32668
rect 18012 32612 18016 32668
rect 17952 32608 18016 32612
rect 18032 32668 18096 32672
rect 18032 32612 18036 32668
rect 18036 32612 18092 32668
rect 18092 32612 18096 32668
rect 18032 32608 18096 32612
rect 18112 32668 18176 32672
rect 18112 32612 18116 32668
rect 18116 32612 18172 32668
rect 18172 32612 18176 32668
rect 18112 32608 18176 32612
rect 18192 32668 18256 32672
rect 18192 32612 18196 32668
rect 18196 32612 18252 32668
rect 18252 32612 18256 32668
rect 18192 32608 18256 32612
rect 2952 32124 3016 32128
rect 2952 32068 2956 32124
rect 2956 32068 3012 32124
rect 3012 32068 3016 32124
rect 2952 32064 3016 32068
rect 3032 32124 3096 32128
rect 3032 32068 3036 32124
rect 3036 32068 3092 32124
rect 3092 32068 3096 32124
rect 3032 32064 3096 32068
rect 3112 32124 3176 32128
rect 3112 32068 3116 32124
rect 3116 32068 3172 32124
rect 3172 32068 3176 32124
rect 3112 32064 3176 32068
rect 3192 32124 3256 32128
rect 3192 32068 3196 32124
rect 3196 32068 3252 32124
rect 3252 32068 3256 32124
rect 3192 32064 3256 32068
rect 12952 32124 13016 32128
rect 12952 32068 12956 32124
rect 12956 32068 13012 32124
rect 13012 32068 13016 32124
rect 12952 32064 13016 32068
rect 13032 32124 13096 32128
rect 13032 32068 13036 32124
rect 13036 32068 13092 32124
rect 13092 32068 13096 32124
rect 13032 32064 13096 32068
rect 13112 32124 13176 32128
rect 13112 32068 13116 32124
rect 13116 32068 13172 32124
rect 13172 32068 13176 32124
rect 13112 32064 13176 32068
rect 13192 32124 13256 32128
rect 13192 32068 13196 32124
rect 13196 32068 13252 32124
rect 13252 32068 13256 32124
rect 13192 32064 13256 32068
rect 22952 32124 23016 32128
rect 22952 32068 22956 32124
rect 22956 32068 23012 32124
rect 23012 32068 23016 32124
rect 22952 32064 23016 32068
rect 23032 32124 23096 32128
rect 23032 32068 23036 32124
rect 23036 32068 23092 32124
rect 23092 32068 23096 32124
rect 23032 32064 23096 32068
rect 23112 32124 23176 32128
rect 23112 32068 23116 32124
rect 23116 32068 23172 32124
rect 23172 32068 23176 32124
rect 23112 32064 23176 32068
rect 23192 32124 23256 32128
rect 23192 32068 23196 32124
rect 23196 32068 23252 32124
rect 23252 32068 23256 32124
rect 23192 32064 23256 32068
rect 7952 31580 8016 31584
rect 7952 31524 7956 31580
rect 7956 31524 8012 31580
rect 8012 31524 8016 31580
rect 7952 31520 8016 31524
rect 8032 31580 8096 31584
rect 8032 31524 8036 31580
rect 8036 31524 8092 31580
rect 8092 31524 8096 31580
rect 8032 31520 8096 31524
rect 8112 31580 8176 31584
rect 8112 31524 8116 31580
rect 8116 31524 8172 31580
rect 8172 31524 8176 31580
rect 8112 31520 8176 31524
rect 8192 31580 8256 31584
rect 8192 31524 8196 31580
rect 8196 31524 8252 31580
rect 8252 31524 8256 31580
rect 8192 31520 8256 31524
rect 17952 31580 18016 31584
rect 17952 31524 17956 31580
rect 17956 31524 18012 31580
rect 18012 31524 18016 31580
rect 17952 31520 18016 31524
rect 18032 31580 18096 31584
rect 18032 31524 18036 31580
rect 18036 31524 18092 31580
rect 18092 31524 18096 31580
rect 18032 31520 18096 31524
rect 18112 31580 18176 31584
rect 18112 31524 18116 31580
rect 18116 31524 18172 31580
rect 18172 31524 18176 31580
rect 18112 31520 18176 31524
rect 18192 31580 18256 31584
rect 18192 31524 18196 31580
rect 18196 31524 18252 31580
rect 18252 31524 18256 31580
rect 18192 31520 18256 31524
rect 2952 31036 3016 31040
rect 2952 30980 2956 31036
rect 2956 30980 3012 31036
rect 3012 30980 3016 31036
rect 2952 30976 3016 30980
rect 3032 31036 3096 31040
rect 3032 30980 3036 31036
rect 3036 30980 3092 31036
rect 3092 30980 3096 31036
rect 3032 30976 3096 30980
rect 3112 31036 3176 31040
rect 3112 30980 3116 31036
rect 3116 30980 3172 31036
rect 3172 30980 3176 31036
rect 3112 30976 3176 30980
rect 3192 31036 3256 31040
rect 3192 30980 3196 31036
rect 3196 30980 3252 31036
rect 3252 30980 3256 31036
rect 3192 30976 3256 30980
rect 12952 31036 13016 31040
rect 12952 30980 12956 31036
rect 12956 30980 13012 31036
rect 13012 30980 13016 31036
rect 12952 30976 13016 30980
rect 13032 31036 13096 31040
rect 13032 30980 13036 31036
rect 13036 30980 13092 31036
rect 13092 30980 13096 31036
rect 13032 30976 13096 30980
rect 13112 31036 13176 31040
rect 13112 30980 13116 31036
rect 13116 30980 13172 31036
rect 13172 30980 13176 31036
rect 13112 30976 13176 30980
rect 13192 31036 13256 31040
rect 13192 30980 13196 31036
rect 13196 30980 13252 31036
rect 13252 30980 13256 31036
rect 13192 30976 13256 30980
rect 22952 31036 23016 31040
rect 22952 30980 22956 31036
rect 22956 30980 23012 31036
rect 23012 30980 23016 31036
rect 22952 30976 23016 30980
rect 23032 31036 23096 31040
rect 23032 30980 23036 31036
rect 23036 30980 23092 31036
rect 23092 30980 23096 31036
rect 23032 30976 23096 30980
rect 23112 31036 23176 31040
rect 23112 30980 23116 31036
rect 23116 30980 23172 31036
rect 23172 30980 23176 31036
rect 23112 30976 23176 30980
rect 23192 31036 23256 31040
rect 23192 30980 23196 31036
rect 23196 30980 23252 31036
rect 23252 30980 23256 31036
rect 23192 30976 23256 30980
rect 7952 30492 8016 30496
rect 7952 30436 7956 30492
rect 7956 30436 8012 30492
rect 8012 30436 8016 30492
rect 7952 30432 8016 30436
rect 8032 30492 8096 30496
rect 8032 30436 8036 30492
rect 8036 30436 8092 30492
rect 8092 30436 8096 30492
rect 8032 30432 8096 30436
rect 8112 30492 8176 30496
rect 8112 30436 8116 30492
rect 8116 30436 8172 30492
rect 8172 30436 8176 30492
rect 8112 30432 8176 30436
rect 8192 30492 8256 30496
rect 8192 30436 8196 30492
rect 8196 30436 8252 30492
rect 8252 30436 8256 30492
rect 8192 30432 8256 30436
rect 17952 30492 18016 30496
rect 17952 30436 17956 30492
rect 17956 30436 18012 30492
rect 18012 30436 18016 30492
rect 17952 30432 18016 30436
rect 18032 30492 18096 30496
rect 18032 30436 18036 30492
rect 18036 30436 18092 30492
rect 18092 30436 18096 30492
rect 18032 30432 18096 30436
rect 18112 30492 18176 30496
rect 18112 30436 18116 30492
rect 18116 30436 18172 30492
rect 18172 30436 18176 30492
rect 18112 30432 18176 30436
rect 18192 30492 18256 30496
rect 18192 30436 18196 30492
rect 18196 30436 18252 30492
rect 18252 30436 18256 30492
rect 18192 30432 18256 30436
rect 2952 29948 3016 29952
rect 2952 29892 2956 29948
rect 2956 29892 3012 29948
rect 3012 29892 3016 29948
rect 2952 29888 3016 29892
rect 3032 29948 3096 29952
rect 3032 29892 3036 29948
rect 3036 29892 3092 29948
rect 3092 29892 3096 29948
rect 3032 29888 3096 29892
rect 3112 29948 3176 29952
rect 3112 29892 3116 29948
rect 3116 29892 3172 29948
rect 3172 29892 3176 29948
rect 3112 29888 3176 29892
rect 3192 29948 3256 29952
rect 3192 29892 3196 29948
rect 3196 29892 3252 29948
rect 3252 29892 3256 29948
rect 3192 29888 3256 29892
rect 12952 29948 13016 29952
rect 12952 29892 12956 29948
rect 12956 29892 13012 29948
rect 13012 29892 13016 29948
rect 12952 29888 13016 29892
rect 13032 29948 13096 29952
rect 13032 29892 13036 29948
rect 13036 29892 13092 29948
rect 13092 29892 13096 29948
rect 13032 29888 13096 29892
rect 13112 29948 13176 29952
rect 13112 29892 13116 29948
rect 13116 29892 13172 29948
rect 13172 29892 13176 29948
rect 13112 29888 13176 29892
rect 13192 29948 13256 29952
rect 13192 29892 13196 29948
rect 13196 29892 13252 29948
rect 13252 29892 13256 29948
rect 13192 29888 13256 29892
rect 22952 29948 23016 29952
rect 22952 29892 22956 29948
rect 22956 29892 23012 29948
rect 23012 29892 23016 29948
rect 22952 29888 23016 29892
rect 23032 29948 23096 29952
rect 23032 29892 23036 29948
rect 23036 29892 23092 29948
rect 23092 29892 23096 29948
rect 23032 29888 23096 29892
rect 23112 29948 23176 29952
rect 23112 29892 23116 29948
rect 23116 29892 23172 29948
rect 23172 29892 23176 29948
rect 23112 29888 23176 29892
rect 23192 29948 23256 29952
rect 23192 29892 23196 29948
rect 23196 29892 23252 29948
rect 23252 29892 23256 29948
rect 23192 29888 23256 29892
rect 7952 29404 8016 29408
rect 7952 29348 7956 29404
rect 7956 29348 8012 29404
rect 8012 29348 8016 29404
rect 7952 29344 8016 29348
rect 8032 29404 8096 29408
rect 8032 29348 8036 29404
rect 8036 29348 8092 29404
rect 8092 29348 8096 29404
rect 8032 29344 8096 29348
rect 8112 29404 8176 29408
rect 8112 29348 8116 29404
rect 8116 29348 8172 29404
rect 8172 29348 8176 29404
rect 8112 29344 8176 29348
rect 8192 29404 8256 29408
rect 8192 29348 8196 29404
rect 8196 29348 8252 29404
rect 8252 29348 8256 29404
rect 8192 29344 8256 29348
rect 17952 29404 18016 29408
rect 17952 29348 17956 29404
rect 17956 29348 18012 29404
rect 18012 29348 18016 29404
rect 17952 29344 18016 29348
rect 18032 29404 18096 29408
rect 18032 29348 18036 29404
rect 18036 29348 18092 29404
rect 18092 29348 18096 29404
rect 18032 29344 18096 29348
rect 18112 29404 18176 29408
rect 18112 29348 18116 29404
rect 18116 29348 18172 29404
rect 18172 29348 18176 29404
rect 18112 29344 18176 29348
rect 18192 29404 18256 29408
rect 18192 29348 18196 29404
rect 18196 29348 18252 29404
rect 18252 29348 18256 29404
rect 18192 29344 18256 29348
rect 21220 29140 21284 29204
rect 22692 29004 22756 29068
rect 2952 28860 3016 28864
rect 2952 28804 2956 28860
rect 2956 28804 3012 28860
rect 3012 28804 3016 28860
rect 2952 28800 3016 28804
rect 3032 28860 3096 28864
rect 3032 28804 3036 28860
rect 3036 28804 3092 28860
rect 3092 28804 3096 28860
rect 3032 28800 3096 28804
rect 3112 28860 3176 28864
rect 3112 28804 3116 28860
rect 3116 28804 3172 28860
rect 3172 28804 3176 28860
rect 3112 28800 3176 28804
rect 3192 28860 3256 28864
rect 3192 28804 3196 28860
rect 3196 28804 3252 28860
rect 3252 28804 3256 28860
rect 3192 28800 3256 28804
rect 12952 28860 13016 28864
rect 12952 28804 12956 28860
rect 12956 28804 13012 28860
rect 13012 28804 13016 28860
rect 12952 28800 13016 28804
rect 13032 28860 13096 28864
rect 13032 28804 13036 28860
rect 13036 28804 13092 28860
rect 13092 28804 13096 28860
rect 13032 28800 13096 28804
rect 13112 28860 13176 28864
rect 13112 28804 13116 28860
rect 13116 28804 13172 28860
rect 13172 28804 13176 28860
rect 13112 28800 13176 28804
rect 13192 28860 13256 28864
rect 13192 28804 13196 28860
rect 13196 28804 13252 28860
rect 13252 28804 13256 28860
rect 13192 28800 13256 28804
rect 22952 28860 23016 28864
rect 22952 28804 22956 28860
rect 22956 28804 23012 28860
rect 23012 28804 23016 28860
rect 22952 28800 23016 28804
rect 23032 28860 23096 28864
rect 23032 28804 23036 28860
rect 23036 28804 23092 28860
rect 23092 28804 23096 28860
rect 23032 28800 23096 28804
rect 23112 28860 23176 28864
rect 23112 28804 23116 28860
rect 23116 28804 23172 28860
rect 23172 28804 23176 28860
rect 23112 28800 23176 28804
rect 23192 28860 23256 28864
rect 23192 28804 23196 28860
rect 23196 28804 23252 28860
rect 23252 28804 23256 28860
rect 23192 28800 23256 28804
rect 7952 28316 8016 28320
rect 7952 28260 7956 28316
rect 7956 28260 8012 28316
rect 8012 28260 8016 28316
rect 7952 28256 8016 28260
rect 8032 28316 8096 28320
rect 8032 28260 8036 28316
rect 8036 28260 8092 28316
rect 8092 28260 8096 28316
rect 8032 28256 8096 28260
rect 8112 28316 8176 28320
rect 8112 28260 8116 28316
rect 8116 28260 8172 28316
rect 8172 28260 8176 28316
rect 8112 28256 8176 28260
rect 8192 28316 8256 28320
rect 8192 28260 8196 28316
rect 8196 28260 8252 28316
rect 8252 28260 8256 28316
rect 8192 28256 8256 28260
rect 17952 28316 18016 28320
rect 17952 28260 17956 28316
rect 17956 28260 18012 28316
rect 18012 28260 18016 28316
rect 17952 28256 18016 28260
rect 18032 28316 18096 28320
rect 18032 28260 18036 28316
rect 18036 28260 18092 28316
rect 18092 28260 18096 28316
rect 18032 28256 18096 28260
rect 18112 28316 18176 28320
rect 18112 28260 18116 28316
rect 18116 28260 18172 28316
rect 18172 28260 18176 28316
rect 18112 28256 18176 28260
rect 18192 28316 18256 28320
rect 18192 28260 18196 28316
rect 18196 28260 18252 28316
rect 18252 28260 18256 28316
rect 18192 28256 18256 28260
rect 2952 27772 3016 27776
rect 2952 27716 2956 27772
rect 2956 27716 3012 27772
rect 3012 27716 3016 27772
rect 2952 27712 3016 27716
rect 3032 27772 3096 27776
rect 3032 27716 3036 27772
rect 3036 27716 3092 27772
rect 3092 27716 3096 27772
rect 3032 27712 3096 27716
rect 3112 27772 3176 27776
rect 3112 27716 3116 27772
rect 3116 27716 3172 27772
rect 3172 27716 3176 27772
rect 3112 27712 3176 27716
rect 3192 27772 3256 27776
rect 3192 27716 3196 27772
rect 3196 27716 3252 27772
rect 3252 27716 3256 27772
rect 3192 27712 3256 27716
rect 12952 27772 13016 27776
rect 12952 27716 12956 27772
rect 12956 27716 13012 27772
rect 13012 27716 13016 27772
rect 12952 27712 13016 27716
rect 13032 27772 13096 27776
rect 13032 27716 13036 27772
rect 13036 27716 13092 27772
rect 13092 27716 13096 27772
rect 13032 27712 13096 27716
rect 13112 27772 13176 27776
rect 13112 27716 13116 27772
rect 13116 27716 13172 27772
rect 13172 27716 13176 27772
rect 13112 27712 13176 27716
rect 13192 27772 13256 27776
rect 13192 27716 13196 27772
rect 13196 27716 13252 27772
rect 13252 27716 13256 27772
rect 13192 27712 13256 27716
rect 22952 27772 23016 27776
rect 22952 27716 22956 27772
rect 22956 27716 23012 27772
rect 23012 27716 23016 27772
rect 22952 27712 23016 27716
rect 23032 27772 23096 27776
rect 23032 27716 23036 27772
rect 23036 27716 23092 27772
rect 23092 27716 23096 27772
rect 23032 27712 23096 27716
rect 23112 27772 23176 27776
rect 23112 27716 23116 27772
rect 23116 27716 23172 27772
rect 23172 27716 23176 27772
rect 23112 27712 23176 27716
rect 23192 27772 23256 27776
rect 23192 27716 23196 27772
rect 23196 27716 23252 27772
rect 23252 27716 23256 27772
rect 23192 27712 23256 27716
rect 17724 27296 17788 27300
rect 17724 27240 17738 27296
rect 17738 27240 17788 27296
rect 17724 27236 17788 27240
rect 7952 27228 8016 27232
rect 7952 27172 7956 27228
rect 7956 27172 8012 27228
rect 8012 27172 8016 27228
rect 7952 27168 8016 27172
rect 8032 27228 8096 27232
rect 8032 27172 8036 27228
rect 8036 27172 8092 27228
rect 8092 27172 8096 27228
rect 8032 27168 8096 27172
rect 8112 27228 8176 27232
rect 8112 27172 8116 27228
rect 8116 27172 8172 27228
rect 8172 27172 8176 27228
rect 8112 27168 8176 27172
rect 8192 27228 8256 27232
rect 8192 27172 8196 27228
rect 8196 27172 8252 27228
rect 8252 27172 8256 27228
rect 8192 27168 8256 27172
rect 17952 27228 18016 27232
rect 17952 27172 17956 27228
rect 17956 27172 18012 27228
rect 18012 27172 18016 27228
rect 17952 27168 18016 27172
rect 18032 27228 18096 27232
rect 18032 27172 18036 27228
rect 18036 27172 18092 27228
rect 18092 27172 18096 27228
rect 18032 27168 18096 27172
rect 18112 27228 18176 27232
rect 18112 27172 18116 27228
rect 18116 27172 18172 27228
rect 18172 27172 18176 27228
rect 18112 27168 18176 27172
rect 18192 27228 18256 27232
rect 18192 27172 18196 27228
rect 18196 27172 18252 27228
rect 18252 27172 18256 27228
rect 18192 27168 18256 27172
rect 2952 26684 3016 26688
rect 2952 26628 2956 26684
rect 2956 26628 3012 26684
rect 3012 26628 3016 26684
rect 2952 26624 3016 26628
rect 3032 26684 3096 26688
rect 3032 26628 3036 26684
rect 3036 26628 3092 26684
rect 3092 26628 3096 26684
rect 3032 26624 3096 26628
rect 3112 26684 3176 26688
rect 3112 26628 3116 26684
rect 3116 26628 3172 26684
rect 3172 26628 3176 26684
rect 3112 26624 3176 26628
rect 3192 26684 3256 26688
rect 3192 26628 3196 26684
rect 3196 26628 3252 26684
rect 3252 26628 3256 26684
rect 3192 26624 3256 26628
rect 12952 26684 13016 26688
rect 12952 26628 12956 26684
rect 12956 26628 13012 26684
rect 13012 26628 13016 26684
rect 12952 26624 13016 26628
rect 13032 26684 13096 26688
rect 13032 26628 13036 26684
rect 13036 26628 13092 26684
rect 13092 26628 13096 26684
rect 13032 26624 13096 26628
rect 13112 26684 13176 26688
rect 13112 26628 13116 26684
rect 13116 26628 13172 26684
rect 13172 26628 13176 26684
rect 13112 26624 13176 26628
rect 13192 26684 13256 26688
rect 13192 26628 13196 26684
rect 13196 26628 13252 26684
rect 13252 26628 13256 26684
rect 13192 26624 13256 26628
rect 22952 26684 23016 26688
rect 22952 26628 22956 26684
rect 22956 26628 23012 26684
rect 23012 26628 23016 26684
rect 22952 26624 23016 26628
rect 23032 26684 23096 26688
rect 23032 26628 23036 26684
rect 23036 26628 23092 26684
rect 23092 26628 23096 26684
rect 23032 26624 23096 26628
rect 23112 26684 23176 26688
rect 23112 26628 23116 26684
rect 23116 26628 23172 26684
rect 23172 26628 23176 26684
rect 23112 26624 23176 26628
rect 23192 26684 23256 26688
rect 23192 26628 23196 26684
rect 23196 26628 23252 26684
rect 23252 26628 23256 26684
rect 23192 26624 23256 26628
rect 18644 26284 18708 26348
rect 7952 26140 8016 26144
rect 7952 26084 7956 26140
rect 7956 26084 8012 26140
rect 8012 26084 8016 26140
rect 7952 26080 8016 26084
rect 8032 26140 8096 26144
rect 8032 26084 8036 26140
rect 8036 26084 8092 26140
rect 8092 26084 8096 26140
rect 8032 26080 8096 26084
rect 8112 26140 8176 26144
rect 8112 26084 8116 26140
rect 8116 26084 8172 26140
rect 8172 26084 8176 26140
rect 8112 26080 8176 26084
rect 8192 26140 8256 26144
rect 8192 26084 8196 26140
rect 8196 26084 8252 26140
rect 8252 26084 8256 26140
rect 8192 26080 8256 26084
rect 17952 26140 18016 26144
rect 17952 26084 17956 26140
rect 17956 26084 18012 26140
rect 18012 26084 18016 26140
rect 17952 26080 18016 26084
rect 18032 26140 18096 26144
rect 18032 26084 18036 26140
rect 18036 26084 18092 26140
rect 18092 26084 18096 26140
rect 18032 26080 18096 26084
rect 18112 26140 18176 26144
rect 18112 26084 18116 26140
rect 18116 26084 18172 26140
rect 18172 26084 18176 26140
rect 18112 26080 18176 26084
rect 18192 26140 18256 26144
rect 18192 26084 18196 26140
rect 18196 26084 18252 26140
rect 18252 26084 18256 26140
rect 18192 26080 18256 26084
rect 22140 25800 22204 25804
rect 22140 25744 22190 25800
rect 22190 25744 22204 25800
rect 22140 25740 22204 25744
rect 2952 25596 3016 25600
rect 2952 25540 2956 25596
rect 2956 25540 3012 25596
rect 3012 25540 3016 25596
rect 2952 25536 3016 25540
rect 3032 25596 3096 25600
rect 3032 25540 3036 25596
rect 3036 25540 3092 25596
rect 3092 25540 3096 25596
rect 3032 25536 3096 25540
rect 3112 25596 3176 25600
rect 3112 25540 3116 25596
rect 3116 25540 3172 25596
rect 3172 25540 3176 25596
rect 3112 25536 3176 25540
rect 3192 25596 3256 25600
rect 3192 25540 3196 25596
rect 3196 25540 3252 25596
rect 3252 25540 3256 25596
rect 3192 25536 3256 25540
rect 12952 25596 13016 25600
rect 12952 25540 12956 25596
rect 12956 25540 13012 25596
rect 13012 25540 13016 25596
rect 12952 25536 13016 25540
rect 13032 25596 13096 25600
rect 13032 25540 13036 25596
rect 13036 25540 13092 25596
rect 13092 25540 13096 25596
rect 13032 25536 13096 25540
rect 13112 25596 13176 25600
rect 13112 25540 13116 25596
rect 13116 25540 13172 25596
rect 13172 25540 13176 25596
rect 13112 25536 13176 25540
rect 13192 25596 13256 25600
rect 13192 25540 13196 25596
rect 13196 25540 13252 25596
rect 13252 25540 13256 25596
rect 13192 25536 13256 25540
rect 22952 25596 23016 25600
rect 22952 25540 22956 25596
rect 22956 25540 23012 25596
rect 23012 25540 23016 25596
rect 22952 25536 23016 25540
rect 23032 25596 23096 25600
rect 23032 25540 23036 25596
rect 23036 25540 23092 25596
rect 23092 25540 23096 25596
rect 23032 25536 23096 25540
rect 23112 25596 23176 25600
rect 23112 25540 23116 25596
rect 23116 25540 23172 25596
rect 23172 25540 23176 25596
rect 23112 25536 23176 25540
rect 23192 25596 23256 25600
rect 23192 25540 23196 25596
rect 23196 25540 23252 25596
rect 23252 25540 23256 25596
rect 23192 25536 23256 25540
rect 15332 25120 15396 25124
rect 15332 25064 15382 25120
rect 15382 25064 15396 25120
rect 15332 25060 15396 25064
rect 19380 25120 19444 25124
rect 19380 25064 19394 25120
rect 19394 25064 19444 25120
rect 19380 25060 19444 25064
rect 7952 25052 8016 25056
rect 7952 24996 7956 25052
rect 7956 24996 8012 25052
rect 8012 24996 8016 25052
rect 7952 24992 8016 24996
rect 8032 25052 8096 25056
rect 8032 24996 8036 25052
rect 8036 24996 8092 25052
rect 8092 24996 8096 25052
rect 8032 24992 8096 24996
rect 8112 25052 8176 25056
rect 8112 24996 8116 25052
rect 8116 24996 8172 25052
rect 8172 24996 8176 25052
rect 8112 24992 8176 24996
rect 8192 25052 8256 25056
rect 8192 24996 8196 25052
rect 8196 24996 8252 25052
rect 8252 24996 8256 25052
rect 8192 24992 8256 24996
rect 17952 25052 18016 25056
rect 17952 24996 17956 25052
rect 17956 24996 18012 25052
rect 18012 24996 18016 25052
rect 17952 24992 18016 24996
rect 18032 25052 18096 25056
rect 18032 24996 18036 25052
rect 18036 24996 18092 25052
rect 18092 24996 18096 25052
rect 18032 24992 18096 24996
rect 18112 25052 18176 25056
rect 18112 24996 18116 25052
rect 18116 24996 18172 25052
rect 18172 24996 18176 25052
rect 18112 24992 18176 24996
rect 18192 25052 18256 25056
rect 18192 24996 18196 25052
rect 18196 24996 18252 25052
rect 18252 24996 18256 25052
rect 18192 24992 18256 24996
rect 21036 24984 21100 24988
rect 21036 24928 21050 24984
rect 21050 24928 21100 24984
rect 21036 24924 21100 24928
rect 2952 24508 3016 24512
rect 2952 24452 2956 24508
rect 2956 24452 3012 24508
rect 3012 24452 3016 24508
rect 2952 24448 3016 24452
rect 3032 24508 3096 24512
rect 3032 24452 3036 24508
rect 3036 24452 3092 24508
rect 3092 24452 3096 24508
rect 3032 24448 3096 24452
rect 3112 24508 3176 24512
rect 3112 24452 3116 24508
rect 3116 24452 3172 24508
rect 3172 24452 3176 24508
rect 3112 24448 3176 24452
rect 3192 24508 3256 24512
rect 3192 24452 3196 24508
rect 3196 24452 3252 24508
rect 3252 24452 3256 24508
rect 3192 24448 3256 24452
rect 12952 24508 13016 24512
rect 12952 24452 12956 24508
rect 12956 24452 13012 24508
rect 13012 24452 13016 24508
rect 12952 24448 13016 24452
rect 13032 24508 13096 24512
rect 13032 24452 13036 24508
rect 13036 24452 13092 24508
rect 13092 24452 13096 24508
rect 13032 24448 13096 24452
rect 13112 24508 13176 24512
rect 13112 24452 13116 24508
rect 13116 24452 13172 24508
rect 13172 24452 13176 24508
rect 13112 24448 13176 24452
rect 13192 24508 13256 24512
rect 13192 24452 13196 24508
rect 13196 24452 13252 24508
rect 13252 24452 13256 24508
rect 13192 24448 13256 24452
rect 22952 24508 23016 24512
rect 22952 24452 22956 24508
rect 22956 24452 23012 24508
rect 23012 24452 23016 24508
rect 22952 24448 23016 24452
rect 23032 24508 23096 24512
rect 23032 24452 23036 24508
rect 23036 24452 23092 24508
rect 23092 24452 23096 24508
rect 23032 24448 23096 24452
rect 23112 24508 23176 24512
rect 23112 24452 23116 24508
rect 23116 24452 23172 24508
rect 23172 24452 23176 24508
rect 23112 24448 23176 24452
rect 23192 24508 23256 24512
rect 23192 24452 23196 24508
rect 23196 24452 23252 24508
rect 23252 24452 23256 24508
rect 23192 24448 23256 24452
rect 7952 23964 8016 23968
rect 7952 23908 7956 23964
rect 7956 23908 8012 23964
rect 8012 23908 8016 23964
rect 7952 23904 8016 23908
rect 8032 23964 8096 23968
rect 8032 23908 8036 23964
rect 8036 23908 8092 23964
rect 8092 23908 8096 23964
rect 8032 23904 8096 23908
rect 8112 23964 8176 23968
rect 8112 23908 8116 23964
rect 8116 23908 8172 23964
rect 8172 23908 8176 23964
rect 8112 23904 8176 23908
rect 8192 23964 8256 23968
rect 8192 23908 8196 23964
rect 8196 23908 8252 23964
rect 8252 23908 8256 23964
rect 8192 23904 8256 23908
rect 17952 23964 18016 23968
rect 17952 23908 17956 23964
rect 17956 23908 18012 23964
rect 18012 23908 18016 23964
rect 17952 23904 18016 23908
rect 18032 23964 18096 23968
rect 18032 23908 18036 23964
rect 18036 23908 18092 23964
rect 18092 23908 18096 23964
rect 18032 23904 18096 23908
rect 18112 23964 18176 23968
rect 18112 23908 18116 23964
rect 18116 23908 18172 23964
rect 18172 23908 18176 23964
rect 18112 23904 18176 23908
rect 18192 23964 18256 23968
rect 18192 23908 18196 23964
rect 18196 23908 18252 23964
rect 18252 23908 18256 23964
rect 18192 23904 18256 23908
rect 17172 23700 17236 23764
rect 22140 23428 22204 23492
rect 2952 23420 3016 23424
rect 2952 23364 2956 23420
rect 2956 23364 3012 23420
rect 3012 23364 3016 23420
rect 2952 23360 3016 23364
rect 3032 23420 3096 23424
rect 3032 23364 3036 23420
rect 3036 23364 3092 23420
rect 3092 23364 3096 23420
rect 3032 23360 3096 23364
rect 3112 23420 3176 23424
rect 3112 23364 3116 23420
rect 3116 23364 3172 23420
rect 3172 23364 3176 23420
rect 3112 23360 3176 23364
rect 3192 23420 3256 23424
rect 3192 23364 3196 23420
rect 3196 23364 3252 23420
rect 3252 23364 3256 23420
rect 3192 23360 3256 23364
rect 12952 23420 13016 23424
rect 12952 23364 12956 23420
rect 12956 23364 13012 23420
rect 13012 23364 13016 23420
rect 12952 23360 13016 23364
rect 13032 23420 13096 23424
rect 13032 23364 13036 23420
rect 13036 23364 13092 23420
rect 13092 23364 13096 23420
rect 13032 23360 13096 23364
rect 13112 23420 13176 23424
rect 13112 23364 13116 23420
rect 13116 23364 13172 23420
rect 13172 23364 13176 23420
rect 13112 23360 13176 23364
rect 13192 23420 13256 23424
rect 13192 23364 13196 23420
rect 13196 23364 13252 23420
rect 13252 23364 13256 23420
rect 13192 23360 13256 23364
rect 22952 23420 23016 23424
rect 22952 23364 22956 23420
rect 22956 23364 23012 23420
rect 23012 23364 23016 23420
rect 22952 23360 23016 23364
rect 23032 23420 23096 23424
rect 23032 23364 23036 23420
rect 23036 23364 23092 23420
rect 23092 23364 23096 23420
rect 23032 23360 23096 23364
rect 23112 23420 23176 23424
rect 23112 23364 23116 23420
rect 23116 23364 23172 23420
rect 23172 23364 23176 23420
rect 23112 23360 23176 23364
rect 23192 23420 23256 23424
rect 23192 23364 23196 23420
rect 23196 23364 23252 23420
rect 23252 23364 23256 23420
rect 23192 23360 23256 23364
rect 7952 22876 8016 22880
rect 7952 22820 7956 22876
rect 7956 22820 8012 22876
rect 8012 22820 8016 22876
rect 7952 22816 8016 22820
rect 8032 22876 8096 22880
rect 8032 22820 8036 22876
rect 8036 22820 8092 22876
rect 8092 22820 8096 22876
rect 8032 22816 8096 22820
rect 8112 22876 8176 22880
rect 8112 22820 8116 22876
rect 8116 22820 8172 22876
rect 8172 22820 8176 22876
rect 8112 22816 8176 22820
rect 8192 22876 8256 22880
rect 8192 22820 8196 22876
rect 8196 22820 8252 22876
rect 8252 22820 8256 22876
rect 8192 22816 8256 22820
rect 17952 22876 18016 22880
rect 17952 22820 17956 22876
rect 17956 22820 18012 22876
rect 18012 22820 18016 22876
rect 17952 22816 18016 22820
rect 18032 22876 18096 22880
rect 18032 22820 18036 22876
rect 18036 22820 18092 22876
rect 18092 22820 18096 22876
rect 18032 22816 18096 22820
rect 18112 22876 18176 22880
rect 18112 22820 18116 22876
rect 18116 22820 18172 22876
rect 18172 22820 18176 22876
rect 18112 22816 18176 22820
rect 18192 22876 18256 22880
rect 18192 22820 18196 22876
rect 18196 22820 18252 22876
rect 18252 22820 18256 22876
rect 18192 22816 18256 22820
rect 2952 22332 3016 22336
rect 2952 22276 2956 22332
rect 2956 22276 3012 22332
rect 3012 22276 3016 22332
rect 2952 22272 3016 22276
rect 3032 22332 3096 22336
rect 3032 22276 3036 22332
rect 3036 22276 3092 22332
rect 3092 22276 3096 22332
rect 3032 22272 3096 22276
rect 3112 22332 3176 22336
rect 3112 22276 3116 22332
rect 3116 22276 3172 22332
rect 3172 22276 3176 22332
rect 3112 22272 3176 22276
rect 3192 22332 3256 22336
rect 3192 22276 3196 22332
rect 3196 22276 3252 22332
rect 3252 22276 3256 22332
rect 3192 22272 3256 22276
rect 12952 22332 13016 22336
rect 12952 22276 12956 22332
rect 12956 22276 13012 22332
rect 13012 22276 13016 22332
rect 12952 22272 13016 22276
rect 13032 22332 13096 22336
rect 13032 22276 13036 22332
rect 13036 22276 13092 22332
rect 13092 22276 13096 22332
rect 13032 22272 13096 22276
rect 13112 22332 13176 22336
rect 13112 22276 13116 22332
rect 13116 22276 13172 22332
rect 13172 22276 13176 22332
rect 13112 22272 13176 22276
rect 13192 22332 13256 22336
rect 13192 22276 13196 22332
rect 13196 22276 13252 22332
rect 13252 22276 13256 22332
rect 13192 22272 13256 22276
rect 22952 22332 23016 22336
rect 22952 22276 22956 22332
rect 22956 22276 23012 22332
rect 23012 22276 23016 22332
rect 22952 22272 23016 22276
rect 23032 22332 23096 22336
rect 23032 22276 23036 22332
rect 23036 22276 23092 22332
rect 23092 22276 23096 22332
rect 23032 22272 23096 22276
rect 23112 22332 23176 22336
rect 23112 22276 23116 22332
rect 23116 22276 23172 22332
rect 23172 22276 23176 22332
rect 23112 22272 23176 22276
rect 23192 22332 23256 22336
rect 23192 22276 23196 22332
rect 23196 22276 23252 22332
rect 23252 22276 23256 22332
rect 23192 22272 23256 22276
rect 7952 21788 8016 21792
rect 7952 21732 7956 21788
rect 7956 21732 8012 21788
rect 8012 21732 8016 21788
rect 7952 21728 8016 21732
rect 8032 21788 8096 21792
rect 8032 21732 8036 21788
rect 8036 21732 8092 21788
rect 8092 21732 8096 21788
rect 8032 21728 8096 21732
rect 8112 21788 8176 21792
rect 8112 21732 8116 21788
rect 8116 21732 8172 21788
rect 8172 21732 8176 21788
rect 8112 21728 8176 21732
rect 8192 21788 8256 21792
rect 8192 21732 8196 21788
rect 8196 21732 8252 21788
rect 8252 21732 8256 21788
rect 8192 21728 8256 21732
rect 17952 21788 18016 21792
rect 17952 21732 17956 21788
rect 17956 21732 18012 21788
rect 18012 21732 18016 21788
rect 17952 21728 18016 21732
rect 18032 21788 18096 21792
rect 18032 21732 18036 21788
rect 18036 21732 18092 21788
rect 18092 21732 18096 21788
rect 18032 21728 18096 21732
rect 18112 21788 18176 21792
rect 18112 21732 18116 21788
rect 18116 21732 18172 21788
rect 18172 21732 18176 21788
rect 18112 21728 18176 21732
rect 18192 21788 18256 21792
rect 18192 21732 18196 21788
rect 18196 21732 18252 21788
rect 18252 21732 18256 21788
rect 18192 21728 18256 21732
rect 2952 21244 3016 21248
rect 2952 21188 2956 21244
rect 2956 21188 3012 21244
rect 3012 21188 3016 21244
rect 2952 21184 3016 21188
rect 3032 21244 3096 21248
rect 3032 21188 3036 21244
rect 3036 21188 3092 21244
rect 3092 21188 3096 21244
rect 3032 21184 3096 21188
rect 3112 21244 3176 21248
rect 3112 21188 3116 21244
rect 3116 21188 3172 21244
rect 3172 21188 3176 21244
rect 3112 21184 3176 21188
rect 3192 21244 3256 21248
rect 3192 21188 3196 21244
rect 3196 21188 3252 21244
rect 3252 21188 3256 21244
rect 3192 21184 3256 21188
rect 12952 21244 13016 21248
rect 12952 21188 12956 21244
rect 12956 21188 13012 21244
rect 13012 21188 13016 21244
rect 12952 21184 13016 21188
rect 13032 21244 13096 21248
rect 13032 21188 13036 21244
rect 13036 21188 13092 21244
rect 13092 21188 13096 21244
rect 13032 21184 13096 21188
rect 13112 21244 13176 21248
rect 13112 21188 13116 21244
rect 13116 21188 13172 21244
rect 13172 21188 13176 21244
rect 13112 21184 13176 21188
rect 13192 21244 13256 21248
rect 13192 21188 13196 21244
rect 13196 21188 13252 21244
rect 13252 21188 13256 21244
rect 13192 21184 13256 21188
rect 22952 21244 23016 21248
rect 22952 21188 22956 21244
rect 22956 21188 23012 21244
rect 23012 21188 23016 21244
rect 22952 21184 23016 21188
rect 23032 21244 23096 21248
rect 23032 21188 23036 21244
rect 23036 21188 23092 21244
rect 23092 21188 23096 21244
rect 23032 21184 23096 21188
rect 23112 21244 23176 21248
rect 23112 21188 23116 21244
rect 23116 21188 23172 21244
rect 23172 21188 23176 21244
rect 23112 21184 23176 21188
rect 23192 21244 23256 21248
rect 23192 21188 23196 21244
rect 23196 21188 23252 21244
rect 23252 21188 23256 21244
rect 23192 21184 23256 21188
rect 7952 20700 8016 20704
rect 7952 20644 7956 20700
rect 7956 20644 8012 20700
rect 8012 20644 8016 20700
rect 7952 20640 8016 20644
rect 8032 20700 8096 20704
rect 8032 20644 8036 20700
rect 8036 20644 8092 20700
rect 8092 20644 8096 20700
rect 8032 20640 8096 20644
rect 8112 20700 8176 20704
rect 8112 20644 8116 20700
rect 8116 20644 8172 20700
rect 8172 20644 8176 20700
rect 8112 20640 8176 20644
rect 8192 20700 8256 20704
rect 8192 20644 8196 20700
rect 8196 20644 8252 20700
rect 8252 20644 8256 20700
rect 8192 20640 8256 20644
rect 17952 20700 18016 20704
rect 17952 20644 17956 20700
rect 17956 20644 18012 20700
rect 18012 20644 18016 20700
rect 17952 20640 18016 20644
rect 18032 20700 18096 20704
rect 18032 20644 18036 20700
rect 18036 20644 18092 20700
rect 18092 20644 18096 20700
rect 18032 20640 18096 20644
rect 18112 20700 18176 20704
rect 18112 20644 18116 20700
rect 18116 20644 18172 20700
rect 18172 20644 18176 20700
rect 18112 20640 18176 20644
rect 18192 20700 18256 20704
rect 18192 20644 18196 20700
rect 18196 20644 18252 20700
rect 18252 20644 18256 20700
rect 18192 20640 18256 20644
rect 2952 20156 3016 20160
rect 2952 20100 2956 20156
rect 2956 20100 3012 20156
rect 3012 20100 3016 20156
rect 2952 20096 3016 20100
rect 3032 20156 3096 20160
rect 3032 20100 3036 20156
rect 3036 20100 3092 20156
rect 3092 20100 3096 20156
rect 3032 20096 3096 20100
rect 3112 20156 3176 20160
rect 3112 20100 3116 20156
rect 3116 20100 3172 20156
rect 3172 20100 3176 20156
rect 3112 20096 3176 20100
rect 3192 20156 3256 20160
rect 3192 20100 3196 20156
rect 3196 20100 3252 20156
rect 3252 20100 3256 20156
rect 3192 20096 3256 20100
rect 12952 20156 13016 20160
rect 12952 20100 12956 20156
rect 12956 20100 13012 20156
rect 13012 20100 13016 20156
rect 12952 20096 13016 20100
rect 13032 20156 13096 20160
rect 13032 20100 13036 20156
rect 13036 20100 13092 20156
rect 13092 20100 13096 20156
rect 13032 20096 13096 20100
rect 13112 20156 13176 20160
rect 13112 20100 13116 20156
rect 13116 20100 13172 20156
rect 13172 20100 13176 20156
rect 13112 20096 13176 20100
rect 13192 20156 13256 20160
rect 13192 20100 13196 20156
rect 13196 20100 13252 20156
rect 13252 20100 13256 20156
rect 13192 20096 13256 20100
rect 22952 20156 23016 20160
rect 22952 20100 22956 20156
rect 22956 20100 23012 20156
rect 23012 20100 23016 20156
rect 22952 20096 23016 20100
rect 23032 20156 23096 20160
rect 23032 20100 23036 20156
rect 23036 20100 23092 20156
rect 23092 20100 23096 20156
rect 23032 20096 23096 20100
rect 23112 20156 23176 20160
rect 23112 20100 23116 20156
rect 23116 20100 23172 20156
rect 23172 20100 23176 20156
rect 23112 20096 23176 20100
rect 23192 20156 23256 20160
rect 23192 20100 23196 20156
rect 23196 20100 23252 20156
rect 23252 20100 23256 20156
rect 23192 20096 23256 20100
rect 7952 19612 8016 19616
rect 7952 19556 7956 19612
rect 7956 19556 8012 19612
rect 8012 19556 8016 19612
rect 7952 19552 8016 19556
rect 8032 19612 8096 19616
rect 8032 19556 8036 19612
rect 8036 19556 8092 19612
rect 8092 19556 8096 19612
rect 8032 19552 8096 19556
rect 8112 19612 8176 19616
rect 8112 19556 8116 19612
rect 8116 19556 8172 19612
rect 8172 19556 8176 19612
rect 8112 19552 8176 19556
rect 8192 19612 8256 19616
rect 8192 19556 8196 19612
rect 8196 19556 8252 19612
rect 8252 19556 8256 19612
rect 8192 19552 8256 19556
rect 17952 19612 18016 19616
rect 17952 19556 17956 19612
rect 17956 19556 18012 19612
rect 18012 19556 18016 19612
rect 17952 19552 18016 19556
rect 18032 19612 18096 19616
rect 18032 19556 18036 19612
rect 18036 19556 18092 19612
rect 18092 19556 18096 19612
rect 18032 19552 18096 19556
rect 18112 19612 18176 19616
rect 18112 19556 18116 19612
rect 18116 19556 18172 19612
rect 18172 19556 18176 19612
rect 18112 19552 18176 19556
rect 18192 19612 18256 19616
rect 18192 19556 18196 19612
rect 18196 19556 18252 19612
rect 18252 19556 18256 19612
rect 18192 19552 18256 19556
rect 19196 19348 19260 19412
rect 2952 19068 3016 19072
rect 2952 19012 2956 19068
rect 2956 19012 3012 19068
rect 3012 19012 3016 19068
rect 2952 19008 3016 19012
rect 3032 19068 3096 19072
rect 3032 19012 3036 19068
rect 3036 19012 3092 19068
rect 3092 19012 3096 19068
rect 3032 19008 3096 19012
rect 3112 19068 3176 19072
rect 3112 19012 3116 19068
rect 3116 19012 3172 19068
rect 3172 19012 3176 19068
rect 3112 19008 3176 19012
rect 3192 19068 3256 19072
rect 3192 19012 3196 19068
rect 3196 19012 3252 19068
rect 3252 19012 3256 19068
rect 3192 19008 3256 19012
rect 12952 19068 13016 19072
rect 12952 19012 12956 19068
rect 12956 19012 13012 19068
rect 13012 19012 13016 19068
rect 12952 19008 13016 19012
rect 13032 19068 13096 19072
rect 13032 19012 13036 19068
rect 13036 19012 13092 19068
rect 13092 19012 13096 19068
rect 13032 19008 13096 19012
rect 13112 19068 13176 19072
rect 13112 19012 13116 19068
rect 13116 19012 13172 19068
rect 13172 19012 13176 19068
rect 13112 19008 13176 19012
rect 13192 19068 13256 19072
rect 13192 19012 13196 19068
rect 13196 19012 13252 19068
rect 13252 19012 13256 19068
rect 13192 19008 13256 19012
rect 22952 19068 23016 19072
rect 22952 19012 22956 19068
rect 22956 19012 23012 19068
rect 23012 19012 23016 19068
rect 22952 19008 23016 19012
rect 23032 19068 23096 19072
rect 23032 19012 23036 19068
rect 23036 19012 23092 19068
rect 23092 19012 23096 19068
rect 23032 19008 23096 19012
rect 23112 19068 23176 19072
rect 23112 19012 23116 19068
rect 23116 19012 23172 19068
rect 23172 19012 23176 19068
rect 23112 19008 23176 19012
rect 23192 19068 23256 19072
rect 23192 19012 23196 19068
rect 23196 19012 23252 19068
rect 23252 19012 23256 19068
rect 23192 19008 23256 19012
rect 7952 18524 8016 18528
rect 7952 18468 7956 18524
rect 7956 18468 8012 18524
rect 8012 18468 8016 18524
rect 7952 18464 8016 18468
rect 8032 18524 8096 18528
rect 8032 18468 8036 18524
rect 8036 18468 8092 18524
rect 8092 18468 8096 18524
rect 8032 18464 8096 18468
rect 8112 18524 8176 18528
rect 8112 18468 8116 18524
rect 8116 18468 8172 18524
rect 8172 18468 8176 18524
rect 8112 18464 8176 18468
rect 8192 18524 8256 18528
rect 8192 18468 8196 18524
rect 8196 18468 8252 18524
rect 8252 18468 8256 18524
rect 8192 18464 8256 18468
rect 17952 18524 18016 18528
rect 17952 18468 17956 18524
rect 17956 18468 18012 18524
rect 18012 18468 18016 18524
rect 17952 18464 18016 18468
rect 18032 18524 18096 18528
rect 18032 18468 18036 18524
rect 18036 18468 18092 18524
rect 18092 18468 18096 18524
rect 18032 18464 18096 18468
rect 18112 18524 18176 18528
rect 18112 18468 18116 18524
rect 18116 18468 18172 18524
rect 18172 18468 18176 18524
rect 18112 18464 18176 18468
rect 18192 18524 18256 18528
rect 18192 18468 18196 18524
rect 18196 18468 18252 18524
rect 18252 18468 18256 18524
rect 18192 18464 18256 18468
rect 18644 18260 18708 18324
rect 18644 18184 18708 18188
rect 18644 18128 18658 18184
rect 18658 18128 18708 18184
rect 18644 18124 18708 18128
rect 21404 18048 21468 18052
rect 21404 17992 21418 18048
rect 21418 17992 21468 18048
rect 21404 17988 21468 17992
rect 2952 17980 3016 17984
rect 2952 17924 2956 17980
rect 2956 17924 3012 17980
rect 3012 17924 3016 17980
rect 2952 17920 3016 17924
rect 3032 17980 3096 17984
rect 3032 17924 3036 17980
rect 3036 17924 3092 17980
rect 3092 17924 3096 17980
rect 3032 17920 3096 17924
rect 3112 17980 3176 17984
rect 3112 17924 3116 17980
rect 3116 17924 3172 17980
rect 3172 17924 3176 17980
rect 3112 17920 3176 17924
rect 3192 17980 3256 17984
rect 3192 17924 3196 17980
rect 3196 17924 3252 17980
rect 3252 17924 3256 17980
rect 3192 17920 3256 17924
rect 12952 17980 13016 17984
rect 12952 17924 12956 17980
rect 12956 17924 13012 17980
rect 13012 17924 13016 17980
rect 12952 17920 13016 17924
rect 13032 17980 13096 17984
rect 13032 17924 13036 17980
rect 13036 17924 13092 17980
rect 13092 17924 13096 17980
rect 13032 17920 13096 17924
rect 13112 17980 13176 17984
rect 13112 17924 13116 17980
rect 13116 17924 13172 17980
rect 13172 17924 13176 17980
rect 13112 17920 13176 17924
rect 13192 17980 13256 17984
rect 13192 17924 13196 17980
rect 13196 17924 13252 17980
rect 13252 17924 13256 17980
rect 13192 17920 13256 17924
rect 22952 17980 23016 17984
rect 22952 17924 22956 17980
rect 22956 17924 23012 17980
rect 23012 17924 23016 17980
rect 22952 17920 23016 17924
rect 23032 17980 23096 17984
rect 23032 17924 23036 17980
rect 23036 17924 23092 17980
rect 23092 17924 23096 17980
rect 23032 17920 23096 17924
rect 23112 17980 23176 17984
rect 23112 17924 23116 17980
rect 23116 17924 23172 17980
rect 23172 17924 23176 17980
rect 23112 17920 23176 17924
rect 23192 17980 23256 17984
rect 23192 17924 23196 17980
rect 23196 17924 23252 17980
rect 23252 17924 23256 17980
rect 23192 17920 23256 17924
rect 7952 17436 8016 17440
rect 7952 17380 7956 17436
rect 7956 17380 8012 17436
rect 8012 17380 8016 17436
rect 7952 17376 8016 17380
rect 8032 17436 8096 17440
rect 8032 17380 8036 17436
rect 8036 17380 8092 17436
rect 8092 17380 8096 17436
rect 8032 17376 8096 17380
rect 8112 17436 8176 17440
rect 8112 17380 8116 17436
rect 8116 17380 8172 17436
rect 8172 17380 8176 17436
rect 8112 17376 8176 17380
rect 8192 17436 8256 17440
rect 8192 17380 8196 17436
rect 8196 17380 8252 17436
rect 8252 17380 8256 17436
rect 8192 17376 8256 17380
rect 17952 17436 18016 17440
rect 17952 17380 17956 17436
rect 17956 17380 18012 17436
rect 18012 17380 18016 17436
rect 17952 17376 18016 17380
rect 18032 17436 18096 17440
rect 18032 17380 18036 17436
rect 18036 17380 18092 17436
rect 18092 17380 18096 17436
rect 18032 17376 18096 17380
rect 18112 17436 18176 17440
rect 18112 17380 18116 17436
rect 18116 17380 18172 17436
rect 18172 17380 18176 17436
rect 18112 17376 18176 17380
rect 18192 17436 18256 17440
rect 18192 17380 18196 17436
rect 18196 17380 18252 17436
rect 18252 17380 18256 17436
rect 18192 17376 18256 17380
rect 21220 17368 21284 17372
rect 21220 17312 21234 17368
rect 21234 17312 21284 17368
rect 21220 17308 21284 17312
rect 16804 17036 16868 17100
rect 22140 17096 22204 17100
rect 22140 17040 22154 17096
rect 22154 17040 22204 17096
rect 22140 17036 22204 17040
rect 2952 16892 3016 16896
rect 2952 16836 2956 16892
rect 2956 16836 3012 16892
rect 3012 16836 3016 16892
rect 2952 16832 3016 16836
rect 3032 16892 3096 16896
rect 3032 16836 3036 16892
rect 3036 16836 3092 16892
rect 3092 16836 3096 16892
rect 3032 16832 3096 16836
rect 3112 16892 3176 16896
rect 3112 16836 3116 16892
rect 3116 16836 3172 16892
rect 3172 16836 3176 16892
rect 3112 16832 3176 16836
rect 3192 16892 3256 16896
rect 3192 16836 3196 16892
rect 3196 16836 3252 16892
rect 3252 16836 3256 16892
rect 3192 16832 3256 16836
rect 12952 16892 13016 16896
rect 12952 16836 12956 16892
rect 12956 16836 13012 16892
rect 13012 16836 13016 16892
rect 12952 16832 13016 16836
rect 13032 16892 13096 16896
rect 13032 16836 13036 16892
rect 13036 16836 13092 16892
rect 13092 16836 13096 16892
rect 13032 16832 13096 16836
rect 13112 16892 13176 16896
rect 13112 16836 13116 16892
rect 13116 16836 13172 16892
rect 13172 16836 13176 16892
rect 13112 16832 13176 16836
rect 13192 16892 13256 16896
rect 13192 16836 13196 16892
rect 13196 16836 13252 16892
rect 13252 16836 13256 16892
rect 13192 16832 13256 16836
rect 22952 16892 23016 16896
rect 22952 16836 22956 16892
rect 22956 16836 23012 16892
rect 23012 16836 23016 16892
rect 22952 16832 23016 16836
rect 23032 16892 23096 16896
rect 23032 16836 23036 16892
rect 23036 16836 23092 16892
rect 23092 16836 23096 16892
rect 23032 16832 23096 16836
rect 23112 16892 23176 16896
rect 23112 16836 23116 16892
rect 23116 16836 23172 16892
rect 23172 16836 23176 16892
rect 23112 16832 23176 16836
rect 23192 16892 23256 16896
rect 23192 16836 23196 16892
rect 23196 16836 23252 16892
rect 23252 16836 23256 16892
rect 23192 16832 23256 16836
rect 13492 16628 13556 16692
rect 19564 16628 19628 16692
rect 13676 16492 13740 16556
rect 7952 16348 8016 16352
rect 7952 16292 7956 16348
rect 7956 16292 8012 16348
rect 8012 16292 8016 16348
rect 7952 16288 8016 16292
rect 8032 16348 8096 16352
rect 8032 16292 8036 16348
rect 8036 16292 8092 16348
rect 8092 16292 8096 16348
rect 8032 16288 8096 16292
rect 8112 16348 8176 16352
rect 8112 16292 8116 16348
rect 8116 16292 8172 16348
rect 8172 16292 8176 16348
rect 8112 16288 8176 16292
rect 8192 16348 8256 16352
rect 8192 16292 8196 16348
rect 8196 16292 8252 16348
rect 8252 16292 8256 16348
rect 8192 16288 8256 16292
rect 17952 16348 18016 16352
rect 17952 16292 17956 16348
rect 17956 16292 18012 16348
rect 18012 16292 18016 16348
rect 17952 16288 18016 16292
rect 18032 16348 18096 16352
rect 18032 16292 18036 16348
rect 18036 16292 18092 16348
rect 18092 16292 18096 16348
rect 18032 16288 18096 16292
rect 18112 16348 18176 16352
rect 18112 16292 18116 16348
rect 18116 16292 18172 16348
rect 18172 16292 18176 16348
rect 18112 16288 18176 16292
rect 18192 16348 18256 16352
rect 18192 16292 18196 16348
rect 18196 16292 18252 16348
rect 18252 16292 18256 16348
rect 18192 16288 18256 16292
rect 17172 16280 17236 16284
rect 17172 16224 17222 16280
rect 17222 16224 17236 16280
rect 17172 16220 17236 16224
rect 2952 15804 3016 15808
rect 2952 15748 2956 15804
rect 2956 15748 3012 15804
rect 3012 15748 3016 15804
rect 2952 15744 3016 15748
rect 3032 15804 3096 15808
rect 3032 15748 3036 15804
rect 3036 15748 3092 15804
rect 3092 15748 3096 15804
rect 3032 15744 3096 15748
rect 3112 15804 3176 15808
rect 3112 15748 3116 15804
rect 3116 15748 3172 15804
rect 3172 15748 3176 15804
rect 3112 15744 3176 15748
rect 3192 15804 3256 15808
rect 3192 15748 3196 15804
rect 3196 15748 3252 15804
rect 3252 15748 3256 15804
rect 3192 15744 3256 15748
rect 12952 15804 13016 15808
rect 12952 15748 12956 15804
rect 12956 15748 13012 15804
rect 13012 15748 13016 15804
rect 12952 15744 13016 15748
rect 13032 15804 13096 15808
rect 13032 15748 13036 15804
rect 13036 15748 13092 15804
rect 13092 15748 13096 15804
rect 13032 15744 13096 15748
rect 13112 15804 13176 15808
rect 13112 15748 13116 15804
rect 13116 15748 13172 15804
rect 13172 15748 13176 15804
rect 13112 15744 13176 15748
rect 13192 15804 13256 15808
rect 13192 15748 13196 15804
rect 13196 15748 13252 15804
rect 13252 15748 13256 15804
rect 13192 15744 13256 15748
rect 22952 15804 23016 15808
rect 22952 15748 22956 15804
rect 22956 15748 23012 15804
rect 23012 15748 23016 15804
rect 22952 15744 23016 15748
rect 23032 15804 23096 15808
rect 23032 15748 23036 15804
rect 23036 15748 23092 15804
rect 23092 15748 23096 15804
rect 23032 15744 23096 15748
rect 23112 15804 23176 15808
rect 23112 15748 23116 15804
rect 23116 15748 23172 15804
rect 23172 15748 23176 15804
rect 23112 15744 23176 15748
rect 23192 15804 23256 15808
rect 23192 15748 23196 15804
rect 23196 15748 23252 15804
rect 23252 15748 23256 15804
rect 23192 15744 23256 15748
rect 13676 15404 13740 15468
rect 17356 15328 17420 15332
rect 17356 15272 17370 15328
rect 17370 15272 17420 15328
rect 17356 15268 17420 15272
rect 7952 15260 8016 15264
rect 7952 15204 7956 15260
rect 7956 15204 8012 15260
rect 8012 15204 8016 15260
rect 7952 15200 8016 15204
rect 8032 15260 8096 15264
rect 8032 15204 8036 15260
rect 8036 15204 8092 15260
rect 8092 15204 8096 15260
rect 8032 15200 8096 15204
rect 8112 15260 8176 15264
rect 8112 15204 8116 15260
rect 8116 15204 8172 15260
rect 8172 15204 8176 15260
rect 8112 15200 8176 15204
rect 8192 15260 8256 15264
rect 8192 15204 8196 15260
rect 8196 15204 8252 15260
rect 8252 15204 8256 15260
rect 8192 15200 8256 15204
rect 17952 15260 18016 15264
rect 17952 15204 17956 15260
rect 17956 15204 18012 15260
rect 18012 15204 18016 15260
rect 17952 15200 18016 15204
rect 18032 15260 18096 15264
rect 18032 15204 18036 15260
rect 18036 15204 18092 15260
rect 18092 15204 18096 15260
rect 18032 15200 18096 15204
rect 18112 15260 18176 15264
rect 18112 15204 18116 15260
rect 18116 15204 18172 15260
rect 18172 15204 18176 15260
rect 18112 15200 18176 15204
rect 18192 15260 18256 15264
rect 18192 15204 18196 15260
rect 18196 15204 18252 15260
rect 18252 15204 18256 15260
rect 18192 15200 18256 15204
rect 2952 14716 3016 14720
rect 2952 14660 2956 14716
rect 2956 14660 3012 14716
rect 3012 14660 3016 14716
rect 2952 14656 3016 14660
rect 3032 14716 3096 14720
rect 3032 14660 3036 14716
rect 3036 14660 3092 14716
rect 3092 14660 3096 14716
rect 3032 14656 3096 14660
rect 3112 14716 3176 14720
rect 3112 14660 3116 14716
rect 3116 14660 3172 14716
rect 3172 14660 3176 14716
rect 3112 14656 3176 14660
rect 3192 14716 3256 14720
rect 3192 14660 3196 14716
rect 3196 14660 3252 14716
rect 3252 14660 3256 14716
rect 3192 14656 3256 14660
rect 12952 14716 13016 14720
rect 12952 14660 12956 14716
rect 12956 14660 13012 14716
rect 13012 14660 13016 14716
rect 12952 14656 13016 14660
rect 13032 14716 13096 14720
rect 13032 14660 13036 14716
rect 13036 14660 13092 14716
rect 13092 14660 13096 14716
rect 13032 14656 13096 14660
rect 13112 14716 13176 14720
rect 13112 14660 13116 14716
rect 13116 14660 13172 14716
rect 13172 14660 13176 14716
rect 13112 14656 13176 14660
rect 13192 14716 13256 14720
rect 13192 14660 13196 14716
rect 13196 14660 13252 14716
rect 13252 14660 13256 14716
rect 13192 14656 13256 14660
rect 22952 14716 23016 14720
rect 22952 14660 22956 14716
rect 22956 14660 23012 14716
rect 23012 14660 23016 14716
rect 22952 14656 23016 14660
rect 23032 14716 23096 14720
rect 23032 14660 23036 14716
rect 23036 14660 23092 14716
rect 23092 14660 23096 14716
rect 23032 14656 23096 14660
rect 23112 14716 23176 14720
rect 23112 14660 23116 14716
rect 23116 14660 23172 14716
rect 23172 14660 23176 14716
rect 23112 14656 23176 14660
rect 23192 14716 23256 14720
rect 23192 14660 23196 14716
rect 23196 14660 23252 14716
rect 23252 14660 23256 14716
rect 23192 14656 23256 14660
rect 16068 14240 16132 14244
rect 16068 14184 16082 14240
rect 16082 14184 16132 14240
rect 16068 14180 16132 14184
rect 7952 14172 8016 14176
rect 7952 14116 7956 14172
rect 7956 14116 8012 14172
rect 8012 14116 8016 14172
rect 7952 14112 8016 14116
rect 8032 14172 8096 14176
rect 8032 14116 8036 14172
rect 8036 14116 8092 14172
rect 8092 14116 8096 14172
rect 8032 14112 8096 14116
rect 8112 14172 8176 14176
rect 8112 14116 8116 14172
rect 8116 14116 8172 14172
rect 8172 14116 8176 14172
rect 8112 14112 8176 14116
rect 8192 14172 8256 14176
rect 8192 14116 8196 14172
rect 8196 14116 8252 14172
rect 8252 14116 8256 14172
rect 8192 14112 8256 14116
rect 17952 14172 18016 14176
rect 17952 14116 17956 14172
rect 17956 14116 18012 14172
rect 18012 14116 18016 14172
rect 17952 14112 18016 14116
rect 18032 14172 18096 14176
rect 18032 14116 18036 14172
rect 18036 14116 18092 14172
rect 18092 14116 18096 14172
rect 18032 14112 18096 14116
rect 18112 14172 18176 14176
rect 18112 14116 18116 14172
rect 18116 14116 18172 14172
rect 18172 14116 18176 14172
rect 18112 14112 18176 14116
rect 18192 14172 18256 14176
rect 18192 14116 18196 14172
rect 18196 14116 18252 14172
rect 18252 14116 18256 14172
rect 18192 14112 18256 14116
rect 2952 13628 3016 13632
rect 2952 13572 2956 13628
rect 2956 13572 3012 13628
rect 3012 13572 3016 13628
rect 2952 13568 3016 13572
rect 3032 13628 3096 13632
rect 3032 13572 3036 13628
rect 3036 13572 3092 13628
rect 3092 13572 3096 13628
rect 3032 13568 3096 13572
rect 3112 13628 3176 13632
rect 3112 13572 3116 13628
rect 3116 13572 3172 13628
rect 3172 13572 3176 13628
rect 3112 13568 3176 13572
rect 3192 13628 3256 13632
rect 3192 13572 3196 13628
rect 3196 13572 3252 13628
rect 3252 13572 3256 13628
rect 3192 13568 3256 13572
rect 12952 13628 13016 13632
rect 12952 13572 12956 13628
rect 12956 13572 13012 13628
rect 13012 13572 13016 13628
rect 12952 13568 13016 13572
rect 13032 13628 13096 13632
rect 13032 13572 13036 13628
rect 13036 13572 13092 13628
rect 13092 13572 13096 13628
rect 13032 13568 13096 13572
rect 13112 13628 13176 13632
rect 13112 13572 13116 13628
rect 13116 13572 13172 13628
rect 13172 13572 13176 13628
rect 13112 13568 13176 13572
rect 13192 13628 13256 13632
rect 13192 13572 13196 13628
rect 13196 13572 13252 13628
rect 13252 13572 13256 13628
rect 13192 13568 13256 13572
rect 22952 13628 23016 13632
rect 22952 13572 22956 13628
rect 22956 13572 23012 13628
rect 23012 13572 23016 13628
rect 22952 13568 23016 13572
rect 23032 13628 23096 13632
rect 23032 13572 23036 13628
rect 23036 13572 23092 13628
rect 23092 13572 23096 13628
rect 23032 13568 23096 13572
rect 23112 13628 23176 13632
rect 23112 13572 23116 13628
rect 23116 13572 23172 13628
rect 23172 13572 23176 13628
rect 23112 13568 23176 13572
rect 23192 13628 23256 13632
rect 23192 13572 23196 13628
rect 23196 13572 23252 13628
rect 23252 13572 23256 13628
rect 23192 13568 23256 13572
rect 19564 13288 19628 13292
rect 19564 13232 19578 13288
rect 19578 13232 19628 13288
rect 19564 13228 19628 13232
rect 7952 13084 8016 13088
rect 7952 13028 7956 13084
rect 7956 13028 8012 13084
rect 8012 13028 8016 13084
rect 7952 13024 8016 13028
rect 8032 13084 8096 13088
rect 8032 13028 8036 13084
rect 8036 13028 8092 13084
rect 8092 13028 8096 13084
rect 8032 13024 8096 13028
rect 8112 13084 8176 13088
rect 8112 13028 8116 13084
rect 8116 13028 8172 13084
rect 8172 13028 8176 13084
rect 8112 13024 8176 13028
rect 8192 13084 8256 13088
rect 8192 13028 8196 13084
rect 8196 13028 8252 13084
rect 8252 13028 8256 13084
rect 8192 13024 8256 13028
rect 17952 13084 18016 13088
rect 17952 13028 17956 13084
rect 17956 13028 18012 13084
rect 18012 13028 18016 13084
rect 17952 13024 18016 13028
rect 18032 13084 18096 13088
rect 18032 13028 18036 13084
rect 18036 13028 18092 13084
rect 18092 13028 18096 13084
rect 18032 13024 18096 13028
rect 18112 13084 18176 13088
rect 18112 13028 18116 13084
rect 18116 13028 18172 13084
rect 18172 13028 18176 13084
rect 18112 13024 18176 13028
rect 18192 13084 18256 13088
rect 18192 13028 18196 13084
rect 18196 13028 18252 13084
rect 18252 13028 18256 13084
rect 18192 13024 18256 13028
rect 22692 12956 22756 13020
rect 18644 12820 18708 12884
rect 20116 12608 20180 12612
rect 20116 12552 20130 12608
rect 20130 12552 20180 12608
rect 20116 12548 20180 12552
rect 2952 12540 3016 12544
rect 2952 12484 2956 12540
rect 2956 12484 3012 12540
rect 3012 12484 3016 12540
rect 2952 12480 3016 12484
rect 3032 12540 3096 12544
rect 3032 12484 3036 12540
rect 3036 12484 3092 12540
rect 3092 12484 3096 12540
rect 3032 12480 3096 12484
rect 3112 12540 3176 12544
rect 3112 12484 3116 12540
rect 3116 12484 3172 12540
rect 3172 12484 3176 12540
rect 3112 12480 3176 12484
rect 3192 12540 3256 12544
rect 3192 12484 3196 12540
rect 3196 12484 3252 12540
rect 3252 12484 3256 12540
rect 3192 12480 3256 12484
rect 12952 12540 13016 12544
rect 12952 12484 12956 12540
rect 12956 12484 13012 12540
rect 13012 12484 13016 12540
rect 12952 12480 13016 12484
rect 13032 12540 13096 12544
rect 13032 12484 13036 12540
rect 13036 12484 13092 12540
rect 13092 12484 13096 12540
rect 13032 12480 13096 12484
rect 13112 12540 13176 12544
rect 13112 12484 13116 12540
rect 13116 12484 13172 12540
rect 13172 12484 13176 12540
rect 13112 12480 13176 12484
rect 13192 12540 13256 12544
rect 13192 12484 13196 12540
rect 13196 12484 13252 12540
rect 13252 12484 13256 12540
rect 13192 12480 13256 12484
rect 22952 12540 23016 12544
rect 22952 12484 22956 12540
rect 22956 12484 23012 12540
rect 23012 12484 23016 12540
rect 22952 12480 23016 12484
rect 23032 12540 23096 12544
rect 23032 12484 23036 12540
rect 23036 12484 23092 12540
rect 23092 12484 23096 12540
rect 23032 12480 23096 12484
rect 23112 12540 23176 12544
rect 23112 12484 23116 12540
rect 23116 12484 23172 12540
rect 23172 12484 23176 12540
rect 23112 12480 23176 12484
rect 23192 12540 23256 12544
rect 23192 12484 23196 12540
rect 23196 12484 23252 12540
rect 23252 12484 23256 12540
rect 23192 12480 23256 12484
rect 7952 11996 8016 12000
rect 7952 11940 7956 11996
rect 7956 11940 8012 11996
rect 8012 11940 8016 11996
rect 7952 11936 8016 11940
rect 8032 11996 8096 12000
rect 8032 11940 8036 11996
rect 8036 11940 8092 11996
rect 8092 11940 8096 11996
rect 8032 11936 8096 11940
rect 8112 11996 8176 12000
rect 8112 11940 8116 11996
rect 8116 11940 8172 11996
rect 8172 11940 8176 11996
rect 8112 11936 8176 11940
rect 8192 11996 8256 12000
rect 8192 11940 8196 11996
rect 8196 11940 8252 11996
rect 8252 11940 8256 11996
rect 8192 11936 8256 11940
rect 17952 11996 18016 12000
rect 17952 11940 17956 11996
rect 17956 11940 18012 11996
rect 18012 11940 18016 11996
rect 17952 11936 18016 11940
rect 18032 11996 18096 12000
rect 18032 11940 18036 11996
rect 18036 11940 18092 11996
rect 18092 11940 18096 11996
rect 18032 11936 18096 11940
rect 18112 11996 18176 12000
rect 18112 11940 18116 11996
rect 18116 11940 18172 11996
rect 18172 11940 18176 11996
rect 18112 11936 18176 11940
rect 18192 11996 18256 12000
rect 18192 11940 18196 11996
rect 18196 11940 18252 11996
rect 18252 11940 18256 11996
rect 18192 11936 18256 11940
rect 13676 11732 13740 11796
rect 14964 11596 15028 11660
rect 18644 11520 18708 11524
rect 18644 11464 18694 11520
rect 18694 11464 18708 11520
rect 18644 11460 18708 11464
rect 2952 11452 3016 11456
rect 2952 11396 2956 11452
rect 2956 11396 3012 11452
rect 3012 11396 3016 11452
rect 2952 11392 3016 11396
rect 3032 11452 3096 11456
rect 3032 11396 3036 11452
rect 3036 11396 3092 11452
rect 3092 11396 3096 11452
rect 3032 11392 3096 11396
rect 3112 11452 3176 11456
rect 3112 11396 3116 11452
rect 3116 11396 3172 11452
rect 3172 11396 3176 11452
rect 3112 11392 3176 11396
rect 3192 11452 3256 11456
rect 3192 11396 3196 11452
rect 3196 11396 3252 11452
rect 3252 11396 3256 11452
rect 3192 11392 3256 11396
rect 12952 11452 13016 11456
rect 12952 11396 12956 11452
rect 12956 11396 13012 11452
rect 13012 11396 13016 11452
rect 12952 11392 13016 11396
rect 13032 11452 13096 11456
rect 13032 11396 13036 11452
rect 13036 11396 13092 11452
rect 13092 11396 13096 11452
rect 13032 11392 13096 11396
rect 13112 11452 13176 11456
rect 13112 11396 13116 11452
rect 13116 11396 13172 11452
rect 13172 11396 13176 11452
rect 13112 11392 13176 11396
rect 13192 11452 13256 11456
rect 13192 11396 13196 11452
rect 13196 11396 13252 11452
rect 13252 11396 13256 11452
rect 13192 11392 13256 11396
rect 22952 11452 23016 11456
rect 22952 11396 22956 11452
rect 22956 11396 23012 11452
rect 23012 11396 23016 11452
rect 22952 11392 23016 11396
rect 23032 11452 23096 11456
rect 23032 11396 23036 11452
rect 23036 11396 23092 11452
rect 23092 11396 23096 11452
rect 23032 11392 23096 11396
rect 23112 11452 23176 11456
rect 23112 11396 23116 11452
rect 23116 11396 23172 11452
rect 23172 11396 23176 11452
rect 23112 11392 23176 11396
rect 23192 11452 23256 11456
rect 23192 11396 23196 11452
rect 23196 11396 23252 11452
rect 23252 11396 23256 11452
rect 23192 11392 23256 11396
rect 7952 10908 8016 10912
rect 7952 10852 7956 10908
rect 7956 10852 8012 10908
rect 8012 10852 8016 10908
rect 7952 10848 8016 10852
rect 8032 10908 8096 10912
rect 8032 10852 8036 10908
rect 8036 10852 8092 10908
rect 8092 10852 8096 10908
rect 8032 10848 8096 10852
rect 8112 10908 8176 10912
rect 8112 10852 8116 10908
rect 8116 10852 8172 10908
rect 8172 10852 8176 10908
rect 8112 10848 8176 10852
rect 8192 10908 8256 10912
rect 8192 10852 8196 10908
rect 8196 10852 8252 10908
rect 8252 10852 8256 10908
rect 8192 10848 8256 10852
rect 17952 10908 18016 10912
rect 17952 10852 17956 10908
rect 17956 10852 18012 10908
rect 18012 10852 18016 10908
rect 17952 10848 18016 10852
rect 18032 10908 18096 10912
rect 18032 10852 18036 10908
rect 18036 10852 18092 10908
rect 18092 10852 18096 10908
rect 18032 10848 18096 10852
rect 18112 10908 18176 10912
rect 18112 10852 18116 10908
rect 18116 10852 18172 10908
rect 18172 10852 18176 10908
rect 18112 10848 18176 10852
rect 18192 10908 18256 10912
rect 18192 10852 18196 10908
rect 18196 10852 18252 10908
rect 18252 10852 18256 10908
rect 18192 10848 18256 10852
rect 17724 10432 17788 10436
rect 17724 10376 17774 10432
rect 17774 10376 17788 10432
rect 17724 10372 17788 10376
rect 2952 10364 3016 10368
rect 2952 10308 2956 10364
rect 2956 10308 3012 10364
rect 3012 10308 3016 10364
rect 2952 10304 3016 10308
rect 3032 10364 3096 10368
rect 3032 10308 3036 10364
rect 3036 10308 3092 10364
rect 3092 10308 3096 10364
rect 3032 10304 3096 10308
rect 3112 10364 3176 10368
rect 3112 10308 3116 10364
rect 3116 10308 3172 10364
rect 3172 10308 3176 10364
rect 3112 10304 3176 10308
rect 3192 10364 3256 10368
rect 3192 10308 3196 10364
rect 3196 10308 3252 10364
rect 3252 10308 3256 10364
rect 3192 10304 3256 10308
rect 12952 10364 13016 10368
rect 12952 10308 12956 10364
rect 12956 10308 13012 10364
rect 13012 10308 13016 10364
rect 12952 10304 13016 10308
rect 13032 10364 13096 10368
rect 13032 10308 13036 10364
rect 13036 10308 13092 10364
rect 13092 10308 13096 10364
rect 13032 10304 13096 10308
rect 13112 10364 13176 10368
rect 13112 10308 13116 10364
rect 13116 10308 13172 10364
rect 13172 10308 13176 10364
rect 13112 10304 13176 10308
rect 13192 10364 13256 10368
rect 13192 10308 13196 10364
rect 13196 10308 13252 10364
rect 13252 10308 13256 10364
rect 13192 10304 13256 10308
rect 22952 10364 23016 10368
rect 22952 10308 22956 10364
rect 22956 10308 23012 10364
rect 23012 10308 23016 10364
rect 22952 10304 23016 10308
rect 23032 10364 23096 10368
rect 23032 10308 23036 10364
rect 23036 10308 23092 10364
rect 23092 10308 23096 10364
rect 23032 10304 23096 10308
rect 23112 10364 23176 10368
rect 23112 10308 23116 10364
rect 23116 10308 23172 10364
rect 23172 10308 23176 10364
rect 23112 10304 23176 10308
rect 23192 10364 23256 10368
rect 23192 10308 23196 10364
rect 23196 10308 23252 10364
rect 23252 10308 23256 10364
rect 23192 10304 23256 10308
rect 16804 10236 16868 10300
rect 14964 9828 15028 9892
rect 7952 9820 8016 9824
rect 7952 9764 7956 9820
rect 7956 9764 8012 9820
rect 8012 9764 8016 9820
rect 7952 9760 8016 9764
rect 8032 9820 8096 9824
rect 8032 9764 8036 9820
rect 8036 9764 8092 9820
rect 8092 9764 8096 9820
rect 8032 9760 8096 9764
rect 8112 9820 8176 9824
rect 8112 9764 8116 9820
rect 8116 9764 8172 9820
rect 8172 9764 8176 9820
rect 8112 9760 8176 9764
rect 8192 9820 8256 9824
rect 8192 9764 8196 9820
rect 8196 9764 8252 9820
rect 8252 9764 8256 9820
rect 8192 9760 8256 9764
rect 17952 9820 18016 9824
rect 17952 9764 17956 9820
rect 17956 9764 18012 9820
rect 18012 9764 18016 9820
rect 17952 9760 18016 9764
rect 18032 9820 18096 9824
rect 18032 9764 18036 9820
rect 18036 9764 18092 9820
rect 18092 9764 18096 9820
rect 18032 9760 18096 9764
rect 18112 9820 18176 9824
rect 18112 9764 18116 9820
rect 18116 9764 18172 9820
rect 18172 9764 18176 9820
rect 18112 9760 18176 9764
rect 18192 9820 18256 9824
rect 18192 9764 18196 9820
rect 18196 9764 18252 9820
rect 18252 9764 18256 9820
rect 18192 9760 18256 9764
rect 19196 9556 19260 9620
rect 2952 9276 3016 9280
rect 2952 9220 2956 9276
rect 2956 9220 3012 9276
rect 3012 9220 3016 9276
rect 2952 9216 3016 9220
rect 3032 9276 3096 9280
rect 3032 9220 3036 9276
rect 3036 9220 3092 9276
rect 3092 9220 3096 9276
rect 3032 9216 3096 9220
rect 3112 9276 3176 9280
rect 3112 9220 3116 9276
rect 3116 9220 3172 9276
rect 3172 9220 3176 9276
rect 3112 9216 3176 9220
rect 3192 9276 3256 9280
rect 3192 9220 3196 9276
rect 3196 9220 3252 9276
rect 3252 9220 3256 9276
rect 3192 9216 3256 9220
rect 12952 9276 13016 9280
rect 12952 9220 12956 9276
rect 12956 9220 13012 9276
rect 13012 9220 13016 9276
rect 12952 9216 13016 9220
rect 13032 9276 13096 9280
rect 13032 9220 13036 9276
rect 13036 9220 13092 9276
rect 13092 9220 13096 9276
rect 13032 9216 13096 9220
rect 13112 9276 13176 9280
rect 13112 9220 13116 9276
rect 13116 9220 13172 9276
rect 13172 9220 13176 9276
rect 13112 9216 13176 9220
rect 13192 9276 13256 9280
rect 13192 9220 13196 9276
rect 13196 9220 13252 9276
rect 13252 9220 13256 9276
rect 13192 9216 13256 9220
rect 22952 9276 23016 9280
rect 22952 9220 22956 9276
rect 22956 9220 23012 9276
rect 23012 9220 23016 9276
rect 22952 9216 23016 9220
rect 23032 9276 23096 9280
rect 23032 9220 23036 9276
rect 23036 9220 23092 9276
rect 23092 9220 23096 9276
rect 23032 9216 23096 9220
rect 23112 9276 23176 9280
rect 23112 9220 23116 9276
rect 23116 9220 23172 9276
rect 23172 9220 23176 9276
rect 23112 9216 23176 9220
rect 23192 9276 23256 9280
rect 23192 9220 23196 9276
rect 23196 9220 23252 9276
rect 23252 9220 23256 9276
rect 23192 9216 23256 9220
rect 7952 8732 8016 8736
rect 7952 8676 7956 8732
rect 7956 8676 8012 8732
rect 8012 8676 8016 8732
rect 7952 8672 8016 8676
rect 8032 8732 8096 8736
rect 8032 8676 8036 8732
rect 8036 8676 8092 8732
rect 8092 8676 8096 8732
rect 8032 8672 8096 8676
rect 8112 8732 8176 8736
rect 8112 8676 8116 8732
rect 8116 8676 8172 8732
rect 8172 8676 8176 8732
rect 8112 8672 8176 8676
rect 8192 8732 8256 8736
rect 8192 8676 8196 8732
rect 8196 8676 8252 8732
rect 8252 8676 8256 8732
rect 8192 8672 8256 8676
rect 17952 8732 18016 8736
rect 17952 8676 17956 8732
rect 17956 8676 18012 8732
rect 18012 8676 18016 8732
rect 17952 8672 18016 8676
rect 18032 8732 18096 8736
rect 18032 8676 18036 8732
rect 18036 8676 18092 8732
rect 18092 8676 18096 8732
rect 18032 8672 18096 8676
rect 18112 8732 18176 8736
rect 18112 8676 18116 8732
rect 18116 8676 18172 8732
rect 18172 8676 18176 8732
rect 18112 8672 18176 8676
rect 18192 8732 18256 8736
rect 18192 8676 18196 8732
rect 18196 8676 18252 8732
rect 18252 8676 18256 8732
rect 18192 8672 18256 8676
rect 19564 8392 19628 8396
rect 19564 8336 19614 8392
rect 19614 8336 19628 8392
rect 19564 8332 19628 8336
rect 2952 8188 3016 8192
rect 2952 8132 2956 8188
rect 2956 8132 3012 8188
rect 3012 8132 3016 8188
rect 2952 8128 3016 8132
rect 3032 8188 3096 8192
rect 3032 8132 3036 8188
rect 3036 8132 3092 8188
rect 3092 8132 3096 8188
rect 3032 8128 3096 8132
rect 3112 8188 3176 8192
rect 3112 8132 3116 8188
rect 3116 8132 3172 8188
rect 3172 8132 3176 8188
rect 3112 8128 3176 8132
rect 3192 8188 3256 8192
rect 3192 8132 3196 8188
rect 3196 8132 3252 8188
rect 3252 8132 3256 8188
rect 3192 8128 3256 8132
rect 12952 8188 13016 8192
rect 12952 8132 12956 8188
rect 12956 8132 13012 8188
rect 13012 8132 13016 8188
rect 12952 8128 13016 8132
rect 13032 8188 13096 8192
rect 13032 8132 13036 8188
rect 13036 8132 13092 8188
rect 13092 8132 13096 8188
rect 13032 8128 13096 8132
rect 13112 8188 13176 8192
rect 13112 8132 13116 8188
rect 13116 8132 13172 8188
rect 13172 8132 13176 8188
rect 13112 8128 13176 8132
rect 13192 8188 13256 8192
rect 13192 8132 13196 8188
rect 13196 8132 13252 8188
rect 13252 8132 13256 8188
rect 13192 8128 13256 8132
rect 22952 8188 23016 8192
rect 22952 8132 22956 8188
rect 22956 8132 23012 8188
rect 23012 8132 23016 8188
rect 22952 8128 23016 8132
rect 23032 8188 23096 8192
rect 23032 8132 23036 8188
rect 23036 8132 23092 8188
rect 23092 8132 23096 8188
rect 23032 8128 23096 8132
rect 23112 8188 23176 8192
rect 23112 8132 23116 8188
rect 23116 8132 23172 8188
rect 23172 8132 23176 8188
rect 23112 8128 23176 8132
rect 23192 8188 23256 8192
rect 23192 8132 23196 8188
rect 23196 8132 23252 8188
rect 23252 8132 23256 8188
rect 23192 8128 23256 8132
rect 15332 7924 15396 7988
rect 7952 7644 8016 7648
rect 7952 7588 7956 7644
rect 7956 7588 8012 7644
rect 8012 7588 8016 7644
rect 7952 7584 8016 7588
rect 8032 7644 8096 7648
rect 8032 7588 8036 7644
rect 8036 7588 8092 7644
rect 8092 7588 8096 7644
rect 8032 7584 8096 7588
rect 8112 7644 8176 7648
rect 8112 7588 8116 7644
rect 8116 7588 8172 7644
rect 8172 7588 8176 7644
rect 8112 7584 8176 7588
rect 8192 7644 8256 7648
rect 8192 7588 8196 7644
rect 8196 7588 8252 7644
rect 8252 7588 8256 7644
rect 8192 7584 8256 7588
rect 17952 7644 18016 7648
rect 17952 7588 17956 7644
rect 17956 7588 18012 7644
rect 18012 7588 18016 7644
rect 17952 7584 18016 7588
rect 18032 7644 18096 7648
rect 18032 7588 18036 7644
rect 18036 7588 18092 7644
rect 18092 7588 18096 7644
rect 18032 7584 18096 7588
rect 18112 7644 18176 7648
rect 18112 7588 18116 7644
rect 18116 7588 18172 7644
rect 18172 7588 18176 7644
rect 18112 7584 18176 7588
rect 18192 7644 18256 7648
rect 18192 7588 18196 7644
rect 18196 7588 18252 7644
rect 18252 7588 18256 7644
rect 18192 7584 18256 7588
rect 15332 7516 15396 7580
rect 2952 7100 3016 7104
rect 2952 7044 2956 7100
rect 2956 7044 3012 7100
rect 3012 7044 3016 7100
rect 2952 7040 3016 7044
rect 3032 7100 3096 7104
rect 3032 7044 3036 7100
rect 3036 7044 3092 7100
rect 3092 7044 3096 7100
rect 3032 7040 3096 7044
rect 3112 7100 3176 7104
rect 3112 7044 3116 7100
rect 3116 7044 3172 7100
rect 3172 7044 3176 7100
rect 3112 7040 3176 7044
rect 3192 7100 3256 7104
rect 3192 7044 3196 7100
rect 3196 7044 3252 7100
rect 3252 7044 3256 7100
rect 3192 7040 3256 7044
rect 12952 7100 13016 7104
rect 12952 7044 12956 7100
rect 12956 7044 13012 7100
rect 13012 7044 13016 7100
rect 12952 7040 13016 7044
rect 13032 7100 13096 7104
rect 13032 7044 13036 7100
rect 13036 7044 13092 7100
rect 13092 7044 13096 7100
rect 13032 7040 13096 7044
rect 13112 7100 13176 7104
rect 13112 7044 13116 7100
rect 13116 7044 13172 7100
rect 13172 7044 13176 7100
rect 13112 7040 13176 7044
rect 13192 7100 13256 7104
rect 13192 7044 13196 7100
rect 13196 7044 13252 7100
rect 13252 7044 13256 7100
rect 13192 7040 13256 7044
rect 22952 7100 23016 7104
rect 22952 7044 22956 7100
rect 22956 7044 23012 7100
rect 23012 7044 23016 7100
rect 22952 7040 23016 7044
rect 23032 7100 23096 7104
rect 23032 7044 23036 7100
rect 23036 7044 23092 7100
rect 23092 7044 23096 7100
rect 23032 7040 23096 7044
rect 23112 7100 23176 7104
rect 23112 7044 23116 7100
rect 23116 7044 23172 7100
rect 23172 7044 23176 7100
rect 23112 7040 23176 7044
rect 23192 7100 23256 7104
rect 23192 7044 23196 7100
rect 23196 7044 23252 7100
rect 23252 7044 23256 7100
rect 23192 7040 23256 7044
rect 23428 7032 23492 7036
rect 23428 6976 23442 7032
rect 23442 6976 23492 7032
rect 23428 6972 23492 6976
rect 7952 6556 8016 6560
rect 7952 6500 7956 6556
rect 7956 6500 8012 6556
rect 8012 6500 8016 6556
rect 7952 6496 8016 6500
rect 8032 6556 8096 6560
rect 8032 6500 8036 6556
rect 8036 6500 8092 6556
rect 8092 6500 8096 6556
rect 8032 6496 8096 6500
rect 8112 6556 8176 6560
rect 8112 6500 8116 6556
rect 8116 6500 8172 6556
rect 8172 6500 8176 6556
rect 8112 6496 8176 6500
rect 8192 6556 8256 6560
rect 8192 6500 8196 6556
rect 8196 6500 8252 6556
rect 8252 6500 8256 6556
rect 8192 6496 8256 6500
rect 17952 6556 18016 6560
rect 17952 6500 17956 6556
rect 17956 6500 18012 6556
rect 18012 6500 18016 6556
rect 17952 6496 18016 6500
rect 18032 6556 18096 6560
rect 18032 6500 18036 6556
rect 18036 6500 18092 6556
rect 18092 6500 18096 6556
rect 18032 6496 18096 6500
rect 18112 6556 18176 6560
rect 18112 6500 18116 6556
rect 18116 6500 18172 6556
rect 18172 6500 18176 6556
rect 18112 6496 18176 6500
rect 18192 6556 18256 6560
rect 18192 6500 18196 6556
rect 18196 6500 18252 6556
rect 18252 6500 18256 6556
rect 18192 6496 18256 6500
rect 2952 6012 3016 6016
rect 2952 5956 2956 6012
rect 2956 5956 3012 6012
rect 3012 5956 3016 6012
rect 2952 5952 3016 5956
rect 3032 6012 3096 6016
rect 3032 5956 3036 6012
rect 3036 5956 3092 6012
rect 3092 5956 3096 6012
rect 3032 5952 3096 5956
rect 3112 6012 3176 6016
rect 3112 5956 3116 6012
rect 3116 5956 3172 6012
rect 3172 5956 3176 6012
rect 3112 5952 3176 5956
rect 3192 6012 3256 6016
rect 3192 5956 3196 6012
rect 3196 5956 3252 6012
rect 3252 5956 3256 6012
rect 3192 5952 3256 5956
rect 12952 6012 13016 6016
rect 12952 5956 12956 6012
rect 12956 5956 13012 6012
rect 13012 5956 13016 6012
rect 12952 5952 13016 5956
rect 13032 6012 13096 6016
rect 13032 5956 13036 6012
rect 13036 5956 13092 6012
rect 13092 5956 13096 6012
rect 13032 5952 13096 5956
rect 13112 6012 13176 6016
rect 13112 5956 13116 6012
rect 13116 5956 13172 6012
rect 13172 5956 13176 6012
rect 13112 5952 13176 5956
rect 13192 6012 13256 6016
rect 13192 5956 13196 6012
rect 13196 5956 13252 6012
rect 13252 5956 13256 6012
rect 13192 5952 13256 5956
rect 22952 6012 23016 6016
rect 22952 5956 22956 6012
rect 22956 5956 23012 6012
rect 23012 5956 23016 6012
rect 22952 5952 23016 5956
rect 23032 6012 23096 6016
rect 23032 5956 23036 6012
rect 23036 5956 23092 6012
rect 23092 5956 23096 6012
rect 23032 5952 23096 5956
rect 23112 6012 23176 6016
rect 23112 5956 23116 6012
rect 23116 5956 23172 6012
rect 23172 5956 23176 6012
rect 23112 5952 23176 5956
rect 23192 6012 23256 6016
rect 23192 5956 23196 6012
rect 23196 5956 23252 6012
rect 23252 5956 23256 6012
rect 23192 5952 23256 5956
rect 21404 5536 21468 5540
rect 21404 5480 21418 5536
rect 21418 5480 21468 5536
rect 21404 5476 21468 5480
rect 23428 5536 23492 5540
rect 23428 5480 23442 5536
rect 23442 5480 23492 5536
rect 23428 5476 23492 5480
rect 7952 5468 8016 5472
rect 7952 5412 7956 5468
rect 7956 5412 8012 5468
rect 8012 5412 8016 5468
rect 7952 5408 8016 5412
rect 8032 5468 8096 5472
rect 8032 5412 8036 5468
rect 8036 5412 8092 5468
rect 8092 5412 8096 5468
rect 8032 5408 8096 5412
rect 8112 5468 8176 5472
rect 8112 5412 8116 5468
rect 8116 5412 8172 5468
rect 8172 5412 8176 5468
rect 8112 5408 8176 5412
rect 8192 5468 8256 5472
rect 8192 5412 8196 5468
rect 8196 5412 8252 5468
rect 8252 5412 8256 5468
rect 8192 5408 8256 5412
rect 17952 5468 18016 5472
rect 17952 5412 17956 5468
rect 17956 5412 18012 5468
rect 18012 5412 18016 5468
rect 17952 5408 18016 5412
rect 18032 5468 18096 5472
rect 18032 5412 18036 5468
rect 18036 5412 18092 5468
rect 18092 5412 18096 5468
rect 18032 5408 18096 5412
rect 18112 5468 18176 5472
rect 18112 5412 18116 5468
rect 18116 5412 18172 5468
rect 18172 5412 18176 5468
rect 18112 5408 18176 5412
rect 18192 5468 18256 5472
rect 18192 5412 18196 5468
rect 18196 5412 18252 5468
rect 18252 5412 18256 5468
rect 18192 5408 18256 5412
rect 2952 4924 3016 4928
rect 2952 4868 2956 4924
rect 2956 4868 3012 4924
rect 3012 4868 3016 4924
rect 2952 4864 3016 4868
rect 3032 4924 3096 4928
rect 3032 4868 3036 4924
rect 3036 4868 3092 4924
rect 3092 4868 3096 4924
rect 3032 4864 3096 4868
rect 3112 4924 3176 4928
rect 3112 4868 3116 4924
rect 3116 4868 3172 4924
rect 3172 4868 3176 4924
rect 3112 4864 3176 4868
rect 3192 4924 3256 4928
rect 3192 4868 3196 4924
rect 3196 4868 3252 4924
rect 3252 4868 3256 4924
rect 3192 4864 3256 4868
rect 12952 4924 13016 4928
rect 12952 4868 12956 4924
rect 12956 4868 13012 4924
rect 13012 4868 13016 4924
rect 12952 4864 13016 4868
rect 13032 4924 13096 4928
rect 13032 4868 13036 4924
rect 13036 4868 13092 4924
rect 13092 4868 13096 4924
rect 13032 4864 13096 4868
rect 13112 4924 13176 4928
rect 13112 4868 13116 4924
rect 13116 4868 13172 4924
rect 13172 4868 13176 4924
rect 13112 4864 13176 4868
rect 13192 4924 13256 4928
rect 13192 4868 13196 4924
rect 13196 4868 13252 4924
rect 13252 4868 13256 4924
rect 13192 4864 13256 4868
rect 22952 4924 23016 4928
rect 22952 4868 22956 4924
rect 22956 4868 23012 4924
rect 23012 4868 23016 4924
rect 22952 4864 23016 4868
rect 23032 4924 23096 4928
rect 23032 4868 23036 4924
rect 23036 4868 23092 4924
rect 23092 4868 23096 4924
rect 23032 4864 23096 4868
rect 23112 4924 23176 4928
rect 23112 4868 23116 4924
rect 23116 4868 23172 4924
rect 23172 4868 23176 4924
rect 23112 4864 23176 4868
rect 23192 4924 23256 4928
rect 23192 4868 23196 4924
rect 23196 4868 23252 4924
rect 23252 4868 23256 4924
rect 23192 4864 23256 4868
rect 7952 4380 8016 4384
rect 7952 4324 7956 4380
rect 7956 4324 8012 4380
rect 8012 4324 8016 4380
rect 7952 4320 8016 4324
rect 8032 4380 8096 4384
rect 8032 4324 8036 4380
rect 8036 4324 8092 4380
rect 8092 4324 8096 4380
rect 8032 4320 8096 4324
rect 8112 4380 8176 4384
rect 8112 4324 8116 4380
rect 8116 4324 8172 4380
rect 8172 4324 8176 4380
rect 8112 4320 8176 4324
rect 8192 4380 8256 4384
rect 8192 4324 8196 4380
rect 8196 4324 8252 4380
rect 8252 4324 8256 4380
rect 8192 4320 8256 4324
rect 17952 4380 18016 4384
rect 17952 4324 17956 4380
rect 17956 4324 18012 4380
rect 18012 4324 18016 4380
rect 17952 4320 18016 4324
rect 18032 4380 18096 4384
rect 18032 4324 18036 4380
rect 18036 4324 18092 4380
rect 18092 4324 18096 4380
rect 18032 4320 18096 4324
rect 18112 4380 18176 4384
rect 18112 4324 18116 4380
rect 18116 4324 18172 4380
rect 18172 4324 18176 4380
rect 18112 4320 18176 4324
rect 18192 4380 18256 4384
rect 18192 4324 18196 4380
rect 18196 4324 18252 4380
rect 18252 4324 18256 4380
rect 18192 4320 18256 4324
rect 20116 3980 20180 4044
rect 22140 4040 22204 4044
rect 22140 3984 22154 4040
rect 22154 3984 22204 4040
rect 22140 3980 22204 3984
rect 2952 3836 3016 3840
rect 2952 3780 2956 3836
rect 2956 3780 3012 3836
rect 3012 3780 3016 3836
rect 2952 3776 3016 3780
rect 3032 3836 3096 3840
rect 3032 3780 3036 3836
rect 3036 3780 3092 3836
rect 3092 3780 3096 3836
rect 3032 3776 3096 3780
rect 3112 3836 3176 3840
rect 3112 3780 3116 3836
rect 3116 3780 3172 3836
rect 3172 3780 3176 3836
rect 3112 3776 3176 3780
rect 3192 3836 3256 3840
rect 3192 3780 3196 3836
rect 3196 3780 3252 3836
rect 3252 3780 3256 3836
rect 3192 3776 3256 3780
rect 12952 3836 13016 3840
rect 12952 3780 12956 3836
rect 12956 3780 13012 3836
rect 13012 3780 13016 3836
rect 12952 3776 13016 3780
rect 13032 3836 13096 3840
rect 13032 3780 13036 3836
rect 13036 3780 13092 3836
rect 13092 3780 13096 3836
rect 13032 3776 13096 3780
rect 13112 3836 13176 3840
rect 13112 3780 13116 3836
rect 13116 3780 13172 3836
rect 13172 3780 13176 3836
rect 13112 3776 13176 3780
rect 13192 3836 13256 3840
rect 13192 3780 13196 3836
rect 13196 3780 13252 3836
rect 13252 3780 13256 3836
rect 13192 3776 13256 3780
rect 22952 3836 23016 3840
rect 22952 3780 22956 3836
rect 22956 3780 23012 3836
rect 23012 3780 23016 3836
rect 22952 3776 23016 3780
rect 23032 3836 23096 3840
rect 23032 3780 23036 3836
rect 23036 3780 23092 3836
rect 23092 3780 23096 3836
rect 23032 3776 23096 3780
rect 23112 3836 23176 3840
rect 23112 3780 23116 3836
rect 23116 3780 23172 3836
rect 23172 3780 23176 3836
rect 23112 3776 23176 3780
rect 23192 3836 23256 3840
rect 23192 3780 23196 3836
rect 23196 3780 23252 3836
rect 23252 3780 23256 3836
rect 23192 3776 23256 3780
rect 17356 3572 17420 3636
rect 19564 3572 19628 3636
rect 19380 3436 19444 3500
rect 7952 3292 8016 3296
rect 7952 3236 7956 3292
rect 7956 3236 8012 3292
rect 8012 3236 8016 3292
rect 7952 3232 8016 3236
rect 8032 3292 8096 3296
rect 8032 3236 8036 3292
rect 8036 3236 8092 3292
rect 8092 3236 8096 3292
rect 8032 3232 8096 3236
rect 8112 3292 8176 3296
rect 8112 3236 8116 3292
rect 8116 3236 8172 3292
rect 8172 3236 8176 3292
rect 8112 3232 8176 3236
rect 8192 3292 8256 3296
rect 8192 3236 8196 3292
rect 8196 3236 8252 3292
rect 8252 3236 8256 3292
rect 8192 3232 8256 3236
rect 17952 3292 18016 3296
rect 17952 3236 17956 3292
rect 17956 3236 18012 3292
rect 18012 3236 18016 3292
rect 17952 3232 18016 3236
rect 18032 3292 18096 3296
rect 18032 3236 18036 3292
rect 18036 3236 18092 3292
rect 18092 3236 18096 3292
rect 18032 3232 18096 3236
rect 18112 3292 18176 3296
rect 18112 3236 18116 3292
rect 18116 3236 18172 3292
rect 18172 3236 18176 3292
rect 18112 3232 18176 3236
rect 18192 3292 18256 3296
rect 18192 3236 18196 3292
rect 18196 3236 18252 3292
rect 18252 3236 18256 3292
rect 18192 3232 18256 3236
rect 13492 3028 13556 3092
rect 2952 2748 3016 2752
rect 2952 2692 2956 2748
rect 2956 2692 3012 2748
rect 3012 2692 3016 2748
rect 2952 2688 3016 2692
rect 3032 2748 3096 2752
rect 3032 2692 3036 2748
rect 3036 2692 3092 2748
rect 3092 2692 3096 2748
rect 3032 2688 3096 2692
rect 3112 2748 3176 2752
rect 3112 2692 3116 2748
rect 3116 2692 3172 2748
rect 3172 2692 3176 2748
rect 3112 2688 3176 2692
rect 3192 2748 3256 2752
rect 3192 2692 3196 2748
rect 3196 2692 3252 2748
rect 3252 2692 3256 2748
rect 3192 2688 3256 2692
rect 12952 2748 13016 2752
rect 12952 2692 12956 2748
rect 12956 2692 13012 2748
rect 13012 2692 13016 2748
rect 12952 2688 13016 2692
rect 13032 2748 13096 2752
rect 13032 2692 13036 2748
rect 13036 2692 13092 2748
rect 13092 2692 13096 2748
rect 13032 2688 13096 2692
rect 13112 2748 13176 2752
rect 13112 2692 13116 2748
rect 13116 2692 13172 2748
rect 13172 2692 13176 2748
rect 13112 2688 13176 2692
rect 13192 2748 13256 2752
rect 13192 2692 13196 2748
rect 13196 2692 13252 2748
rect 13252 2692 13256 2748
rect 13192 2688 13256 2692
rect 22952 2748 23016 2752
rect 22952 2692 22956 2748
rect 22956 2692 23012 2748
rect 23012 2692 23016 2748
rect 22952 2688 23016 2692
rect 23032 2748 23096 2752
rect 23032 2692 23036 2748
rect 23036 2692 23092 2748
rect 23092 2692 23096 2748
rect 23032 2688 23096 2692
rect 23112 2748 23176 2752
rect 23112 2692 23116 2748
rect 23116 2692 23172 2748
rect 23172 2692 23176 2748
rect 23112 2688 23176 2692
rect 23192 2748 23256 2752
rect 23192 2692 23196 2748
rect 23196 2692 23252 2748
rect 23252 2692 23256 2748
rect 23192 2688 23256 2692
rect 14964 2484 15028 2548
rect 21036 2484 21100 2548
rect 16068 2348 16132 2412
rect 7952 2204 8016 2208
rect 7952 2148 7956 2204
rect 7956 2148 8012 2204
rect 8012 2148 8016 2204
rect 7952 2144 8016 2148
rect 8032 2204 8096 2208
rect 8032 2148 8036 2204
rect 8036 2148 8092 2204
rect 8092 2148 8096 2204
rect 8032 2144 8096 2148
rect 8112 2204 8176 2208
rect 8112 2148 8116 2204
rect 8116 2148 8172 2204
rect 8172 2148 8176 2204
rect 8112 2144 8176 2148
rect 8192 2204 8256 2208
rect 8192 2148 8196 2204
rect 8196 2148 8252 2204
rect 8252 2148 8256 2204
rect 8192 2144 8256 2148
rect 17952 2204 18016 2208
rect 17952 2148 17956 2204
rect 17956 2148 18012 2204
rect 18012 2148 18016 2204
rect 17952 2144 18016 2148
rect 18032 2204 18096 2208
rect 18032 2148 18036 2204
rect 18036 2148 18092 2204
rect 18092 2148 18096 2204
rect 18032 2144 18096 2148
rect 18112 2204 18176 2208
rect 18112 2148 18116 2204
rect 18116 2148 18172 2204
rect 18172 2148 18176 2204
rect 18112 2144 18176 2148
rect 18192 2204 18256 2208
rect 18192 2148 18196 2204
rect 18196 2148 18252 2204
rect 18252 2148 18256 2204
rect 18192 2144 18256 2148
<< metal4 >>
rect 2944 53888 3264 54448
rect 2944 53824 2952 53888
rect 3016 53824 3032 53888
rect 3096 53824 3112 53888
rect 3176 53824 3192 53888
rect 3256 53824 3264 53888
rect 2944 52800 3264 53824
rect 2944 52736 2952 52800
rect 3016 52736 3032 52800
rect 3096 52736 3112 52800
rect 3176 52736 3192 52800
rect 3256 52736 3264 52800
rect 2944 51712 3264 52736
rect 2944 51648 2952 51712
rect 3016 51648 3032 51712
rect 3096 51648 3112 51712
rect 3176 51648 3192 51712
rect 3256 51648 3264 51712
rect 2944 50624 3264 51648
rect 2944 50560 2952 50624
rect 3016 50560 3032 50624
rect 3096 50560 3112 50624
rect 3176 50560 3192 50624
rect 3256 50560 3264 50624
rect 2944 49536 3264 50560
rect 2944 49472 2952 49536
rect 3016 49472 3032 49536
rect 3096 49472 3112 49536
rect 3176 49472 3192 49536
rect 3256 49472 3264 49536
rect 2944 48448 3264 49472
rect 2944 48384 2952 48448
rect 3016 48384 3032 48448
rect 3096 48384 3112 48448
rect 3176 48384 3192 48448
rect 3256 48384 3264 48448
rect 2944 47360 3264 48384
rect 2944 47296 2952 47360
rect 3016 47296 3032 47360
rect 3096 47296 3112 47360
rect 3176 47296 3192 47360
rect 3256 47296 3264 47360
rect 2944 46272 3264 47296
rect 2944 46208 2952 46272
rect 3016 46208 3032 46272
rect 3096 46208 3112 46272
rect 3176 46208 3192 46272
rect 3256 46208 3264 46272
rect 2944 45184 3264 46208
rect 2944 45120 2952 45184
rect 3016 45120 3032 45184
rect 3096 45120 3112 45184
rect 3176 45120 3192 45184
rect 3256 45120 3264 45184
rect 2944 44096 3264 45120
rect 2944 44032 2952 44096
rect 3016 44032 3032 44096
rect 3096 44032 3112 44096
rect 3176 44032 3192 44096
rect 3256 44032 3264 44096
rect 2944 43008 3264 44032
rect 2944 42944 2952 43008
rect 3016 42944 3032 43008
rect 3096 42944 3112 43008
rect 3176 42944 3192 43008
rect 3256 42944 3264 43008
rect 2944 41920 3264 42944
rect 2944 41856 2952 41920
rect 3016 41856 3032 41920
rect 3096 41856 3112 41920
rect 3176 41856 3192 41920
rect 3256 41856 3264 41920
rect 2944 40832 3264 41856
rect 2944 40768 2952 40832
rect 3016 40768 3032 40832
rect 3096 40768 3112 40832
rect 3176 40768 3192 40832
rect 3256 40768 3264 40832
rect 2944 39744 3264 40768
rect 2944 39680 2952 39744
rect 3016 39680 3032 39744
rect 3096 39680 3112 39744
rect 3176 39680 3192 39744
rect 3256 39680 3264 39744
rect 2944 38656 3264 39680
rect 2944 38592 2952 38656
rect 3016 38592 3032 38656
rect 3096 38592 3112 38656
rect 3176 38592 3192 38656
rect 3256 38592 3264 38656
rect 2944 37568 3264 38592
rect 2944 37504 2952 37568
rect 3016 37504 3032 37568
rect 3096 37504 3112 37568
rect 3176 37504 3192 37568
rect 3256 37504 3264 37568
rect 2944 36480 3264 37504
rect 2944 36416 2952 36480
rect 3016 36416 3032 36480
rect 3096 36416 3112 36480
rect 3176 36416 3192 36480
rect 3256 36416 3264 36480
rect 2944 35392 3264 36416
rect 2944 35328 2952 35392
rect 3016 35328 3032 35392
rect 3096 35328 3112 35392
rect 3176 35328 3192 35392
rect 3256 35328 3264 35392
rect 2944 34304 3264 35328
rect 2944 34240 2952 34304
rect 3016 34240 3032 34304
rect 3096 34240 3112 34304
rect 3176 34240 3192 34304
rect 3256 34240 3264 34304
rect 2944 33216 3264 34240
rect 2944 33152 2952 33216
rect 3016 33152 3032 33216
rect 3096 33152 3112 33216
rect 3176 33152 3192 33216
rect 3256 33152 3264 33216
rect 2944 32128 3264 33152
rect 2944 32064 2952 32128
rect 3016 32064 3032 32128
rect 3096 32064 3112 32128
rect 3176 32064 3192 32128
rect 3256 32064 3264 32128
rect 2944 31040 3264 32064
rect 2944 30976 2952 31040
rect 3016 30976 3032 31040
rect 3096 30976 3112 31040
rect 3176 30976 3192 31040
rect 3256 30976 3264 31040
rect 2944 29952 3264 30976
rect 2944 29888 2952 29952
rect 3016 29888 3032 29952
rect 3096 29888 3112 29952
rect 3176 29888 3192 29952
rect 3256 29888 3264 29952
rect 2944 28864 3264 29888
rect 2944 28800 2952 28864
rect 3016 28800 3032 28864
rect 3096 28800 3112 28864
rect 3176 28800 3192 28864
rect 3256 28800 3264 28864
rect 2944 27776 3264 28800
rect 2944 27712 2952 27776
rect 3016 27712 3032 27776
rect 3096 27712 3112 27776
rect 3176 27712 3192 27776
rect 3256 27712 3264 27776
rect 2944 26688 3264 27712
rect 2944 26624 2952 26688
rect 3016 26624 3032 26688
rect 3096 26624 3112 26688
rect 3176 26624 3192 26688
rect 3256 26624 3264 26688
rect 2944 25600 3264 26624
rect 2944 25536 2952 25600
rect 3016 25536 3032 25600
rect 3096 25536 3112 25600
rect 3176 25536 3192 25600
rect 3256 25536 3264 25600
rect 2944 24512 3264 25536
rect 2944 24448 2952 24512
rect 3016 24448 3032 24512
rect 3096 24448 3112 24512
rect 3176 24448 3192 24512
rect 3256 24448 3264 24512
rect 2944 23424 3264 24448
rect 2944 23360 2952 23424
rect 3016 23360 3032 23424
rect 3096 23360 3112 23424
rect 3176 23360 3192 23424
rect 3256 23360 3264 23424
rect 2944 22336 3264 23360
rect 2944 22272 2952 22336
rect 3016 22272 3032 22336
rect 3096 22272 3112 22336
rect 3176 22272 3192 22336
rect 3256 22272 3264 22336
rect 2944 21248 3264 22272
rect 2944 21184 2952 21248
rect 3016 21184 3032 21248
rect 3096 21184 3112 21248
rect 3176 21184 3192 21248
rect 3256 21184 3264 21248
rect 2944 20160 3264 21184
rect 2944 20096 2952 20160
rect 3016 20096 3032 20160
rect 3096 20096 3112 20160
rect 3176 20096 3192 20160
rect 3256 20096 3264 20160
rect 2944 19072 3264 20096
rect 2944 19008 2952 19072
rect 3016 19008 3032 19072
rect 3096 19008 3112 19072
rect 3176 19008 3192 19072
rect 3256 19008 3264 19072
rect 2944 17984 3264 19008
rect 2944 17920 2952 17984
rect 3016 17920 3032 17984
rect 3096 17920 3112 17984
rect 3176 17920 3192 17984
rect 3256 17920 3264 17984
rect 2944 16896 3264 17920
rect 2944 16832 2952 16896
rect 3016 16832 3032 16896
rect 3096 16832 3112 16896
rect 3176 16832 3192 16896
rect 3256 16832 3264 16896
rect 2944 15808 3264 16832
rect 2944 15744 2952 15808
rect 3016 15744 3032 15808
rect 3096 15744 3112 15808
rect 3176 15744 3192 15808
rect 3256 15744 3264 15808
rect 2944 14720 3264 15744
rect 2944 14656 2952 14720
rect 3016 14656 3032 14720
rect 3096 14656 3112 14720
rect 3176 14656 3192 14720
rect 3256 14656 3264 14720
rect 2944 13632 3264 14656
rect 2944 13568 2952 13632
rect 3016 13568 3032 13632
rect 3096 13568 3112 13632
rect 3176 13568 3192 13632
rect 3256 13568 3264 13632
rect 2944 12544 3264 13568
rect 2944 12480 2952 12544
rect 3016 12480 3032 12544
rect 3096 12480 3112 12544
rect 3176 12480 3192 12544
rect 3256 12480 3264 12544
rect 2944 11456 3264 12480
rect 2944 11392 2952 11456
rect 3016 11392 3032 11456
rect 3096 11392 3112 11456
rect 3176 11392 3192 11456
rect 3256 11392 3264 11456
rect 2944 10368 3264 11392
rect 2944 10304 2952 10368
rect 3016 10304 3032 10368
rect 3096 10304 3112 10368
rect 3176 10304 3192 10368
rect 3256 10304 3264 10368
rect 2944 9280 3264 10304
rect 2944 9216 2952 9280
rect 3016 9216 3032 9280
rect 3096 9216 3112 9280
rect 3176 9216 3192 9280
rect 3256 9216 3264 9280
rect 2944 8192 3264 9216
rect 2944 8128 2952 8192
rect 3016 8128 3032 8192
rect 3096 8128 3112 8192
rect 3176 8128 3192 8192
rect 3256 8128 3264 8192
rect 2944 7104 3264 8128
rect 2944 7040 2952 7104
rect 3016 7040 3032 7104
rect 3096 7040 3112 7104
rect 3176 7040 3192 7104
rect 3256 7040 3264 7104
rect 2944 6016 3264 7040
rect 2944 5952 2952 6016
rect 3016 5952 3032 6016
rect 3096 5952 3112 6016
rect 3176 5952 3192 6016
rect 3256 5952 3264 6016
rect 2944 4928 3264 5952
rect 2944 4864 2952 4928
rect 3016 4864 3032 4928
rect 3096 4864 3112 4928
rect 3176 4864 3192 4928
rect 3256 4864 3264 4928
rect 2944 3840 3264 4864
rect 2944 3776 2952 3840
rect 3016 3776 3032 3840
rect 3096 3776 3112 3840
rect 3176 3776 3192 3840
rect 3256 3776 3264 3840
rect 2944 2752 3264 3776
rect 2944 2688 2952 2752
rect 3016 2688 3032 2752
rect 3096 2688 3112 2752
rect 3176 2688 3192 2752
rect 3256 2688 3264 2752
rect 2944 2128 3264 2688
rect 7944 54432 8264 54448
rect 7944 54368 7952 54432
rect 8016 54368 8032 54432
rect 8096 54368 8112 54432
rect 8176 54368 8192 54432
rect 8256 54368 8264 54432
rect 7944 53344 8264 54368
rect 7944 53280 7952 53344
rect 8016 53280 8032 53344
rect 8096 53280 8112 53344
rect 8176 53280 8192 53344
rect 8256 53280 8264 53344
rect 7944 52256 8264 53280
rect 7944 52192 7952 52256
rect 8016 52192 8032 52256
rect 8096 52192 8112 52256
rect 8176 52192 8192 52256
rect 8256 52192 8264 52256
rect 7944 51168 8264 52192
rect 7944 51104 7952 51168
rect 8016 51104 8032 51168
rect 8096 51104 8112 51168
rect 8176 51104 8192 51168
rect 8256 51104 8264 51168
rect 7944 50080 8264 51104
rect 7944 50016 7952 50080
rect 8016 50016 8032 50080
rect 8096 50016 8112 50080
rect 8176 50016 8192 50080
rect 8256 50016 8264 50080
rect 7944 48992 8264 50016
rect 7944 48928 7952 48992
rect 8016 48928 8032 48992
rect 8096 48928 8112 48992
rect 8176 48928 8192 48992
rect 8256 48928 8264 48992
rect 7944 47904 8264 48928
rect 7944 47840 7952 47904
rect 8016 47840 8032 47904
rect 8096 47840 8112 47904
rect 8176 47840 8192 47904
rect 8256 47840 8264 47904
rect 7944 46816 8264 47840
rect 7944 46752 7952 46816
rect 8016 46752 8032 46816
rect 8096 46752 8112 46816
rect 8176 46752 8192 46816
rect 8256 46752 8264 46816
rect 7944 45728 8264 46752
rect 7944 45664 7952 45728
rect 8016 45664 8032 45728
rect 8096 45664 8112 45728
rect 8176 45664 8192 45728
rect 8256 45664 8264 45728
rect 7944 44640 8264 45664
rect 7944 44576 7952 44640
rect 8016 44576 8032 44640
rect 8096 44576 8112 44640
rect 8176 44576 8192 44640
rect 8256 44576 8264 44640
rect 7944 43552 8264 44576
rect 7944 43488 7952 43552
rect 8016 43488 8032 43552
rect 8096 43488 8112 43552
rect 8176 43488 8192 43552
rect 8256 43488 8264 43552
rect 7944 42464 8264 43488
rect 7944 42400 7952 42464
rect 8016 42400 8032 42464
rect 8096 42400 8112 42464
rect 8176 42400 8192 42464
rect 8256 42400 8264 42464
rect 7944 41376 8264 42400
rect 7944 41312 7952 41376
rect 8016 41312 8032 41376
rect 8096 41312 8112 41376
rect 8176 41312 8192 41376
rect 8256 41312 8264 41376
rect 7944 40288 8264 41312
rect 7944 40224 7952 40288
rect 8016 40224 8032 40288
rect 8096 40224 8112 40288
rect 8176 40224 8192 40288
rect 8256 40224 8264 40288
rect 7944 39200 8264 40224
rect 7944 39136 7952 39200
rect 8016 39136 8032 39200
rect 8096 39136 8112 39200
rect 8176 39136 8192 39200
rect 8256 39136 8264 39200
rect 7944 38112 8264 39136
rect 7944 38048 7952 38112
rect 8016 38048 8032 38112
rect 8096 38048 8112 38112
rect 8176 38048 8192 38112
rect 8256 38048 8264 38112
rect 7944 37024 8264 38048
rect 7944 36960 7952 37024
rect 8016 36960 8032 37024
rect 8096 36960 8112 37024
rect 8176 36960 8192 37024
rect 8256 36960 8264 37024
rect 7944 35936 8264 36960
rect 7944 35872 7952 35936
rect 8016 35872 8032 35936
rect 8096 35872 8112 35936
rect 8176 35872 8192 35936
rect 8256 35872 8264 35936
rect 7944 34848 8264 35872
rect 7944 34784 7952 34848
rect 8016 34784 8032 34848
rect 8096 34784 8112 34848
rect 8176 34784 8192 34848
rect 8256 34784 8264 34848
rect 7944 33760 8264 34784
rect 7944 33696 7952 33760
rect 8016 33696 8032 33760
rect 8096 33696 8112 33760
rect 8176 33696 8192 33760
rect 8256 33696 8264 33760
rect 7944 32672 8264 33696
rect 7944 32608 7952 32672
rect 8016 32608 8032 32672
rect 8096 32608 8112 32672
rect 8176 32608 8192 32672
rect 8256 32608 8264 32672
rect 7944 31584 8264 32608
rect 7944 31520 7952 31584
rect 8016 31520 8032 31584
rect 8096 31520 8112 31584
rect 8176 31520 8192 31584
rect 8256 31520 8264 31584
rect 7944 30496 8264 31520
rect 7944 30432 7952 30496
rect 8016 30432 8032 30496
rect 8096 30432 8112 30496
rect 8176 30432 8192 30496
rect 8256 30432 8264 30496
rect 7944 29408 8264 30432
rect 7944 29344 7952 29408
rect 8016 29344 8032 29408
rect 8096 29344 8112 29408
rect 8176 29344 8192 29408
rect 8256 29344 8264 29408
rect 7944 28320 8264 29344
rect 7944 28256 7952 28320
rect 8016 28256 8032 28320
rect 8096 28256 8112 28320
rect 8176 28256 8192 28320
rect 8256 28256 8264 28320
rect 7944 27232 8264 28256
rect 7944 27168 7952 27232
rect 8016 27168 8032 27232
rect 8096 27168 8112 27232
rect 8176 27168 8192 27232
rect 8256 27168 8264 27232
rect 7944 26144 8264 27168
rect 7944 26080 7952 26144
rect 8016 26080 8032 26144
rect 8096 26080 8112 26144
rect 8176 26080 8192 26144
rect 8256 26080 8264 26144
rect 7944 25056 8264 26080
rect 7944 24992 7952 25056
rect 8016 24992 8032 25056
rect 8096 24992 8112 25056
rect 8176 24992 8192 25056
rect 8256 24992 8264 25056
rect 7944 23968 8264 24992
rect 7944 23904 7952 23968
rect 8016 23904 8032 23968
rect 8096 23904 8112 23968
rect 8176 23904 8192 23968
rect 8256 23904 8264 23968
rect 7944 22880 8264 23904
rect 7944 22816 7952 22880
rect 8016 22816 8032 22880
rect 8096 22816 8112 22880
rect 8176 22816 8192 22880
rect 8256 22816 8264 22880
rect 7944 21792 8264 22816
rect 7944 21728 7952 21792
rect 8016 21728 8032 21792
rect 8096 21728 8112 21792
rect 8176 21728 8192 21792
rect 8256 21728 8264 21792
rect 7944 20704 8264 21728
rect 7944 20640 7952 20704
rect 8016 20640 8032 20704
rect 8096 20640 8112 20704
rect 8176 20640 8192 20704
rect 8256 20640 8264 20704
rect 7944 19616 8264 20640
rect 7944 19552 7952 19616
rect 8016 19552 8032 19616
rect 8096 19552 8112 19616
rect 8176 19552 8192 19616
rect 8256 19552 8264 19616
rect 7944 18528 8264 19552
rect 7944 18464 7952 18528
rect 8016 18464 8032 18528
rect 8096 18464 8112 18528
rect 8176 18464 8192 18528
rect 8256 18464 8264 18528
rect 7944 17440 8264 18464
rect 7944 17376 7952 17440
rect 8016 17376 8032 17440
rect 8096 17376 8112 17440
rect 8176 17376 8192 17440
rect 8256 17376 8264 17440
rect 7944 16352 8264 17376
rect 7944 16288 7952 16352
rect 8016 16288 8032 16352
rect 8096 16288 8112 16352
rect 8176 16288 8192 16352
rect 8256 16288 8264 16352
rect 7944 15264 8264 16288
rect 7944 15200 7952 15264
rect 8016 15200 8032 15264
rect 8096 15200 8112 15264
rect 8176 15200 8192 15264
rect 8256 15200 8264 15264
rect 7944 14176 8264 15200
rect 7944 14112 7952 14176
rect 8016 14112 8032 14176
rect 8096 14112 8112 14176
rect 8176 14112 8192 14176
rect 8256 14112 8264 14176
rect 7944 13088 8264 14112
rect 7944 13024 7952 13088
rect 8016 13024 8032 13088
rect 8096 13024 8112 13088
rect 8176 13024 8192 13088
rect 8256 13024 8264 13088
rect 7944 12000 8264 13024
rect 7944 11936 7952 12000
rect 8016 11936 8032 12000
rect 8096 11936 8112 12000
rect 8176 11936 8192 12000
rect 8256 11936 8264 12000
rect 7944 10912 8264 11936
rect 7944 10848 7952 10912
rect 8016 10848 8032 10912
rect 8096 10848 8112 10912
rect 8176 10848 8192 10912
rect 8256 10848 8264 10912
rect 7944 9824 8264 10848
rect 7944 9760 7952 9824
rect 8016 9760 8032 9824
rect 8096 9760 8112 9824
rect 8176 9760 8192 9824
rect 8256 9760 8264 9824
rect 7944 8736 8264 9760
rect 7944 8672 7952 8736
rect 8016 8672 8032 8736
rect 8096 8672 8112 8736
rect 8176 8672 8192 8736
rect 8256 8672 8264 8736
rect 7944 7648 8264 8672
rect 7944 7584 7952 7648
rect 8016 7584 8032 7648
rect 8096 7584 8112 7648
rect 8176 7584 8192 7648
rect 8256 7584 8264 7648
rect 7944 6560 8264 7584
rect 7944 6496 7952 6560
rect 8016 6496 8032 6560
rect 8096 6496 8112 6560
rect 8176 6496 8192 6560
rect 8256 6496 8264 6560
rect 7944 5472 8264 6496
rect 7944 5408 7952 5472
rect 8016 5408 8032 5472
rect 8096 5408 8112 5472
rect 8176 5408 8192 5472
rect 8256 5408 8264 5472
rect 7944 4384 8264 5408
rect 7944 4320 7952 4384
rect 8016 4320 8032 4384
rect 8096 4320 8112 4384
rect 8176 4320 8192 4384
rect 8256 4320 8264 4384
rect 7944 3296 8264 4320
rect 7944 3232 7952 3296
rect 8016 3232 8032 3296
rect 8096 3232 8112 3296
rect 8176 3232 8192 3296
rect 8256 3232 8264 3296
rect 7944 2208 8264 3232
rect 7944 2144 7952 2208
rect 8016 2144 8032 2208
rect 8096 2144 8112 2208
rect 8176 2144 8192 2208
rect 8256 2144 8264 2208
rect 7944 2128 8264 2144
rect 12944 53888 13264 54448
rect 12944 53824 12952 53888
rect 13016 53824 13032 53888
rect 13096 53824 13112 53888
rect 13176 53824 13192 53888
rect 13256 53824 13264 53888
rect 12944 52800 13264 53824
rect 12944 52736 12952 52800
rect 13016 52736 13032 52800
rect 13096 52736 13112 52800
rect 13176 52736 13192 52800
rect 13256 52736 13264 52800
rect 12944 51712 13264 52736
rect 12944 51648 12952 51712
rect 13016 51648 13032 51712
rect 13096 51648 13112 51712
rect 13176 51648 13192 51712
rect 13256 51648 13264 51712
rect 12944 50624 13264 51648
rect 12944 50560 12952 50624
rect 13016 50560 13032 50624
rect 13096 50560 13112 50624
rect 13176 50560 13192 50624
rect 13256 50560 13264 50624
rect 12944 49536 13264 50560
rect 12944 49472 12952 49536
rect 13016 49472 13032 49536
rect 13096 49472 13112 49536
rect 13176 49472 13192 49536
rect 13256 49472 13264 49536
rect 12944 48448 13264 49472
rect 12944 48384 12952 48448
rect 13016 48384 13032 48448
rect 13096 48384 13112 48448
rect 13176 48384 13192 48448
rect 13256 48384 13264 48448
rect 12944 47360 13264 48384
rect 12944 47296 12952 47360
rect 13016 47296 13032 47360
rect 13096 47296 13112 47360
rect 13176 47296 13192 47360
rect 13256 47296 13264 47360
rect 12944 46272 13264 47296
rect 12944 46208 12952 46272
rect 13016 46208 13032 46272
rect 13096 46208 13112 46272
rect 13176 46208 13192 46272
rect 13256 46208 13264 46272
rect 12944 45184 13264 46208
rect 12944 45120 12952 45184
rect 13016 45120 13032 45184
rect 13096 45120 13112 45184
rect 13176 45120 13192 45184
rect 13256 45120 13264 45184
rect 12944 44096 13264 45120
rect 12944 44032 12952 44096
rect 13016 44032 13032 44096
rect 13096 44032 13112 44096
rect 13176 44032 13192 44096
rect 13256 44032 13264 44096
rect 12944 43008 13264 44032
rect 12944 42944 12952 43008
rect 13016 42944 13032 43008
rect 13096 42944 13112 43008
rect 13176 42944 13192 43008
rect 13256 42944 13264 43008
rect 12944 41920 13264 42944
rect 12944 41856 12952 41920
rect 13016 41856 13032 41920
rect 13096 41856 13112 41920
rect 13176 41856 13192 41920
rect 13256 41856 13264 41920
rect 12944 40832 13264 41856
rect 12944 40768 12952 40832
rect 13016 40768 13032 40832
rect 13096 40768 13112 40832
rect 13176 40768 13192 40832
rect 13256 40768 13264 40832
rect 12944 39744 13264 40768
rect 12944 39680 12952 39744
rect 13016 39680 13032 39744
rect 13096 39680 13112 39744
rect 13176 39680 13192 39744
rect 13256 39680 13264 39744
rect 12944 38656 13264 39680
rect 12944 38592 12952 38656
rect 13016 38592 13032 38656
rect 13096 38592 13112 38656
rect 13176 38592 13192 38656
rect 13256 38592 13264 38656
rect 12944 37568 13264 38592
rect 12944 37504 12952 37568
rect 13016 37504 13032 37568
rect 13096 37504 13112 37568
rect 13176 37504 13192 37568
rect 13256 37504 13264 37568
rect 12944 36480 13264 37504
rect 12944 36416 12952 36480
rect 13016 36416 13032 36480
rect 13096 36416 13112 36480
rect 13176 36416 13192 36480
rect 13256 36416 13264 36480
rect 12944 35392 13264 36416
rect 12944 35328 12952 35392
rect 13016 35328 13032 35392
rect 13096 35328 13112 35392
rect 13176 35328 13192 35392
rect 13256 35328 13264 35392
rect 12944 34304 13264 35328
rect 12944 34240 12952 34304
rect 13016 34240 13032 34304
rect 13096 34240 13112 34304
rect 13176 34240 13192 34304
rect 13256 34240 13264 34304
rect 12944 33216 13264 34240
rect 12944 33152 12952 33216
rect 13016 33152 13032 33216
rect 13096 33152 13112 33216
rect 13176 33152 13192 33216
rect 13256 33152 13264 33216
rect 12944 32128 13264 33152
rect 12944 32064 12952 32128
rect 13016 32064 13032 32128
rect 13096 32064 13112 32128
rect 13176 32064 13192 32128
rect 13256 32064 13264 32128
rect 12944 31040 13264 32064
rect 12944 30976 12952 31040
rect 13016 30976 13032 31040
rect 13096 30976 13112 31040
rect 13176 30976 13192 31040
rect 13256 30976 13264 31040
rect 12944 29952 13264 30976
rect 12944 29888 12952 29952
rect 13016 29888 13032 29952
rect 13096 29888 13112 29952
rect 13176 29888 13192 29952
rect 13256 29888 13264 29952
rect 12944 28864 13264 29888
rect 12944 28800 12952 28864
rect 13016 28800 13032 28864
rect 13096 28800 13112 28864
rect 13176 28800 13192 28864
rect 13256 28800 13264 28864
rect 12944 27776 13264 28800
rect 12944 27712 12952 27776
rect 13016 27712 13032 27776
rect 13096 27712 13112 27776
rect 13176 27712 13192 27776
rect 13256 27712 13264 27776
rect 12944 26688 13264 27712
rect 17944 54432 18264 54448
rect 17944 54368 17952 54432
rect 18016 54368 18032 54432
rect 18096 54368 18112 54432
rect 18176 54368 18192 54432
rect 18256 54368 18264 54432
rect 17944 53344 18264 54368
rect 17944 53280 17952 53344
rect 18016 53280 18032 53344
rect 18096 53280 18112 53344
rect 18176 53280 18192 53344
rect 18256 53280 18264 53344
rect 17944 52256 18264 53280
rect 17944 52192 17952 52256
rect 18016 52192 18032 52256
rect 18096 52192 18112 52256
rect 18176 52192 18192 52256
rect 18256 52192 18264 52256
rect 17944 51168 18264 52192
rect 17944 51104 17952 51168
rect 18016 51104 18032 51168
rect 18096 51104 18112 51168
rect 18176 51104 18192 51168
rect 18256 51104 18264 51168
rect 17944 50080 18264 51104
rect 17944 50016 17952 50080
rect 18016 50016 18032 50080
rect 18096 50016 18112 50080
rect 18176 50016 18192 50080
rect 18256 50016 18264 50080
rect 17944 48992 18264 50016
rect 17944 48928 17952 48992
rect 18016 48928 18032 48992
rect 18096 48928 18112 48992
rect 18176 48928 18192 48992
rect 18256 48928 18264 48992
rect 17944 47904 18264 48928
rect 17944 47840 17952 47904
rect 18016 47840 18032 47904
rect 18096 47840 18112 47904
rect 18176 47840 18192 47904
rect 18256 47840 18264 47904
rect 17944 46816 18264 47840
rect 17944 46752 17952 46816
rect 18016 46752 18032 46816
rect 18096 46752 18112 46816
rect 18176 46752 18192 46816
rect 18256 46752 18264 46816
rect 17944 45728 18264 46752
rect 17944 45664 17952 45728
rect 18016 45664 18032 45728
rect 18096 45664 18112 45728
rect 18176 45664 18192 45728
rect 18256 45664 18264 45728
rect 17944 44640 18264 45664
rect 17944 44576 17952 44640
rect 18016 44576 18032 44640
rect 18096 44576 18112 44640
rect 18176 44576 18192 44640
rect 18256 44576 18264 44640
rect 17944 43552 18264 44576
rect 17944 43488 17952 43552
rect 18016 43488 18032 43552
rect 18096 43488 18112 43552
rect 18176 43488 18192 43552
rect 18256 43488 18264 43552
rect 17944 42464 18264 43488
rect 17944 42400 17952 42464
rect 18016 42400 18032 42464
rect 18096 42400 18112 42464
rect 18176 42400 18192 42464
rect 18256 42400 18264 42464
rect 17944 41376 18264 42400
rect 17944 41312 17952 41376
rect 18016 41312 18032 41376
rect 18096 41312 18112 41376
rect 18176 41312 18192 41376
rect 18256 41312 18264 41376
rect 17944 40288 18264 41312
rect 17944 40224 17952 40288
rect 18016 40224 18032 40288
rect 18096 40224 18112 40288
rect 18176 40224 18192 40288
rect 18256 40224 18264 40288
rect 17944 39200 18264 40224
rect 17944 39136 17952 39200
rect 18016 39136 18032 39200
rect 18096 39136 18112 39200
rect 18176 39136 18192 39200
rect 18256 39136 18264 39200
rect 17944 38112 18264 39136
rect 17944 38048 17952 38112
rect 18016 38048 18032 38112
rect 18096 38048 18112 38112
rect 18176 38048 18192 38112
rect 18256 38048 18264 38112
rect 17944 37024 18264 38048
rect 17944 36960 17952 37024
rect 18016 36960 18032 37024
rect 18096 36960 18112 37024
rect 18176 36960 18192 37024
rect 18256 36960 18264 37024
rect 17944 35936 18264 36960
rect 17944 35872 17952 35936
rect 18016 35872 18032 35936
rect 18096 35872 18112 35936
rect 18176 35872 18192 35936
rect 18256 35872 18264 35936
rect 17944 34848 18264 35872
rect 17944 34784 17952 34848
rect 18016 34784 18032 34848
rect 18096 34784 18112 34848
rect 18176 34784 18192 34848
rect 18256 34784 18264 34848
rect 17944 33760 18264 34784
rect 17944 33696 17952 33760
rect 18016 33696 18032 33760
rect 18096 33696 18112 33760
rect 18176 33696 18192 33760
rect 18256 33696 18264 33760
rect 17944 32672 18264 33696
rect 17944 32608 17952 32672
rect 18016 32608 18032 32672
rect 18096 32608 18112 32672
rect 18176 32608 18192 32672
rect 18256 32608 18264 32672
rect 17944 31584 18264 32608
rect 17944 31520 17952 31584
rect 18016 31520 18032 31584
rect 18096 31520 18112 31584
rect 18176 31520 18192 31584
rect 18256 31520 18264 31584
rect 17944 30496 18264 31520
rect 17944 30432 17952 30496
rect 18016 30432 18032 30496
rect 18096 30432 18112 30496
rect 18176 30432 18192 30496
rect 18256 30432 18264 30496
rect 17944 29408 18264 30432
rect 17944 29344 17952 29408
rect 18016 29344 18032 29408
rect 18096 29344 18112 29408
rect 18176 29344 18192 29408
rect 18256 29344 18264 29408
rect 17944 28320 18264 29344
rect 22944 53888 23264 54448
rect 22944 53824 22952 53888
rect 23016 53824 23032 53888
rect 23096 53824 23112 53888
rect 23176 53824 23192 53888
rect 23256 53824 23264 53888
rect 22944 52800 23264 53824
rect 22944 52736 22952 52800
rect 23016 52736 23032 52800
rect 23096 52736 23112 52800
rect 23176 52736 23192 52800
rect 23256 52736 23264 52800
rect 22944 51712 23264 52736
rect 22944 51648 22952 51712
rect 23016 51648 23032 51712
rect 23096 51648 23112 51712
rect 23176 51648 23192 51712
rect 23256 51648 23264 51712
rect 22944 50624 23264 51648
rect 22944 50560 22952 50624
rect 23016 50560 23032 50624
rect 23096 50560 23112 50624
rect 23176 50560 23192 50624
rect 23256 50560 23264 50624
rect 22944 49536 23264 50560
rect 22944 49472 22952 49536
rect 23016 49472 23032 49536
rect 23096 49472 23112 49536
rect 23176 49472 23192 49536
rect 23256 49472 23264 49536
rect 22944 48448 23264 49472
rect 22944 48384 22952 48448
rect 23016 48384 23032 48448
rect 23096 48384 23112 48448
rect 23176 48384 23192 48448
rect 23256 48384 23264 48448
rect 22944 47360 23264 48384
rect 22944 47296 22952 47360
rect 23016 47296 23032 47360
rect 23096 47296 23112 47360
rect 23176 47296 23192 47360
rect 23256 47296 23264 47360
rect 22944 46272 23264 47296
rect 22944 46208 22952 46272
rect 23016 46208 23032 46272
rect 23096 46208 23112 46272
rect 23176 46208 23192 46272
rect 23256 46208 23264 46272
rect 22944 45184 23264 46208
rect 22944 45120 22952 45184
rect 23016 45120 23032 45184
rect 23096 45120 23112 45184
rect 23176 45120 23192 45184
rect 23256 45120 23264 45184
rect 22944 44096 23264 45120
rect 22944 44032 22952 44096
rect 23016 44032 23032 44096
rect 23096 44032 23112 44096
rect 23176 44032 23192 44096
rect 23256 44032 23264 44096
rect 22944 43008 23264 44032
rect 22944 42944 22952 43008
rect 23016 42944 23032 43008
rect 23096 42944 23112 43008
rect 23176 42944 23192 43008
rect 23256 42944 23264 43008
rect 22944 41920 23264 42944
rect 22944 41856 22952 41920
rect 23016 41856 23032 41920
rect 23096 41856 23112 41920
rect 23176 41856 23192 41920
rect 23256 41856 23264 41920
rect 22944 40832 23264 41856
rect 22944 40768 22952 40832
rect 23016 40768 23032 40832
rect 23096 40768 23112 40832
rect 23176 40768 23192 40832
rect 23256 40768 23264 40832
rect 22944 39744 23264 40768
rect 22944 39680 22952 39744
rect 23016 39680 23032 39744
rect 23096 39680 23112 39744
rect 23176 39680 23192 39744
rect 23256 39680 23264 39744
rect 22944 38656 23264 39680
rect 22944 38592 22952 38656
rect 23016 38592 23032 38656
rect 23096 38592 23112 38656
rect 23176 38592 23192 38656
rect 23256 38592 23264 38656
rect 22944 37568 23264 38592
rect 22944 37504 22952 37568
rect 23016 37504 23032 37568
rect 23096 37504 23112 37568
rect 23176 37504 23192 37568
rect 23256 37504 23264 37568
rect 22944 36480 23264 37504
rect 22944 36416 22952 36480
rect 23016 36416 23032 36480
rect 23096 36416 23112 36480
rect 23176 36416 23192 36480
rect 23256 36416 23264 36480
rect 22944 35392 23264 36416
rect 22944 35328 22952 35392
rect 23016 35328 23032 35392
rect 23096 35328 23112 35392
rect 23176 35328 23192 35392
rect 23256 35328 23264 35392
rect 22944 34304 23264 35328
rect 22944 34240 22952 34304
rect 23016 34240 23032 34304
rect 23096 34240 23112 34304
rect 23176 34240 23192 34304
rect 23256 34240 23264 34304
rect 22944 33216 23264 34240
rect 22944 33152 22952 33216
rect 23016 33152 23032 33216
rect 23096 33152 23112 33216
rect 23176 33152 23192 33216
rect 23256 33152 23264 33216
rect 22944 32128 23264 33152
rect 22944 32064 22952 32128
rect 23016 32064 23032 32128
rect 23096 32064 23112 32128
rect 23176 32064 23192 32128
rect 23256 32064 23264 32128
rect 22944 31040 23264 32064
rect 22944 30976 22952 31040
rect 23016 30976 23032 31040
rect 23096 30976 23112 31040
rect 23176 30976 23192 31040
rect 23256 30976 23264 31040
rect 22944 29952 23264 30976
rect 22944 29888 22952 29952
rect 23016 29888 23032 29952
rect 23096 29888 23112 29952
rect 23176 29888 23192 29952
rect 23256 29888 23264 29952
rect 21219 29204 21285 29205
rect 21219 29140 21220 29204
rect 21284 29140 21285 29204
rect 21219 29139 21285 29140
rect 17944 28256 17952 28320
rect 18016 28256 18032 28320
rect 18096 28256 18112 28320
rect 18176 28256 18192 28320
rect 18256 28256 18264 28320
rect 17723 27300 17789 27301
rect 17723 27236 17724 27300
rect 17788 27236 17789 27300
rect 17723 27235 17789 27236
rect 12944 26624 12952 26688
rect 13016 26624 13032 26688
rect 13096 26624 13112 26688
rect 13176 26624 13192 26688
rect 13256 26624 13264 26688
rect 12944 25600 13264 26624
rect 12944 25536 12952 25600
rect 13016 25536 13032 25600
rect 13096 25536 13112 25600
rect 13176 25536 13192 25600
rect 13256 25536 13264 25600
rect 12944 24512 13264 25536
rect 15331 25124 15397 25125
rect 15331 25060 15332 25124
rect 15396 25060 15397 25124
rect 15331 25059 15397 25060
rect 12944 24448 12952 24512
rect 13016 24448 13032 24512
rect 13096 24448 13112 24512
rect 13176 24448 13192 24512
rect 13256 24448 13264 24512
rect 12944 23424 13264 24448
rect 12944 23360 12952 23424
rect 13016 23360 13032 23424
rect 13096 23360 13112 23424
rect 13176 23360 13192 23424
rect 13256 23360 13264 23424
rect 12944 22336 13264 23360
rect 12944 22272 12952 22336
rect 13016 22272 13032 22336
rect 13096 22272 13112 22336
rect 13176 22272 13192 22336
rect 13256 22272 13264 22336
rect 12944 21248 13264 22272
rect 12944 21184 12952 21248
rect 13016 21184 13032 21248
rect 13096 21184 13112 21248
rect 13176 21184 13192 21248
rect 13256 21184 13264 21248
rect 12944 20160 13264 21184
rect 12944 20096 12952 20160
rect 13016 20096 13032 20160
rect 13096 20096 13112 20160
rect 13176 20096 13192 20160
rect 13256 20096 13264 20160
rect 12944 19072 13264 20096
rect 12944 19008 12952 19072
rect 13016 19008 13032 19072
rect 13096 19008 13112 19072
rect 13176 19008 13192 19072
rect 13256 19008 13264 19072
rect 12944 17984 13264 19008
rect 12944 17920 12952 17984
rect 13016 17920 13032 17984
rect 13096 17920 13112 17984
rect 13176 17920 13192 17984
rect 13256 17920 13264 17984
rect 12944 16896 13264 17920
rect 12944 16832 12952 16896
rect 13016 16832 13032 16896
rect 13096 16832 13112 16896
rect 13176 16832 13192 16896
rect 13256 16832 13264 16896
rect 12944 15808 13264 16832
rect 13491 16692 13557 16693
rect 13491 16628 13492 16692
rect 13556 16628 13557 16692
rect 13491 16627 13557 16628
rect 12944 15744 12952 15808
rect 13016 15744 13032 15808
rect 13096 15744 13112 15808
rect 13176 15744 13192 15808
rect 13256 15744 13264 15808
rect 12944 14720 13264 15744
rect 12944 14656 12952 14720
rect 13016 14656 13032 14720
rect 13096 14656 13112 14720
rect 13176 14656 13192 14720
rect 13256 14656 13264 14720
rect 12944 13632 13264 14656
rect 12944 13568 12952 13632
rect 13016 13568 13032 13632
rect 13096 13568 13112 13632
rect 13176 13568 13192 13632
rect 13256 13568 13264 13632
rect 12944 12544 13264 13568
rect 12944 12480 12952 12544
rect 13016 12480 13032 12544
rect 13096 12480 13112 12544
rect 13176 12480 13192 12544
rect 13256 12480 13264 12544
rect 12944 11456 13264 12480
rect 12944 11392 12952 11456
rect 13016 11392 13032 11456
rect 13096 11392 13112 11456
rect 13176 11392 13192 11456
rect 13256 11392 13264 11456
rect 12944 10368 13264 11392
rect 12944 10304 12952 10368
rect 13016 10304 13032 10368
rect 13096 10304 13112 10368
rect 13176 10304 13192 10368
rect 13256 10304 13264 10368
rect 12944 9280 13264 10304
rect 12944 9216 12952 9280
rect 13016 9216 13032 9280
rect 13096 9216 13112 9280
rect 13176 9216 13192 9280
rect 13256 9216 13264 9280
rect 12944 8192 13264 9216
rect 12944 8128 12952 8192
rect 13016 8128 13032 8192
rect 13096 8128 13112 8192
rect 13176 8128 13192 8192
rect 13256 8128 13264 8192
rect 12944 7104 13264 8128
rect 12944 7040 12952 7104
rect 13016 7040 13032 7104
rect 13096 7040 13112 7104
rect 13176 7040 13192 7104
rect 13256 7040 13264 7104
rect 12944 6016 13264 7040
rect 12944 5952 12952 6016
rect 13016 5952 13032 6016
rect 13096 5952 13112 6016
rect 13176 5952 13192 6016
rect 13256 5952 13264 6016
rect 12944 4928 13264 5952
rect 12944 4864 12952 4928
rect 13016 4864 13032 4928
rect 13096 4864 13112 4928
rect 13176 4864 13192 4928
rect 13256 4864 13264 4928
rect 12944 3840 13264 4864
rect 12944 3776 12952 3840
rect 13016 3776 13032 3840
rect 13096 3776 13112 3840
rect 13176 3776 13192 3840
rect 13256 3776 13264 3840
rect 12944 2752 13264 3776
rect 13494 3093 13554 16627
rect 13675 16556 13741 16557
rect 13675 16492 13676 16556
rect 13740 16492 13741 16556
rect 13675 16491 13741 16492
rect 13678 15469 13738 16491
rect 13675 15468 13741 15469
rect 13675 15404 13676 15468
rect 13740 15404 13741 15468
rect 13675 15403 13741 15404
rect 13678 11797 13738 15403
rect 13675 11796 13741 11797
rect 13675 11732 13676 11796
rect 13740 11732 13741 11796
rect 13675 11731 13741 11732
rect 14963 11660 15029 11661
rect 14963 11596 14964 11660
rect 15028 11596 15029 11660
rect 14963 11595 15029 11596
rect 14966 9893 15026 11595
rect 14963 9892 15029 9893
rect 14963 9828 14964 9892
rect 15028 9828 15029 9892
rect 14963 9827 15029 9828
rect 13491 3092 13557 3093
rect 13491 3028 13492 3092
rect 13556 3028 13557 3092
rect 13491 3027 13557 3028
rect 12944 2688 12952 2752
rect 13016 2688 13032 2752
rect 13096 2688 13112 2752
rect 13176 2688 13192 2752
rect 13256 2688 13264 2752
rect 12944 2128 13264 2688
rect 14966 2549 15026 9827
rect 15334 7989 15394 25059
rect 17171 23764 17237 23765
rect 17171 23700 17172 23764
rect 17236 23700 17237 23764
rect 17171 23699 17237 23700
rect 16803 17100 16869 17101
rect 16803 17036 16804 17100
rect 16868 17036 16869 17100
rect 16803 17035 16869 17036
rect 16067 14244 16133 14245
rect 16067 14180 16068 14244
rect 16132 14180 16133 14244
rect 16067 14179 16133 14180
rect 15331 7988 15397 7989
rect 15331 7924 15332 7988
rect 15396 7924 15397 7988
rect 15331 7923 15397 7924
rect 15334 7581 15394 7923
rect 15331 7580 15397 7581
rect 15331 7516 15332 7580
rect 15396 7516 15397 7580
rect 15331 7515 15397 7516
rect 14963 2548 15029 2549
rect 14963 2484 14964 2548
rect 15028 2484 15029 2548
rect 14963 2483 15029 2484
rect 16070 2413 16130 14179
rect 16806 10301 16866 17035
rect 17174 16285 17234 23699
rect 17171 16284 17237 16285
rect 17171 16220 17172 16284
rect 17236 16220 17237 16284
rect 17171 16219 17237 16220
rect 17355 15332 17421 15333
rect 17355 15268 17356 15332
rect 17420 15268 17421 15332
rect 17355 15267 17421 15268
rect 16803 10300 16869 10301
rect 16803 10236 16804 10300
rect 16868 10236 16869 10300
rect 16803 10235 16869 10236
rect 17358 3637 17418 15267
rect 17726 10437 17786 27235
rect 17944 27232 18264 28256
rect 17944 27168 17952 27232
rect 18016 27168 18032 27232
rect 18096 27168 18112 27232
rect 18176 27168 18192 27232
rect 18256 27168 18264 27232
rect 17944 26144 18264 27168
rect 18643 26348 18709 26349
rect 18643 26284 18644 26348
rect 18708 26284 18709 26348
rect 18643 26283 18709 26284
rect 17944 26080 17952 26144
rect 18016 26080 18032 26144
rect 18096 26080 18112 26144
rect 18176 26080 18192 26144
rect 18256 26080 18264 26144
rect 17944 25056 18264 26080
rect 17944 24992 17952 25056
rect 18016 24992 18032 25056
rect 18096 24992 18112 25056
rect 18176 24992 18192 25056
rect 18256 24992 18264 25056
rect 17944 23968 18264 24992
rect 17944 23904 17952 23968
rect 18016 23904 18032 23968
rect 18096 23904 18112 23968
rect 18176 23904 18192 23968
rect 18256 23904 18264 23968
rect 17944 22880 18264 23904
rect 17944 22816 17952 22880
rect 18016 22816 18032 22880
rect 18096 22816 18112 22880
rect 18176 22816 18192 22880
rect 18256 22816 18264 22880
rect 17944 21792 18264 22816
rect 17944 21728 17952 21792
rect 18016 21728 18032 21792
rect 18096 21728 18112 21792
rect 18176 21728 18192 21792
rect 18256 21728 18264 21792
rect 17944 20704 18264 21728
rect 17944 20640 17952 20704
rect 18016 20640 18032 20704
rect 18096 20640 18112 20704
rect 18176 20640 18192 20704
rect 18256 20640 18264 20704
rect 17944 19616 18264 20640
rect 17944 19552 17952 19616
rect 18016 19552 18032 19616
rect 18096 19552 18112 19616
rect 18176 19552 18192 19616
rect 18256 19552 18264 19616
rect 17944 18528 18264 19552
rect 17944 18464 17952 18528
rect 18016 18464 18032 18528
rect 18096 18464 18112 18528
rect 18176 18464 18192 18528
rect 18256 18464 18264 18528
rect 17944 17440 18264 18464
rect 18646 18325 18706 26283
rect 19379 25124 19445 25125
rect 19379 25060 19380 25124
rect 19444 25060 19445 25124
rect 19379 25059 19445 25060
rect 19195 19412 19261 19413
rect 19195 19348 19196 19412
rect 19260 19348 19261 19412
rect 19195 19347 19261 19348
rect 18643 18324 18709 18325
rect 18643 18260 18644 18324
rect 18708 18260 18709 18324
rect 18643 18259 18709 18260
rect 18643 18188 18709 18189
rect 18643 18124 18644 18188
rect 18708 18124 18709 18188
rect 18643 18123 18709 18124
rect 17944 17376 17952 17440
rect 18016 17376 18032 17440
rect 18096 17376 18112 17440
rect 18176 17376 18192 17440
rect 18256 17376 18264 17440
rect 17944 16352 18264 17376
rect 17944 16288 17952 16352
rect 18016 16288 18032 16352
rect 18096 16288 18112 16352
rect 18176 16288 18192 16352
rect 18256 16288 18264 16352
rect 17944 15264 18264 16288
rect 17944 15200 17952 15264
rect 18016 15200 18032 15264
rect 18096 15200 18112 15264
rect 18176 15200 18192 15264
rect 18256 15200 18264 15264
rect 17944 14176 18264 15200
rect 17944 14112 17952 14176
rect 18016 14112 18032 14176
rect 18096 14112 18112 14176
rect 18176 14112 18192 14176
rect 18256 14112 18264 14176
rect 17944 13088 18264 14112
rect 17944 13024 17952 13088
rect 18016 13024 18032 13088
rect 18096 13024 18112 13088
rect 18176 13024 18192 13088
rect 18256 13024 18264 13088
rect 17944 12000 18264 13024
rect 18646 12885 18706 18123
rect 18643 12884 18709 12885
rect 18643 12820 18644 12884
rect 18708 12820 18709 12884
rect 18643 12819 18709 12820
rect 17944 11936 17952 12000
rect 18016 11936 18032 12000
rect 18096 11936 18112 12000
rect 18176 11936 18192 12000
rect 18256 11936 18264 12000
rect 17944 10912 18264 11936
rect 18646 11525 18706 12819
rect 18643 11524 18709 11525
rect 18643 11460 18644 11524
rect 18708 11460 18709 11524
rect 18643 11459 18709 11460
rect 17944 10848 17952 10912
rect 18016 10848 18032 10912
rect 18096 10848 18112 10912
rect 18176 10848 18192 10912
rect 18256 10848 18264 10912
rect 17723 10436 17789 10437
rect 17723 10372 17724 10436
rect 17788 10372 17789 10436
rect 17723 10371 17789 10372
rect 17944 9824 18264 10848
rect 17944 9760 17952 9824
rect 18016 9760 18032 9824
rect 18096 9760 18112 9824
rect 18176 9760 18192 9824
rect 18256 9760 18264 9824
rect 17944 8736 18264 9760
rect 19198 9621 19258 19347
rect 19195 9620 19261 9621
rect 19195 9556 19196 9620
rect 19260 9556 19261 9620
rect 19195 9555 19261 9556
rect 17944 8672 17952 8736
rect 18016 8672 18032 8736
rect 18096 8672 18112 8736
rect 18176 8672 18192 8736
rect 18256 8672 18264 8736
rect 17944 7648 18264 8672
rect 17944 7584 17952 7648
rect 18016 7584 18032 7648
rect 18096 7584 18112 7648
rect 18176 7584 18192 7648
rect 18256 7584 18264 7648
rect 17944 6560 18264 7584
rect 17944 6496 17952 6560
rect 18016 6496 18032 6560
rect 18096 6496 18112 6560
rect 18176 6496 18192 6560
rect 18256 6496 18264 6560
rect 17944 5472 18264 6496
rect 17944 5408 17952 5472
rect 18016 5408 18032 5472
rect 18096 5408 18112 5472
rect 18176 5408 18192 5472
rect 18256 5408 18264 5472
rect 17944 4384 18264 5408
rect 17944 4320 17952 4384
rect 18016 4320 18032 4384
rect 18096 4320 18112 4384
rect 18176 4320 18192 4384
rect 18256 4320 18264 4384
rect 17355 3636 17421 3637
rect 17355 3572 17356 3636
rect 17420 3572 17421 3636
rect 17355 3571 17421 3572
rect 17944 3296 18264 4320
rect 19382 3501 19442 25059
rect 21035 24988 21101 24989
rect 21035 24924 21036 24988
rect 21100 24924 21101 24988
rect 21035 24923 21101 24924
rect 19563 16692 19629 16693
rect 19563 16628 19564 16692
rect 19628 16628 19629 16692
rect 19563 16627 19629 16628
rect 19566 13293 19626 16627
rect 19563 13292 19629 13293
rect 19563 13228 19564 13292
rect 19628 13228 19629 13292
rect 19563 13227 19629 13228
rect 20115 12612 20181 12613
rect 20115 12548 20116 12612
rect 20180 12548 20181 12612
rect 20115 12547 20181 12548
rect 19563 8396 19629 8397
rect 19563 8332 19564 8396
rect 19628 8332 19629 8396
rect 19563 8331 19629 8332
rect 19566 3637 19626 8331
rect 20118 4045 20178 12547
rect 20115 4044 20181 4045
rect 20115 3980 20116 4044
rect 20180 3980 20181 4044
rect 20115 3979 20181 3980
rect 19563 3636 19629 3637
rect 19563 3572 19564 3636
rect 19628 3572 19629 3636
rect 19563 3571 19629 3572
rect 19379 3500 19445 3501
rect 19379 3436 19380 3500
rect 19444 3436 19445 3500
rect 19379 3435 19445 3436
rect 17944 3232 17952 3296
rect 18016 3232 18032 3296
rect 18096 3232 18112 3296
rect 18176 3232 18192 3296
rect 18256 3232 18264 3296
rect 16067 2412 16133 2413
rect 16067 2348 16068 2412
rect 16132 2348 16133 2412
rect 16067 2347 16133 2348
rect 17944 2208 18264 3232
rect 21038 2549 21098 24923
rect 21222 17373 21282 29139
rect 22691 29068 22757 29069
rect 22691 29004 22692 29068
rect 22756 29004 22757 29068
rect 22691 29003 22757 29004
rect 22139 25804 22205 25805
rect 22139 25740 22140 25804
rect 22204 25740 22205 25804
rect 22139 25739 22205 25740
rect 22142 23493 22202 25739
rect 22139 23492 22205 23493
rect 22139 23428 22140 23492
rect 22204 23428 22205 23492
rect 22139 23427 22205 23428
rect 21403 18052 21469 18053
rect 21403 17988 21404 18052
rect 21468 17988 21469 18052
rect 21403 17987 21469 17988
rect 21219 17372 21285 17373
rect 21219 17308 21220 17372
rect 21284 17308 21285 17372
rect 21219 17307 21285 17308
rect 21406 5541 21466 17987
rect 22139 17100 22205 17101
rect 22139 17036 22140 17100
rect 22204 17036 22205 17100
rect 22139 17035 22205 17036
rect 21403 5540 21469 5541
rect 21403 5476 21404 5540
rect 21468 5476 21469 5540
rect 21403 5475 21469 5476
rect 22142 4045 22202 17035
rect 22694 13021 22754 29003
rect 22944 28864 23264 29888
rect 22944 28800 22952 28864
rect 23016 28800 23032 28864
rect 23096 28800 23112 28864
rect 23176 28800 23192 28864
rect 23256 28800 23264 28864
rect 22944 27776 23264 28800
rect 22944 27712 22952 27776
rect 23016 27712 23032 27776
rect 23096 27712 23112 27776
rect 23176 27712 23192 27776
rect 23256 27712 23264 27776
rect 22944 26688 23264 27712
rect 22944 26624 22952 26688
rect 23016 26624 23032 26688
rect 23096 26624 23112 26688
rect 23176 26624 23192 26688
rect 23256 26624 23264 26688
rect 22944 25600 23264 26624
rect 22944 25536 22952 25600
rect 23016 25536 23032 25600
rect 23096 25536 23112 25600
rect 23176 25536 23192 25600
rect 23256 25536 23264 25600
rect 22944 24512 23264 25536
rect 22944 24448 22952 24512
rect 23016 24448 23032 24512
rect 23096 24448 23112 24512
rect 23176 24448 23192 24512
rect 23256 24448 23264 24512
rect 22944 23424 23264 24448
rect 22944 23360 22952 23424
rect 23016 23360 23032 23424
rect 23096 23360 23112 23424
rect 23176 23360 23192 23424
rect 23256 23360 23264 23424
rect 22944 22336 23264 23360
rect 22944 22272 22952 22336
rect 23016 22272 23032 22336
rect 23096 22272 23112 22336
rect 23176 22272 23192 22336
rect 23256 22272 23264 22336
rect 22944 21248 23264 22272
rect 22944 21184 22952 21248
rect 23016 21184 23032 21248
rect 23096 21184 23112 21248
rect 23176 21184 23192 21248
rect 23256 21184 23264 21248
rect 22944 20160 23264 21184
rect 22944 20096 22952 20160
rect 23016 20096 23032 20160
rect 23096 20096 23112 20160
rect 23176 20096 23192 20160
rect 23256 20096 23264 20160
rect 22944 19072 23264 20096
rect 22944 19008 22952 19072
rect 23016 19008 23032 19072
rect 23096 19008 23112 19072
rect 23176 19008 23192 19072
rect 23256 19008 23264 19072
rect 22944 17984 23264 19008
rect 22944 17920 22952 17984
rect 23016 17920 23032 17984
rect 23096 17920 23112 17984
rect 23176 17920 23192 17984
rect 23256 17920 23264 17984
rect 22944 16896 23264 17920
rect 22944 16832 22952 16896
rect 23016 16832 23032 16896
rect 23096 16832 23112 16896
rect 23176 16832 23192 16896
rect 23256 16832 23264 16896
rect 22944 15808 23264 16832
rect 22944 15744 22952 15808
rect 23016 15744 23032 15808
rect 23096 15744 23112 15808
rect 23176 15744 23192 15808
rect 23256 15744 23264 15808
rect 22944 14720 23264 15744
rect 22944 14656 22952 14720
rect 23016 14656 23032 14720
rect 23096 14656 23112 14720
rect 23176 14656 23192 14720
rect 23256 14656 23264 14720
rect 22944 13632 23264 14656
rect 22944 13568 22952 13632
rect 23016 13568 23032 13632
rect 23096 13568 23112 13632
rect 23176 13568 23192 13632
rect 23256 13568 23264 13632
rect 22691 13020 22757 13021
rect 22691 12956 22692 13020
rect 22756 12956 22757 13020
rect 22691 12955 22757 12956
rect 22944 12544 23264 13568
rect 22944 12480 22952 12544
rect 23016 12480 23032 12544
rect 23096 12480 23112 12544
rect 23176 12480 23192 12544
rect 23256 12480 23264 12544
rect 22944 11456 23264 12480
rect 22944 11392 22952 11456
rect 23016 11392 23032 11456
rect 23096 11392 23112 11456
rect 23176 11392 23192 11456
rect 23256 11392 23264 11456
rect 22944 10368 23264 11392
rect 22944 10304 22952 10368
rect 23016 10304 23032 10368
rect 23096 10304 23112 10368
rect 23176 10304 23192 10368
rect 23256 10304 23264 10368
rect 22944 9280 23264 10304
rect 22944 9216 22952 9280
rect 23016 9216 23032 9280
rect 23096 9216 23112 9280
rect 23176 9216 23192 9280
rect 23256 9216 23264 9280
rect 22944 8192 23264 9216
rect 22944 8128 22952 8192
rect 23016 8128 23032 8192
rect 23096 8128 23112 8192
rect 23176 8128 23192 8192
rect 23256 8128 23264 8192
rect 22944 7104 23264 8128
rect 22944 7040 22952 7104
rect 23016 7040 23032 7104
rect 23096 7040 23112 7104
rect 23176 7040 23192 7104
rect 23256 7040 23264 7104
rect 22944 6016 23264 7040
rect 23427 7036 23493 7037
rect 23427 6972 23428 7036
rect 23492 6972 23493 7036
rect 23427 6971 23493 6972
rect 22944 5952 22952 6016
rect 23016 5952 23032 6016
rect 23096 5952 23112 6016
rect 23176 5952 23192 6016
rect 23256 5952 23264 6016
rect 22944 4928 23264 5952
rect 23430 5541 23490 6971
rect 23427 5540 23493 5541
rect 23427 5476 23428 5540
rect 23492 5476 23493 5540
rect 23427 5475 23493 5476
rect 22944 4864 22952 4928
rect 23016 4864 23032 4928
rect 23096 4864 23112 4928
rect 23176 4864 23192 4928
rect 23256 4864 23264 4928
rect 22139 4044 22205 4045
rect 22139 3980 22140 4044
rect 22204 3980 22205 4044
rect 22139 3979 22205 3980
rect 22944 3840 23264 4864
rect 22944 3776 22952 3840
rect 23016 3776 23032 3840
rect 23096 3776 23112 3840
rect 23176 3776 23192 3840
rect 23256 3776 23264 3840
rect 22944 2752 23264 3776
rect 22944 2688 22952 2752
rect 23016 2688 23032 2752
rect 23096 2688 23112 2752
rect 23176 2688 23192 2752
rect 23256 2688 23264 2752
rect 21035 2548 21101 2549
rect 21035 2484 21036 2548
rect 21100 2484 21101 2548
rect 21035 2483 21101 2484
rect 17944 2144 17952 2208
rect 18016 2144 18032 2208
rect 18096 2144 18112 2208
rect 18176 2144 18192 2208
rect 18256 2144 18264 2208
rect 17944 2128 18264 2144
rect 22944 2128 23264 2688
use sky130_fd_sc_hd__clkbuf_2  _104_ pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1679235063
transform 1 0 23460 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  _105_ pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1679235063
transform 1 0 12972 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _106_ pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1679235063
transform 1 0 11040 0 1 3264
box -38 -48 958 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _107_
timestamp 1679235063
transform 1 0 12880 0 1 4352
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_1  _108_
timestamp 1679235063
transform 1 0 16468 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _109_
timestamp 1679235063
transform 1 0 14260 0 -1 8704
box -38 -48 958 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _110_
timestamp 1679235063
transform 1 0 21988 0 -1 10880
box -38 -48 958 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _111_
timestamp 1679235063
transform 1 0 10304 0 1 8704
box -38 -48 958 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _112_
timestamp 1679235063
transform 1 0 11592 0 1 4352
box -38 -48 958 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _113_
timestamp 1679235063
transform 1 0 10304 0 -1 4352
box -38 -48 958 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _114_
timestamp 1679235063
transform 1 0 11684 0 -1 5440
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_1  _115_
timestamp 1679235063
transform 1 0 8372 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _116_
timestamp 1679235063
transform 1 0 9108 0 1 10880
box -38 -48 958 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _117_
timestamp 1679235063
transform 1 0 16836 0 -1 15232
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_1  _118_
timestamp 1679235063
transform 1 0 23828 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _119_
timestamp 1679235063
transform 1 0 18676 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _120_
timestamp 1679235063
transform 1 0 17204 0 1 14144
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_2  _121_
timestamp 1679235063
transform 1 0 21160 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  _122_
timestamp 1679235063
transform 1 0 23276 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  _123_
timestamp 1679235063
transform 1 0 21528 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  _124_
timestamp 1679235063
transform 1 0 20884 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _125_
timestamp 1679235063
transform 1 0 15456 0 -1 18496
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_1  _126_
timestamp 1679235063
transform 1 0 14352 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _127_
timestamp 1679235063
transform 1 0 18676 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _128_
timestamp 1679235063
transform 1 0 21988 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _129_
timestamp 1679235063
transform 1 0 20792 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _130_
timestamp 1679235063
transform 1 0 17388 0 1 20672
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_1  _131_
timestamp 1679235063
transform 1 0 23828 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  _132_
timestamp 1679235063
transform 1 0 21804 0 1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _133_
timestamp 1679235063
transform 1 0 18584 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _134_
timestamp 1679235063
transform 1 0 19872 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _135_
timestamp 1679235063
transform 1 0 20792 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _136_
timestamp 1679235063
transform 1 0 16836 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _137_
timestamp 1679235063
transform 1 0 17112 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  _138_
timestamp 1679235063
transform 1 0 14444 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  _139_
timestamp 1679235063
transform 1 0 14260 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _140_
timestamp 1679235063
transform 1 0 16836 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _141_
timestamp 1679235063
transform 1 0 17940 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _142_
timestamp 1679235063
transform 1 0 19412 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _143_
timestamp 1679235063
transform 1 0 18492 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _144_
timestamp 1679235063
transform 1 0 19412 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _145_
timestamp 1679235063
transform 1 0 19412 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _146_
timestamp 1679235063
transform 1 0 18952 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _147_
timestamp 1679235063
transform 1 0 21068 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _148_
timestamp 1679235063
transform 1 0 16008 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _149_
timestamp 1679235063
transform 1 0 15548 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _150_
timestamp 1679235063
transform 1 0 20792 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _151_
timestamp 1679235063
transform 1 0 20148 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _152_
timestamp 1679235063
transform 1 0 21160 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _153_
timestamp 1679235063
transform 1 0 21896 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  _154_
timestamp 1679235063
transform 1 0 18676 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  _155_
timestamp 1679235063
transform 1 0 19412 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _156_
timestamp 1679235063
transform 1 0 19412 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _157_
timestamp 1679235063
transform 1 0 20516 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _158_
timestamp 1679235063
transform 1 0 24564 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _159_
timestamp 1679235063
transform 1 0 21988 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _160_
timestamp 1679235063
transform 1 0 16008 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _161_
timestamp 1679235063
transform 1 0 22724 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _162_
timestamp 1679235063
transform 1 0 24564 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _163_
timestamp 1679235063
transform 1 0 24564 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  _164_
timestamp 1679235063
transform 1 0 4968 0 -1 53312
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _165_
timestamp 1679235063
transform 1 0 6532 0 -1 53312
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _166_
timestamp 1679235063
transform 1 0 7636 0 1 52224
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  _167_
timestamp 1679235063
transform 1 0 8648 0 -1 52224
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA_1 pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1679235063
transform 1 0 10764 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_2
timestamp 1679235063
transform 1 0 10120 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_3
timestamp 1679235063
transform 1 0 23276 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_4
timestamp 1679235063
transform 1 0 10212 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__134__A
timestamp 1679235063
transform 1 0 20792 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__135__A
timestamp 1679235063
transform 1 0 21436 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__136__A
timestamp 1679235063
transform 1 0 18032 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__137__A
timestamp 1679235063
transform 1 0 16744 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__138__A
timestamp 1679235063
transform 1 0 14076 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__139__A
timestamp 1679235063
transform 1 0 14812 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__142__A
timestamp 1679235063
transform 1 0 20424 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__143__A
timestamp 1679235063
transform 1 0 19228 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__144__A
timestamp 1679235063
transform 1 0 20332 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__145__A
timestamp 1679235063
transform 1 0 19964 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__150__A
timestamp 1679235063
transform 1 0 21528 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__151__A
timestamp 1679235063
transform 1 0 21344 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__152__A
timestamp 1679235063
transform 1 0 21528 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__153__A
timestamp 1679235063
transform 1 0 20608 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__154__A
timestamp 1679235063
transform 1 0 18860 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__158__A
timestamp 1679235063
transform 1 0 25116 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__162__A
timestamp 1679235063
transform 1 0 25116 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__163__A
timestamp 1679235063
transform 1 0 25116 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_cby_0__8_.cby_0__1_.mem_right_ipin_0.sky130_fd_sc_hd__dfrtp_1_0__RESET_B
timestamp 1679235063
transform 1 0 7360 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_cby_0__8_.cby_0__1_.mem_right_ipin_0.sky130_fd_sc_hd__dfrtp_1_1__D
timestamp 1679235063
transform 1 0 7820 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_cby_0__8_.cby_0__1_.mem_right_ipin_0.sky130_fd_sc_hd__dfrtp_1_1__RESET_B
timestamp 1679235063
transform 1 0 11224 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_cby_0__8_.cby_0__1_.mem_right_ipin_0.sky130_fd_sc_hd__dfrtp_1_2__RESET_B
timestamp 1679235063
transform 1 0 8556 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_cby_0__8_.cby_0__1_.mem_right_ipin_0.sky130_fd_sc_hd__dfrtp_1_3__RESET_B
timestamp 1679235063
transform 1 0 7912 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_cby_0__8_.cby_0__1_.mem_right_ipin_1.sky130_fd_sc_hd__dfrtp_1_0__RESET_B
timestamp 1679235063
transform 1 0 9844 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_cby_0__8_.cby_0__1_.mem_right_ipin_1.sky130_fd_sc_hd__dfrtp_1_1__RESET_B
timestamp 1679235063
transform 1 0 11132 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_cby_0__8_.cby_0__1_.mem_right_ipin_1.sky130_fd_sc_hd__dfrtp_1_2__RESET_B
timestamp 1679235063
transform 1 0 9200 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_cby_0__8_.cby_0__1_.mem_right_ipin_1.sky130_fd_sc_hd__dfrtp_1_3__RESET_B
timestamp 1679235063
transform 1 0 8372 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_cby_0__8_.cby_0__1_.mem_right_ipin_2.sky130_fd_sc_hd__dfrtp_1_0__RESET_B
timestamp 1679235063
transform 1 0 9568 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_cby_0__8_.cby_0__1_.mem_right_ipin_2.sky130_fd_sc_hd__dfrtp_1_1__RESET_B
timestamp 1679235063
transform 1 0 12236 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_cby_0__8_.cby_0__1_.mem_right_ipin_2.sky130_fd_sc_hd__dfrtp_1_2__RESET_B
timestamp 1679235063
transform 1 0 9476 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_cby_0__8_.cby_0__1_.mem_right_ipin_2.sky130_fd_sc_hd__dfrtp_1_3__RESET_B
timestamp 1679235063
transform 1 0 8924 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_cby_0__8_.cby_0__1_.mem_right_ipin_3.sky130_fd_sc_hd__dfrtp_1_0__RESET_B
timestamp 1679235063
transform 1 0 9844 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_cby_0__8_.cby_0__1_.mem_right_ipin_3.sky130_fd_sc_hd__dfrtp_1_1__RESET_B
timestamp 1679235063
transform 1 0 11408 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_cby_0__8_.cby_0__1_.mem_right_ipin_3.sky130_fd_sc_hd__dfrtp_1_2__D
timestamp 1679235063
transform 1 0 9108 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_cby_0__8_.cby_0__1_.mem_right_ipin_3.sky130_fd_sc_hd__dfrtp_1_2__RESET_B
timestamp 1679235063
transform 1 0 8924 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_cby_0__8_.cby_0__1_.mem_right_ipin_3.sky130_fd_sc_hd__dfrtp_1_3__RESET_B
timestamp 1679235063
transform 1 0 11132 0 1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_cby_0__8_.cby_0__1_.mux_right_ipin_0.mux_l1_in_0__A0
timestamp 1679235063
transform 1 0 16560 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_cby_0__8_.cby_0__1_.mux_right_ipin_0.mux_l1_in_0__S
timestamp 1679235063
transform 1 0 15640 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_cby_0__8_.cby_0__1_.mux_right_ipin_0.mux_l1_in_1__A1
timestamp 1679235063
transform 1 0 13616 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_cby_0__8_.cby_0__1_.mux_right_ipin_0.mux_l1_in_1__S
timestamp 1679235063
transform 1 0 13524 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_cby_0__8_.cby_0__1_.mux_right_ipin_0.mux_l1_in_2__A1
timestamp 1679235063
transform 1 0 13800 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_cby_0__8_.cby_0__1_.mux_right_ipin_0.mux_l1_in_2__S
timestamp 1679235063
transform 1 0 14076 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_cby_0__8_.cby_0__1_.mux_right_ipin_0.mux_l1_in_3__A0
timestamp 1679235063
transform 1 0 16192 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_cby_0__8_.cby_0__1_.mux_right_ipin_0.mux_l1_in_3__A1
timestamp 1679235063
transform 1 0 16008 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_cby_0__8_.cby_0__1_.mux_right_ipin_0.mux_l1_in_3__S
timestamp 1679235063
transform 1 0 15548 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_cby_0__8_.cby_0__1_.mux_right_ipin_0.mux_l1_in_4__A0
timestamp 1679235063
transform 1 0 13616 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_cby_0__8_.cby_0__1_.mux_right_ipin_0.mux_l1_in_4__A1
timestamp 1679235063
transform 1 0 13616 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_cby_0__8_.cby_0__1_.mux_right_ipin_0.mux_l1_in_4__S
timestamp 1679235063
transform 1 0 11592 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_cby_0__8_.cby_0__1_.mux_right_ipin_0.mux_l2_in_2__A0
timestamp 1679235063
transform 1 0 8924 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_cby_0__8_.cby_0__1_.mux_right_ipin_0.mux_l2_in_3__A1
timestamp 1679235063
transform 1 0 12604 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_cby_0__8_.cby_0__1_.mux_right_ipin_1.mux_l1_in_0__A0
timestamp 1679235063
transform 1 0 16744 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_cby_0__8_.cby_0__1_.mux_right_ipin_1.mux_l1_in_1__A1
timestamp 1679235063
transform 1 0 15180 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_cby_0__8_.cby_0__1_.mux_right_ipin_1.mux_l1_in_3__A0
timestamp 1679235063
transform 1 0 16836 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_cby_0__8_.cby_0__1_.mux_right_ipin_1.mux_l1_in_3__A1
timestamp 1679235063
transform 1 0 15088 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_cby_0__8_.cby_0__1_.mux_right_ipin_1.mux_l1_in_4__A0
timestamp 1679235063
transform 1 0 13064 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_cby_0__8_.cby_0__1_.mux_right_ipin_1.mux_l1_in_4__A1
timestamp 1679235063
transform 1 0 12788 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_cby_0__8_.cby_0__1_.mux_right_ipin_1.mux_l2_in_2__A0
timestamp 1679235063
transform 1 0 9384 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_cby_0__8_.cby_0__1_.mux_right_ipin_1.mux_l2_in_3__A1
timestamp 1679235063
transform 1 0 11132 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_cby_0__8_.cby_0__1_.mux_right_ipin_2.mux_l1_in_1__A0
timestamp 1679235063
transform 1 0 14904 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_cby_0__8_.cby_0__1_.mux_right_ipin_2.mux_l1_in_1__A1
timestamp 1679235063
transform 1 0 15088 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_cby_0__8_.cby_0__1_.mux_right_ipin_2.mux_l1_in_3__A1
timestamp 1679235063
transform 1 0 13800 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_cby_0__8_.cby_0__1_.mux_right_ipin_2.mux_l1_in_4__A0
timestamp 1679235063
transform 1 0 14076 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_cby_0__8_.cby_0__1_.mux_right_ipin_2.mux_l1_in_4__A1
timestamp 1679235063
transform 1 0 14260 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_cby_0__8_.cby_0__1_.mux_right_ipin_2.mux_l2_in_2__A0
timestamp 1679235063
transform 1 0 9844 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_cby_0__8_.cby_0__1_.mux_right_ipin_2.mux_l2_in_3__A1
timestamp 1679235063
transform 1 0 16284 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_cby_0__8_.cby_0__1_.mux_right_ipin_3.mux_l1_in_0__A0
timestamp 1679235063
transform 1 0 14260 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_cby_0__8_.cby_0__1_.mux_right_ipin_3.mux_l1_in_1__A1
timestamp 1679235063
transform 1 0 13800 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_cby_0__8_.cby_0__1_.mux_right_ipin_3.mux_l1_in_2__A0
timestamp 1679235063
transform 1 0 14076 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_cby_0__8_.cby_0__1_.mux_right_ipin_3.mux_l1_in_4__A0
timestamp 1679235063
transform 1 0 13800 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_cby_0__8_.cby_0__1_.mux_right_ipin_3.mux_l1_in_4__A1
timestamp 1679235063
transform 1 0 12788 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_cby_0__8_.cby_0__1_.mux_right_ipin_3.mux_l2_in_0__S
timestamp 1679235063
transform 1 0 11408 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_cby_0__8_.cby_0__1_.mux_right_ipin_3.mux_l2_in_1__S
timestamp 1679235063
transform 1 0 11776 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_cby_0__8_.cby_0__1_.mux_right_ipin_3.mux_l2_in_2__A0
timestamp 1679235063
transform 1 0 9752 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_cby_0__8_.cby_0__1_.mux_right_ipin_3.mux_l2_in_2__S
timestamp 1679235063
transform 1 0 11132 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_cby_0__8_.cby_0__1_.mux_right_ipin_3.mux_l2_in_3__A1
timestamp 1679235063
transform 1 0 16836 0 1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_cby_0__8_.cby_0__1_.mux_right_ipin_3.mux_l2_in_3__S
timestamp 1679235063
transform 1 0 16652 0 1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_cby_0__8_.grid_io_left_left_0__1_.logical_tile_io_mode_io__0.logical_tile_io_mode_physical__iopad_0.io_0_.ISOL_EN_GATE_B_N
timestamp 1679235063
transform 1 0 11868 0 1 44608
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_cby_0__8_.grid_io_left_left_0__1_.logical_tile_io_mode_io__0.logical_tile_io_mode_physical__iopad_0.io_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_0__CLK
timestamp 1679235063
transform 1 0 11500 0 -1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_cby_0__8_.grid_io_left_left_0__1_.logical_tile_io_mode_io__0.logical_tile_io_mode_physical__iopad_0.io_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_0__RESET_B
timestamp 1679235063
transform 1 0 11684 0 -1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_cby_0__8_.grid_io_left_left_0__1_.logical_tile_io_mode_io__1.logical_tile_io_mode_physical__iopad_0.io_0_.ISOL_EN_GATE_B_N
timestamp 1679235063
transform 1 0 11132 0 1 46784
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_cby_0__8_.grid_io_left_left_0__1_.logical_tile_io_mode_io__1.logical_tile_io_mode_physical__iopad_0.io_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_0__CLK
timestamp 1679235063
transform 1 0 11500 0 -1 43520
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_cby_0__8_.grid_io_left_left_0__1_.logical_tile_io_mode_io__1.logical_tile_io_mode_physical__iopad_0.io_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_0__RESET_B
timestamp 1679235063
transform 1 0 11684 0 -1 43520
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_cby_0__8_.grid_io_left_left_0__1_.logical_tile_io_mode_io__2.logical_tile_io_mode_physical__iopad_0.io_0_.ISOL_EN_GATE_B_N
timestamp 1679235063
transform 1 0 10120 0 1 48960
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_cby_0__8_.grid_io_left_left_0__1_.logical_tile_io_mode_io__2.logical_tile_io_mode_physical__iopad_0.io_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_0__CLK
timestamp 1679235063
transform 1 0 10856 0 -1 46784
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_cby_0__8_.grid_io_left_left_0__1_.logical_tile_io_mode_io__2.logical_tile_io_mode_physical__iopad_0.io_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_0__RESET_B
timestamp 1679235063
transform 1 0 11040 0 -1 46784
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_cby_0__8_.grid_io_left_left_0__1_.logical_tile_io_mode_io__3.logical_tile_io_mode_physical__iopad_0.io_0_.ISOL_EN_GATE_B_N
timestamp 1679235063
transform 1 0 8372 0 1 51136
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_cby_0__8_.grid_io_left_left_0__1_.logical_tile_io_mode_io__3.logical_tile_io_mode_physical__iopad_0.io_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_0__CLK
timestamp 1679235063
transform 1 0 8648 0 1 48960
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_cby_0__8_.grid_io_left_left_0__1_.logical_tile_io_mode_io__3.logical_tile_io_mode_physical__iopad_0.io_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_0__RESET_B
timestamp 1679235063
transform 1 0 8924 0 1 48960
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_0_prog_clk_A
timestamp 1679235063
transform 1 0 19228 0 1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_4_0_0_prog_clk_A
timestamp 1679235063
transform 1 0 11224 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_4_1_0_prog_clk_A
timestamp 1679235063
transform 1 0 13156 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_4_2_0_prog_clk_A
timestamp 1679235063
transform 1 0 11592 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_4_3_0_prog_clk_A
timestamp 1679235063
transform 1 0 13340 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_4_4_0_prog_clk_A
timestamp 1679235063
transform 1 0 17848 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_4_5_0_prog_clk_A
timestamp 1679235063
transform 1 0 18308 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_4_6_0_prog_clk_A
timestamp 1679235063
transform 1 0 16928 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_4_7_0_prog_clk_A
timestamp 1679235063
transform 1 0 18952 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_4_8_0_prog_clk_A
timestamp 1679235063
transform 1 0 15548 0 -1 31552
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_4_9_0_prog_clk_A
timestamp 1679235063
transform 1 0 15640 0 1 30464
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_4_10_0_prog_clk_A
timestamp 1679235063
transform 1 0 16284 0 -1 34816
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_4_11_0_prog_clk_A
timestamp 1679235063
transform 1 0 16836 0 1 33728
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_4_12_0_prog_clk_A
timestamp 1679235063
transform 1 0 20148 0 -1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_4_13_0_prog_clk_A
timestamp 1679235063
transform 1 0 21988 0 1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_4_14_0_prog_clk_A
timestamp 1679235063
transform 1 0 19688 0 -1 32640
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_4_15_0_prog_clk_A
timestamp 1679235063
transform 1 0 21528 0 -1 32640
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_hold97_A
timestamp 1679235063
transform 1 0 11500 0 -1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input1_A
timestamp 1679235063
transform 1 0 23368 0 1 53312
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input2_A
timestamp 1679235063
transform 1 0 1380 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input3_A
timestamp 1679235063
transform 1 0 22172 0 1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input4_A
timestamp 1679235063
transform 1 0 24748 0 -1 35904
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input5_A
timestamp 1679235063
transform 1 0 24748 0 1 35904
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input6_A
timestamp 1679235063
transform 1 0 24748 0 1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input7_A
timestamp 1679235063
transform 1 0 24656 0 -1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input8_A
timestamp 1679235063
transform 1 0 24656 0 -1 38080
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input9_A
timestamp 1679235063
transform 1 0 25392 0 -1 39168
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input10_A
timestamp 1679235063
transform 1 0 24748 0 1 39168
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input11_A
timestamp 1679235063
transform 1 0 25392 0 1 40256
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input12_A
timestamp 1679235063
transform 1 0 24748 0 -1 41344
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input13_A
timestamp 1679235063
transform 1 0 25392 0 -1 42432
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input14_A
timestamp 1679235063
transform 1 0 16192 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input15_A
timestamp 1679235063
transform 1 0 24656 0 1 42432
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input16_A
timestamp 1679235063
transform 1 0 25392 0 1 43520
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input17_A
timestamp 1679235063
transform 1 0 24656 0 -1 44608
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input18_A
timestamp 1679235063
transform 1 0 25392 0 -1 45696
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input19_A
timestamp 1679235063
transform 1 0 24748 0 1 45696
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input20_A
timestamp 1679235063
transform 1 0 25392 0 1 46784
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input21_A
timestamp 1679235063
transform 1 0 24748 0 -1 47872
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input22_A
timestamp 1679235063
transform 1 0 25392 0 -1 48960
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input23_A
timestamp 1679235063
transform 1 0 24656 0 1 48960
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input24_A
timestamp 1679235063
transform 1 0 25392 0 1 50048
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input25_A
timestamp 1679235063
transform 1 0 18860 0 1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input26_A
timestamp 1679235063
transform 1 0 19228 0 1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input27_A
timestamp 1679235063
transform 1 0 24380 0 1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input28_A
timestamp 1679235063
transform 1 0 25208 0 -1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input29_A
timestamp 1679235063
transform 1 0 24748 0 1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input30_A
timestamp 1679235063
transform 1 0 24104 0 -1 34816
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input31_A
timestamp 1679235063
transform 1 0 24564 0 1 34816
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input32_A
timestamp 1679235063
transform 1 0 24380 0 1 34816
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input33_A
timestamp 1679235063
transform 1 0 2668 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input34_A
timestamp 1679235063
transform 1 0 6072 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input35_A
timestamp 1679235063
transform 1 0 4140 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input36_A
timestamp 1679235063
transform 1 0 5980 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input37_A
timestamp 1679235063
transform 1 0 6992 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input38_A
timestamp 1679235063
transform 1 0 7176 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input39_A
timestamp 1679235063
transform 1 0 7452 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input40_A
timestamp 1679235063
transform 1 0 7636 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input41_A
timestamp 1679235063
transform 1 0 6716 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input42_A
timestamp 1679235063
transform 1 0 7820 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input43_A
timestamp 1679235063
transform 1 0 6532 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input44_A
timestamp 1679235063
transform 1 0 3496 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input45_A
timestamp 1679235063
transform 1 0 9752 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input46_A
timestamp 1679235063
transform 1 0 8004 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input47_A
timestamp 1679235063
transform 1 0 9936 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input48_A
timestamp 1679235063
transform 1 0 9108 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input49_A
timestamp 1679235063
transform 1 0 8924 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input50_A
timestamp 1679235063
transform 1 0 8924 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input51_A
timestamp 1679235063
transform 1 0 11500 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input52_A
timestamp 1679235063
transform 1 0 9292 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input53_A
timestamp 1679235063
transform 1 0 9108 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input54_A
timestamp 1679235063
transform 1 0 9292 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input55_A
timestamp 1679235063
transform 1 0 3772 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input56_A
timestamp 1679235063
transform 1 0 3956 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input57_A
timestamp 1679235063
transform 1 0 3312 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input58_A
timestamp 1679235063
transform 1 0 2852 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input59_A
timestamp 1679235063
transform 1 0 4600 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input60_A
timestamp 1679235063
transform 1 0 4508 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input61_A
timestamp 1679235063
transform 1 0 4692 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input62_A
timestamp 1679235063
transform 1 0 6348 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input63_A
timestamp 1679235063
transform 1 0 14076 0 -1 54400
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input64_A
timestamp 1679235063
transform 1 0 15364 0 -1 54400
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input65_A
timestamp 1679235063
transform 1 0 17296 0 -1 54400
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input66_A
timestamp 1679235063
transform 1 0 18124 0 -1 54400
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input67_A
timestamp 1679235063
transform 1 0 18952 0 -1 54400
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input68_A
timestamp 1679235063
transform 1 0 25392 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input69_A
timestamp 1679235063
transform 1 0 24472 0 -1 51136
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input70_A
timestamp 1679235063
transform 1 0 25392 0 -1 52224
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input71_A
timestamp 1679235063
transform 1 0 24472 0 1 52224
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input72_A
timestamp 1679235063
transform 1 0 24656 0 -1 53312
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input73_A
timestamp 1679235063
transform 1 0 24656 0 -1 54400
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input74_A
timestamp 1679235063
transform 1 0 24656 0 1 53312
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input75_A
timestamp 1679235063
transform 1 0 24380 0 -1 54400
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input76_A
timestamp 1679235063
transform 1 0 24380 0 1 53312
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output77_A
timestamp 1679235063
transform 1 0 14076 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output120_A
timestamp 1679235063
transform 1 0 16100 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__8_.mem_bottom_track_1.sky130_fd_sc_hd__dfrtp_1_0__RESET_B
timestamp 1679235063
transform 1 0 20792 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__8_.mem_bottom_track_1.sky130_fd_sc_hd__dfrtp_1_1__RESET_B
timestamp 1679235063
transform 1 0 22264 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__8_.mem_bottom_track_3.sky130_fd_sc_hd__dfrtp_1_0__RESET_B
timestamp 1679235063
transform 1 0 19504 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__8_.mem_bottom_track_3.sky130_fd_sc_hd__dfrtp_1_1__RESET_B
timestamp 1679235063
transform 1 0 20332 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__8_.mem_bottom_track_5.sky130_fd_sc_hd__dfrtp_1_0__RESET_B
timestamp 1679235063
transform 1 0 19320 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__8_.mem_bottom_track_5.sky130_fd_sc_hd__dfrtp_1_1__RESET_B
timestamp 1679235063
transform 1 0 22908 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__8_.mem_bottom_track_7.sky130_fd_sc_hd__dfrtp_1_0__RESET_B
timestamp 1679235063
transform 1 0 25300 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__8_.mem_bottom_track_7.sky130_fd_sc_hd__dfrtp_1_1__RESET_B
timestamp 1679235063
transform 1 0 21436 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__8_.mem_bottom_track_9.sky130_fd_sc_hd__dfrtp_1_0__RESET_B
timestamp 1679235063
transform 1 0 23092 0 -1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__8_.mem_bottom_track_9.sky130_fd_sc_hd__dfrtp_1_1__RESET_B
timestamp 1679235063
transform 1 0 24104 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__8_.mem_bottom_track_11.sky130_fd_sc_hd__dfrtp_1_0__RESET_B
timestamp 1679235063
transform 1 0 25392 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__8_.mem_bottom_track_11.sky130_fd_sc_hd__dfrtp_1_1__RESET_B
timestamp 1679235063
transform 1 0 25208 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__8_.mem_bottom_track_13.sky130_fd_sc_hd__dfrtp_1_0__RESET_B
timestamp 1679235063
transform 1 0 25392 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__8_.mem_bottom_track_13.sky130_fd_sc_hd__dfrtp_1_1__RESET_B
timestamp 1679235063
transform 1 0 25208 0 -1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__8_.mem_bottom_track_15.sky130_fd_sc_hd__dfrtp_1_0__RESET_B
timestamp 1679235063
transform 1 0 25392 0 -1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__8_.mem_bottom_track_15.sky130_fd_sc_hd__dfrtp_1_1__RESET_B
timestamp 1679235063
transform 1 0 21436 0 1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__8_.mem_bottom_track_17.sky130_fd_sc_hd__dfrtp_1_0__RESET_B
timestamp 1679235063
transform 1 0 20424 0 -1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__8_.mem_bottom_track_17.sky130_fd_sc_hd__dfrtp_1_1__RESET_B
timestamp 1679235063
transform 1 0 19964 0 -1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__8_.mem_bottom_track_19.sky130_fd_sc_hd__dfrtp_1_0__RESET_B
timestamp 1679235063
transform 1 0 18676 0 -1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__8_.mem_bottom_track_19.sky130_fd_sc_hd__dfrtp_1_1__RESET_B
timestamp 1679235063
transform 1 0 18860 0 -1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__8_.mem_bottom_track_29.sky130_fd_sc_hd__dfrtp_1_0__RESET_B
timestamp 1679235063
transform 1 0 18860 0 1 30464
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__8_.mem_bottom_track_29.sky130_fd_sc_hd__dfrtp_1_1__RESET_B
timestamp 1679235063
transform 1 0 18860 0 1 31552
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__8_.mem_bottom_track_31.sky130_fd_sc_hd__dfrtp_1_0__RESET_B
timestamp 1679235063
transform 1 0 19412 0 -1 32640
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__8_.mem_bottom_track_31.sky130_fd_sc_hd__dfrtp_1_1__RESET_B
timestamp 1679235063
transform 1 0 21252 0 -1 31552
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__8_.mem_bottom_track_33.sky130_fd_sc_hd__dfrtp_1_0__RESET_B
timestamp 1679235063
transform 1 0 23828 0 1 30464
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__8_.mem_bottom_track_33.sky130_fd_sc_hd__dfrtp_1_1__RESET_B
timestamp 1679235063
transform 1 0 24104 0 1 30464
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__8_.mem_bottom_track_35.sky130_fd_sc_hd__dfrtp_1_0__RESET_B
timestamp 1679235063
transform 1 0 25300 0 -1 30464
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__8_.mem_bottom_track_35.sky130_fd_sc_hd__dfrtp_1_1__RESET_B
timestamp 1679235063
transform 1 0 25300 0 -1 33728
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__8_.mem_bottom_track_45.sky130_fd_sc_hd__dfrtp_1_0__RESET_B
timestamp 1679235063
transform 1 0 24104 0 1 31552
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__8_.mem_bottom_track_45.sky130_fd_sc_hd__dfrtp_1_1__RESET_B
timestamp 1679235063
transform 1 0 23828 0 1 33728
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__8_.mem_bottom_track_47.sky130_fd_sc_hd__dfrtp_1_0__RESET_B
timestamp 1679235063
transform 1 0 23644 0 1 33728
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__8_.mem_bottom_track_47.sky130_fd_sc_hd__dfrtp_1_1__RESET_B
timestamp 1679235063
transform 1 0 21436 0 -1 33728
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__8_.mem_bottom_track_49.sky130_fd_sc_hd__dfrtp_1_0__RESET_B
timestamp 1679235063
transform 1 0 21252 0 1 34816
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__8_.mem_bottom_track_49.sky130_fd_sc_hd__dfrtp_1_1__RESET_B
timestamp 1679235063
transform 1 0 21436 0 1 32640
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__8_.mem_bottom_track_51.sky130_fd_sc_hd__dfrtp_1_0__RESET_B
timestamp 1679235063
transform 1 0 24012 0 1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__8_.mem_bottom_track_51.sky130_fd_sc_hd__dfrtp_1_1__RESET_B
timestamp 1679235063
transform 1 0 24104 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__8_.mem_right_track_0.sky130_fd_sc_hd__dfrtp_1_0__RESET_B
timestamp 1679235063
transform 1 0 22448 0 1 44608
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__8_.mem_right_track_0.sky130_fd_sc_hd__dfrtp_1_1__RESET_B
timestamp 1679235063
transform 1 0 15364 0 -1 31552
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__8_.mem_right_track_0.sky130_fd_sc_hd__dfrtp_1_2__RESET_B
timestamp 1679235063
transform 1 0 11132 0 1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__8_.mem_right_track_2.sky130_fd_sc_hd__dfrtp_1_0__RESET_B
timestamp 1679235063
transform 1 0 12052 0 -1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__8_.mem_right_track_2.sky130_fd_sc_hd__dfrtp_1_1__RESET_B
timestamp 1679235063
transform 1 0 12604 0 -1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__8_.mem_right_track_2.sky130_fd_sc_hd__dfrtp_1_2__RESET_B
timestamp 1679235063
transform 1 0 11500 0 -1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__8_.mem_right_track_4.sky130_fd_sc_hd__dfrtp_1_0__RESET_B
timestamp 1679235063
transform 1 0 13524 0 1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__8_.mem_right_track_4.sky130_fd_sc_hd__dfrtp_1_1__RESET_B
timestamp 1679235063
transform 1 0 14076 0 1 30464
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__8_.mem_right_track_4.sky130_fd_sc_hd__dfrtp_1_2__RESET_B
timestamp 1679235063
transform 1 0 14076 0 1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__8_.mem_right_track_6.sky130_fd_sc_hd__dfrtp_1_0__RESET_B
timestamp 1679235063
transform 1 0 16284 0 1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__8_.mem_right_track_6.sky130_fd_sc_hd__dfrtp_1_1__RESET_B
timestamp 1679235063
transform 1 0 14536 0 1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__8_.mem_right_track_6.sky130_fd_sc_hd__dfrtp_1_2__RESET_B
timestamp 1679235063
transform 1 0 13708 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__8_.mem_right_track_8.sky130_fd_sc_hd__dfrtp_1_0__RESET_B
timestamp 1679235063
transform 1 0 14076 0 1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__8_.mem_right_track_8.sky130_fd_sc_hd__dfrtp_1_1__RESET_B
timestamp 1679235063
transform 1 0 12420 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__8_.mem_right_track_8.sky130_fd_sc_hd__dfrtp_1_2__RESET_B
timestamp 1679235063
transform 1 0 10580 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__8_.mem_right_track_10.sky130_fd_sc_hd__dfrtp_1_0__RESET_B
timestamp 1679235063
transform 1 0 11224 0 -1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__8_.mem_right_track_10.sky130_fd_sc_hd__dfrtp_1_1__RESET_B
timestamp 1679235063
transform 1 0 10212 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__8_.mem_right_track_10.sky130_fd_sc_hd__dfrtp_1_2__RESET_B
timestamp 1679235063
transform 1 0 8372 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__8_.mem_right_track_12.sky130_fd_sc_hd__dfrtp_1_0__RESET_B
timestamp 1679235063
transform 1 0 8648 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__8_.mem_right_track_12.sky130_fd_sc_hd__dfrtp_1_1__RESET_B
timestamp 1679235063
transform 1 0 11132 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__8_.mem_right_track_14.sky130_fd_sc_hd__dfrtp_1_0__RESET_B
timestamp 1679235063
transform 1 0 13800 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__8_.mem_right_track_14.sky130_fd_sc_hd__dfrtp_1_1__RESET_B
timestamp 1679235063
transform 1 0 14628 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__8_.mem_right_track_16.sky130_fd_sc_hd__dfrtp_1_0__RESET_B
timestamp 1679235063
transform 1 0 15272 0 1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__8_.mem_right_track_16.sky130_fd_sc_hd__dfrtp_1_1__RESET_B
timestamp 1679235063
transform 1 0 14812 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__8_.mem_right_track_18.sky130_fd_sc_hd__dfrtp_1_0__RESET_B
timestamp 1679235063
transform 1 0 13800 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__8_.mem_right_track_18.sky130_fd_sc_hd__dfrtp_1_1__RESET_B
timestamp 1679235063
transform 1 0 13708 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__8_.mem_right_track_20.sky130_fd_sc_hd__dfrtp_1_0__RESET_B
timestamp 1679235063
transform 1 0 14076 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__8_.mem_right_track_20.sky130_fd_sc_hd__dfrtp_1_1__RESET_B
timestamp 1679235063
transform 1 0 11040 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__8_.mem_right_track_22.sky130_fd_sc_hd__dfrtp_1_0__RESET_B
timestamp 1679235063
transform 1 0 10580 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__8_.mem_right_track_22.sky130_fd_sc_hd__dfrtp_1_1__RESET_B
timestamp 1679235063
transform 1 0 11040 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__8_.mem_right_track_24.sky130_fd_sc_hd__dfrtp_1_0__RESET_B
timestamp 1679235063
transform 1 0 11960 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__8_.mem_right_track_24.sky130_fd_sc_hd__dfrtp_1_1__RESET_B
timestamp 1679235063
transform 1 0 12604 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__8_.mem_right_track_26.sky130_fd_sc_hd__dfrtp_1_0__RESET_B
timestamp 1679235063
transform 1 0 13800 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__8_.mem_right_track_26.sky130_fd_sc_hd__dfrtp_1_1__RESET_B
timestamp 1679235063
transform 1 0 15732 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__8_.mem_right_track_28.sky130_fd_sc_hd__dfrtp_1_0__RESET_B
timestamp 1679235063
transform 1 0 16652 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__8_.mem_right_track_28.sky130_fd_sc_hd__dfrtp_1_1__RESET_B
timestamp 1679235063
transform 1 0 16284 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__8_.mem_right_track_30.sky130_fd_sc_hd__dfrtp_1_0__RESET_B
timestamp 1679235063
transform 1 0 17756 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__8_.mem_right_track_30.sky130_fd_sc_hd__dfrtp_1_1__RESET_B
timestamp 1679235063
transform 1 0 18124 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__8_.mem_right_track_32.sky130_fd_sc_hd__dfrtp_1_0__RESET_B
timestamp 1679235063
transform 1 0 19504 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__8_.mem_right_track_32.sky130_fd_sc_hd__dfrtp_1_1__RESET_B
timestamp 1679235063
transform 1 0 18952 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__8_.mem_right_track_34.sky130_fd_sc_hd__dfrtp_1_0__RESET_B
timestamp 1679235063
transform 1 0 18032 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__8_.mem_right_track_34.sky130_fd_sc_hd__dfrtp_1_1__RESET_B
timestamp 1679235063
transform 1 0 17296 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__8_.mem_right_track_36.sky130_fd_sc_hd__dfrtp_1_0__RESET_B
timestamp 1679235063
transform 1 0 16100 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__8_.mem_right_track_36.sky130_fd_sc_hd__dfrtp_1_1__RESET_B
timestamp 1679235063
transform 1 0 15180 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__8_.mem_right_track_38.sky130_fd_sc_hd__dfrtp_1_0__RESET_B
timestamp 1679235063
transform 1 0 15272 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__8_.mem_right_track_38.sky130_fd_sc_hd__dfrtp_1_1__RESET_B
timestamp 1679235063
transform 1 0 16376 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__8_.mem_right_track_40.sky130_fd_sc_hd__dfrtp_1_0__RESET_B
timestamp 1679235063
transform 1 0 19964 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__8_.mem_right_track_40.sky130_fd_sc_hd__dfrtp_1_1__RESET_B
timestamp 1679235063
transform 1 0 19504 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__8_.mem_right_track_42.sky130_fd_sc_hd__dfrtp_1_0__RESET_B
timestamp 1679235063
transform 1 0 19964 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__8_.mem_right_track_42.sky130_fd_sc_hd__dfrtp_1_1__RESET_B
timestamp 1679235063
transform 1 0 21804 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__8_.mem_right_track_44.sky130_fd_sc_hd__dfrtp_1_0__RESET_B
timestamp 1679235063
transform 1 0 22632 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__8_.mem_right_track_44.sky130_fd_sc_hd__dfrtp_1_1__RESET_B
timestamp 1679235063
transform 1 0 21988 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__8_.mem_right_track_46.sky130_fd_sc_hd__dfrtp_1_0__RESET_B
timestamp 1679235063
transform 1 0 21804 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__8_.mem_right_track_46.sky130_fd_sc_hd__dfrtp_1_1__RESET_B
timestamp 1679235063
transform 1 0 23552 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__8_.mem_right_track_48.sky130_fd_sc_hd__dfrtp_1_0__RESET_B
timestamp 1679235063
transform 1 0 23368 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__8_.mem_right_track_48.sky130_fd_sc_hd__dfrtp_1_1__RESET_B
timestamp 1679235063
transform 1 0 25024 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__8_.mem_right_track_50.sky130_fd_sc_hd__dfrtp_1_0__RESET_B
timestamp 1679235063
transform 1 0 25024 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__8_.mem_right_track_50.sky130_fd_sc_hd__dfrtp_1_1__RESET_B
timestamp 1679235063
transform 1 0 25116 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__8_.mem_right_track_52.sky130_fd_sc_hd__dfrtp_1_0__RESET_B
timestamp 1679235063
transform 1 0 25024 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__8_.mem_right_track_52.sky130_fd_sc_hd__dfrtp_1_1__RESET_B
timestamp 1679235063
transform 1 0 24104 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__8_.mem_right_track_54.sky130_fd_sc_hd__dfrtp_1_0__RESET_B
timestamp 1679235063
transform 1 0 23828 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__8_.mem_right_track_54.sky130_fd_sc_hd__dfrtp_1_1__RESET_B
timestamp 1679235063
transform 1 0 21528 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__8_.mem_right_track_56.sky130_fd_sc_hd__dfrtp_1_0__RESET_B
timestamp 1679235063
transform 1 0 24012 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__8_.mem_right_track_56.sky130_fd_sc_hd__dfrtp_1_1__RESET_B
timestamp 1679235063
transform 1 0 21988 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__8_.mem_right_track_58.sky130_fd_sc_hd__dfrtp_1_0__RESET_B
timestamp 1679235063
transform 1 0 19228 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__8_.mem_right_track_58.sky130_fd_sc_hd__dfrtp_1_1__RESET_B
timestamp 1679235063
transform 1 0 20240 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__8_.mux_bottom_track_1.mux_l1_in_0__A0
timestamp 1679235063
transform 1 0 19228 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__8_.mux_bottom_track_1.mux_l1_in_1__A1
timestamp 1679235063
transform 1 0 18308 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__8_.mux_bottom_track_3.mux_l1_in_0__A0
timestamp 1679235063
transform 1 0 25392 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__8_.mux_bottom_track_5.mux_l1_in_0__A0
timestamp 1679235063
transform 1 0 24104 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__8_.mux_bottom_track_7.mux_l1_in_0__A0
timestamp 1679235063
transform 1 0 23184 0 -1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__8_.mux_bottom_track_7.mux_l1_in_1__A1
timestamp 1679235063
transform 1 0 18860 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__8_.mux_bottom_track_9.mux_l1_in_0__A0
timestamp 1679235063
transform 1 0 23920 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__8_.mux_bottom_track_11.mux_l1_in_0__A0
timestamp 1679235063
transform 1 0 25392 0 -1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__8_.mux_bottom_track_13.mux_l1_in_0__A0
timestamp 1679235063
transform 1 0 24564 0 1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__8_.mux_bottom_track_15.mux_l1_in_0__A0
timestamp 1679235063
transform 1 0 23000 0 -1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__8_.mux_bottom_track_17.mux_l1_in_0__A0
timestamp 1679235063
transform 1 0 20332 0 -1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__8_.mux_bottom_track_19.mux_l1_in_0__A0
timestamp 1679235063
transform 1 0 20424 0 -1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__8_.mux_bottom_track_29.mux_l1_in_0__A0
timestamp 1679235063
transform 1 0 20332 0 1 30464
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__8_.mux_bottom_track_31.mux_l1_in_0__A0
timestamp 1679235063
transform 1 0 21436 0 -1 31552
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__8_.mux_bottom_track_33.mux_l1_in_0__A0
timestamp 1679235063
transform 1 0 24748 0 1 34816
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__8_.mux_bottom_track_35.mux_l1_in_0__A0
timestamp 1679235063
transform 1 0 24012 0 1 33728
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__8_.mux_bottom_track_45.mux_l1_in_0__A0
timestamp 1679235063
transform 1 0 22356 0 1 34816
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__8_.mux_bottom_track_47.mux_l1_in_0__A0
timestamp 1679235063
transform 1 0 21804 0 1 34816
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__8_.mux_bottom_track_49.mux_l1_in_0__A0
timestamp 1679235063
transform 1 0 20332 0 -1 35904
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__8_.mux_bottom_track_51.mux_l1_in_0__A0
timestamp 1679235063
transform 1 0 21528 0 -1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__8_.mux_bottom_track_51.mux_l1_in_0__A1
timestamp 1679235063
transform 1 0 24748 0 -1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__8_.mux_bottom_track_51.mux_l2_in_0__S
timestamp 1679235063
transform 1 0 20332 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__8_.mux_right_track_0.mux_l1_in_0__A0
timestamp 1679235063
transform 1 0 17020 0 -1 32640
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__8_.mux_right_track_0.mux_l1_in_0__A1
timestamp 1679235063
transform 1 0 16836 0 -1 32640
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__8_.mux_right_track_0.mux_l1_in_1__A0
timestamp 1679235063
transform 1 0 16652 0 -1 32640
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__8_.mux_right_track_0.mux_l1_in_1__A1
timestamp 1679235063
transform 1 0 16652 0 -1 31552
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__8_.mux_right_track_0.mux_l2_in_0__S
timestamp 1679235063
transform 1 0 13800 0 1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__8_.mux_right_track_0.mux_l2_in_1__A1
timestamp 1679235063
transform 1 0 7268 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__8_.mux_right_track_0.mux_l2_in_1__S
timestamp 1679235063
transform 1 0 8924 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__8_.mux_right_track_2.mux_l1_in_0__A0
timestamp 1679235063
transform 1 0 16376 0 -1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__8_.mux_right_track_2.mux_l1_in_0__A1
timestamp 1679235063
transform 1 0 16468 0 1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__8_.mux_right_track_2.mux_l1_in_1__A0
timestamp 1679235063
transform 1 0 16928 0 1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__8_.mux_right_track_2.mux_l1_in_1__A1
timestamp 1679235063
transform 1 0 16744 0 1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__8_.mux_right_track_2.mux_l2_in_1__A1
timestamp 1679235063
transform 1 0 9292 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__8_.mux_right_track_4.mux_l1_in_0__A0
timestamp 1679235063
transform 1 0 16376 0 -1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__8_.mux_right_track_4.mux_l1_in_0__A1
timestamp 1679235063
transform 1 0 16468 0 1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__8_.mux_right_track_4.mux_l1_in_1__A0
timestamp 1679235063
transform 1 0 16836 0 -1 30464
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__8_.mux_right_track_4.mux_l1_in_1__A1
timestamp 1679235063
transform 1 0 16652 0 -1 30464
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__8_.mux_right_track_4.mux_l2_in_1__A1
timestamp 1679235063
transform 1 0 12788 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__8_.mux_right_track_6.mux_l1_in_0__A0
timestamp 1679235063
transform 1 0 18032 0 -1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__8_.mux_right_track_6.mux_l1_in_0__A1
timestamp 1679235063
transform 1 0 17848 0 -1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__8_.mux_right_track_6.mux_l1_in_1__A0
timestamp 1679235063
transform 1 0 17480 0 1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__8_.mux_right_track_6.mux_l1_in_1__A1
timestamp 1679235063
transform 1 0 17664 0 1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__8_.mux_right_track_6.mux_l2_in_1__A1
timestamp 1679235063
transform 1 0 11500 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__8_.mux_right_track_8.mux_l1_in_0__A0
timestamp 1679235063
transform 1 0 16008 0 -1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__8_.mux_right_track_8.mux_l1_in_0__A1
timestamp 1679235063
transform 1 0 16192 0 -1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__8_.mux_right_track_8.mux_l1_in_1__A0
timestamp 1679235063
transform 1 0 17296 0 1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__8_.mux_right_track_8.mux_l1_in_1__A1
timestamp 1679235063
transform 1 0 17112 0 1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__8_.mux_right_track_8.mux_l2_in_1__A1
timestamp 1679235063
transform 1 0 8740 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__8_.mux_right_track_10.mux_l1_in_0__A0
timestamp 1679235063
transform 1 0 15272 0 1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__8_.mux_right_track_10.mux_l1_in_0__A1
timestamp 1679235063
transform 1 0 15180 0 -1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__8_.mux_right_track_10.mux_l1_in_1__A0
timestamp 1679235063
transform 1 0 16376 0 -1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__8_.mux_right_track_10.mux_l1_in_1__A1
timestamp 1679235063
transform 1 0 16192 0 -1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__8_.mux_right_track_12.mux_l1_in_0__A0
timestamp 1679235063
transform 1 0 14260 0 1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__8_.mux_right_track_12.mux_l1_in_0__A1
timestamp 1679235063
transform 1 0 14076 0 1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__8_.mux_right_track_14.mux_l1_in_0__A0
timestamp 1679235063
transform 1 0 16376 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__8_.mux_right_track_14.mux_l1_in_0__A1
timestamp 1679235063
transform 1 0 16008 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__8_.mux_right_track_14.mux_l1_in_1__A1
timestamp 1679235063
transform 1 0 13616 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__8_.mux_right_track_16.mux_l1_in_0__A0
timestamp 1679235063
transform 1 0 19044 0 -1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__8_.mux_right_track_16.mux_l1_in_0__A1
timestamp 1679235063
transform 1 0 18860 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__8_.mux_right_track_16.mux_l1_in_1__A1
timestamp 1679235063
transform 1 0 13892 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__8_.mux_right_track_18.mux_l1_in_0__A0
timestamp 1679235063
transform 1 0 12604 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__8_.mux_right_track_18.mux_l1_in_0__A1
timestamp 1679235063
transform 1 0 14720 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__8_.mux_right_track_20.mux_l1_in_0__A0
timestamp 1679235063
transform 1 0 10304 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__8_.mux_right_track_20.mux_l1_in_0__A1
timestamp 1679235063
transform 1 0 12144 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__8_.mux_right_track_22.mux_l1_in_0__A1
timestamp 1679235063
transform 1 0 11408 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__8_.mux_right_track_24.mux_l1_in_0__A1
timestamp 1679235063
transform 1 0 12696 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__8_.mux_right_track_26.mux_l1_in_0__A1
timestamp 1679235063
transform 1 0 16652 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__8_.mux_right_track_28.mux_l1_in_0__A0
timestamp 1679235063
transform 1 0 18492 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__8_.mux_right_track_28.mux_l1_in_0__A1
timestamp 1679235063
transform 1 0 18676 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__8_.mux_right_track_28.mux_l1_in_1__A1
timestamp 1679235063
transform 1 0 13248 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__8_.mux_right_track_30.mux_l1_in_0__A0
timestamp 1679235063
transform 1 0 19228 0 -1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__8_.mux_right_track_30.mux_l1_in_0__A1
timestamp 1679235063
transform 1 0 18676 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__8_.mux_right_track_30.mux_l1_in_1__A1
timestamp 1679235063
transform 1 0 14904 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__8_.mux_right_track_32.mux_l1_in_0__A0
timestamp 1679235063
transform 1 0 18492 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__8_.mux_right_track_32.mux_l1_in_0__A1
timestamp 1679235063
transform 1 0 18308 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__8_.mux_right_track_32.mux_l1_in_1__A1
timestamp 1679235063
transform 1 0 15732 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__8_.mux_right_track_34.mux_l1_in_0__A0
timestamp 1679235063
transform 1 0 18952 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__8_.mux_right_track_34.mux_l1_in_0__A1
timestamp 1679235063
transform 1 0 19044 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__8_.mux_right_track_36.mux_l1_in_0__A1
timestamp 1679235063
transform 1 0 12604 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__8_.mux_right_track_38.mux_l1_in_0__A1
timestamp 1679235063
transform 1 0 16284 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__8_.mux_right_track_40.mux_l1_in_0__A1
timestamp 1679235063
transform 1 0 17848 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__8_.mux_right_track_42.mux_l1_in_0__A1
timestamp 1679235063
transform 1 0 18768 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__8_.mux_right_track_44.mux_l1_in_0__A0
timestamp 1679235063
transform 1 0 19688 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__8_.mux_right_track_44.mux_l1_in_0__A1
timestamp 1679235063
transform 1 0 21988 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__8_.mux_right_track_44.mux_l1_in_1__A1
timestamp 1679235063
transform 1 0 19044 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__8_.mux_right_track_46.mux_l1_in_0__A0
timestamp 1679235063
transform 1 0 21620 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__8_.mux_right_track_46.mux_l1_in_0__A1
timestamp 1679235063
transform 1 0 18124 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__8_.mux_right_track_46.mux_l1_in_1__A1
timestamp 1679235063
transform 1 0 18124 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__8_.mux_right_track_48.mux_l1_in_0__A0
timestamp 1679235063
transform 1 0 21804 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__8_.mux_right_track_48.mux_l1_in_0__A1
timestamp 1679235063
transform 1 0 21804 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__8_.mux_right_track_48.mux_l1_in_1__A1
timestamp 1679235063
transform 1 0 18952 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__8_.mux_right_track_48.sky130_fd_sc_hd__buf_4_0__A
timestamp 1679235063
transform 1 0 8924 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__8_.mux_right_track_50.mux_l1_in_0__A0
timestamp 1679235063
transform 1 0 20608 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__8_.mux_right_track_50.mux_l1_in_0__A1
timestamp 1679235063
transform 1 0 22448 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__8_.mux_right_track_50.mux_l2_in_0__A0
timestamp 1679235063
transform 1 0 22356 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__8_.mux_right_track_52.mux_l1_in_0__A1
timestamp 1679235063
transform 1 0 21804 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__8_.mux_right_track_52.mux_l2_in_0__A0
timestamp 1679235063
transform 1 0 24104 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__8_.mux_right_track_54.mux_l1_in_0__A1
timestamp 1679235063
transform 1 0 19320 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__8_.mux_right_track_56.mux_l1_in_0__A1
timestamp 1679235063
transform 1 0 18584 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__8_.mux_right_track_58.mux_l1_in_0__A0
timestamp 1679235063
transform 1 0 19688 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__8_.mux_right_track_58.mux_l1_in_0__A1
timestamp 1679235063
transform 1 0 18860 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__dfrtp_4  cby_0__8_.cby_0__1_.mem_right_ipin_0.sky130_fd_sc_hd__dfrtp_1_0_ pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1679235063
transform 1 0 5060 0 1 4352
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_2  cby_0__8_.cby_0__1_.mem_right_ipin_0.sky130_fd_sc_hd__dfrtp_1_1_ pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1679235063
transform 1 0 8188 0 -1 9792
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_1  cby_0__8_.cby_0__1_.mem_right_ipin_0.sky130_fd_sc_hd__dfrtp_1_2_ pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1679235063
transform 1 0 6532 0 -1 14144
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  cby_0__8_.cby_0__1_.mem_right_ipin_0.sky130_fd_sc_hd__dfrtp_1_3_
timestamp 1679235063
transform 1 0 5888 0 1 16320
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_4  cby_0__8_.cby_0__1_.mem_right_ipin_1.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1679235063
transform 1 0 7544 0 -1 16320
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_2  cby_0__8_.cby_0__1_.mem_right_ipin_1.sky130_fd_sc_hd__dfrtp_1_1_
timestamp 1679235063
transform 1 0 9200 0 -1 10880
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_1  cby_0__8_.cby_0__1_.mem_right_ipin_1.sky130_fd_sc_hd__dfrtp_1_2_
timestamp 1679235063
transform 1 0 7176 0 -1 13056
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  cby_0__8_.cby_0__1_.mem_right_ipin_1.sky130_fd_sc_hd__dfrtp_1_3_
timestamp 1679235063
transform 1 0 6348 0 1 15232
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_4  cby_0__8_.cby_0__1_.mem_right_ipin_2.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1679235063
transform 1 0 7728 0 -1 15232
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_4  cby_0__8_.cby_0__1_.mem_right_ipin_2.sky130_fd_sc_hd__dfrtp_1_1_
timestamp 1679235063
transform 1 0 9936 0 1 15232
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_1  cby_0__8_.cby_0__1_.mem_right_ipin_2.sky130_fd_sc_hd__dfrtp_1_2_
timestamp 1679235063
transform 1 0 7452 0 -1 19584
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  cby_0__8_.cby_0__1_.mem_right_ipin_2.sky130_fd_sc_hd__dfrtp_1_3_
timestamp 1679235063
transform 1 0 6808 0 1 21760
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_4  cby_0__8_.cby_0__1_.mem_right_ipin_3.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1679235063
transform 1 0 7544 0 -1 21760
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_4  cby_0__8_.cby_0__1_.mem_right_ipin_3.sky130_fd_sc_hd__dfrtp_1_1_
timestamp 1679235063
transform 1 0 9108 0 -1 18496
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_1  cby_0__8_.cby_0__1_.mem_right_ipin_3.sky130_fd_sc_hd__dfrtp_1_2_
timestamp 1679235063
transform 1 0 6808 0 1 23936
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  cby_0__8_.cby_0__1_.mem_right_ipin_3.sky130_fd_sc_hd__dfrtp_1_3_
timestamp 1679235063
transform 1 0 9108 0 1 29376
box -38 -48 1878 592
use sky130_fd_sc_hd__mux2_1  cby_0__8_.cby_0__1_.mux_right_ipin_0.mux_l1_in_0_ pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1679235063
transform 1 0 15640 0 1 9792
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  cby_0__8_.cby_0__1_.mux_right_ipin_0.mux_l1_in_1_
timestamp 1679235063
transform 1 0 13892 0 -1 10880
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  cby_0__8_.cby_0__1_.mux_right_ipin_0.mux_l1_in_2_
timestamp 1679235063
transform 1 0 14444 0 1 9792
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  cby_0__8_.cby_0__1_.mux_right_ipin_0.mux_l1_in_3_
timestamp 1679235063
transform 1 0 14996 0 1 14144
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  cby_0__8_.cby_0__1_.mux_right_ipin_0.mux_l1_in_4_
timestamp 1679235063
transform 1 0 12604 0 -1 13056
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  cby_0__8_.cby_0__1_.mux_right_ipin_0.mux_l2_in_0_
timestamp 1679235063
transform 1 0 11408 0 1 11968
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  cby_0__8_.cby_0__1_.mux_right_ipin_0.mux_l2_in_1_
timestamp 1679235063
transform 1 0 11960 0 -1 11968
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  cby_0__8_.cby_0__1_.mux_right_ipin_0.mux_l2_in_2_
timestamp 1679235063
transform 1 0 8924 0 -1 11968
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  cby_0__8_.cby_0__1_.mux_right_ipin_0.mux_l2_in_3__186 pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1679235063
transform 1 0 11684 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  cby_0__8_.cby_0__1_.mux_right_ipin_0.mux_l2_in_3_
timestamp 1679235063
transform 1 0 10396 0 -1 14144
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  cby_0__8_.cby_0__1_.mux_right_ipin_0.mux_l3_in_0_
timestamp 1679235063
transform 1 0 10212 0 -1 15232
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  cby_0__8_.cby_0__1_.mux_right_ipin_0.mux_l3_in_1_
timestamp 1679235063
transform 1 0 9108 0 1 14144
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  cby_0__8_.cby_0__1_.mux_right_ipin_0.mux_l4_in_0_
timestamp 1679235063
transform 1 0 8004 0 -1 20672
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  cby_0__8_.cby_0__1_.mux_right_ipin_0.sky130_fd_sc_hd__buf_4_0_
timestamp 1679235063
transform 1 0 9108 0 1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  cby_0__8_.cby_0__1_.mux_right_ipin_1.mux_l1_in_0_
timestamp 1679235063
transform 1 0 15548 0 -1 8704
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  cby_0__8_.cby_0__1_.mux_right_ipin_1.mux_l1_in_1_
timestamp 1679235063
transform 1 0 15548 0 1 8704
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  cby_0__8_.cby_0__1_.mux_right_ipin_1.mux_l1_in_2_
timestamp 1679235063
transform 1 0 14628 0 -1 9792
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  cby_0__8_.cby_0__1_.mux_right_ipin_1.mux_l1_in_3_
timestamp 1679235063
transform 1 0 15180 0 1 13056
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  cby_0__8_.cby_0__1_.mux_right_ipin_1.mux_l1_in_4_
timestamp 1679235063
transform 1 0 12972 0 1 14144
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  cby_0__8_.cby_0__1_.mux_right_ipin_1.mux_l2_in_0_
timestamp 1679235063
transform 1 0 12972 0 1 8704
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  cby_0__8_.cby_0__1_.mux_right_ipin_1.mux_l2_in_1_
timestamp 1679235063
transform 1 0 12604 0 1 10880
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  cby_0__8_.cby_0__1_.mux_right_ipin_1.mux_l2_in_2_
timestamp 1679235063
transform 1 0 9752 0 1 11968
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  cby_0__8_.cby_0__1_.mux_right_ipin_1.mux_l2_in_3_
timestamp 1679235063
transform 1 0 10120 0 -1 11968
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  cby_0__8_.cby_0__1_.mux_right_ipin_1.mux_l2_in_3__187
timestamp 1679235063
transform 1 0 11684 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  cby_0__8_.cby_0__1_.mux_right_ipin_1.mux_l3_in_0_
timestamp 1679235063
transform 1 0 10304 0 -1 13056
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  cby_0__8_.cby_0__1_.mux_right_ipin_1.mux_l3_in_1_
timestamp 1679235063
transform 1 0 9108 0 -1 14144
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  cby_0__8_.cby_0__1_.mux_right_ipin_1.mux_l4_in_0_
timestamp 1679235063
transform 1 0 7912 0 -1 18496
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  cby_0__8_.cby_0__1_.mux_right_ipin_1.sky130_fd_sc_hd__buf_4_0_
timestamp 1679235063
transform 1 0 8924 0 -1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  cby_0__8_.cby_0__1_.mux_right_ipin_2.mux_l1_in_0_
timestamp 1679235063
transform 1 0 16836 0 1 9792
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  cby_0__8_.cby_0__1_.mux_right_ipin_2.mux_l1_in_1_
timestamp 1679235063
transform 1 0 15456 0 -1 10880
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  cby_0__8_.cby_0__1_.mux_right_ipin_2.mux_l1_in_2_
timestamp 1679235063
transform 1 0 12696 0 1 9792
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  cby_0__8_.cby_0__1_.mux_right_ipin_2.mux_l1_in_3_
timestamp 1679235063
transform 1 0 12512 0 -1 10880
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  cby_0__8_.cby_0__1_.mux_right_ipin_2.mux_l1_in_4_
timestamp 1679235063
transform 1 0 12972 0 1 16320
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  cby_0__8_.cby_0__1_.mux_right_ipin_2.mux_l2_in_0_
timestamp 1679235063
transform 1 0 12328 0 -1 14144
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  cby_0__8_.cby_0__1_.mux_right_ipin_2.mux_l2_in_1_
timestamp 1679235063
transform 1 0 11684 0 1 14144
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  cby_0__8_.cby_0__1_.mux_right_ipin_2.mux_l2_in_2_
timestamp 1679235063
transform 1 0 10212 0 1 16320
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  cby_0__8_.cby_0__1_.mux_right_ipin_2.mux_l2_in_3__188
timestamp 1679235063
transform 1 0 15824 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  cby_0__8_.cby_0__1_.mux_right_ipin_2.mux_l2_in_3_
timestamp 1679235063
transform 1 0 14628 0 -1 23936
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  cby_0__8_.cby_0__1_.mux_right_ipin_2.mux_l3_in_0_
timestamp 1679235063
transform 1 0 10304 0 -1 17408
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  cby_0__8_.cby_0__1_.mux_right_ipin_2.mux_l3_in_1_
timestamp 1679235063
transform 1 0 10304 0 -1 21760
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  cby_0__8_.cby_0__1_.mux_right_ipin_2.mux_l4_in_0_
timestamp 1679235063
transform 1 0 8004 0 -1 25024
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  cby_0__8_.cby_0__1_.mux_right_ipin_2.sky130_fd_sc_hd__buf_4_0_
timestamp 1679235063
transform 1 0 9108 0 1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  cby_0__8_.cby_0__1_.mux_right_ipin_3.mux_l1_in_0_
timestamp 1679235063
transform 1 0 14352 0 -1 11968
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  cby_0__8_.cby_0__1_.mux_right_ipin_3.mux_l1_in_1_
timestamp 1679235063
transform 1 0 14352 0 1 11968
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  cby_0__8_.cby_0__1_.mux_right_ipin_3.mux_l1_in_2_
timestamp 1679235063
transform 1 0 13156 0 -1 11968
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  cby_0__8_.cby_0__1_.mux_right_ipin_3.mux_l1_in_3_
timestamp 1679235063
transform 1 0 12604 0 1 11968
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  cby_0__8_.cby_0__1_.mux_right_ipin_3.mux_l1_in_4_
timestamp 1679235063
transform 1 0 13156 0 -1 18496
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  cby_0__8_.cby_0__1_.mux_right_ipin_3.mux_l2_in_0_
timestamp 1679235063
transform 1 0 11776 0 1 16320
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  cby_0__8_.cby_0__1_.mux_right_ipin_3.mux_l2_in_1_
timestamp 1679235063
transform 1 0 11684 0 -1 17408
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  cby_0__8_.cby_0__1_.mux_right_ipin_3.mux_l2_in_2_
timestamp 1679235063
transform 1 0 10120 0 -1 19584
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  cby_0__8_.cby_0__1_.mux_right_ipin_3.mux_l2_in_3_
timestamp 1679235063
transform 1 0 15640 0 1 26112
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  cby_0__8_.cby_0__1_.mux_right_ipin_3.mux_l2_in_3__189
timestamp 1679235063
transform 1 0 15732 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  cby_0__8_.cby_0__1_.mux_right_ipin_3.mux_l3_in_0_
timestamp 1679235063
transform 1 0 10120 0 1 21760
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  cby_0__8_.cby_0__1_.mux_right_ipin_3.mux_l3_in_1_
timestamp 1679235063
transform 1 0 10304 0 1 25024
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  cby_0__8_.cby_0__1_.mux_right_ipin_3.mux_l4_in_0_
timestamp 1679235063
transform 1 0 9660 0 -1 30464
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  cby_0__8_.cby_0__1_.mux_right_ipin_3.sky130_fd_sc_hd__buf_4_0_
timestamp 1679235063
transform 1 0 9108 0 1 39168
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_8  cby_0__8_.grid_io_left_left_0__1_.logical_tile_io_mode_io__0.logical_tile_io_mode_physical__iopad_0.io_0_.IN_PROTECT_GATE pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1679235063
transform 1 0 15640 0 1 45696
box -38 -48 1970 592
use sky130_fd_sc_hd__inv_1  cby_0__8_.grid_io_left_left_0__1_.logical_tile_io_mode_io__0.logical_tile_io_mode_physical__iopad_0.io_0_.INV_SOC_DIR pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1679235063
transform 1 0 13340 0 1 46784
box -38 -48 314 592
use sky130_fd_sc_hd__or2b_2  cby_0__8_.grid_io_left_left_0__1_.logical_tile_io_mode_io__0.logical_tile_io_mode_physical__iopad_0.io_0_.ISOL_EN_GATE pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1679235063
transform 1 0 11040 0 1 44608
box -38 -48 682 592
use sky130_fd_sc_hd__ebufn_8  cby_0__8_.grid_io_left_left_0__1_.logical_tile_io_mode_io__0.logical_tile_io_mode_physical__iopad_0.io_0_.OUT_PROTECT_GATE
timestamp 1679235063
transform 1 0 10396 0 1 45696
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_1  cby_0__8_.grid_io_left_left_0__1_.logical_tile_io_mode_io__0.logical_tile_io_mode_physical__iopad_0.io_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1679235063
transform 1 0 9384 0 -1 36992
box -38 -48 1878 592
use sky130_fd_sc_hd__ebufn_8  cby_0__8_.grid_io_left_left_0__1_.logical_tile_io_mode_io__1.logical_tile_io_mode_physical__iopad_0.io_0_.IN_PROTECT_GATE
timestamp 1679235063
transform 1 0 14444 0 -1 46784
box -38 -48 1970 592
use sky130_fd_sc_hd__inv_1  cby_0__8_.grid_io_left_left_0__1_.logical_tile_io_mode_io__1.logical_tile_io_mode_physical__iopad_0.io_0_.INV_SOC_DIR
timestamp 1679235063
transform 1 0 12512 0 1 46784
box -38 -48 314 592
use sky130_fd_sc_hd__or2b_2  cby_0__8_.grid_io_left_left_0__1_.logical_tile_io_mode_io__1.logical_tile_io_mode_physical__iopad_0.io_0_.ISOL_EN_GATE
timestamp 1679235063
transform 1 0 10304 0 1 46784
box -38 -48 682 592
use sky130_fd_sc_hd__ebufn_8  cby_0__8_.grid_io_left_left_0__1_.logical_tile_io_mode_io__1.logical_tile_io_mode_physical__iopad_0.io_0_.OUT_PROTECT_GATE
timestamp 1679235063
transform 1 0 9292 0 -1 45696
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_1  cby_0__8_.grid_io_left_left_0__1_.logical_tile_io_mode_io__1.logical_tile_io_mode_physical__iopad_0.io_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1679235063
transform 1 0 9384 0 -1 43520
box -38 -48 1878 592
use sky130_fd_sc_hd__ebufn_8  cby_0__8_.grid_io_left_left_0__1_.logical_tile_io_mode_io__2.logical_tile_io_mode_physical__iopad_0.io_0_.IN_PROTECT_GATE
timestamp 1679235063
transform 1 0 14260 0 1 46784
box -38 -48 1970 592
use sky130_fd_sc_hd__inv_1  cby_0__8_.grid_io_left_left_0__1_.logical_tile_io_mode_io__2.logical_tile_io_mode_physical__iopad_0.io_0_.INV_SOC_DIR
timestamp 1679235063
transform 1 0 11500 0 1 47872
box -38 -48 314 592
use sky130_fd_sc_hd__or2b_2  cby_0__8_.grid_io_left_left_0__1_.logical_tile_io_mode_io__2.logical_tile_io_mode_physical__iopad_0.io_0_.ISOL_EN_GATE
timestamp 1679235063
transform 1 0 9292 0 1 48960
box -38 -48 682 592
use sky130_fd_sc_hd__ebufn_8  cby_0__8_.grid_io_left_left_0__1_.logical_tile_io_mode_io__2.logical_tile_io_mode_physical__iopad_0.io_0_.OUT_PROTECT_GATE
timestamp 1679235063
transform 1 0 8648 0 -1 47872
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_1  cby_0__8_.grid_io_left_left_0__1_.logical_tile_io_mode_io__2.logical_tile_io_mode_physical__iopad_0.io_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1679235063
transform 1 0 8832 0 -1 46784
box -38 -48 1878 592
use sky130_fd_sc_hd__ebufn_8  cby_0__8_.grid_io_left_left_0__1_.logical_tile_io_mode_io__3.logical_tile_io_mode_physical__iopad_0.io_0_.IN_PROTECT_GATE
timestamp 1679235063
transform 1 0 12604 0 -1 47872
box -38 -48 1970 592
use sky130_fd_sc_hd__inv_1  cby_0__8_.grid_io_left_left_0__1_.logical_tile_io_mode_io__3.logical_tile_io_mode_physical__iopad_0.io_0_.INV_SOC_DIR
timestamp 1679235063
transform 1 0 10212 0 -1 48960
box -38 -48 314 592
use sky130_fd_sc_hd__or2b_2  cby_0__8_.grid_io_left_left_0__1_.logical_tile_io_mode_io__3.logical_tile_io_mode_physical__iopad_0.io_0_.ISOL_EN_GATE
timestamp 1679235063
transform 1 0 7544 0 1 51136
box -38 -48 682 592
use sky130_fd_sc_hd__ebufn_8  cby_0__8_.grid_io_left_left_0__1_.logical_tile_io_mode_io__3.logical_tile_io_mode_physical__iopad_0.io_0_.OUT_PROTECT_GATE
timestamp 1679235063
transform 1 0 7728 0 -1 48960
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_1  cby_0__8_.grid_io_left_left_0__1_.logical_tile_io_mode_io__3.logical_tile_io_mode_physical__iopad_0.io_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1679235063
transform 1 0 6624 0 1 48960
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_0_prog_clk pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1679235063
transform 1 0 15640 0 1 25024
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_8  clkbuf_4_0_0_prog_clk pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1679235063
transform 1 0 10304 0 1 14144
box -38 -48 1050 592
use sky130_fd_sc_hd__clkbuf_8  clkbuf_4_1_0_prog_clk
timestamp 1679235063
transform 1 0 11960 0 1 13056
box -38 -48 1050 592
use sky130_fd_sc_hd__clkbuf_8  clkbuf_4_2_0_prog_clk
timestamp 1679235063
transform 1 0 10212 0 1 17408
box -38 -48 1050 592
use sky130_fd_sc_hd__clkbuf_8  clkbuf_4_3_0_prog_clk
timestamp 1679235063
transform 1 0 12144 0 1 18496
box -38 -48 1050 592
use sky130_fd_sc_hd__clkbuf_8  clkbuf_4_4_0_prog_clk
timestamp 1679235063
transform 1 0 17204 0 -1 13056
box -38 -48 1050 592
use sky130_fd_sc_hd__clkbuf_8  clkbuf_4_5_0_prog_clk
timestamp 1679235063
transform 1 0 19044 0 -1 14144
box -38 -48 1050 592
use sky130_fd_sc_hd__clkbuf_8  clkbuf_4_6_0_prog_clk
timestamp 1679235063
transform 1 0 17296 0 -1 17408
box -38 -48 1050 592
use sky130_fd_sc_hd__clkbuf_8  clkbuf_4_7_0_prog_clk
timestamp 1679235063
transform 1 0 19412 0 1 16320
box -38 -48 1050 592
use sky130_fd_sc_hd__clkbuf_8  clkbuf_4_8_0_prog_clk
timestamp 1679235063
transform 1 0 14260 0 1 31552
box -38 -48 1050 592
use sky130_fd_sc_hd__clkbuf_8  clkbuf_4_9_0_prog_clk
timestamp 1679235063
transform 1 0 14444 0 1 30464
box -38 -48 1050 592
use sky130_fd_sc_hd__clkbuf_8  clkbuf_4_10_0_prog_clk
timestamp 1679235063
transform 1 0 15088 0 -1 34816
box -38 -48 1050 592
use sky130_fd_sc_hd__clkbuf_8  clkbuf_4_11_0_prog_clk
timestamp 1679235063
transform 1 0 17204 0 1 33728
box -38 -48 1050 592
use sky130_fd_sc_hd__clkbuf_8  clkbuf_4_12_0_prog_clk
timestamp 1679235063
transform 1 0 20516 0 -1 28288
box -38 -48 1050 592
use sky130_fd_sc_hd__clkbuf_8  clkbuf_4_13_0_prog_clk
timestamp 1679235063
transform 1 0 22816 0 1 28288
box -38 -48 1050 592
use sky130_fd_sc_hd__clkbuf_8  clkbuf_4_14_0_prog_clk
timestamp 1679235063
transform 1 0 20056 0 -1 32640
box -38 -48 1050 592
use sky130_fd_sc_hd__clkbuf_8  clkbuf_4_15_0_prog_clk
timestamp 1679235063
transform 1 0 22080 0 -1 32640
box -38 -48 1050 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3 pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1679235063
transform 1 0 1380 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_15 pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1679235063
transform 1 0 2484 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_26 pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1679235063
transform 1 0 3496 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_35
timestamp 1679235063
transform 1 0 4324 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_40 pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1679235063
transform 1 0 4784 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_54
timestamp 1679235063
transform 1 0 6072 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_63
timestamp 1679235063
transform 1 0 6900 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_68
timestamp 1679235063
transform 1 0 7360 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_75
timestamp 1679235063
transform 1 0 8004 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_82
timestamp 1679235063
transform 1 0 8648 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_91
timestamp 1679235063
transform 1 0 9476 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_96
timestamp 1679235063
transform 1 0 9936 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_110
timestamp 1679235063
transform 1 0 11224 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_113
timestamp 1679235063
transform 1 0 11500 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_118
timestamp 1679235063
transform 1 0 11960 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_138
timestamp 1679235063
transform 1 0 13800 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_143
timestamp 1679235063
transform 1 0 14260 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_161
timestamp 1679235063
transform 1 0 15916 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_165 pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1679235063
transform 1 0 16284 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_169
timestamp 1679235063
transform 1 0 16652 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_187
timestamp 1679235063
transform 1 0 18308 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_194
timestamp 1679235063
transform 1 0 18952 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_197
timestamp 1679235063
transform 1 0 19228 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_215
timestamp 1679235063
transform 1 0 20884 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_222
timestamp 1679235063
transform 1 0 21528 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_225
timestamp 1679235063
transform 1 0 21804 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_243
timestamp 1679235063
transform 1 0 23460 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_250
timestamp 1679235063
transform 1 0 24104 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_253
timestamp 1679235063
transform 1 0 24380 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_259
timestamp 1679235063
transform 1 0 24932 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_263
timestamp 1679235063
transform 1 0 25300 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_1_3 pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1679235063
transform 1 0 1380 0 -1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_1_21
timestamp 1679235063
transform 1 0 3036 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_1_35
timestamp 1679235063
transform 1 0 4324 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_1_41
timestamp 1679235063
transform 1 0 4876 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_1_54
timestamp 1679235063
transform 1 0 6072 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_1_57
timestamp 1679235063
transform 1 0 6348 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_1_62
timestamp 1679235063
transform 1 0 6808 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_69
timestamp 1679235063
transform 1 0 7452 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_1_83
timestamp 1679235063
transform 1 0 8740 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_1_91
timestamp 1679235063
transform 1 0 9476 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_1_96
timestamp 1679235063
transform 1 0 9936 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_103
timestamp 1679235063
transform 1 0 10580 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_1_110
timestamp 1679235063
transform 1 0 11224 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_1_113
timestamp 1679235063
transform 1 0 11500 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_1_125
timestamp 1679235063
transform 1 0 12604 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_145
timestamp 1679235063
transform 1 0 14444 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_1_165
timestamp 1679235063
transform 1 0 16284 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_1_169
timestamp 1679235063
transform 1 0 16652 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_1_187
timestamp 1679235063
transform 1 0 18308 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_207
timestamp 1679235063
transform 1 0 20148 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_215
timestamp 1679235063
transform 1 0 20884 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_1_222
timestamp 1679235063
transform 1 0 21528 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_1_225
timestamp 1679235063
transform 1 0 21804 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_1_231
timestamp 1679235063
transform 1 0 22356 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_239
timestamp 1679235063
transform 1 0 23092 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_1_243
timestamp 1679235063
transform 1 0 23460 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_1_264
timestamp 1679235063
transform 1 0 25392 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_2_3
timestamp 1679235063
transform 1 0 1380 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_2_15
timestamp 1679235063
transform 1 0 2484 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_2_22
timestamp 1679235063
transform 1 0 3128 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_2_29
timestamp 1679235063
transform 1 0 3772 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_2_33
timestamp 1679235063
transform 1 0 4140 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_2_37
timestamp 1679235063
transform 1 0 4508 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_2_51
timestamp 1679235063
transform 1 0 5796 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_2_55
timestamp 1679235063
transform 1 0 6164 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_2_60
timestamp 1679235063
transform 1 0 6624 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_2_64
timestamp 1679235063
transform 1 0 6992 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_2_68
timestamp 1679235063
transform 1 0 7360 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_2_77
timestamp 1679235063
transform 1 0 8188 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_2_82
timestamp 1679235063
transform 1 0 8648 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_2_85
timestamp 1679235063
transform 1 0 8924 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_2_90
timestamp 1679235063
transform 1 0 9384 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_2_97
timestamp 1679235063
transform 1 0 10028 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_2_104
timestamp 1679235063
transform 1 0 10672 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_2_118
timestamp 1679235063
transform 1 0 11960 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_2_138
timestamp 1679235063
transform 1 0 13800 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_2_141
timestamp 1679235063
transform 1 0 14076 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_2_159
timestamp 1679235063
transform 1 0 15732 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_2_179
timestamp 1679235063
transform 1 0 17572 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_2_191
timestamp 1679235063
transform 1 0 18676 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_2_195
timestamp 1679235063
transform 1 0 19044 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_2_197
timestamp 1679235063
transform 1 0 19228 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_2_215
timestamp 1679235063
transform 1 0 20884 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_2_235 pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1679235063
transform 1 0 22724 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_2_247
timestamp 1679235063
transform 1 0 23828 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_2_251
timestamp 1679235063
transform 1 0 24196 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_2_253
timestamp 1679235063
transform 1 0 24380 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_2_259
timestamp 1679235063
transform 1 0 24932 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_2_263
timestamp 1679235063
transform 1 0 25300 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_3_3
timestamp 1679235063
transform 1 0 1380 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_3_8
timestamp 1679235063
transform 1 0 1840 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_3_15
timestamp 1679235063
transform 1 0 2484 0 -1 4352
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_3_21
timestamp 1679235063
transform 1 0 3036 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_3_36
timestamp 1679235063
transform 1 0 4416 0 -1 4352
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_3_40
timestamp 1679235063
transform 1 0 4784 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_3_52
timestamp 1679235063
transform 1 0 5888 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_3_57
timestamp 1679235063
transform 1 0 6348 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_3_62
timestamp 1679235063
transform 1 0 6808 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_3_68
timestamp 1679235063
transform 1 0 7360 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_3_71
timestamp 1679235063
transform 1 0 7636 0 -1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_3_79
timestamp 1679235063
transform 1 0 8372 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_3_85
timestamp 1679235063
transform 1 0 8924 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_3_92
timestamp 1679235063
transform 1 0 9568 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_3_98
timestamp 1679235063
transform 1 0 10120 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_3_110
timestamp 1679235063
transform 1 0 11224 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_3_115
timestamp 1679235063
transform 1 0 11684 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_3_125
timestamp 1679235063
transform 1 0 12604 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_3_145
timestamp 1679235063
transform 1 0 14444 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_3_149
timestamp 1679235063
transform 1 0 14812 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_3_166
timestamp 1679235063
transform 1 0 16376 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_3_169
timestamp 1679235063
transform 1 0 16652 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_3_187
timestamp 1679235063
transform 1 0 18308 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_3_207
timestamp 1679235063
transform 1 0 20148 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_3_220
timestamp 1679235063
transform 1 0 21344 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_3_225
timestamp 1679235063
transform 1 0 21804 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_3_243
timestamp 1679235063
transform 1 0 23460 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_3_263
timestamp 1679235063
transform 1 0 25300 0 -1 4352
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_4_5
timestamp 1679235063
transform 1 0 1564 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_4_17
timestamp 1679235063
transform 1 0 2668 0 1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_4_25
timestamp 1679235063
transform 1 0 3404 0 1 4352
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_4_29
timestamp 1679235063
transform 1 0 3772 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_4_41
timestamp 1679235063
transform 1 0 4876 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_4_66
timestamp 1679235063
transform 1 0 7176 0 1 4352
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_4_70
timestamp 1679235063
transform 1 0 7544 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_4_82
timestamp 1679235063
transform 1 0 8648 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_4_87
timestamp 1679235063
transform 1 0 9108 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_4_96
timestamp 1679235063
transform 1 0 9936 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_4_103
timestamp 1679235063
transform 1 0 10580 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_4_110
timestamp 1679235063
transform 1 0 11224 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_4_124
timestamp 1679235063
transform 1 0 12512 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_4_138
timestamp 1679235063
transform 1 0 13800 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_4_143
timestamp 1679235063
transform 1 0 14260 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_4_148
timestamp 1679235063
transform 1 0 14720 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_4_172
timestamp 1679235063
transform 1 0 16928 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_4_176
timestamp 1679235063
transform 1 0 17296 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_4_193
timestamp 1679235063
transform 1 0 18860 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_4_197
timestamp 1679235063
transform 1 0 19228 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_4_215
timestamp 1679235063
transform 1 0 20884 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_4_235
timestamp 1679235063
transform 1 0 22724 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_4_247
timestamp 1679235063
transform 1 0 23828 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_4_251
timestamp 1679235063
transform 1 0 24196 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_4_253
timestamp 1679235063
transform 1 0 24380 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_4_259
timestamp 1679235063
transform 1 0 24932 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_4_263
timestamp 1679235063
transform 1 0 25300 0 1 4352
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_5_3
timestamp 1679235063
transform 1 0 1380 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_15
timestamp 1679235063
transform 1 0 2484 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_27
timestamp 1679235063
transform 1 0 3588 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_39
timestamp 1679235063
transform 1 0 4692 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_5_51
timestamp 1679235063
transform 1 0 5796 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_5_55
timestamp 1679235063
transform 1 0 6164 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_5_57
timestamp 1679235063
transform 1 0 6348 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_69
timestamp 1679235063
transform 1 0 7452 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_81
timestamp 1679235063
transform 1 0 8556 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_5_93
timestamp 1679235063
transform 1 0 9660 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_99
timestamp 1679235063
transform 1 0 10212 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_5_103
timestamp 1679235063
transform 1 0 10580 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_5_110
timestamp 1679235063
transform 1 0 11224 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_5_113
timestamp 1679235063
transform 1 0 11500 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_5_125
timestamp 1679235063
transform 1 0 12604 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_5_132
timestamp 1679235063
transform 1 0 13248 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_5_136
timestamp 1679235063
transform 1 0 13616 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_5_157
timestamp 1679235063
transform 1 0 15548 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_5_161
timestamp 1679235063
transform 1 0 15916 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_5_166
timestamp 1679235063
transform 1 0 16376 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_5_169
timestamp 1679235063
transform 1 0 16652 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_5_191
timestamp 1679235063
transform 1 0 18676 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_5_198
timestamp 1679235063
transform 1 0 19320 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_5_222
timestamp 1679235063
transform 1 0 21528 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_5_225
timestamp 1679235063
transform 1 0 21804 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_5_243
timestamp 1679235063
transform 1 0 23460 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_5_247
timestamp 1679235063
transform 1 0 23828 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_5_264
timestamp 1679235063
transform 1 0 25392 0 -1 5440
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_6_3
timestamp 1679235063
transform 1 0 1380 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_15
timestamp 1679235063
transform 1 0 2484 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_6_27
timestamp 1679235063
transform 1 0 3588 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_6_29
timestamp 1679235063
transform 1 0 3772 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_41
timestamp 1679235063
transform 1 0 4876 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_53
timestamp 1679235063
transform 1 0 5980 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_65
timestamp 1679235063
transform 1 0 7084 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_6_77
timestamp 1679235063
transform 1 0 8188 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_83
timestamp 1679235063
transform 1 0 8740 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_6_85
timestamp 1679235063
transform 1 0 8924 0 1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_6_93
timestamp 1679235063
transform 1 0 9660 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_6_116
timestamp 1679235063
transform 1 0 11776 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_6_120
timestamp 1679235063
transform 1 0 12144 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_6_125
timestamp 1679235063
transform 1 0 12604 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_6_129
timestamp 1679235063
transform 1 0 12972 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_6_138
timestamp 1679235063
transform 1 0 13800 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_6_141
timestamp 1679235063
transform 1 0 14076 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_6_152
timestamp 1679235063
transform 1 0 15088 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_6_156
timestamp 1679235063
transform 1 0 15456 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_6_174
timestamp 1679235063
transform 1 0 17112 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_6_194
timestamp 1679235063
transform 1 0 18952 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_6_197
timestamp 1679235063
transform 1 0 19228 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_6_203
timestamp 1679235063
transform 1 0 19780 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_6_207
timestamp 1679235063
transform 1 0 20148 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_6_225
timestamp 1679235063
transform 1 0 21804 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_6_245
timestamp 1679235063
transform 1 0 23644 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_6_249
timestamp 1679235063
transform 1 0 24012 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_6_253
timestamp 1679235063
transform 1 0 24380 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_6_263
timestamp 1679235063
transform 1 0 25300 0 1 5440
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_7_3
timestamp 1679235063
transform 1 0 1380 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_15
timestamp 1679235063
transform 1 0 2484 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_27
timestamp 1679235063
transform 1 0 3588 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_39
timestamp 1679235063
transform 1 0 4692 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_7_51
timestamp 1679235063
transform 1 0 5796 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_7_55
timestamp 1679235063
transform 1 0 6164 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_7_57
timestamp 1679235063
transform 1 0 6348 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_69
timestamp 1679235063
transform 1 0 7452 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_81
timestamp 1679235063
transform 1 0 8556 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_7_93
timestamp 1679235063
transform 1 0 9660 0 -1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_7_101
timestamp 1679235063
transform 1 0 10396 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_7_110
timestamp 1679235063
transform 1 0 11224 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_7_113
timestamp 1679235063
transform 1 0 11500 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_7_123
timestamp 1679235063
transform 1 0 12420 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_7_127
timestamp 1679235063
transform 1 0 12788 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_7_149
timestamp 1679235063
transform 1 0 14812 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_7_162
timestamp 1679235063
transform 1 0 16008 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_7_169
timestamp 1679235063
transform 1 0 16652 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_7_191
timestamp 1679235063
transform 1 0 18676 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_7_198
timestamp 1679235063
transform 1 0 19320 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_7_202
timestamp 1679235063
transform 1 0 19688 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_7_222
timestamp 1679235063
transform 1 0 21528 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_7_225
timestamp 1679235063
transform 1 0 21804 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_7_243
timestamp 1679235063
transform 1 0 23460 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_7_247
timestamp 1679235063
transform 1 0 23828 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_7_264
timestamp 1679235063
transform 1 0 25392 0 -1 6528
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_8_3
timestamp 1679235063
transform 1 0 1380 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_15
timestamp 1679235063
transform 1 0 2484 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_8_27
timestamp 1679235063
transform 1 0 3588 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_8_29
timestamp 1679235063
transform 1 0 3772 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_41
timestamp 1679235063
transform 1 0 4876 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_53
timestamp 1679235063
transform 1 0 5980 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_65
timestamp 1679235063
transform 1 0 7084 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_8_77
timestamp 1679235063
transform 1 0 8188 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_83
timestamp 1679235063
transform 1 0 8740 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_8_85
timestamp 1679235063
transform 1 0 8924 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_8_97
timestamp 1679235063
transform 1 0 10028 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_8_123
timestamp 1679235063
transform 1 0 12420 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_8_127
timestamp 1679235063
transform 1 0 12788 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_8_138
timestamp 1679235063
transform 1 0 13800 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_8_141
timestamp 1679235063
transform 1 0 14076 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_8_151
timestamp 1679235063
transform 1 0 14996 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_8_155
timestamp 1679235063
transform 1 0 15364 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_8_161
timestamp 1679235063
transform 1 0 15916 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_8_174
timestamp 1679235063
transform 1 0 17112 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_8_194
timestamp 1679235063
transform 1 0 18952 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_8_197
timestamp 1679235063
transform 1 0 19228 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_8_223
timestamp 1679235063
transform 1 0 21620 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_8_247
timestamp 1679235063
transform 1 0 23828 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_8_251
timestamp 1679235063
transform 1 0 24196 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_8_253
timestamp 1679235063
transform 1 0 24380 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_8_264
timestamp 1679235063
transform 1 0 25392 0 1 6528
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_9_3
timestamp 1679235063
transform 1 0 1380 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_15
timestamp 1679235063
transform 1 0 2484 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_27
timestamp 1679235063
transform 1 0 3588 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_39
timestamp 1679235063
transform 1 0 4692 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_9_51
timestamp 1679235063
transform 1 0 5796 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_9_55
timestamp 1679235063
transform 1 0 6164 0 -1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_9_57
timestamp 1679235063
transform 1 0 6348 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_69
timestamp 1679235063
transform 1 0 7452 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_9_81
timestamp 1679235063
transform 1 0 8556 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_9_85
timestamp 1679235063
transform 1 0 8924 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_9_106
timestamp 1679235063
transform 1 0 10856 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_9_110
timestamp 1679235063
transform 1 0 11224 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_9_113
timestamp 1679235063
transform 1 0 11500 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_9_124
timestamp 1679235063
transform 1 0 12512 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_9_128
timestamp 1679235063
transform 1 0 12880 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_9_139
timestamp 1679235063
transform 1 0 13892 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_9_146
timestamp 1679235063
transform 1 0 14536 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_9_150
timestamp 1679235063
transform 1 0 14904 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_9_160
timestamp 1679235063
transform 1 0 15824 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_9_167
timestamp 1679235063
transform 1 0 16468 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_9_169
timestamp 1679235063
transform 1 0 16652 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_9_182
timestamp 1679235063
transform 1 0 17848 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_9_202
timestamp 1679235063
transform 1 0 19688 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_9_222
timestamp 1679235063
transform 1 0 21528 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_9_225
timestamp 1679235063
transform 1 0 21804 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_9_244
timestamp 1679235063
transform 1 0 23552 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_9_264
timestamp 1679235063
transform 1 0 25392 0 -1 7616
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_10_3
timestamp 1679235063
transform 1 0 1380 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_15
timestamp 1679235063
transform 1 0 2484 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_10_27
timestamp 1679235063
transform 1 0 3588 0 1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_10_29
timestamp 1679235063
transform 1 0 3772 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_41
timestamp 1679235063
transform 1 0 4876 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_53
timestamp 1679235063
transform 1 0 5980 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_65
timestamp 1679235063
transform 1 0 7084 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_10_77
timestamp 1679235063
transform 1 0 8188 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_10_83
timestamp 1679235063
transform 1 0 8740 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_10_85
timestamp 1679235063
transform 1 0 8924 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_10_97
timestamp 1679235063
transform 1 0 10028 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_10_110
timestamp 1679235063
transform 1 0 11224 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_10_114
timestamp 1679235063
transform 1 0 11592 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_10_125
timestamp 1679235063
transform 1 0 12604 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_10_138
timestamp 1679235063
transform 1 0 13800 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_10_141
timestamp 1679235063
transform 1 0 14076 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_10_163
timestamp 1679235063
transform 1 0 16100 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_10_170
timestamp 1679235063
transform 1 0 16744 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_10_194
timestamp 1679235063
transform 1 0 18952 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_10_197
timestamp 1679235063
transform 1 0 19228 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_10_203
timestamp 1679235063
transform 1 0 19780 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_10_207
timestamp 1679235063
transform 1 0 20148 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_10_225
timestamp 1679235063
transform 1 0 21804 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_10_245
timestamp 1679235063
transform 1 0 23644 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_10_249
timestamp 1679235063
transform 1 0 24012 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_10_253
timestamp 1679235063
transform 1 0 24380 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_10_263
timestamp 1679235063
transform 1 0 25300 0 1 7616
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_11_3
timestamp 1679235063
transform 1 0 1380 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_15
timestamp 1679235063
transform 1 0 2484 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_27
timestamp 1679235063
transform 1 0 3588 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_39
timestamp 1679235063
transform 1 0 4692 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_11_51
timestamp 1679235063
transform 1 0 5796 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_11_55
timestamp 1679235063
transform 1 0 6164 0 -1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_11_57
timestamp 1679235063
transform 1 0 6348 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_11_69
timestamp 1679235063
transform 1 0 7452 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_11_73
timestamp 1679235063
transform 1 0 7820 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_11_77
timestamp 1679235063
transform 1 0 8188 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_11_101
timestamp 1679235063
transform 1 0 10396 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_11_105
timestamp 1679235063
transform 1 0 10764 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_11_110
timestamp 1679235063
transform 1 0 11224 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_11_113
timestamp 1679235063
transform 1 0 11500 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_11_124
timestamp 1679235063
transform 1 0 12512 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_11_136
timestamp 1679235063
transform 1 0 13616 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_11_140
timestamp 1679235063
transform 1 0 13984 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_11_153
timestamp 1679235063
transform 1 0 15180 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_11_166
timestamp 1679235063
transform 1 0 16376 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_11_169
timestamp 1679235063
transform 1 0 16652 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_11_180
timestamp 1679235063
transform 1 0 17664 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_11_184
timestamp 1679235063
transform 1 0 18032 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_11_196
timestamp 1679235063
transform 1 0 19136 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_11_200
timestamp 1679235063
transform 1 0 19504 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_11_222
timestamp 1679235063
transform 1 0 21528 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_11_229
timestamp 1679235063
transform 1 0 22172 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_11_251
timestamp 1679235063
transform 1 0 24196 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_11_263
timestamp 1679235063
transform 1 0 25300 0 -1 8704
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_12_3
timestamp 1679235063
transform 1 0 1380 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_15
timestamp 1679235063
transform 1 0 2484 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_12_27
timestamp 1679235063
transform 1 0 3588 0 1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_12_29
timestamp 1679235063
transform 1 0 3772 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_41
timestamp 1679235063
transform 1 0 4876 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_53
timestamp 1679235063
transform 1 0 5980 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_65
timestamp 1679235063
transform 1 0 7084 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_12_77
timestamp 1679235063
transform 1 0 8188 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_12_83
timestamp 1679235063
transform 1 0 8740 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_12_85
timestamp 1679235063
transform 1 0 8924 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_12_95
timestamp 1679235063
transform 1 0 9844 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_12_99
timestamp 1679235063
transform 1 0 10212 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_12_110
timestamp 1679235063
transform 1 0 11224 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_12_114
timestamp 1679235063
transform 1 0 11592 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_12_118
timestamp 1679235063
transform 1 0 11960 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_12_125
timestamp 1679235063
transform 1 0 12604 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_12_138
timestamp 1679235063
transform 1 0 13800 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_12_141
timestamp 1679235063
transform 1 0 14076 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_12_147
timestamp 1679235063
transform 1 0 14628 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_12_151
timestamp 1679235063
transform 1 0 14996 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_12_155
timestamp 1679235063
transform 1 0 15364 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_12_166
timestamp 1679235063
transform 1 0 16376 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_12_172
timestamp 1679235063
transform 1 0 16928 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_12_182
timestamp 1679235063
transform 1 0 17848 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_12_194
timestamp 1679235063
transform 1 0 18952 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_12_199
timestamp 1679235063
transform 1 0 19412 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_12_210
timestamp 1679235063
transform 1 0 20424 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_12_230
timestamp 1679235063
transform 1 0 22264 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_12_250
timestamp 1679235063
transform 1 0 24104 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_12_253
timestamp 1679235063
transform 1 0 24380 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_12_263
timestamp 1679235063
transform 1 0 25300 0 1 8704
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_13_3
timestamp 1679235063
transform 1 0 1380 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_15
timestamp 1679235063
transform 1 0 2484 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_27
timestamp 1679235063
transform 1 0 3588 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_39
timestamp 1679235063
transform 1 0 4692 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_13_51
timestamp 1679235063
transform 1 0 5796 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_13_55
timestamp 1679235063
transform 1 0 6164 0 -1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_13_57
timestamp 1679235063
transform 1 0 6348 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_13_69
timestamp 1679235063
transform 1 0 7452 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_13_75
timestamp 1679235063
transform 1 0 8004 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_13_98
timestamp 1679235063
transform 1 0 10120 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_13_102
timestamp 1679235063
transform 1 0 10488 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_13_106
timestamp 1679235063
transform 1 0 10856 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_13_113
timestamp 1679235063
transform 1 0 11500 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_13_135
timestamp 1679235063
transform 1 0 13524 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_13_142
timestamp 1679235063
transform 1 0 14168 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_13_146
timestamp 1679235063
transform 1 0 14536 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_13_156
timestamp 1679235063
transform 1 0 15456 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_13_160
timestamp 1679235063
transform 1 0 15824 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_13_166
timestamp 1679235063
transform 1 0 16376 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_13_169
timestamp 1679235063
transform 1 0 16652 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_13_175
timestamp 1679235063
transform 1 0 17204 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_13_179
timestamp 1679235063
transform 1 0 17572 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_13_200
timestamp 1679235063
transform 1 0 19504 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_13_213
timestamp 1679235063
transform 1 0 20700 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_13_221
timestamp 1679235063
transform 1 0 21436 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_13_225
timestamp 1679235063
transform 1 0 21804 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_13_244
timestamp 1679235063
transform 1 0 23552 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_13_264
timestamp 1679235063
transform 1 0 25392 0 -1 9792
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_14_3
timestamp 1679235063
transform 1 0 1380 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_15
timestamp 1679235063
transform 1 0 2484 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_14_27
timestamp 1679235063
transform 1 0 3588 0 1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_14_29
timestamp 1679235063
transform 1 0 3772 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_41
timestamp 1679235063
transform 1 0 4876 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_53
timestamp 1679235063
transform 1 0 5980 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_65
timestamp 1679235063
transform 1 0 7084 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_14_77
timestamp 1679235063
transform 1 0 8188 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_14_82
timestamp 1679235063
transform 1 0 8648 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_14_85
timestamp 1679235063
transform 1 0 8924 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_14_107
timestamp 1679235063
transform 1 0 10948 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_14_111
timestamp 1679235063
transform 1 0 11316 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_14_122
timestamp 1679235063
transform 1 0 12328 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_14_135
timestamp 1679235063
transform 1 0 13524 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_14_143
timestamp 1679235063
transform 1 0 14260 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_14_154
timestamp 1679235063
transform 1 0 15272 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_14_167
timestamp 1679235063
transform 1 0 16468 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_14_180
timestamp 1679235063
transform 1 0 17664 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_14_184
timestamp 1679235063
transform 1 0 18032 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_14_194
timestamp 1679235063
transform 1 0 18952 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_14_197
timestamp 1679235063
transform 1 0 19228 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_14_207
timestamp 1679235063
transform 1 0 20148 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_14_211
timestamp 1679235063
transform 1 0 20516 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_14_223
timestamp 1679235063
transform 1 0 21620 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_14_227
timestamp 1679235063
transform 1 0 21988 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_14_250
timestamp 1679235063
transform 1 0 24104 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_14_253
timestamp 1679235063
transform 1 0 24380 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_14_258
timestamp 1679235063
transform 1 0 24840 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_14_262
timestamp 1679235063
transform 1 0 25208 0 1 9792
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_15_3
timestamp 1679235063
transform 1 0 1380 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_15
timestamp 1679235063
transform 1 0 2484 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_27
timestamp 1679235063
transform 1 0 3588 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_39
timestamp 1679235063
transform 1 0 4692 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_15_51
timestamp 1679235063
transform 1 0 5796 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_15_55
timestamp 1679235063
transform 1 0 6164 0 -1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_15_57
timestamp 1679235063
transform 1 0 6348 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_69
timestamp 1679235063
transform 1 0 7452 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_15_81
timestamp 1679235063
transform 1 0 8556 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_15_87
timestamp 1679235063
transform 1 0 9108 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_15_109
timestamp 1679235063
transform 1 0 11132 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_15_113
timestamp 1679235063
transform 1 0 11500 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_15_118
timestamp 1679235063
transform 1 0 11960 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_15_122
timestamp 1679235063
transform 1 0 12328 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_15_133
timestamp 1679235063
transform 1 0 13340 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_15_137
timestamp 1679235063
transform 1 0 13708 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_15_148
timestamp 1679235063
transform 1 0 14720 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_15_154
timestamp 1679235063
transform 1 0 15272 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_15_165
timestamp 1679235063
transform 1 0 16284 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_15_169
timestamp 1679235063
transform 1 0 16652 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_15_179
timestamp 1679235063
transform 1 0 17572 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_15_187
timestamp 1679235063
transform 1 0 18308 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_15_192
timestamp 1679235063
transform 1 0 18768 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_15_198
timestamp 1679235063
transform 1 0 19320 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_15_222
timestamp 1679235063
transform 1 0 21528 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_15_225
timestamp 1679235063
transform 1 0 21804 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_15_237
timestamp 1679235063
transform 1 0 22908 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_15_244
timestamp 1679235063
transform 1 0 23552 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_15_264
timestamp 1679235063
transform 1 0 25392 0 -1 10880
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_16_3
timestamp 1679235063
transform 1 0 1380 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_15
timestamp 1679235063
transform 1 0 2484 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_16_27
timestamp 1679235063
transform 1 0 3588 0 1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_16_29
timestamp 1679235063
transform 1 0 3772 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_41
timestamp 1679235063
transform 1 0 4876 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_53
timestamp 1679235063
transform 1 0 5980 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_16_65
timestamp 1679235063
transform 1 0 7084 0 1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_16_73
timestamp 1679235063
transform 1 0 7820 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_16_82
timestamp 1679235063
transform 1 0 8648 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_16_85
timestamp 1679235063
transform 1 0 8924 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_16_97
timestamp 1679235063
transform 1 0 10028 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_16_102
timestamp 1679235063
transform 1 0 10488 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_16_107
timestamp 1679235063
transform 1 0 10948 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_16_120
timestamp 1679235063
transform 1 0 12144 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_16_124
timestamp 1679235063
transform 1 0 12512 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_16_134
timestamp 1679235063
transform 1 0 13432 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_16_145
timestamp 1679235063
transform 1 0 14444 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_16_167
timestamp 1679235063
transform 1 0 16468 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_16_174
timestamp 1679235063
transform 1 0 17112 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_16_178
timestamp 1679235063
transform 1 0 17480 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_16_190
timestamp 1679235063
transform 1 0 18584 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_16_197
timestamp 1679235063
transform 1 0 19228 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_16_203
timestamp 1679235063
transform 1 0 19780 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_16_211
timestamp 1679235063
transform 1 0 20516 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_16_218
timestamp 1679235063
transform 1 0 21160 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_16_225
timestamp 1679235063
transform 1 0 21804 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_16_233
timestamp 1679235063
transform 1 0 22540 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_16_244
timestamp 1679235063
transform 1 0 23552 0 1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_16_253
timestamp 1679235063
transform 1 0 24380 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_16_263
timestamp 1679235063
transform 1 0 25300 0 1 10880
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_17_3
timestamp 1679235063
transform 1 0 1380 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_15
timestamp 1679235063
transform 1 0 2484 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_27
timestamp 1679235063
transform 1 0 3588 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_39
timestamp 1679235063
transform 1 0 4692 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_17_51
timestamp 1679235063
transform 1 0 5796 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_17_55
timestamp 1679235063
transform 1 0 6164 0 -1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_17_57
timestamp 1679235063
transform 1 0 6348 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_17_69
timestamp 1679235063
transform 1 0 7452 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_17_81
timestamp 1679235063
transform 1 0 8556 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_17_94
timestamp 1679235063
transform 1 0 9752 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_17_107
timestamp 1679235063
transform 1 0 10948 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_17_111
timestamp 1679235063
transform 1 0 11316 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_17_113
timestamp 1679235063
transform 1 0 11500 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_17_117
timestamp 1679235063
transform 1 0 11868 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_17_127
timestamp 1679235063
transform 1 0 12788 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_17_140
timestamp 1679235063
transform 1 0 13984 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_17_153
timestamp 1679235063
transform 1 0 15180 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_17_165
timestamp 1679235063
transform 1 0 16284 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_17_169
timestamp 1679235063
transform 1 0 16652 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_17_180
timestamp 1679235063
transform 1 0 17664 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_17_193
timestamp 1679235063
transform 1 0 18860 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_17_199
timestamp 1679235063
transform 1 0 19412 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_17_210
timestamp 1679235063
transform 1 0 20424 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_17_218
timestamp 1679235063
transform 1 0 21160 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_17_225
timestamp 1679235063
transform 1 0 21804 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_17_235
timestamp 1679235063
transform 1 0 22724 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_17_259
timestamp 1679235063
transform 1 0 24932 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_17_263
timestamp 1679235063
transform 1 0 25300 0 -1 11968
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_18_3
timestamp 1679235063
transform 1 0 1380 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_15
timestamp 1679235063
transform 1 0 2484 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_18_27
timestamp 1679235063
transform 1 0 3588 0 1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_18_29
timestamp 1679235063
transform 1 0 3772 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_41
timestamp 1679235063
transform 1 0 4876 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_53
timestamp 1679235063
transform 1 0 5980 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_18_65
timestamp 1679235063
transform 1 0 7084 0 1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_18_82
timestamp 1679235063
transform 1 0 8648 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_18_87
timestamp 1679235063
transform 1 0 9108 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_18_92
timestamp 1679235063
transform 1 0 9568 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_18_103
timestamp 1679235063
transform 1 0 10580 0 1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_18_111
timestamp 1679235063
transform 1 0 11316 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_18_121
timestamp 1679235063
transform 1 0 12236 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_18_134
timestamp 1679235063
transform 1 0 13432 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_18_141
timestamp 1679235063
transform 1 0 14076 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_18_153
timestamp 1679235063
transform 1 0 15180 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_18_160
timestamp 1679235063
transform 1 0 15824 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_18_167
timestamp 1679235063
transform 1 0 16468 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_18_180
timestamp 1679235063
transform 1 0 17664 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_18_184
timestamp 1679235063
transform 1 0 18032 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_18_187
timestamp 1679235063
transform 1 0 18308 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_18_193
timestamp 1679235063
transform 1 0 18860 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_18_197
timestamp 1679235063
transform 1 0 19228 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_18_203
timestamp 1679235063
transform 1 0 19780 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_18_207
timestamp 1679235063
transform 1 0 20148 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_18_229
timestamp 1679235063
transform 1 0 22172 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_18_233
timestamp 1679235063
transform 1 0 22540 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_18_250
timestamp 1679235063
transform 1 0 24104 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_18_253
timestamp 1679235063
transform 1 0 24380 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_18_264
timestamp 1679235063
transform 1 0 25392 0 1 11968
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_19_3
timestamp 1679235063
transform 1 0 1380 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_15
timestamp 1679235063
transform 1 0 2484 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_27
timestamp 1679235063
transform 1 0 3588 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_39
timestamp 1679235063
transform 1 0 4692 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_19_51
timestamp 1679235063
transform 1 0 5796 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_19_55
timestamp 1679235063
transform 1 0 6164 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_19_57
timestamp 1679235063
transform 1 0 6348 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_19_62
timestamp 1679235063
transform 1 0 6808 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_19_86
timestamp 1679235063
transform 1 0 9016 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_19_90
timestamp 1679235063
transform 1 0 9384 0 -1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_19_98
timestamp 1679235063
transform 1 0 10120 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_19_109
timestamp 1679235063
transform 1 0 11132 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_19_113
timestamp 1679235063
transform 1 0 11500 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_19_116
timestamp 1679235063
transform 1 0 11776 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_19_121
timestamp 1679235063
transform 1 0 12236 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_19_134
timestamp 1679235063
transform 1 0 13432 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_19_138
timestamp 1679235063
transform 1 0 13800 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_19_150
timestamp 1679235063
transform 1 0 14904 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_19_154
timestamp 1679235063
transform 1 0 15272 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_19_159
timestamp 1679235063
transform 1 0 15732 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_19_166
timestamp 1679235063
transform 1 0 16376 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_19_173
timestamp 1679235063
transform 1 0 17020 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_19_186
timestamp 1679235063
transform 1 0 18216 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_19_190
timestamp 1679235063
transform 1 0 18584 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_19_200
timestamp 1679235063
transform 1 0 19504 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_19_208
timestamp 1679235063
transform 1 0 20240 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_19_216
timestamp 1679235063
transform 1 0 20976 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_19_222
timestamp 1679235063
transform 1 0 21528 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_19_225
timestamp 1679235063
transform 1 0 21804 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_19_230
timestamp 1679235063
transform 1 0 22264 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_19_236
timestamp 1679235063
transform 1 0 22816 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_19_258
timestamp 1679235063
transform 1 0 24840 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_19_262
timestamp 1679235063
transform 1 0 25208 0 -1 13056
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_20_3
timestamp 1679235063
transform 1 0 1380 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_15
timestamp 1679235063
transform 1 0 2484 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_20_27
timestamp 1679235063
transform 1 0 3588 0 1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_20_29
timestamp 1679235063
transform 1 0 3772 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_41
timestamp 1679235063
transform 1 0 4876 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_20_53
timestamp 1679235063
transform 1 0 5980 0 1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_20_61
timestamp 1679235063
transform 1 0 6716 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_20_73
timestamp 1679235063
transform 1 0 7820 0 1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_20_81
timestamp 1679235063
transform 1 0 8556 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_20_85
timestamp 1679235063
transform 1 0 8924 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_20_90
timestamp 1679235063
transform 1 0 9384 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_20_114
timestamp 1679235063
transform 1 0 11592 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_20_129
timestamp 1679235063
transform 1 0 12972 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_20_133
timestamp 1679235063
transform 1 0 13340 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_20_138
timestamp 1679235063
transform 1 0 13800 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_20_143
timestamp 1679235063
transform 1 0 14260 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_20_149
timestamp 1679235063
transform 1 0 14812 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_20_162
timestamp 1679235063
transform 1 0 16008 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_20_175
timestamp 1679235063
transform 1 0 17204 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_20_187
timestamp 1679235063
transform 1 0 18308 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_20_194
timestamp 1679235063
transform 1 0 18952 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_20_197
timestamp 1679235063
transform 1 0 19228 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_20_203
timestamp 1679235063
transform 1 0 19780 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_20_216
timestamp 1679235063
transform 1 0 20976 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_20_220
timestamp 1679235063
transform 1 0 21344 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_20_230
timestamp 1679235063
transform 1 0 22264 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_20_250
timestamp 1679235063
transform 1 0 24104 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_20_253
timestamp 1679235063
transform 1 0 24380 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_20_263
timestamp 1679235063
transform 1 0 25300 0 1 13056
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_21_3
timestamp 1679235063
transform 1 0 1380 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_15
timestamp 1679235063
transform 1 0 2484 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_27
timestamp 1679235063
transform 1 0 3588 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_39
timestamp 1679235063
transform 1 0 4692 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_21_51
timestamp 1679235063
transform 1 0 5796 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_21_55
timestamp 1679235063
transform 1 0 6164 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_21_57
timestamp 1679235063
transform 1 0 6348 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_21_79
timestamp 1679235063
transform 1 0 8372 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_21_83
timestamp 1679235063
transform 1 0 8740 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_21_96
timestamp 1679235063
transform 1 0 9936 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_21_100
timestamp 1679235063
transform 1 0 10304 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_21_110
timestamp 1679235063
transform 1 0 11224 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_21_113
timestamp 1679235063
transform 1 0 11500 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_21_118
timestamp 1679235063
transform 1 0 11960 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_21_131
timestamp 1679235063
transform 1 0 13156 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_21_155
timestamp 1679235063
transform 1 0 15364 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_21_161
timestamp 1679235063
transform 1 0 15916 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_21_166
timestamp 1679235063
transform 1 0 16376 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_21_169
timestamp 1679235063
transform 1 0 16652 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_21_191
timestamp 1679235063
transform 1 0 18676 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_21_206
timestamp 1679235063
transform 1 0 20056 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_21_210
timestamp 1679235063
transform 1 0 20424 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_21_215
timestamp 1679235063
transform 1 0 20884 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_21_222
timestamp 1679235063
transform 1 0 21528 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_21_225
timestamp 1679235063
transform 1 0 21804 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_21_244
timestamp 1679235063
transform 1 0 23552 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_21_264
timestamp 1679235063
transform 1 0 25392 0 -1 14144
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_22_3
timestamp 1679235063
transform 1 0 1380 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_15
timestamp 1679235063
transform 1 0 2484 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_22_27
timestamp 1679235063
transform 1 0 3588 0 1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_22_29
timestamp 1679235063
transform 1 0 3772 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_41
timestamp 1679235063
transform 1 0 4876 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_53
timestamp 1679235063
transform 1 0 5980 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_22_65
timestamp 1679235063
transform 1 0 7084 0 1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_22_73
timestamp 1679235063
transform 1 0 7820 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_22_82
timestamp 1679235063
transform 1 0 8648 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_22_85
timestamp 1679235063
transform 1 0 8924 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_22_96
timestamp 1679235063
transform 1 0 9936 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_22_111
timestamp 1679235063
transform 1 0 11316 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_22_124
timestamp 1679235063
transform 1 0 12512 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_22_128
timestamp 1679235063
transform 1 0 12880 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_22_138
timestamp 1679235063
transform 1 0 13800 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_22_141
timestamp 1679235063
transform 1 0 14076 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_22_147
timestamp 1679235063
transform 1 0 14628 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_22_160
timestamp 1679235063
transform 1 0 15824 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_22_166
timestamp 1679235063
transform 1 0 16376 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_22_171
timestamp 1679235063
transform 1 0 16836 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_22_185
timestamp 1679235063
transform 1 0 18124 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_22_189
timestamp 1679235063
transform 1 0 18492 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_22_194
timestamp 1679235063
transform 1 0 18952 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_22_197
timestamp 1679235063
transform 1 0 19228 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_22_203
timestamp 1679235063
transform 1 0 19780 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_22_210
timestamp 1679235063
transform 1 0 20424 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_22_214
timestamp 1679235063
transform 1 0 20792 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_22_218
timestamp 1679235063
transform 1 0 21160 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_22_226
timestamp 1679235063
transform 1 0 21896 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_22_250
timestamp 1679235063
transform 1 0 24104 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_22_253
timestamp 1679235063
transform 1 0 24380 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_22_258
timestamp 1679235063
transform 1 0 24840 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_22_262
timestamp 1679235063
transform 1 0 25208 0 1 14144
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_23_3
timestamp 1679235063
transform 1 0 1380 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_15
timestamp 1679235063
transform 1 0 2484 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_27
timestamp 1679235063
transform 1 0 3588 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_39
timestamp 1679235063
transform 1 0 4692 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_23_51
timestamp 1679235063
transform 1 0 5796 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_23_55
timestamp 1679235063
transform 1 0 6164 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_23_57
timestamp 1679235063
transform 1 0 6348 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_23_68
timestamp 1679235063
transform 1 0 7360 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_23_95
timestamp 1679235063
transform 1 0 9844 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_23_108
timestamp 1679235063
transform 1 0 11040 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_23_113
timestamp 1679235063
transform 1 0 11500 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_23_123
timestamp 1679235063
transform 1 0 12420 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_23_129
timestamp 1679235063
transform 1 0 12972 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_23_134
timestamp 1679235063
transform 1 0 13432 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_23_145
timestamp 1679235063
transform 1 0 14444 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_23_149
timestamp 1679235063
transform 1 0 14812 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_23_153
timestamp 1679235063
transform 1 0 15180 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_23_166
timestamp 1679235063
transform 1 0 16376 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_23_169
timestamp 1679235063
transform 1 0 16652 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_23_181
timestamp 1679235063
transform 1 0 17756 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_23_186
timestamp 1679235063
transform 1 0 18216 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_23_193
timestamp 1679235063
transform 1 0 18860 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_23_199
timestamp 1679235063
transform 1 0 19412 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_23_209
timestamp 1679235063
transform 1 0 20332 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_23_222
timestamp 1679235063
transform 1 0 21528 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_23_229
timestamp 1679235063
transform 1 0 22172 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_23_240
timestamp 1679235063
transform 1 0 23184 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_23_246
timestamp 1679235063
transform 1 0 23736 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_23_264
timestamp 1679235063
transform 1 0 25392 0 -1 15232
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_24_3
timestamp 1679235063
transform 1 0 1380 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_15
timestamp 1679235063
transform 1 0 2484 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_24_27
timestamp 1679235063
transform 1 0 3588 0 1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_24_29
timestamp 1679235063
transform 1 0 3772 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_41
timestamp 1679235063
transform 1 0 4876 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_24_53
timestamp 1679235063
transform 1 0 5980 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_24_77
timestamp 1679235063
transform 1 0 8188 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_24_81
timestamp 1679235063
transform 1 0 8556 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_24_85
timestamp 1679235063
transform 1 0 8924 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_24_91
timestamp 1679235063
transform 1 0 9476 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_24_94
timestamp 1679235063
transform 1 0 9752 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_24_119
timestamp 1679235063
transform 1 0 12052 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_24_123
timestamp 1679235063
transform 1 0 12420 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_24_127
timestamp 1679235063
transform 1 0 12788 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_24_138
timestamp 1679235063
transform 1 0 13800 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_24_141
timestamp 1679235063
transform 1 0 14076 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_24_146
timestamp 1679235063
transform 1 0 14536 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_24_150
timestamp 1679235063
transform 1 0 14904 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_24_157
timestamp 1679235063
transform 1 0 15548 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_24_161
timestamp 1679235063
transform 1 0 15916 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_24_184
timestamp 1679235063
transform 1 0 18032 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_24_188
timestamp 1679235063
transform 1 0 18400 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_24_192
timestamp 1679235063
transform 1 0 18768 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_24_197
timestamp 1679235063
transform 1 0 19228 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_24_219
timestamp 1679235063
transform 1 0 21252 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_24_226
timestamp 1679235063
transform 1 0 21896 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_24_250
timestamp 1679235063
transform 1 0 24104 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_24_253
timestamp 1679235063
transform 1 0 24380 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_24_263
timestamp 1679235063
transform 1 0 25300 0 1 15232
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_25_3
timestamp 1679235063
transform 1 0 1380 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_15
timestamp 1679235063
transform 1 0 2484 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_27
timestamp 1679235063
transform 1 0 3588 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_39
timestamp 1679235063
transform 1 0 4692 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_25_51
timestamp 1679235063
transform 1 0 5796 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_25_55
timestamp 1679235063
transform 1 0 6164 0 -1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_25_57
timestamp 1679235063
transform 1 0 6348 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_25_69
timestamp 1679235063
transform 1 0 7452 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_25_93
timestamp 1679235063
transform 1 0 9660 0 -1 16320
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_25_97
timestamp 1679235063
transform 1 0 10028 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_25_109
timestamp 1679235063
transform 1 0 11132 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_25_113
timestamp 1679235063
transform 1 0 11500 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_25_135
timestamp 1679235063
transform 1 0 13524 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_25_139
timestamp 1679235063
transform 1 0 13892 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_25_150
timestamp 1679235063
transform 1 0 14904 0 -1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_25_166
timestamp 1679235063
transform 1 0 16376 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_25_169
timestamp 1679235063
transform 1 0 16652 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_25_172
timestamp 1679235063
transform 1 0 16928 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_25_178
timestamp 1679235063
transform 1 0 17480 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_25_182
timestamp 1679235063
transform 1 0 17848 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_25_186
timestamp 1679235063
transform 1 0 18216 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_25_198
timestamp 1679235063
transform 1 0 19320 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_25_222
timestamp 1679235063
transform 1 0 21528 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_25_225
timestamp 1679235063
transform 1 0 21804 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_25_247
timestamp 1679235063
transform 1 0 23828 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_25_252
timestamp 1679235063
transform 1 0 24288 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_25_262
timestamp 1679235063
transform 1 0 25208 0 -1 16320
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_26_3
timestamp 1679235063
transform 1 0 1380 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_15
timestamp 1679235063
transform 1 0 2484 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_26_27
timestamp 1679235063
transform 1 0 3588 0 1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_26_29
timestamp 1679235063
transform 1 0 3772 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_26_41
timestamp 1679235063
transform 1 0 4876 0 1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_26_49
timestamp 1679235063
transform 1 0 5612 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_26_72
timestamp 1679235063
transform 1 0 7728 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_26_76
timestamp 1679235063
transform 1 0 8096 0 1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_26_85
timestamp 1679235063
transform 1 0 8924 0 1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_26_93
timestamp 1679235063
transform 1 0 9660 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_26_97
timestamp 1679235063
transform 1 0 10028 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_26_108
timestamp 1679235063
transform 1 0 11040 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_26_114
timestamp 1679235063
transform 1 0 11592 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_26_125
timestamp 1679235063
transform 1 0 12604 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_26_138
timestamp 1679235063
transform 1 0 13800 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_26_145
timestamp 1679235063
transform 1 0 14444 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_26_149
timestamp 1679235063
transform 1 0 14812 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_26_152
timestamp 1679235063
transform 1 0 15088 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_26_163
timestamp 1679235063
transform 1 0 16100 0 1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_26_175
timestamp 1679235063
transform 1 0 17204 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_26_182
timestamp 1679235063
transform 1 0 17848 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_26_186
timestamp 1679235063
transform 1 0 18216 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_26_191
timestamp 1679235063
transform 1 0 18676 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_26_197
timestamp 1679235063
transform 1 0 19228 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_26_210
timestamp 1679235063
transform 1 0 20424 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_26_222
timestamp 1679235063
transform 1 0 21528 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_26_229
timestamp 1679235063
transform 1 0 22172 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_26_233
timestamp 1679235063
transform 1 0 22540 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_26_250
timestamp 1679235063
transform 1 0 24104 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_26_253
timestamp 1679235063
transform 1 0 24380 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_26_263
timestamp 1679235063
transform 1 0 25300 0 1 16320
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_27_3
timestamp 1679235063
transform 1 0 1380 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_15
timestamp 1679235063
transform 1 0 2484 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_27
timestamp 1679235063
transform 1 0 3588 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_39
timestamp 1679235063
transform 1 0 4692 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_27_51
timestamp 1679235063
transform 1 0 5796 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_27_55
timestamp 1679235063
transform 1 0 6164 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_27_57
timestamp 1679235063
transform 1 0 6348 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_27_71
timestamp 1679235063
transform 1 0 7636 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_27_78
timestamp 1679235063
transform 1 0 8280 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_27_82
timestamp 1679235063
transform 1 0 8648 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_27_85
timestamp 1679235063
transform 1 0 8924 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_27_96
timestamp 1679235063
transform 1 0 9936 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_27_109
timestamp 1679235063
transform 1 0 11132 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_27_113
timestamp 1679235063
transform 1 0 11500 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_27_124
timestamp 1679235063
transform 1 0 12512 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_27_137
timestamp 1679235063
transform 1 0 13708 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_27_141
timestamp 1679235063
transform 1 0 14076 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_27_165
timestamp 1679235063
transform 1 0 16284 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_27_171
timestamp 1679235063
transform 1 0 16836 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_27_174
timestamp 1679235063
transform 1 0 17112 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_27_187
timestamp 1679235063
transform 1 0 18308 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_27_199
timestamp 1679235063
transform 1 0 19412 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_27_207
timestamp 1679235063
transform 1 0 20148 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_27_211
timestamp 1679235063
transform 1 0 20516 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_27_222
timestamp 1679235063
transform 1 0 21528 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_27_225
timestamp 1679235063
transform 1 0 21804 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_27_244
timestamp 1679235063
transform 1 0 23552 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_27_264
timestamp 1679235063
transform 1 0 25392 0 -1 17408
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_28_3
timestamp 1679235063
transform 1 0 1380 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_15
timestamp 1679235063
transform 1 0 2484 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_28_27
timestamp 1679235063
transform 1 0 3588 0 1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_28_29
timestamp 1679235063
transform 1 0 3772 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_41
timestamp 1679235063
transform 1 0 4876 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_53
timestamp 1679235063
transform 1 0 5980 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_28_65
timestamp 1679235063
transform 1 0 7084 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_28_69
timestamp 1679235063
transform 1 0 7452 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_28_80
timestamp 1679235063
transform 1 0 8464 0 1 17408
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_28_87
timestamp 1679235063
transform 1 0 9108 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_28_110
timestamp 1679235063
transform 1 0 11224 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_28_118
timestamp 1679235063
transform 1 0 11960 0 1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_28_126
timestamp 1679235063
transform 1 0 12696 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_28_135
timestamp 1679235063
transform 1 0 13524 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_28_141
timestamp 1679235063
transform 1 0 14076 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_28_147
timestamp 1679235063
transform 1 0 14628 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_28_154
timestamp 1679235063
transform 1 0 15272 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_28_161
timestamp 1679235063
transform 1 0 15916 0 1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_28_172
timestamp 1679235063
transform 1 0 16928 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_28_179
timestamp 1679235063
transform 1 0 17572 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_28_192
timestamp 1679235063
transform 1 0 18768 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_28_197
timestamp 1679235063
transform 1 0 19228 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_28_219
timestamp 1679235063
transform 1 0 21252 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_28_224
timestamp 1679235063
transform 1 0 21712 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_28_230
timestamp 1679235063
transform 1 0 22264 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_28_250
timestamp 1679235063
transform 1 0 24104 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_28_253
timestamp 1679235063
transform 1 0 24380 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_28_264
timestamp 1679235063
transform 1 0 25392 0 1 17408
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_29_3
timestamp 1679235063
transform 1 0 1380 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_15
timestamp 1679235063
transform 1 0 2484 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_27
timestamp 1679235063
transform 1 0 3588 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_39
timestamp 1679235063
transform 1 0 4692 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_29_51
timestamp 1679235063
transform 1 0 5796 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_29_55
timestamp 1679235063
transform 1 0 6164 0 -1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_29_57
timestamp 1679235063
transform 1 0 6348 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_29_69
timestamp 1679235063
transform 1 0 7452 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_29_73
timestamp 1679235063
transform 1 0 7820 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_29_83
timestamp 1679235063
transform 1 0 8740 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_29_110
timestamp 1679235063
transform 1 0 11224 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_29_113
timestamp 1679235063
transform 1 0 11500 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_29_118
timestamp 1679235063
transform 1 0 11960 0 -1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_29_126
timestamp 1679235063
transform 1 0 12696 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_29_129
timestamp 1679235063
transform 1 0 12972 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_29_140
timestamp 1679235063
transform 1 0 13984 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_29_152
timestamp 1679235063
transform 1 0 15088 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_29_166
timestamp 1679235063
transform 1 0 16376 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_29_169
timestamp 1679235063
transform 1 0 16652 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_29_191
timestamp 1679235063
transform 1 0 18676 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_29_197
timestamp 1679235063
transform 1 0 19228 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_29_202
timestamp 1679235063
transform 1 0 19688 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_29_209
timestamp 1679235063
transform 1 0 20332 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_29_216
timestamp 1679235063
transform 1 0 20976 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_29_222
timestamp 1679235063
transform 1 0 21528 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_29_225
timestamp 1679235063
transform 1 0 21804 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_29_235
timestamp 1679235063
transform 1 0 22724 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_29_239
timestamp 1679235063
transform 1 0 23092 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_29_264
timestamp 1679235063
transform 1 0 25392 0 -1 18496
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_30_3
timestamp 1679235063
transform 1 0 1380 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_15
timestamp 1679235063
transform 1 0 2484 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_30_27
timestamp 1679235063
transform 1 0 3588 0 1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_30_29
timestamp 1679235063
transform 1 0 3772 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_41
timestamp 1679235063
transform 1 0 4876 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_30_53
timestamp 1679235063
transform 1 0 5980 0 1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_30_61
timestamp 1679235063
transform 1 0 6716 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_30_82
timestamp 1679235063
transform 1 0 8648 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_30_85
timestamp 1679235063
transform 1 0 8924 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_30_90
timestamp 1679235063
transform 1 0 9384 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_30_103
timestamp 1679235063
transform 1 0 10580 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_30_116
timestamp 1679235063
transform 1 0 11776 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_30_131
timestamp 1679235063
transform 1 0 13156 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_30_135
timestamp 1679235063
transform 1 0 13524 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_30_141
timestamp 1679235063
transform 1 0 14076 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_30_152
timestamp 1679235063
transform 1 0 15088 0 1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_30_160
timestamp 1679235063
transform 1 0 15824 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_30_165
timestamp 1679235063
transform 1 0 16284 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_30_169
timestamp 1679235063
transform 1 0 16652 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_30_179
timestamp 1679235063
transform 1 0 17572 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_30_192
timestamp 1679235063
transform 1 0 18768 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_30_197
timestamp 1679235063
transform 1 0 19228 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_30_207
timestamp 1679235063
transform 1 0 20148 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_30_211
timestamp 1679235063
transform 1 0 20516 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_30_221
timestamp 1679235063
transform 1 0 21436 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_30_228
timestamp 1679235063
transform 1 0 22080 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_30_232
timestamp 1679235063
transform 1 0 22448 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_30_250
timestamp 1679235063
transform 1 0 24104 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_30_253
timestamp 1679235063
transform 1 0 24380 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_30_264
timestamp 1679235063
transform 1 0 25392 0 1 18496
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_31_3
timestamp 1679235063
transform 1 0 1380 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_15
timestamp 1679235063
transform 1 0 2484 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_27
timestamp 1679235063
transform 1 0 3588 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_39
timestamp 1679235063
transform 1 0 4692 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_31_51
timestamp 1679235063
transform 1 0 5796 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_31_55
timestamp 1679235063
transform 1 0 6164 0 -1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_31_57
timestamp 1679235063
transform 1 0 6348 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_31_89
timestamp 1679235063
transform 1 0 9292 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_31_93
timestamp 1679235063
transform 1 0 9660 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_31_96
timestamp 1679235063
transform 1 0 9936 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_31_107
timestamp 1679235063
transform 1 0 10948 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_31_111
timestamp 1679235063
transform 1 0 11316 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_31_115
timestamp 1679235063
transform 1 0 11684 0 -1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_31_121
timestamp 1679235063
transform 1 0 12236 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_31_142
timestamp 1679235063
transform 1 0 14168 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_31_154
timestamp 1679235063
transform 1 0 15272 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_31_161
timestamp 1679235063
transform 1 0 15916 0 -1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_31_167
timestamp 1679235063
transform 1 0 16468 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_31_169
timestamp 1679235063
transform 1 0 16652 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_31_180
timestamp 1679235063
transform 1 0 17664 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_31_184
timestamp 1679235063
transform 1 0 18032 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_31_193
timestamp 1679235063
transform 1 0 18860 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_31_200
timestamp 1679235063
transform 1 0 19504 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_31_204
timestamp 1679235063
transform 1 0 19872 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_31_215
timestamp 1679235063
transform 1 0 20884 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_31_222
timestamp 1679235063
transform 1 0 21528 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_31_227
timestamp 1679235063
transform 1 0 21988 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_31_238
timestamp 1679235063
transform 1 0 23000 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_31_262
timestamp 1679235063
transform 1 0 25208 0 -1 19584
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_32_3
timestamp 1679235063
transform 1 0 1380 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_15
timestamp 1679235063
transform 1 0 2484 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_32_27
timestamp 1679235063
transform 1 0 3588 0 1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_32_29
timestamp 1679235063
transform 1 0 3772 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_41
timestamp 1679235063
transform 1 0 4876 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_32_53
timestamp 1679235063
transform 1 0 5980 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_32_77
timestamp 1679235063
transform 1 0 8188 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_32_81
timestamp 1679235063
transform 1 0 8556 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_32_85
timestamp 1679235063
transform 1 0 8924 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_32_107
timestamp 1679235063
transform 1 0 10948 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_32_111
timestamp 1679235063
transform 1 0 11316 0 1 19584
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_32_126
timestamp 1679235063
transform 1 0 12696 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_32_138
timestamp 1679235063
transform 1 0 13800 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_32_141
timestamp 1679235063
transform 1 0 14076 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_32_163
timestamp 1679235063
transform 1 0 16100 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_32_167
timestamp 1679235063
transform 1 0 16468 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_32_172
timestamp 1679235063
transform 1 0 16928 0 1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_32_187
timestamp 1679235063
transform 1 0 18308 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_32_194
timestamp 1679235063
transform 1 0 18952 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_32_197
timestamp 1679235063
transform 1 0 19228 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_32_202
timestamp 1679235063
transform 1 0 19688 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_32_224
timestamp 1679235063
transform 1 0 21712 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_32_248
timestamp 1679235063
transform 1 0 23920 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_32_253
timestamp 1679235063
transform 1 0 24380 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_32_263
timestamp 1679235063
transform 1 0 25300 0 1 19584
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_33_3
timestamp 1679235063
transform 1 0 1380 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_15
timestamp 1679235063
transform 1 0 2484 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_27
timestamp 1679235063
transform 1 0 3588 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_39
timestamp 1679235063
transform 1 0 4692 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_33_51
timestamp 1679235063
transform 1 0 5796 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_33_55
timestamp 1679235063
transform 1 0 6164 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_33_57
timestamp 1679235063
transform 1 0 6348 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_33_69
timestamp 1679235063
transform 1 0 7452 0 -1 20672
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_33_84
timestamp 1679235063
transform 1 0 8832 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_96
timestamp 1679235063
transform 1 0 9936 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_33_108
timestamp 1679235063
transform 1 0 11040 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_33_113
timestamp 1679235063
transform 1 0 11500 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_33_123
timestamp 1679235063
transform 1 0 12420 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_33_147
timestamp 1679235063
transform 1 0 14628 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_33_160
timestamp 1679235063
transform 1 0 15824 0 -1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_33_169
timestamp 1679235063
transform 1 0 16652 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_33_191
timestamp 1679235063
transform 1 0 18676 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_33_198
timestamp 1679235063
transform 1 0 19320 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_33_204
timestamp 1679235063
transform 1 0 19872 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_33_222
timestamp 1679235063
transform 1 0 21528 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_33_229
timestamp 1679235063
transform 1 0 22172 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_33_240
timestamp 1679235063
transform 1 0 23184 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_33_264
timestamp 1679235063
transform 1 0 25392 0 -1 20672
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_34_3
timestamp 1679235063
transform 1 0 1380 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_15
timestamp 1679235063
transform 1 0 2484 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_34_27
timestamp 1679235063
transform 1 0 3588 0 1 20672
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_34_29
timestamp 1679235063
transform 1 0 3772 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_41
timestamp 1679235063
transform 1 0 4876 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_53
timestamp 1679235063
transform 1 0 5980 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_34_65
timestamp 1679235063
transform 1 0 7084 0 1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_34_73
timestamp 1679235063
transform 1 0 7820 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_34_82
timestamp 1679235063
transform 1 0 8648 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_34_85
timestamp 1679235063
transform 1 0 8924 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_34_91
timestamp 1679235063
transform 1 0 9476 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_34_102
timestamp 1679235063
transform 1 0 10488 0 1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_34_108
timestamp 1679235063
transform 1 0 11040 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_34_129
timestamp 1679235063
transform 1 0 12972 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_34_136
timestamp 1679235063
transform 1 0 13616 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_34_141
timestamp 1679235063
transform 1 0 14076 0 1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_34_151
timestamp 1679235063
transform 1 0 14996 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_34_173
timestamp 1679235063
transform 1 0 17020 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_34_187
timestamp 1679235063
transform 1 0 18308 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_34_194
timestamp 1679235063
transform 1 0 18952 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_34_197
timestamp 1679235063
transform 1 0 19228 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_34_208
timestamp 1679235063
transform 1 0 20240 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_34_221
timestamp 1679235063
transform 1 0 21436 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_34_225
timestamp 1679235063
transform 1 0 21804 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_34_230
timestamp 1679235063
transform 1 0 22264 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_34_250
timestamp 1679235063
transform 1 0 24104 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_34_253
timestamp 1679235063
transform 1 0 24380 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_34_264
timestamp 1679235063
transform 1 0 25392 0 1 20672
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_35_3
timestamp 1679235063
transform 1 0 1380 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_15
timestamp 1679235063
transform 1 0 2484 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_27
timestamp 1679235063
transform 1 0 3588 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_39
timestamp 1679235063
transform 1 0 4692 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_35_51
timestamp 1679235063
transform 1 0 5796 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_35_55
timestamp 1679235063
transform 1 0 6164 0 -1 21760
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_35_57
timestamp 1679235063
transform 1 0 6348 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_35_69
timestamp 1679235063
transform 1 0 7452 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_35_93
timestamp 1679235063
transform 1 0 9660 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_35_97
timestamp 1679235063
transform 1 0 10028 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_35_109
timestamp 1679235063
transform 1 0 11132 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_35_113
timestamp 1679235063
transform 1 0 11500 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_35_123
timestamp 1679235063
transform 1 0 12420 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_35_147
timestamp 1679235063
transform 1 0 14628 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_35_159
timestamp 1679235063
transform 1 0 15732 0 -1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_35_167
timestamp 1679235063
transform 1 0 16468 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_35_169
timestamp 1679235063
transform 1 0 16652 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_35_179
timestamp 1679235063
transform 1 0 17572 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_35_183
timestamp 1679235063
transform 1 0 17940 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_35_189
timestamp 1679235063
transform 1 0 18492 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_35_202
timestamp 1679235063
transform 1 0 19688 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_35_222
timestamp 1679235063
transform 1 0 21528 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_35_225
timestamp 1679235063
transform 1 0 21804 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_35_236
timestamp 1679235063
transform 1 0 22816 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_35_240
timestamp 1679235063
transform 1 0 23184 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_35_261
timestamp 1679235063
transform 1 0 25116 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_35_265
timestamp 1679235063
transform 1 0 25484 0 -1 21760
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_36_3
timestamp 1679235063
transform 1 0 1380 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_15
timestamp 1679235063
transform 1 0 2484 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_36_27
timestamp 1679235063
transform 1 0 3588 0 1 21760
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_36_29
timestamp 1679235063
transform 1 0 3772 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_41
timestamp 1679235063
transform 1 0 4876 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_36_53
timestamp 1679235063
transform 1 0 5980 0 1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_36_61
timestamp 1679235063
transform 1 0 6716 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_36_82
timestamp 1679235063
transform 1 0 8648 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_36_87
timestamp 1679235063
transform 1 0 9108 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_36_94
timestamp 1679235063
transform 1 0 9752 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_36_107
timestamp 1679235063
transform 1 0 10948 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_36_120
timestamp 1679235063
transform 1 0 12144 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_36_133
timestamp 1679235063
transform 1 0 13340 0 1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_36_139
timestamp 1679235063
transform 1 0 13892 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_36_141
timestamp 1679235063
transform 1 0 14076 0 1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_36_149
timestamp 1679235063
transform 1 0 14812 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_36_159
timestamp 1679235063
transform 1 0 15732 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_36_183
timestamp 1679235063
transform 1 0 17940 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_36_189
timestamp 1679235063
transform 1 0 18492 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_36_194
timestamp 1679235063
transform 1 0 18952 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_36_199
timestamp 1679235063
transform 1 0 19412 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_36_211
timestamp 1679235063
transform 1 0 20516 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_36_218
timestamp 1679235063
transform 1 0 21160 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_36_242
timestamp 1679235063
transform 1 0 23368 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_36_246
timestamp 1679235063
transform 1 0 23736 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_36_250
timestamp 1679235063
transform 1 0 24104 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_36_253
timestamp 1679235063
transform 1 0 24380 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_36_264
timestamp 1679235063
transform 1 0 25392 0 1 21760
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_37_3
timestamp 1679235063
transform 1 0 1380 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_15
timestamp 1679235063
transform 1 0 2484 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_27
timestamp 1679235063
transform 1 0 3588 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_39
timestamp 1679235063
transform 1 0 4692 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_37_51
timestamp 1679235063
transform 1 0 5796 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_37_55
timestamp 1679235063
transform 1 0 6164 0 -1 22848
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_37_57
timestamp 1679235063
transform 1 0 6348 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_37_69
timestamp 1679235063
transform 1 0 7452 0 -1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_37_97
timestamp 1679235063
transform 1 0 10028 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_37_101
timestamp 1679235063
transform 1 0 10396 0 -1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_37_109
timestamp 1679235063
transform 1 0 11132 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_37_113
timestamp 1679235063
transform 1 0 11500 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_37_125
timestamp 1679235063
transform 1 0 12604 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_37_129
timestamp 1679235063
transform 1 0 12972 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_37_133
timestamp 1679235063
transform 1 0 13340 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_37_154
timestamp 1679235063
transform 1 0 15272 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_37_162
timestamp 1679235063
transform 1 0 16008 0 -1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_37_169
timestamp 1679235063
transform 1 0 16652 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_37_174
timestamp 1679235063
transform 1 0 17112 0 -1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_37_182
timestamp 1679235063
transform 1 0 17848 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_37_195
timestamp 1679235063
transform 1 0 19044 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_37_201
timestamp 1679235063
transform 1 0 19596 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_37_208
timestamp 1679235063
transform 1 0 20240 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_37_212
timestamp 1679235063
transform 1 0 20608 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_37_222
timestamp 1679235063
transform 1 0 21528 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_37_225
timestamp 1679235063
transform 1 0 21804 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_37_244
timestamp 1679235063
transform 1 0 23552 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_37_264
timestamp 1679235063
transform 1 0 25392 0 -1 22848
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_38_3
timestamp 1679235063
transform 1 0 1380 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_15
timestamp 1679235063
transform 1 0 2484 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_38_27
timestamp 1679235063
transform 1 0 3588 0 1 22848
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_38_29
timestamp 1679235063
transform 1 0 3772 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_41
timestamp 1679235063
transform 1 0 4876 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_53
timestamp 1679235063
transform 1 0 5980 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_65
timestamp 1679235063
transform 1 0 7084 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_38_77
timestamp 1679235063
transform 1 0 8188 0 1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_38_83
timestamp 1679235063
transform 1 0 8740 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_38_85
timestamp 1679235063
transform 1 0 8924 0 1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_38_99
timestamp 1679235063
transform 1 0 10212 0 1 22848
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_38_111
timestamp 1679235063
transform 1 0 11316 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_38_123
timestamp 1679235063
transform 1 0 12420 0 1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_38_138
timestamp 1679235063
transform 1 0 13800 0 1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_38_145
timestamp 1679235063
transform 1 0 14444 0 1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_38_153
timestamp 1679235063
transform 1 0 15180 0 1 22848
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_38_156
timestamp 1679235063
transform 1 0 15456 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_168
timestamp 1679235063
transform 1 0 16560 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_38_180
timestamp 1679235063
transform 1 0 17664 0 1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_38_191
timestamp 1679235063
transform 1 0 18676 0 1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_38_195
timestamp 1679235063
transform 1 0 19044 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_38_197
timestamp 1679235063
transform 1 0 19228 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_38_209
timestamp 1679235063
transform 1 0 20332 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_38_213
timestamp 1679235063
transform 1 0 20700 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_38_217
timestamp 1679235063
transform 1 0 21068 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_38_221
timestamp 1679235063
transform 1 0 21436 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_38_230
timestamp 1679235063
transform 1 0 22264 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_38_250
timestamp 1679235063
transform 1 0 24104 0 1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_38_253
timestamp 1679235063
transform 1 0 24380 0 1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_38_264
timestamp 1679235063
transform 1 0 25392 0 1 22848
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_39_3
timestamp 1679235063
transform 1 0 1380 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_15
timestamp 1679235063
transform 1 0 2484 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_27
timestamp 1679235063
transform 1 0 3588 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_39
timestamp 1679235063
transform 1 0 4692 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_39_51
timestamp 1679235063
transform 1 0 5796 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_39_55
timestamp 1679235063
transform 1 0 6164 0 -1 23936
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_39_57
timestamp 1679235063
transform 1 0 6348 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_69
timestamp 1679235063
transform 1 0 7452 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_39_101
timestamp 1679235063
transform 1 0 10396 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_39_105
timestamp 1679235063
transform 1 0 10764 0 -1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_39_111
timestamp 1679235063
transform 1 0 11316 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_39_113
timestamp 1679235063
transform 1 0 11500 0 -1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_39_121
timestamp 1679235063
transform 1 0 12236 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_39_125
timestamp 1679235063
transform 1 0 12604 0 -1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_39_133
timestamp 1679235063
transform 1 0 13340 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_39_143
timestamp 1679235063
transform 1 0 14260 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_39_156
timestamp 1679235063
transform 1 0 15456 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_39_163
timestamp 1679235063
transform 1 0 16100 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_39_167
timestamp 1679235063
transform 1 0 16468 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_39_169
timestamp 1679235063
transform 1 0 16652 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_39_180
timestamp 1679235063
transform 1 0 17664 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_39_187
timestamp 1679235063
transform 1 0 18308 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_39_195
timestamp 1679235063
transform 1 0 19044 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_39_206
timestamp 1679235063
transform 1 0 20056 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_39_219
timestamp 1679235063
transform 1 0 21252 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_39_223
timestamp 1679235063
transform 1 0 21620 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_39_225
timestamp 1679235063
transform 1 0 21804 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_39_235
timestamp 1679235063
transform 1 0 22724 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_39_239
timestamp 1679235063
transform 1 0 23092 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_39_260
timestamp 1679235063
transform 1 0 25024 0 -1 23936
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_40_3
timestamp 1679235063
transform 1 0 1380 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_15
timestamp 1679235063
transform 1 0 2484 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_40_27
timestamp 1679235063
transform 1 0 3588 0 1 23936
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_40_29
timestamp 1679235063
transform 1 0 3772 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_41
timestamp 1679235063
transform 1 0 4876 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_40_53
timestamp 1679235063
transform 1 0 5980 0 1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_40_61
timestamp 1679235063
transform 1 0 6716 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_40_82
timestamp 1679235063
transform 1 0 8648 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_40_89
timestamp 1679235063
transform 1 0 9292 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_40_99
timestamp 1679235063
transform 1 0 10212 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_40_123
timestamp 1679235063
transform 1 0 12420 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_40_135
timestamp 1679235063
transform 1 0 13524 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_40_139
timestamp 1679235063
transform 1 0 13892 0 1 23936
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_40_141
timestamp 1679235063
transform 1 0 14076 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_40_153
timestamp 1679235063
transform 1 0 15180 0 1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_40_161
timestamp 1679235063
transform 1 0 15916 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_40_168
timestamp 1679235063
transform 1 0 16560 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_40_174
timestamp 1679235063
transform 1 0 17112 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_40_181
timestamp 1679235063
transform 1 0 17756 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_40_194
timestamp 1679235063
transform 1 0 18952 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_40_197
timestamp 1679235063
transform 1 0 19228 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_40_219
timestamp 1679235063
transform 1 0 21252 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_40_223
timestamp 1679235063
transform 1 0 21620 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_40_246
timestamp 1679235063
transform 1 0 23736 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_40_253
timestamp 1679235063
transform 1 0 24380 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_40_263
timestamp 1679235063
transform 1 0 25300 0 1 23936
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_41_3
timestamp 1679235063
transform 1 0 1380 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_15
timestamp 1679235063
transform 1 0 2484 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_27
timestamp 1679235063
transform 1 0 3588 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_39
timestamp 1679235063
transform 1 0 4692 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_41_51
timestamp 1679235063
transform 1 0 5796 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_41_55
timestamp 1679235063
transform 1 0 6164 0 -1 25024
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_41_57
timestamp 1679235063
transform 1 0 6348 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_41_69
timestamp 1679235063
transform 1 0 7452 0 -1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_41_84
timestamp 1679235063
transform 1 0 8832 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_41_108
timestamp 1679235063
transform 1 0 11040 0 -1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_41_113
timestamp 1679235063
transform 1 0 11500 0 -1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_41_135
timestamp 1679235063
transform 1 0 13524 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_41_148
timestamp 1679235063
transform 1 0 14720 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_41_152
timestamp 1679235063
transform 1 0 15088 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_41_155
timestamp 1679235063
transform 1 0 15364 0 -1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_41_166
timestamp 1679235063
transform 1 0 16376 0 -1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_41_169
timestamp 1679235063
transform 1 0 16652 0 -1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_41_180
timestamp 1679235063
transform 1 0 17664 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_41_193
timestamp 1679235063
transform 1 0 18860 0 -1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_41_199
timestamp 1679235063
transform 1 0 19412 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_41_222
timestamp 1679235063
transform 1 0 21528 0 -1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_41_225
timestamp 1679235063
transform 1 0 21804 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_41_237
timestamp 1679235063
transform 1 0 22908 0 -1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_41_241
timestamp 1679235063
transform 1 0 23276 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_41_264
timestamp 1679235063
transform 1 0 25392 0 -1 25024
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_42_3
timestamp 1679235063
transform 1 0 1380 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_15
timestamp 1679235063
transform 1 0 2484 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_42_27
timestamp 1679235063
transform 1 0 3588 0 1 25024
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_42_29
timestamp 1679235063
transform 1 0 3772 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_41
timestamp 1679235063
transform 1 0 4876 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_53
timestamp 1679235063
transform 1 0 5980 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_65
timestamp 1679235063
transform 1 0 7084 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_42_77
timestamp 1679235063
transform 1 0 8188 0 1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_42_83
timestamp 1679235063
transform 1 0 8740 0 1 25024
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_42_85
timestamp 1679235063
transform 1 0 8924 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_42_97
timestamp 1679235063
transform 1 0 10028 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_42_109
timestamp 1679235063
transform 1 0 11132 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_42_122
timestamp 1679235063
transform 1 0 12328 0 1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_42_138
timestamp 1679235063
transform 1 0 13800 0 1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_42_141
timestamp 1679235063
transform 1 0 14076 0 1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_42_152
timestamp 1679235063
transform 1 0 15088 0 1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_42_156
timestamp 1679235063
transform 1 0 15456 0 1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_42_178
timestamp 1679235063
transform 1 0 17480 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_42_185
timestamp 1679235063
transform 1 0 18124 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_42_189
timestamp 1679235063
transform 1 0 18492 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_42_194
timestamp 1679235063
transform 1 0 18952 0 1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_42_199
timestamp 1679235063
transform 1 0 19412 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_42_210
timestamp 1679235063
transform 1 0 20424 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_42_218
timestamp 1679235063
transform 1 0 21160 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_42_230
timestamp 1679235063
transform 1 0 22264 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_42_250
timestamp 1679235063
transform 1 0 24104 0 1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_42_253
timestamp 1679235063
transform 1 0 24380 0 1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_42_263
timestamp 1679235063
transform 1 0 25300 0 1 25024
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_43_3
timestamp 1679235063
transform 1 0 1380 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_15
timestamp 1679235063
transform 1 0 2484 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_27
timestamp 1679235063
transform 1 0 3588 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_39
timestamp 1679235063
transform 1 0 4692 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_43_51
timestamp 1679235063
transform 1 0 5796 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_43_55
timestamp 1679235063
transform 1 0 6164 0 -1 26112
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_43_57
timestamp 1679235063
transform 1 0 6348 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_69
timestamp 1679235063
transform 1 0 7452 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_81
timestamp 1679235063
transform 1 0 8556 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_43_93
timestamp 1679235063
transform 1 0 9660 0 -1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_43_101
timestamp 1679235063
transform 1 0 10396 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_43_110
timestamp 1679235063
transform 1 0 11224 0 -1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_43_113
timestamp 1679235063
transform 1 0 11500 0 -1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_43_121
timestamp 1679235063
transform 1 0 12236 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_43_142
timestamp 1679235063
transform 1 0 14168 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_43_155
timestamp 1679235063
transform 1 0 15364 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_43_162
timestamp 1679235063
transform 1 0 16008 0 -1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_43_169
timestamp 1679235063
transform 1 0 16652 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_43_175
timestamp 1679235063
transform 1 0 17204 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_43_182
timestamp 1679235063
transform 1 0 17848 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_43_189
timestamp 1679235063
transform 1 0 18492 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_43_196
timestamp 1679235063
transform 1 0 19136 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_43_208
timestamp 1679235063
transform 1 0 20240 0 -1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_43_212
timestamp 1679235063
transform 1 0 20608 0 -1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_43_222
timestamp 1679235063
transform 1 0 21528 0 -1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_43_225
timestamp 1679235063
transform 1 0 21804 0 -1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_43_236
timestamp 1679235063
transform 1 0 22816 0 -1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_43_242
timestamp 1679235063
transform 1 0 23368 0 -1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_43_264
timestamp 1679235063
transform 1 0 25392 0 -1 26112
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_44_3
timestamp 1679235063
transform 1 0 1380 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_15
timestamp 1679235063
transform 1 0 2484 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_44_27
timestamp 1679235063
transform 1 0 3588 0 1 26112
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_44_29
timestamp 1679235063
transform 1 0 3772 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_41
timestamp 1679235063
transform 1 0 4876 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_53
timestamp 1679235063
transform 1 0 5980 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_65
timestamp 1679235063
transform 1 0 7084 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_44_77
timestamp 1679235063
transform 1 0 8188 0 1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_44_83
timestamp 1679235063
transform 1 0 8740 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_44_85
timestamp 1679235063
transform 1 0 8924 0 1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_44_107
timestamp 1679235063
transform 1 0 10948 0 1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_44_111
timestamp 1679235063
transform 1 0 11316 0 1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_44_115
timestamp 1679235063
transform 1 0 11684 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_44_125
timestamp 1679235063
transform 1 0 12604 0 1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_44_138
timestamp 1679235063
transform 1 0 13800 0 1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_44_143
timestamp 1679235063
transform 1 0 14260 0 1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_44_154
timestamp 1679235063
transform 1 0 15272 0 1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_44_167
timestamp 1679235063
transform 1 0 16468 0 1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_44_173
timestamp 1679235063
transform 1 0 17020 0 1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_44_181
timestamp 1679235063
transform 1 0 17756 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_44_191
timestamp 1679235063
transform 1 0 18676 0 1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_44_195
timestamp 1679235063
transform 1 0 19044 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_44_197
timestamp 1679235063
transform 1 0 19228 0 1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_44_219
timestamp 1679235063
transform 1 0 21252 0 1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_44_223
timestamp 1679235063
transform 1 0 21620 0 1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_44_229
timestamp 1679235063
transform 1 0 22172 0 1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_44_233
timestamp 1679235063
transform 1 0 22540 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_44_243
timestamp 1679235063
transform 1 0 23460 0 1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_44_250
timestamp 1679235063
transform 1 0 24104 0 1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_44_253
timestamp 1679235063
transform 1 0 24380 0 1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_44_264
timestamp 1679235063
transform 1 0 25392 0 1 26112
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_45_3
timestamp 1679235063
transform 1 0 1380 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_15
timestamp 1679235063
transform 1 0 2484 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_27
timestamp 1679235063
transform 1 0 3588 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_39
timestamp 1679235063
transform 1 0 4692 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_45_51
timestamp 1679235063
transform 1 0 5796 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_45_55
timestamp 1679235063
transform 1 0 6164 0 -1 27200
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_45_57
timestamp 1679235063
transform 1 0 6348 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_69
timestamp 1679235063
transform 1 0 7452 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_45_81
timestamp 1679235063
transform 1 0 8556 0 -1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_45_89
timestamp 1679235063
transform 1 0 9292 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_45_110
timestamp 1679235063
transform 1 0 11224 0 -1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_45_115
timestamp 1679235063
transform 1 0 11684 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_45_121
timestamp 1679235063
transform 1 0 12236 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_45_125
timestamp 1679235063
transform 1 0 12604 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_45_146
timestamp 1679235063
transform 1 0 14536 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_45_150
timestamp 1679235063
transform 1 0 14904 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_45_160
timestamp 1679235063
transform 1 0 15824 0 -1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_45_166
timestamp 1679235063
transform 1 0 16376 0 -1 27200
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_45_169
timestamp 1679235063
transform 1 0 16652 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_45_181
timestamp 1679235063
transform 1 0 17756 0 -1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_45_203
timestamp 1679235063
transform 1 0 19780 0 -1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_45_207
timestamp 1679235063
transform 1 0 20148 0 -1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_45_211
timestamp 1679235063
transform 1 0 20516 0 -1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_45_222
timestamp 1679235063
transform 1 0 21528 0 -1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_45_225
timestamp 1679235063
transform 1 0 21804 0 -1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_45_235
timestamp 1679235063
transform 1 0 22724 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_45_239
timestamp 1679235063
transform 1 0 23092 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_45_260
timestamp 1679235063
transform 1 0 25024 0 -1 27200
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_46_3
timestamp 1679235063
transform 1 0 1380 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_15
timestamp 1679235063
transform 1 0 2484 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_46_27
timestamp 1679235063
transform 1 0 3588 0 1 27200
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_46_29
timestamp 1679235063
transform 1 0 3772 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_41
timestamp 1679235063
transform 1 0 4876 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_53
timestamp 1679235063
transform 1 0 5980 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_65
timestamp 1679235063
transform 1 0 7084 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_46_77
timestamp 1679235063
transform 1 0 8188 0 1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_46_83
timestamp 1679235063
transform 1 0 8740 0 1 27200
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_46_85
timestamp 1679235063
transform 1 0 8924 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_46_97
timestamp 1679235063
transform 1 0 10028 0 1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_46_119
timestamp 1679235063
transform 1 0 12052 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_46_131
timestamp 1679235063
transform 1 0 13156 0 1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_46_139
timestamp 1679235063
transform 1 0 13892 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_46_141
timestamp 1679235063
transform 1 0 14076 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_46_145
timestamp 1679235063
transform 1 0 14444 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_46_148
timestamp 1679235063
transform 1 0 14720 0 1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_46_165
timestamp 1679235063
transform 1 0 16284 0 1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_46_169
timestamp 1679235063
transform 1 0 16652 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_46_182
timestamp 1679235063
transform 1 0 17848 0 1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_46_187
timestamp 1679235063
transform 1 0 18308 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_46_194
timestamp 1679235063
transform 1 0 18952 0 1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_46_199
timestamp 1679235063
transform 1 0 19412 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_46_203
timestamp 1679235063
transform 1 0 19780 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_46_224
timestamp 1679235063
transform 1 0 21712 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_46_237
timestamp 1679235063
transform 1 0 22908 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_46_250
timestamp 1679235063
transform 1 0 24104 0 1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_46_253
timestamp 1679235063
transform 1 0 24380 0 1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_46_263
timestamp 1679235063
transform 1 0 25300 0 1 27200
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_47_3
timestamp 1679235063
transform 1 0 1380 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_15
timestamp 1679235063
transform 1 0 2484 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_27
timestamp 1679235063
transform 1 0 3588 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_39
timestamp 1679235063
transform 1 0 4692 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_47_51
timestamp 1679235063
transform 1 0 5796 0 -1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_47_55
timestamp 1679235063
transform 1 0 6164 0 -1 28288
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_47_57
timestamp 1679235063
transform 1 0 6348 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_69
timestamp 1679235063
transform 1 0 7452 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_81
timestamp 1679235063
transform 1 0 8556 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_47_93
timestamp 1679235063
transform 1 0 9660 0 -1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_47_101
timestamp 1679235063
transform 1 0 10396 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_47_110
timestamp 1679235063
transform 1 0 11224 0 -1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_47_113
timestamp 1679235063
transform 1 0 11500 0 -1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_47_123
timestamp 1679235063
transform 1 0 12420 0 -1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_47_127
timestamp 1679235063
transform 1 0 12788 0 -1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_47_140
timestamp 1679235063
transform 1 0 13984 0 -1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_47_152
timestamp 1679235063
transform 1 0 15088 0 -1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_47_164
timestamp 1679235063
transform 1 0 16192 0 -1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_47_169
timestamp 1679235063
transform 1 0 16652 0 -1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_47_180
timestamp 1679235063
transform 1 0 17664 0 -1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_47_193
timestamp 1679235063
transform 1 0 18860 0 -1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_47_205
timestamp 1679235063
transform 1 0 19964 0 -1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_47_209
timestamp 1679235063
transform 1 0 20332 0 -1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_47_222
timestamp 1679235063
transform 1 0 21528 0 -1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_47_225
timestamp 1679235063
transform 1 0 21804 0 -1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_47_247
timestamp 1679235063
transform 1 0 23828 0 -1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_47_260
timestamp 1679235063
transform 1 0 25024 0 -1 28288
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_48_3
timestamp 1679235063
transform 1 0 1380 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_15
timestamp 1679235063
transform 1 0 2484 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_48_27
timestamp 1679235063
transform 1 0 3588 0 1 28288
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_48_29
timestamp 1679235063
transform 1 0 3772 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_41
timestamp 1679235063
transform 1 0 4876 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_53
timestamp 1679235063
transform 1 0 5980 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_65
timestamp 1679235063
transform 1 0 7084 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_48_77
timestamp 1679235063
transform 1 0 8188 0 1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_48_83
timestamp 1679235063
transform 1 0 8740 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_48_85
timestamp 1679235063
transform 1 0 8924 0 1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_48_111
timestamp 1679235063
transform 1 0 11316 0 1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_48_135
timestamp 1679235063
transform 1 0 13524 0 1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_48_143
timestamp 1679235063
transform 1 0 14260 0 1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_48_147
timestamp 1679235063
transform 1 0 14628 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_48_157
timestamp 1679235063
transform 1 0 15548 0 1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_48_170
timestamp 1679235063
transform 1 0 16744 0 1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_48_194
timestamp 1679235063
transform 1 0 18952 0 1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_48_197
timestamp 1679235063
transform 1 0 19228 0 1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_48_208
timestamp 1679235063
transform 1 0 20240 0 1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_48_232
timestamp 1679235063
transform 1 0 22448 0 1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_48_247
timestamp 1679235063
transform 1 0 23828 0 1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_48_251
timestamp 1679235063
transform 1 0 24196 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_48_253
timestamp 1679235063
transform 1 0 24380 0 1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_48_264
timestamp 1679235063
transform 1 0 25392 0 1 28288
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_49_3
timestamp 1679235063
transform 1 0 1380 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_15
timestamp 1679235063
transform 1 0 2484 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_27
timestamp 1679235063
transform 1 0 3588 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_39
timestamp 1679235063
transform 1 0 4692 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_49_51
timestamp 1679235063
transform 1 0 5796 0 -1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_49_55
timestamp 1679235063
transform 1 0 6164 0 -1 29376
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_49_57
timestamp 1679235063
transform 1 0 6348 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_69
timestamp 1679235063
transform 1 0 7452 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_81
timestamp 1679235063
transform 1 0 8556 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_49_93
timestamp 1679235063
transform 1 0 9660 0 -1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_49_101
timestamp 1679235063
transform 1 0 10396 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_49_110
timestamp 1679235063
transform 1 0 11224 0 -1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_49_115
timestamp 1679235063
transform 1 0 11684 0 -1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_49_125
timestamp 1679235063
transform 1 0 12604 0 -1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_49_138
timestamp 1679235063
transform 1 0 13800 0 -1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_49_151
timestamp 1679235063
transform 1 0 14996 0 -1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_49_164
timestamp 1679235063
transform 1 0 16192 0 -1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_49_169
timestamp 1679235063
transform 1 0 16652 0 -1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_49_180
timestamp 1679235063
transform 1 0 17664 0 -1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_49_186
timestamp 1679235063
transform 1 0 18216 0 -1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_49_190
timestamp 1679235063
transform 1 0 18584 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_49_195
timestamp 1679235063
transform 1 0 19044 0 -1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_49_200
timestamp 1679235063
transform 1 0 19504 0 -1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_49_207
timestamp 1679235063
transform 1 0 20148 0 -1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_49_212
timestamp 1679235063
transform 1 0 20608 0 -1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_49_220
timestamp 1679235063
transform 1 0 21344 0 -1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_49_225
timestamp 1679235063
transform 1 0 21804 0 -1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_49_235
timestamp 1679235063
transform 1 0 22724 0 -1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_49_248
timestamp 1679235063
transform 1 0 23920 0 -1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_49_255
timestamp 1679235063
transform 1 0 24564 0 -1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_49_259
timestamp 1679235063
transform 1 0 24932 0 -1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_49_264
timestamp 1679235063
transform 1 0 25392 0 -1 29376
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_50_3
timestamp 1679235063
transform 1 0 1380 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_15
timestamp 1679235063
transform 1 0 2484 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_50_27
timestamp 1679235063
transform 1 0 3588 0 1 29376
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_50_29
timestamp 1679235063
transform 1 0 3772 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_41
timestamp 1679235063
transform 1 0 4876 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_53
timestamp 1679235063
transform 1 0 5980 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_65
timestamp 1679235063
transform 1 0 7084 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_50_77
timestamp 1679235063
transform 1 0 8188 0 1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_50_83
timestamp 1679235063
transform 1 0 8740 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_50_85
timestamp 1679235063
transform 1 0 8924 0 1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_50_107
timestamp 1679235063
transform 1 0 10948 0 1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_50_111
timestamp 1679235063
transform 1 0 11316 0 1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_50_133
timestamp 1679235063
transform 1 0 13340 0 1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_50_137
timestamp 1679235063
transform 1 0 13708 0 1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_50_141
timestamp 1679235063
transform 1 0 14076 0 1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_50_163
timestamp 1679235063
transform 1 0 16100 0 1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_50_169
timestamp 1679235063
transform 1 0 16652 0 1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_50_173
timestamp 1679235063
transform 1 0 17020 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_50_194
timestamp 1679235063
transform 1 0 18952 0 1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_50_197
timestamp 1679235063
transform 1 0 19228 0 1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_50_208
timestamp 1679235063
transform 1 0 20240 0 1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_50_221
timestamp 1679235063
transform 1 0 21436 0 1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_50_231
timestamp 1679235063
transform 1 0 22356 0 1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_50_236
timestamp 1679235063
transform 1 0 22816 0 1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_50_243
timestamp 1679235063
transform 1 0 23460 0 1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_50_250
timestamp 1679235063
transform 1 0 24104 0 1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_50_259
timestamp 1679235063
transform 1 0 24932 0 1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_50_264
timestamp 1679235063
transform 1 0 25392 0 1 29376
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_51_3
timestamp 1679235063
transform 1 0 1380 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_15
timestamp 1679235063
transform 1 0 2484 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_27
timestamp 1679235063
transform 1 0 3588 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_39
timestamp 1679235063
transform 1 0 4692 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_51_51
timestamp 1679235063
transform 1 0 5796 0 -1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_51_55
timestamp 1679235063
transform 1 0 6164 0 -1 30464
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_51_57
timestamp 1679235063
transform 1 0 6348 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_69
timestamp 1679235063
transform 1 0 7452 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_81
timestamp 1679235063
transform 1 0 8556 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_51_102
timestamp 1679235063
transform 1 0 10488 0 -1 30464
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_51_110
timestamp 1679235063
transform 1 0 11224 0 -1 30464
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_51_113
timestamp 1679235063
transform 1 0 11500 0 -1 30464
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_51_141
timestamp 1679235063
transform 1 0 14076 0 -1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_51_153
timestamp 1679235063
transform 1 0 15180 0 -1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_51_166
timestamp 1679235063
transform 1 0 16376 0 -1 30464
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_51_173
timestamp 1679235063
transform 1 0 17020 0 -1 30464
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_51_184
timestamp 1679235063
transform 1 0 18032 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_51_196
timestamp 1679235063
transform 1 0 19136 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_51_200
timestamp 1679235063
transform 1 0 19504 0 -1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_51_213
timestamp 1679235063
transform 1 0 20700 0 -1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_51_222
timestamp 1679235063
transform 1 0 21528 0 -1 30464
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_51_225
timestamp 1679235063
transform 1 0 21804 0 -1 30464
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_51_236
timestamp 1679235063
transform 1 0 22816 0 -1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_51_240
timestamp 1679235063
transform 1 0 23184 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_51_261
timestamp 1679235063
transform 1 0 25116 0 -1 30464
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_51_265
timestamp 1679235063
transform 1 0 25484 0 -1 30464
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_52_3
timestamp 1679235063
transform 1 0 1380 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_15
timestamp 1679235063
transform 1 0 2484 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_52_27
timestamp 1679235063
transform 1 0 3588 0 1 30464
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_52_29
timestamp 1679235063
transform 1 0 3772 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_41
timestamp 1679235063
transform 1 0 4876 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_53
timestamp 1679235063
transform 1 0 5980 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_65
timestamp 1679235063
transform 1 0 7084 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_52_77
timestamp 1679235063
transform 1 0 8188 0 1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_52_83
timestamp 1679235063
transform 1 0 8740 0 1 30464
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_52_85
timestamp 1679235063
transform 1 0 8924 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_97
timestamp 1679235063
transform 1 0 10028 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_109
timestamp 1679235063
transform 1 0 11132 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_121
timestamp 1679235063
transform 1 0 12236 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_52_133
timestamp 1679235063
transform 1 0 13340 0 1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_52_139
timestamp 1679235063
transform 1 0 13892 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_52_143
timestamp 1679235063
transform 1 0 14260 0 1 30464
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_52_156
timestamp 1679235063
transform 1 0 15456 0 1 30464
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_52_160
timestamp 1679235063
transform 1 0 15824 0 1 30464
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_52_168
timestamp 1679235063
transform 1 0 16560 0 1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_52_191
timestamp 1679235063
transform 1 0 18676 0 1 30464
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_52_195
timestamp 1679235063
transform 1 0 19044 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_52_197
timestamp 1679235063
transform 1 0 19228 0 1 30464
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_52_207
timestamp 1679235063
transform 1 0 20148 0 1 30464
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_52_211
timestamp 1679235063
transform 1 0 20516 0 1 30464
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_52_233
timestamp 1679235063
transform 1 0 22540 0 1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_52_245
timestamp 1679235063
transform 1 0 23644 0 1 30464
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_52_249
timestamp 1679235063
transform 1 0 24012 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_52_253
timestamp 1679235063
transform 1 0 24380 0 1 30464
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_52_263
timestamp 1679235063
transform 1 0 25300 0 1 30464
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_53_3
timestamp 1679235063
transform 1 0 1380 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_15
timestamp 1679235063
transform 1 0 2484 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_27
timestamp 1679235063
transform 1 0 3588 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_39
timestamp 1679235063
transform 1 0 4692 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_53_51
timestamp 1679235063
transform 1 0 5796 0 -1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_53_55
timestamp 1679235063
transform 1 0 6164 0 -1 31552
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_53_57
timestamp 1679235063
transform 1 0 6348 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_69
timestamp 1679235063
transform 1 0 7452 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_81
timestamp 1679235063
transform 1 0 8556 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_93
timestamp 1679235063
transform 1 0 9660 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_53_105
timestamp 1679235063
transform 1 0 10764 0 -1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_53_111
timestamp 1679235063
transform 1 0 11316 0 -1 31552
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_53_113
timestamp 1679235063
transform 1 0 11500 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_53_125
timestamp 1679235063
transform 1 0 12604 0 -1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_53_131
timestamp 1679235063
transform 1 0 13156 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_53_153
timestamp 1679235063
transform 1 0 15180 0 -1 31552
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_53_159
timestamp 1679235063
transform 1 0 15732 0 -1 31552
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_53_167
timestamp 1679235063
transform 1 0 16468 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_53_171
timestamp 1679235063
transform 1 0 16836 0 -1 31552
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_53_181
timestamp 1679235063
transform 1 0 17756 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_53_193
timestamp 1679235063
transform 1 0 18860 0 -1 31552
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_53_203
timestamp 1679235063
transform 1 0 19780 0 -1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_53_216
timestamp 1679235063
transform 1 0 20976 0 -1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_53_223
timestamp 1679235063
transform 1 0 21620 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_53_225
timestamp 1679235063
transform 1 0 21804 0 -1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_53_231
timestamp 1679235063
transform 1 0 22356 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_53_252
timestamp 1679235063
transform 1 0 24288 0 -1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_53_264
timestamp 1679235063
transform 1 0 25392 0 -1 31552
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_54_3
timestamp 1679235063
transform 1 0 1380 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_15
timestamp 1679235063
transform 1 0 2484 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_54_27
timestamp 1679235063
transform 1 0 3588 0 1 31552
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_54_29
timestamp 1679235063
transform 1 0 3772 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_41
timestamp 1679235063
transform 1 0 4876 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_53
timestamp 1679235063
transform 1 0 5980 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_65
timestamp 1679235063
transform 1 0 7084 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_54_77
timestamp 1679235063
transform 1 0 8188 0 1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_54_83
timestamp 1679235063
transform 1 0 8740 0 1 31552
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_54_85
timestamp 1679235063
transform 1 0 8924 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_97
timestamp 1679235063
transform 1 0 10028 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_109
timestamp 1679235063
transform 1 0 11132 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_121
timestamp 1679235063
transform 1 0 12236 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_54_133
timestamp 1679235063
transform 1 0 13340 0 1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_54_139
timestamp 1679235063
transform 1 0 13892 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_54_141
timestamp 1679235063
transform 1 0 14076 0 1 31552
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_54_154
timestamp 1679235063
transform 1 0 15272 0 1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_54_167
timestamp 1679235063
transform 1 0 16468 0 1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_54_191
timestamp 1679235063
transform 1 0 18676 0 1 31552
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_54_195
timestamp 1679235063
transform 1 0 19044 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_54_197
timestamp 1679235063
transform 1 0 19228 0 1 31552
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_54_219
timestamp 1679235063
transform 1 0 21252 0 1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_54_232
timestamp 1679235063
transform 1 0 22448 0 1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_54_244
timestamp 1679235063
transform 1 0 23552 0 1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_54_253
timestamp 1679235063
transform 1 0 24380 0 1 31552
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_54_263
timestamp 1679235063
transform 1 0 25300 0 1 31552
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_55_3
timestamp 1679235063
transform 1 0 1380 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_15
timestamp 1679235063
transform 1 0 2484 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_27
timestamp 1679235063
transform 1 0 3588 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_39
timestamp 1679235063
transform 1 0 4692 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_55_51
timestamp 1679235063
transform 1 0 5796 0 -1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_55_55
timestamp 1679235063
transform 1 0 6164 0 -1 32640
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_55_57
timestamp 1679235063
transform 1 0 6348 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_69
timestamp 1679235063
transform 1 0 7452 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_55_81
timestamp 1679235063
transform 1 0 8556 0 -1 32640
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_55_88
timestamp 1679235063
transform 1 0 9200 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_100
timestamp 1679235063
transform 1 0 10304 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_113
timestamp 1679235063
transform 1 0 11500 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_125
timestamp 1679235063
transform 1 0 12604 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_137
timestamp 1679235063
transform 1 0 13708 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_55_149
timestamp 1679235063
transform 1 0 14812 0 -1 32640
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_55_166
timestamp 1679235063
transform 1 0 16376 0 -1 32640
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_55_175
timestamp 1679235063
transform 1 0 17204 0 -1 32640
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_55_197
timestamp 1679235063
transform 1 0 19228 0 -1 32640
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_55_201
timestamp 1679235063
transform 1 0 19596 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_55_204
timestamp 1679235063
transform 1 0 19872 0 -1 32640
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_55_217
timestamp 1679235063
transform 1 0 21068 0 -1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_55_221
timestamp 1679235063
transform 1 0 21436 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_55_225
timestamp 1679235063
transform 1 0 21804 0 -1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_55_239
timestamp 1679235063
transform 1 0 23092 0 -1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_55_263
timestamp 1679235063
transform 1 0 25300 0 -1 32640
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_56_3
timestamp 1679235063
transform 1 0 1380 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_15
timestamp 1679235063
transform 1 0 2484 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_56_27
timestamp 1679235063
transform 1 0 3588 0 1 32640
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_56_29
timestamp 1679235063
transform 1 0 3772 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_41
timestamp 1679235063
transform 1 0 4876 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_53
timestamp 1679235063
transform 1 0 5980 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_65
timestamp 1679235063
transform 1 0 7084 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_56_77
timestamp 1679235063
transform 1 0 8188 0 1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_56_83
timestamp 1679235063
transform 1 0 8740 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_56_85
timestamp 1679235063
transform 1 0 8924 0 1 32640
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_56_90
timestamp 1679235063
transform 1 0 9384 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_102
timestamp 1679235063
transform 1 0 10488 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_114
timestamp 1679235063
transform 1 0 11592 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_126
timestamp 1679235063
transform 1 0 12696 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_56_138
timestamp 1679235063
transform 1 0 13800 0 1 32640
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_56_141
timestamp 1679235063
transform 1 0 14076 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_153
timestamp 1679235063
transform 1 0 15180 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_165
timestamp 1679235063
transform 1 0 16284 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_56_177
timestamp 1679235063
transform 1 0 17388 0 1 32640
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_56_193
timestamp 1679235063
transform 1 0 18860 0 1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_56_197
timestamp 1679235063
transform 1 0 19228 0 1 32640
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_56_219
timestamp 1679235063
transform 1 0 21252 0 1 32640
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_56_223
timestamp 1679235063
transform 1 0 21620 0 1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_56_229
timestamp 1679235063
transform 1 0 22172 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_56_250
timestamp 1679235063
transform 1 0 24104 0 1 32640
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_56_253
timestamp 1679235063
transform 1 0 24380 0 1 32640
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_56_264
timestamp 1679235063
transform 1 0 25392 0 1 32640
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_57_3
timestamp 1679235063
transform 1 0 1380 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_15
timestamp 1679235063
transform 1 0 2484 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_27
timestamp 1679235063
transform 1 0 3588 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_39
timestamp 1679235063
transform 1 0 4692 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_57_51
timestamp 1679235063
transform 1 0 5796 0 -1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_57_55
timestamp 1679235063
transform 1 0 6164 0 -1 33728
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_57_57
timestamp 1679235063
transform 1 0 6348 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_69
timestamp 1679235063
transform 1 0 7452 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_57_81
timestamp 1679235063
transform 1 0 8556 0 -1 33728
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_57_89
timestamp 1679235063
transform 1 0 9292 0 -1 33728
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_57_98
timestamp 1679235063
transform 1 0 10120 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_57_110
timestamp 1679235063
transform 1 0 11224 0 -1 33728
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_57_113
timestamp 1679235063
transform 1 0 11500 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_125
timestamp 1679235063
transform 1 0 12604 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_137
timestamp 1679235063
transform 1 0 13708 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_149
timestamp 1679235063
transform 1 0 14812 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_57_161
timestamp 1679235063
transform 1 0 15916 0 -1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_57_167
timestamp 1679235063
transform 1 0 16468 0 -1 33728
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_57_169
timestamp 1679235063
transform 1 0 16652 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_181
timestamp 1679235063
transform 1 0 17756 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_57_193
timestamp 1679235063
transform 1 0 18860 0 -1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_57_219
timestamp 1679235063
transform 1 0 21252 0 -1 33728
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_57_223
timestamp 1679235063
transform 1 0 21620 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_57_225
timestamp 1679235063
transform 1 0 21804 0 -1 33728
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_57_247
timestamp 1679235063
transform 1 0 23828 0 -1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_57_260
timestamp 1679235063
transform 1 0 25024 0 -1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_57_265
timestamp 1679235063
transform 1 0 25484 0 -1 33728
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_58_3
timestamp 1679235063
transform 1 0 1380 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_15
timestamp 1679235063
transform 1 0 2484 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_58_27
timestamp 1679235063
transform 1 0 3588 0 1 33728
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_58_29
timestamp 1679235063
transform 1 0 3772 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_41
timestamp 1679235063
transform 1 0 4876 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_53
timestamp 1679235063
transform 1 0 5980 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_65
timestamp 1679235063
transform 1 0 7084 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_58_77
timestamp 1679235063
transform 1 0 8188 0 1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_58_83
timestamp 1679235063
transform 1 0 8740 0 1 33728
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_58_85
timestamp 1679235063
transform 1 0 8924 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_97
timestamp 1679235063
transform 1 0 10028 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_109
timestamp 1679235063
transform 1 0 11132 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_121
timestamp 1679235063
transform 1 0 12236 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_58_133
timestamp 1679235063
transform 1 0 13340 0 1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_58_139
timestamp 1679235063
transform 1 0 13892 0 1 33728
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_58_141
timestamp 1679235063
transform 1 0 14076 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_153
timestamp 1679235063
transform 1 0 15180 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_58_165
timestamp 1679235063
transform 1 0 16284 0 1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_58_173
timestamp 1679235063
transform 1 0 17020 0 1 33728
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_58_186
timestamp 1679235063
transform 1 0 18216 0 1 33728
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_58_194
timestamp 1679235063
transform 1 0 18952 0 1 33728
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_58_197
timestamp 1679235063
transform 1 0 19228 0 1 33728
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_58_219
timestamp 1679235063
transform 1 0 21252 0 1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_58_243
timestamp 1679235063
transform 1 0 23460 0 1 33728
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_58_251
timestamp 1679235063
transform 1 0 24196 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_58_253
timestamp 1679235063
transform 1 0 24380 0 1 33728
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_58_263
timestamp 1679235063
transform 1 0 25300 0 1 33728
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_59_3
timestamp 1679235063
transform 1 0 1380 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_15
timestamp 1679235063
transform 1 0 2484 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_27
timestamp 1679235063
transform 1 0 3588 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_39
timestamp 1679235063
transform 1 0 4692 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_59_51
timestamp 1679235063
transform 1 0 5796 0 -1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_59_55
timestamp 1679235063
transform 1 0 6164 0 -1 34816
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_59_57
timestamp 1679235063
transform 1 0 6348 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_69
timestamp 1679235063
transform 1 0 7452 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_81
timestamp 1679235063
transform 1 0 8556 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_93
timestamp 1679235063
transform 1 0 9660 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_59_105
timestamp 1679235063
transform 1 0 10764 0 -1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_59_111
timestamp 1679235063
transform 1 0 11316 0 -1 34816
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_59_113
timestamp 1679235063
transform 1 0 11500 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_125
timestamp 1679235063
transform 1 0 12604 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_137
timestamp 1679235063
transform 1 0 13708 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_59_149
timestamp 1679235063
transform 1 0 14812 0 -1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_59_163
timestamp 1679235063
transform 1 0 16100 0 -1 34816
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_59_167
timestamp 1679235063
transform 1 0 16468 0 -1 34816
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_59_169
timestamp 1679235063
transform 1 0 16652 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_181
timestamp 1679235063
transform 1 0 17756 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_59_193
timestamp 1679235063
transform 1 0 18860 0 -1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_59_207
timestamp 1679235063
transform 1 0 20148 0 -1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_59_213
timestamp 1679235063
transform 1 0 20700 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_59_222
timestamp 1679235063
transform 1 0 21528 0 -1 34816
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_59_225
timestamp 1679235063
transform 1 0 21804 0 -1 34816
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_59_235
timestamp 1679235063
transform 1 0 22724 0 -1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_59_247
timestamp 1679235063
transform 1 0 23828 0 -1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_59_252
timestamp 1679235063
transform 1 0 24288 0 -1 34816
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_59_257
timestamp 1679235063
transform 1 0 24748 0 -1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_59_264
timestamp 1679235063
transform 1 0 25392 0 -1 34816
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_60_3
timestamp 1679235063
transform 1 0 1380 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_15
timestamp 1679235063
transform 1 0 2484 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_60_27
timestamp 1679235063
transform 1 0 3588 0 1 34816
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_60_29
timestamp 1679235063
transform 1 0 3772 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_41
timestamp 1679235063
transform 1 0 4876 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_53
timestamp 1679235063
transform 1 0 5980 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_65
timestamp 1679235063
transform 1 0 7084 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_60_77
timestamp 1679235063
transform 1 0 8188 0 1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_60_83
timestamp 1679235063
transform 1 0 8740 0 1 34816
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_60_85
timestamp 1679235063
transform 1 0 8924 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_97
timestamp 1679235063
transform 1 0 10028 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_109
timestamp 1679235063
transform 1 0 11132 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_121
timestamp 1679235063
transform 1 0 12236 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_60_133
timestamp 1679235063
transform 1 0 13340 0 1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_60_139
timestamp 1679235063
transform 1 0 13892 0 1 34816
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_60_141
timestamp 1679235063
transform 1 0 14076 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_153
timestamp 1679235063
transform 1 0 15180 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_165
timestamp 1679235063
transform 1 0 16284 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_177
timestamp 1679235063
transform 1 0 17388 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_60_189
timestamp 1679235063
transform 1 0 18492 0 1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_60_195
timestamp 1679235063
transform 1 0 19044 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_60_197
timestamp 1679235063
transform 1 0 19228 0 1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_60_209
timestamp 1679235063
transform 1 0 20332 0 1 34816
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_60_217
timestamp 1679235063
transform 1 0 21068 0 1 34816
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_60_221
timestamp 1679235063
transform 1 0 21436 0 1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_60_227
timestamp 1679235063
transform 1 0 21988 0 1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_60_233
timestamp 1679235063
transform 1 0 22540 0 1 34816
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_60_244
timestamp 1679235063
transform 1 0 23552 0 1 34816
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_60_259
timestamp 1679235063
transform 1 0 24932 0 1 34816
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_60_264
timestamp 1679235063
transform 1 0 25392 0 1 34816
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_61_3
timestamp 1679235063
transform 1 0 1380 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_15
timestamp 1679235063
transform 1 0 2484 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_27
timestamp 1679235063
transform 1 0 3588 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_39
timestamp 1679235063
transform 1 0 4692 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_61_51
timestamp 1679235063
transform 1 0 5796 0 -1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_61_55
timestamp 1679235063
transform 1 0 6164 0 -1 35904
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_61_57
timestamp 1679235063
transform 1 0 6348 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_69
timestamp 1679235063
transform 1 0 7452 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_81
timestamp 1679235063
transform 1 0 8556 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_93
timestamp 1679235063
transform 1 0 9660 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_61_105
timestamp 1679235063
transform 1 0 10764 0 -1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_61_111
timestamp 1679235063
transform 1 0 11316 0 -1 35904
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_61_113
timestamp 1679235063
transform 1 0 11500 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_125
timestamp 1679235063
transform 1 0 12604 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_137
timestamp 1679235063
transform 1 0 13708 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_149
timestamp 1679235063
transform 1 0 14812 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_61_161
timestamp 1679235063
transform 1 0 15916 0 -1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_61_167
timestamp 1679235063
transform 1 0 16468 0 -1 35904
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_61_169
timestamp 1679235063
transform 1 0 16652 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_181
timestamp 1679235063
transform 1 0 17756 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_193
timestamp 1679235063
transform 1 0 18860 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_61_205
timestamp 1679235063
transform 1 0 19964 0 -1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_61_211
timestamp 1679235063
transform 1 0 20516 0 -1 35904
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_61_222
timestamp 1679235063
transform 1 0 21528 0 -1 35904
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_61_225
timestamp 1679235063
transform 1 0 21804 0 -1 35904
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_61_236
timestamp 1679235063
transform 1 0 22816 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_61_248
timestamp 1679235063
transform 1 0 23920 0 -1 35904
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_61_256
timestamp 1679235063
transform 1 0 24656 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_61_259
timestamp 1679235063
transform 1 0 24932 0 -1 35904
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_61_264
timestamp 1679235063
transform 1 0 25392 0 -1 35904
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_62_3
timestamp 1679235063
transform 1 0 1380 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_15
timestamp 1679235063
transform 1 0 2484 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_62_27
timestamp 1679235063
transform 1 0 3588 0 1 35904
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_62_29
timestamp 1679235063
transform 1 0 3772 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_41
timestamp 1679235063
transform 1 0 4876 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_53
timestamp 1679235063
transform 1 0 5980 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_65
timestamp 1679235063
transform 1 0 7084 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_62_77
timestamp 1679235063
transform 1 0 8188 0 1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_62_83
timestamp 1679235063
transform 1 0 8740 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_62_85
timestamp 1679235063
transform 1 0 8924 0 1 35904
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_62_90
timestamp 1679235063
transform 1 0 9384 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_102
timestamp 1679235063
transform 1 0 10488 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_114
timestamp 1679235063
transform 1 0 11592 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_126
timestamp 1679235063
transform 1 0 12696 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_62_138
timestamp 1679235063
transform 1 0 13800 0 1 35904
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_62_141
timestamp 1679235063
transform 1 0 14076 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_153
timestamp 1679235063
transform 1 0 15180 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_165
timestamp 1679235063
transform 1 0 16284 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_177
timestamp 1679235063
transform 1 0 17388 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_62_189
timestamp 1679235063
transform 1 0 18492 0 1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_62_195
timestamp 1679235063
transform 1 0 19044 0 1 35904
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_62_197
timestamp 1679235063
transform 1 0 19228 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_209
timestamp 1679235063
transform 1 0 20332 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_221
timestamp 1679235063
transform 1 0 21436 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_233
timestamp 1679235063
transform 1 0 22540 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_62_245
timestamp 1679235063
transform 1 0 23644 0 1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_62_251
timestamp 1679235063
transform 1 0 24196 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_62_253
timestamp 1679235063
transform 1 0 24380 0 1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_62_259
timestamp 1679235063
transform 1 0 24932 0 1 35904
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_62_264
timestamp 1679235063
transform 1 0 25392 0 1 35904
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_63_3
timestamp 1679235063
transform 1 0 1380 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_63_15
timestamp 1679235063
transform 1 0 2484 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_63_27
timestamp 1679235063
transform 1 0 3588 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_63_39
timestamp 1679235063
transform 1 0 4692 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_63_51
timestamp 1679235063
transform 1 0 5796 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_63_55
timestamp 1679235063
transform 1 0 6164 0 -1 36992
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_63_57
timestamp 1679235063
transform 1 0 6348 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_63_69
timestamp 1679235063
transform 1 0 7452 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_63_81
timestamp 1679235063
transform 1 0 8556 0 -1 36992
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_63_89
timestamp 1679235063
transform 1 0 9292 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_63_110
timestamp 1679235063
transform 1 0 11224 0 -1 36992
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_63_117
timestamp 1679235063
transform 1 0 11868 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_63_129
timestamp 1679235063
transform 1 0 12972 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_63_141
timestamp 1679235063
transform 1 0 14076 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_63_153
timestamp 1679235063
transform 1 0 15180 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_63_165
timestamp 1679235063
transform 1 0 16284 0 -1 36992
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_63_169
timestamp 1679235063
transform 1 0 16652 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_63_181
timestamp 1679235063
transform 1 0 17756 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_63_193
timestamp 1679235063
transform 1 0 18860 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_63_205
timestamp 1679235063
transform 1 0 19964 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_63_217
timestamp 1679235063
transform 1 0 21068 0 -1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_63_223
timestamp 1679235063
transform 1 0 21620 0 -1 36992
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_63_225
timestamp 1679235063
transform 1 0 21804 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_63_237
timestamp 1679235063
transform 1 0 22908 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_63_249
timestamp 1679235063
transform 1 0 24012 0 -1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_63_255
timestamp 1679235063
transform 1 0 24564 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_63_258
timestamp 1679235063
transform 1 0 24840 0 -1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_63_264
timestamp 1679235063
transform 1 0 25392 0 -1 36992
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_64_3
timestamp 1679235063
transform 1 0 1380 0 1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_64_15
timestamp 1679235063
transform 1 0 2484 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_64_27
timestamp 1679235063
transform 1 0 3588 0 1 36992
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_64_29
timestamp 1679235063
transform 1 0 3772 0 1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_64_41
timestamp 1679235063
transform 1 0 4876 0 1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_64_53
timestamp 1679235063
transform 1 0 5980 0 1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_64_65
timestamp 1679235063
transform 1 0 7084 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_64_77
timestamp 1679235063
transform 1 0 8188 0 1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_64_83
timestamp 1679235063
transform 1 0 8740 0 1 36992
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_64_85
timestamp 1679235063
transform 1 0 8924 0 1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_64_97
timestamp 1679235063
transform 1 0 10028 0 1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_64_109
timestamp 1679235063
transform 1 0 11132 0 1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_64_121
timestamp 1679235063
transform 1 0 12236 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_64_133
timestamp 1679235063
transform 1 0 13340 0 1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_64_139
timestamp 1679235063
transform 1 0 13892 0 1 36992
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_64_141
timestamp 1679235063
transform 1 0 14076 0 1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_64_153
timestamp 1679235063
transform 1 0 15180 0 1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_64_165
timestamp 1679235063
transform 1 0 16284 0 1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_64_177
timestamp 1679235063
transform 1 0 17388 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_64_189
timestamp 1679235063
transform 1 0 18492 0 1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_64_195
timestamp 1679235063
transform 1 0 19044 0 1 36992
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_64_197
timestamp 1679235063
transform 1 0 19228 0 1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_64_209
timestamp 1679235063
transform 1 0 20332 0 1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_64_221
timestamp 1679235063
transform 1 0 21436 0 1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_64_233
timestamp 1679235063
transform 1 0 22540 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_64_245
timestamp 1679235063
transform 1 0 23644 0 1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_64_251
timestamp 1679235063
transform 1 0 24196 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_64_253
timestamp 1679235063
transform 1 0 24380 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_64_259
timestamp 1679235063
transform 1 0 24932 0 1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_64_264
timestamp 1679235063
transform 1 0 25392 0 1 36992
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_65_3
timestamp 1679235063
transform 1 0 1380 0 -1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_65_15
timestamp 1679235063
transform 1 0 2484 0 -1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_65_27
timestamp 1679235063
transform 1 0 3588 0 -1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_65_39
timestamp 1679235063
transform 1 0 4692 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_65_51
timestamp 1679235063
transform 1 0 5796 0 -1 38080
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_65_55
timestamp 1679235063
transform 1 0 6164 0 -1 38080
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_65_57
timestamp 1679235063
transform 1 0 6348 0 -1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_65_69
timestamp 1679235063
transform 1 0 7452 0 -1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_65_81
timestamp 1679235063
transform 1 0 8556 0 -1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_65_93
timestamp 1679235063
transform 1 0 9660 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_65_105
timestamp 1679235063
transform 1 0 10764 0 -1 38080
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_65_111
timestamp 1679235063
transform 1 0 11316 0 -1 38080
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_65_113
timestamp 1679235063
transform 1 0 11500 0 -1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_65_125
timestamp 1679235063
transform 1 0 12604 0 -1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_65_137
timestamp 1679235063
transform 1 0 13708 0 -1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_65_149
timestamp 1679235063
transform 1 0 14812 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_65_161
timestamp 1679235063
transform 1 0 15916 0 -1 38080
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_65_167
timestamp 1679235063
transform 1 0 16468 0 -1 38080
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_65_169
timestamp 1679235063
transform 1 0 16652 0 -1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_65_181
timestamp 1679235063
transform 1 0 17756 0 -1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_65_193
timestamp 1679235063
transform 1 0 18860 0 -1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_65_205
timestamp 1679235063
transform 1 0 19964 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_65_217
timestamp 1679235063
transform 1 0 21068 0 -1 38080
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_65_223
timestamp 1679235063
transform 1 0 21620 0 -1 38080
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_65_225
timestamp 1679235063
transform 1 0 21804 0 -1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_65_237
timestamp 1679235063
transform 1 0 22908 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_65_249
timestamp 1679235063
transform 1 0 24012 0 -1 38080
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_65_255
timestamp 1679235063
transform 1 0 24564 0 -1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_65_258
timestamp 1679235063
transform 1 0 24840 0 -1 38080
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_65_264
timestamp 1679235063
transform 1 0 25392 0 -1 38080
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_66_3
timestamp 1679235063
transform 1 0 1380 0 1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_66_15
timestamp 1679235063
transform 1 0 2484 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_66_27
timestamp 1679235063
transform 1 0 3588 0 1 38080
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_66_29
timestamp 1679235063
transform 1 0 3772 0 1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_66_41
timestamp 1679235063
transform 1 0 4876 0 1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_66_53
timestamp 1679235063
transform 1 0 5980 0 1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_66_65
timestamp 1679235063
transform 1 0 7084 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_66_77
timestamp 1679235063
transform 1 0 8188 0 1 38080
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_66_83
timestamp 1679235063
transform 1 0 8740 0 1 38080
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_66_85
timestamp 1679235063
transform 1 0 8924 0 1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_66_97
timestamp 1679235063
transform 1 0 10028 0 1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_66_109
timestamp 1679235063
transform 1 0 11132 0 1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_66_121
timestamp 1679235063
transform 1 0 12236 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_66_133
timestamp 1679235063
transform 1 0 13340 0 1 38080
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_66_139
timestamp 1679235063
transform 1 0 13892 0 1 38080
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_66_141
timestamp 1679235063
transform 1 0 14076 0 1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_66_153
timestamp 1679235063
transform 1 0 15180 0 1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_66_165
timestamp 1679235063
transform 1 0 16284 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_66_177
timestamp 1679235063
transform 1 0 17388 0 1 38080
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_66_188
timestamp 1679235063
transform 1 0 18400 0 1 38080
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_66_197
timestamp 1679235063
transform 1 0 19228 0 1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_66_209
timestamp 1679235063
transform 1 0 20332 0 1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_66_221
timestamp 1679235063
transform 1 0 21436 0 1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_66_233
timestamp 1679235063
transform 1 0 22540 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_66_245
timestamp 1679235063
transform 1 0 23644 0 1 38080
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_66_251
timestamp 1679235063
transform 1 0 24196 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_66_253
timestamp 1679235063
transform 1 0 24380 0 1 38080
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_66_264
timestamp 1679235063
transform 1 0 25392 0 1 38080
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_67_3
timestamp 1679235063
transform 1 0 1380 0 -1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_67_15
timestamp 1679235063
transform 1 0 2484 0 -1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_67_27
timestamp 1679235063
transform 1 0 3588 0 -1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_67_39
timestamp 1679235063
transform 1 0 4692 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_67_51
timestamp 1679235063
transform 1 0 5796 0 -1 39168
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_67_55
timestamp 1679235063
transform 1 0 6164 0 -1 39168
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_67_57
timestamp 1679235063
transform 1 0 6348 0 -1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_67_69
timestamp 1679235063
transform 1 0 7452 0 -1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_67_81
timestamp 1679235063
transform 1 0 8556 0 -1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_67_93
timestamp 1679235063
transform 1 0 9660 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_67_105
timestamp 1679235063
transform 1 0 10764 0 -1 39168
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_67_111
timestamp 1679235063
transform 1 0 11316 0 -1 39168
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_67_113
timestamp 1679235063
transform 1 0 11500 0 -1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_67_125
timestamp 1679235063
transform 1 0 12604 0 -1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_67_137
timestamp 1679235063
transform 1 0 13708 0 -1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_67_149
timestamp 1679235063
transform 1 0 14812 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_67_161
timestamp 1679235063
transform 1 0 15916 0 -1 39168
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_67_167
timestamp 1679235063
transform 1 0 16468 0 -1 39168
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_67_169
timestamp 1679235063
transform 1 0 16652 0 -1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_67_181
timestamp 1679235063
transform 1 0 17756 0 -1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_67_193
timestamp 1679235063
transform 1 0 18860 0 -1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_67_205
timestamp 1679235063
transform 1 0 19964 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_67_217
timestamp 1679235063
transform 1 0 21068 0 -1 39168
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_67_223
timestamp 1679235063
transform 1 0 21620 0 -1 39168
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_67_225
timestamp 1679235063
transform 1 0 21804 0 -1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_67_237
timestamp 1679235063
transform 1 0 22908 0 -1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_67_249
timestamp 1679235063
transform 1 0 24012 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_67_261
timestamp 1679235063
transform 1 0 25116 0 -1 39168
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_68_3
timestamp 1679235063
transform 1 0 1380 0 1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_68_15
timestamp 1679235063
transform 1 0 2484 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_68_27
timestamp 1679235063
transform 1 0 3588 0 1 39168
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_68_29
timestamp 1679235063
transform 1 0 3772 0 1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_68_41
timestamp 1679235063
transform 1 0 4876 0 1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_68_53
timestamp 1679235063
transform 1 0 5980 0 1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_68_65
timestamp 1679235063
transform 1 0 7084 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_68_77
timestamp 1679235063
transform 1 0 8188 0 1 39168
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_68_83
timestamp 1679235063
transform 1 0 8740 0 1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_68_85
timestamp 1679235063
transform 1 0 8924 0 1 39168
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_68_90
timestamp 1679235063
transform 1 0 9384 0 1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_68_102
timestamp 1679235063
transform 1 0 10488 0 1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_68_114
timestamp 1679235063
transform 1 0 11592 0 1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_68_126
timestamp 1679235063
transform 1 0 12696 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_68_138
timestamp 1679235063
transform 1 0 13800 0 1 39168
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_68_141
timestamp 1679235063
transform 1 0 14076 0 1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_68_153
timestamp 1679235063
transform 1 0 15180 0 1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_68_165
timestamp 1679235063
transform 1 0 16284 0 1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_68_177
timestamp 1679235063
transform 1 0 17388 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_68_189
timestamp 1679235063
transform 1 0 18492 0 1 39168
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_68_195
timestamp 1679235063
transform 1 0 19044 0 1 39168
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_68_197
timestamp 1679235063
transform 1 0 19228 0 1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_68_209
timestamp 1679235063
transform 1 0 20332 0 1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_68_221
timestamp 1679235063
transform 1 0 21436 0 1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_68_233
timestamp 1679235063
transform 1 0 22540 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_68_245
timestamp 1679235063
transform 1 0 23644 0 1 39168
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_68_251
timestamp 1679235063
transform 1 0 24196 0 1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_68_253
timestamp 1679235063
transform 1 0 24380 0 1 39168
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_68_259
timestamp 1679235063
transform 1 0 24932 0 1 39168
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_68_264
timestamp 1679235063
transform 1 0 25392 0 1 39168
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_69_3
timestamp 1679235063
transform 1 0 1380 0 -1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_69_15
timestamp 1679235063
transform 1 0 2484 0 -1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_69_27
timestamp 1679235063
transform 1 0 3588 0 -1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_69_39
timestamp 1679235063
transform 1 0 4692 0 -1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_69_51
timestamp 1679235063
transform 1 0 5796 0 -1 40256
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_69_55
timestamp 1679235063
transform 1 0 6164 0 -1 40256
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_69_57
timestamp 1679235063
transform 1 0 6348 0 -1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_69_69
timestamp 1679235063
transform 1 0 7452 0 -1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_69_81
timestamp 1679235063
transform 1 0 8556 0 -1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_69_93
timestamp 1679235063
transform 1 0 9660 0 -1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_69_105
timestamp 1679235063
transform 1 0 10764 0 -1 40256
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_69_111
timestamp 1679235063
transform 1 0 11316 0 -1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_69_113
timestamp 1679235063
transform 1 0 11500 0 -1 40256
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_69_123
timestamp 1679235063
transform 1 0 12420 0 -1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_69_135
timestamp 1679235063
transform 1 0 13524 0 -1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_69_147
timestamp 1679235063
transform 1 0 14628 0 -1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_69_159
timestamp 1679235063
transform 1 0 15732 0 -1 40256
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_69_167
timestamp 1679235063
transform 1 0 16468 0 -1 40256
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_69_169
timestamp 1679235063
transform 1 0 16652 0 -1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_69_181
timestamp 1679235063
transform 1 0 17756 0 -1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_69_193
timestamp 1679235063
transform 1 0 18860 0 -1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_69_205
timestamp 1679235063
transform 1 0 19964 0 -1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_69_217
timestamp 1679235063
transform 1 0 21068 0 -1 40256
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_69_223
timestamp 1679235063
transform 1 0 21620 0 -1 40256
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_69_225
timestamp 1679235063
transform 1 0 21804 0 -1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_69_237
timestamp 1679235063
transform 1 0 22908 0 -1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_69_249
timestamp 1679235063
transform 1 0 24012 0 -1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_69_264
timestamp 1679235063
transform 1 0 25392 0 -1 40256
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_70_3
timestamp 1679235063
transform 1 0 1380 0 1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_70_15
timestamp 1679235063
transform 1 0 2484 0 1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_70_27
timestamp 1679235063
transform 1 0 3588 0 1 40256
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_70_29
timestamp 1679235063
transform 1 0 3772 0 1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_70_41
timestamp 1679235063
transform 1 0 4876 0 1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_70_53
timestamp 1679235063
transform 1 0 5980 0 1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_70_65
timestamp 1679235063
transform 1 0 7084 0 1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_70_77
timestamp 1679235063
transform 1 0 8188 0 1 40256
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_70_83
timestamp 1679235063
transform 1 0 8740 0 1 40256
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_70_85
timestamp 1679235063
transform 1 0 8924 0 1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_70_97
timestamp 1679235063
transform 1 0 10028 0 1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_70_109
timestamp 1679235063
transform 1 0 11132 0 1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_70_121
timestamp 1679235063
transform 1 0 12236 0 1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_70_133
timestamp 1679235063
transform 1 0 13340 0 1 40256
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_70_139
timestamp 1679235063
transform 1 0 13892 0 1 40256
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_70_141
timestamp 1679235063
transform 1 0 14076 0 1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_70_153
timestamp 1679235063
transform 1 0 15180 0 1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_70_165
timestamp 1679235063
transform 1 0 16284 0 1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_70_177
timestamp 1679235063
transform 1 0 17388 0 1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_70_189
timestamp 1679235063
transform 1 0 18492 0 1 40256
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_70_195
timestamp 1679235063
transform 1 0 19044 0 1 40256
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_70_197
timestamp 1679235063
transform 1 0 19228 0 1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_70_209
timestamp 1679235063
transform 1 0 20332 0 1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_70_221
timestamp 1679235063
transform 1 0 21436 0 1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_70_233
timestamp 1679235063
transform 1 0 22540 0 1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_70_245
timestamp 1679235063
transform 1 0 23644 0 1 40256
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_70_251
timestamp 1679235063
transform 1 0 24196 0 1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_70_253
timestamp 1679235063
transform 1 0 24380 0 1 40256
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_70_261
timestamp 1679235063
transform 1 0 25116 0 1 40256
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_71_3
timestamp 1679235063
transform 1 0 1380 0 -1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_71_15
timestamp 1679235063
transform 1 0 2484 0 -1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_71_27
timestamp 1679235063
transform 1 0 3588 0 -1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_71_39
timestamp 1679235063
transform 1 0 4692 0 -1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_71_51
timestamp 1679235063
transform 1 0 5796 0 -1 41344
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_71_55
timestamp 1679235063
transform 1 0 6164 0 -1 41344
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_71_57
timestamp 1679235063
transform 1 0 6348 0 -1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_71_69
timestamp 1679235063
transform 1 0 7452 0 -1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_71_81
timestamp 1679235063
transform 1 0 8556 0 -1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_71_93
timestamp 1679235063
transform 1 0 9660 0 -1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_71_105
timestamp 1679235063
transform 1 0 10764 0 -1 41344
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_71_111
timestamp 1679235063
transform 1 0 11316 0 -1 41344
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_71_113
timestamp 1679235063
transform 1 0 11500 0 -1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_71_125
timestamp 1679235063
transform 1 0 12604 0 -1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_71_137
timestamp 1679235063
transform 1 0 13708 0 -1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_71_149
timestamp 1679235063
transform 1 0 14812 0 -1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_71_161
timestamp 1679235063
transform 1 0 15916 0 -1 41344
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_71_167
timestamp 1679235063
transform 1 0 16468 0 -1 41344
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_71_169
timestamp 1679235063
transform 1 0 16652 0 -1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_71_181
timestamp 1679235063
transform 1 0 17756 0 -1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_71_193
timestamp 1679235063
transform 1 0 18860 0 -1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_71_205
timestamp 1679235063
transform 1 0 19964 0 -1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_71_217
timestamp 1679235063
transform 1 0 21068 0 -1 41344
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_71_223
timestamp 1679235063
transform 1 0 21620 0 -1 41344
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_71_225
timestamp 1679235063
transform 1 0 21804 0 -1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_71_237
timestamp 1679235063
transform 1 0 22908 0 -1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_71_249
timestamp 1679235063
transform 1 0 24012 0 -1 41344
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_71_259
timestamp 1679235063
transform 1 0 24932 0 -1 41344
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_71_264
timestamp 1679235063
transform 1 0 25392 0 -1 41344
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_72_3
timestamp 1679235063
transform 1 0 1380 0 1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_72_15
timestamp 1679235063
transform 1 0 2484 0 1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_72_27
timestamp 1679235063
transform 1 0 3588 0 1 41344
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_72_29
timestamp 1679235063
transform 1 0 3772 0 1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_72_41
timestamp 1679235063
transform 1 0 4876 0 1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_72_53
timestamp 1679235063
transform 1 0 5980 0 1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_72_65
timestamp 1679235063
transform 1 0 7084 0 1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_72_77
timestamp 1679235063
transform 1 0 8188 0 1 41344
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_72_83
timestamp 1679235063
transform 1 0 8740 0 1 41344
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_72_85
timestamp 1679235063
transform 1 0 8924 0 1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_72_97
timestamp 1679235063
transform 1 0 10028 0 1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_72_109
timestamp 1679235063
transform 1 0 11132 0 1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_72_121
timestamp 1679235063
transform 1 0 12236 0 1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_72_133
timestamp 1679235063
transform 1 0 13340 0 1 41344
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_72_139
timestamp 1679235063
transform 1 0 13892 0 1 41344
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_72_141
timestamp 1679235063
transform 1 0 14076 0 1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_72_153
timestamp 1679235063
transform 1 0 15180 0 1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_72_165
timestamp 1679235063
transform 1 0 16284 0 1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_72_177
timestamp 1679235063
transform 1 0 17388 0 1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_72_189
timestamp 1679235063
transform 1 0 18492 0 1 41344
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_72_195
timestamp 1679235063
transform 1 0 19044 0 1 41344
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_72_197
timestamp 1679235063
transform 1 0 19228 0 1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_72_209
timestamp 1679235063
transform 1 0 20332 0 1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_72_221
timestamp 1679235063
transform 1 0 21436 0 1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_72_233
timestamp 1679235063
transform 1 0 22540 0 1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_72_245
timestamp 1679235063
transform 1 0 23644 0 1 41344
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_72_251
timestamp 1679235063
transform 1 0 24196 0 1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_72_253
timestamp 1679235063
transform 1 0 24380 0 1 41344
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_72_259
timestamp 1679235063
transform 1 0 24932 0 1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_72_264
timestamp 1679235063
transform 1 0 25392 0 1 41344
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_73_3
timestamp 1679235063
transform 1 0 1380 0 -1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_73_15
timestamp 1679235063
transform 1 0 2484 0 -1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_73_27
timestamp 1679235063
transform 1 0 3588 0 -1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_73_39
timestamp 1679235063
transform 1 0 4692 0 -1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_73_51
timestamp 1679235063
transform 1 0 5796 0 -1 42432
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_73_55
timestamp 1679235063
transform 1 0 6164 0 -1 42432
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_73_57
timestamp 1679235063
transform 1 0 6348 0 -1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_73_69
timestamp 1679235063
transform 1 0 7452 0 -1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_73_81
timestamp 1679235063
transform 1 0 8556 0 -1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_73_93
timestamp 1679235063
transform 1 0 9660 0 -1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_73_105
timestamp 1679235063
transform 1 0 10764 0 -1 42432
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_73_111
timestamp 1679235063
transform 1 0 11316 0 -1 42432
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_73_113
timestamp 1679235063
transform 1 0 11500 0 -1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_73_125
timestamp 1679235063
transform 1 0 12604 0 -1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_73_137
timestamp 1679235063
transform 1 0 13708 0 -1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_73_149
timestamp 1679235063
transform 1 0 14812 0 -1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_73_161
timestamp 1679235063
transform 1 0 15916 0 -1 42432
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_73_167
timestamp 1679235063
transform 1 0 16468 0 -1 42432
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_73_169
timestamp 1679235063
transform 1 0 16652 0 -1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_73_181
timestamp 1679235063
transform 1 0 17756 0 -1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_73_193
timestamp 1679235063
transform 1 0 18860 0 -1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_73_205
timestamp 1679235063
transform 1 0 19964 0 -1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_73_217
timestamp 1679235063
transform 1 0 21068 0 -1 42432
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_73_223
timestamp 1679235063
transform 1 0 21620 0 -1 42432
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_73_225
timestamp 1679235063
transform 1 0 21804 0 -1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_73_237
timestamp 1679235063
transform 1 0 22908 0 -1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_73_249
timestamp 1679235063
transform 1 0 24012 0 -1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_73_261
timestamp 1679235063
transform 1 0 25116 0 -1 42432
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_74_3
timestamp 1679235063
transform 1 0 1380 0 1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_74_15
timestamp 1679235063
transform 1 0 2484 0 1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_74_27
timestamp 1679235063
transform 1 0 3588 0 1 42432
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_74_29
timestamp 1679235063
transform 1 0 3772 0 1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_74_41
timestamp 1679235063
transform 1 0 4876 0 1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_74_53
timestamp 1679235063
transform 1 0 5980 0 1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_74_65
timestamp 1679235063
transform 1 0 7084 0 1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_74_77
timestamp 1679235063
transform 1 0 8188 0 1 42432
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_74_83
timestamp 1679235063
transform 1 0 8740 0 1 42432
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_74_85
timestamp 1679235063
transform 1 0 8924 0 1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_74_97
timestamp 1679235063
transform 1 0 10028 0 1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_74_109
timestamp 1679235063
transform 1 0 11132 0 1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_74_121
timestamp 1679235063
transform 1 0 12236 0 1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_74_133
timestamp 1679235063
transform 1 0 13340 0 1 42432
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_74_139
timestamp 1679235063
transform 1 0 13892 0 1 42432
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_74_141
timestamp 1679235063
transform 1 0 14076 0 1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_74_153
timestamp 1679235063
transform 1 0 15180 0 1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_74_165
timestamp 1679235063
transform 1 0 16284 0 1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_74_177
timestamp 1679235063
transform 1 0 17388 0 1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_74_189
timestamp 1679235063
transform 1 0 18492 0 1 42432
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_74_195
timestamp 1679235063
transform 1 0 19044 0 1 42432
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_74_197
timestamp 1679235063
transform 1 0 19228 0 1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_74_209
timestamp 1679235063
transform 1 0 20332 0 1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_74_221
timestamp 1679235063
transform 1 0 21436 0 1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_74_233
timestamp 1679235063
transform 1 0 22540 0 1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_74_245
timestamp 1679235063
transform 1 0 23644 0 1 42432
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_74_251
timestamp 1679235063
transform 1 0 24196 0 1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_74_253
timestamp 1679235063
transform 1 0 24380 0 1 42432
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_74_258
timestamp 1679235063
transform 1 0 24840 0 1 42432
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_74_264
timestamp 1679235063
transform 1 0 25392 0 1 42432
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_75_3
timestamp 1679235063
transform 1 0 1380 0 -1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_75_15
timestamp 1679235063
transform 1 0 2484 0 -1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_75_27
timestamp 1679235063
transform 1 0 3588 0 -1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_75_39
timestamp 1679235063
transform 1 0 4692 0 -1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_75_51
timestamp 1679235063
transform 1 0 5796 0 -1 43520
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_75_55
timestamp 1679235063
transform 1 0 6164 0 -1 43520
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_75_57
timestamp 1679235063
transform 1 0 6348 0 -1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_75_69
timestamp 1679235063
transform 1 0 7452 0 -1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_75_81
timestamp 1679235063
transform 1 0 8556 0 -1 43520
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_75_89
timestamp 1679235063
transform 1 0 9292 0 -1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_75_110
timestamp 1679235063
transform 1 0 11224 0 -1 43520
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_75_117
timestamp 1679235063
transform 1 0 11868 0 -1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_75_129
timestamp 1679235063
transform 1 0 12972 0 -1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_75_141
timestamp 1679235063
transform 1 0 14076 0 -1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_75_153
timestamp 1679235063
transform 1 0 15180 0 -1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_75_165
timestamp 1679235063
transform 1 0 16284 0 -1 43520
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_75_169
timestamp 1679235063
transform 1 0 16652 0 -1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_75_181
timestamp 1679235063
transform 1 0 17756 0 -1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_75_193
timestamp 1679235063
transform 1 0 18860 0 -1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_75_205
timestamp 1679235063
transform 1 0 19964 0 -1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_75_217
timestamp 1679235063
transform 1 0 21068 0 -1 43520
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_75_223
timestamp 1679235063
transform 1 0 21620 0 -1 43520
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_75_225
timestamp 1679235063
transform 1 0 21804 0 -1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_75_237
timestamp 1679235063
transform 1 0 22908 0 -1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_75_249
timestamp 1679235063
transform 1 0 24012 0 -1 43520
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_75_257
timestamp 1679235063
transform 1 0 24748 0 -1 43520
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_75_264
timestamp 1679235063
transform 1 0 25392 0 -1 43520
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_76_3
timestamp 1679235063
transform 1 0 1380 0 1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_76_15
timestamp 1679235063
transform 1 0 2484 0 1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_76_27
timestamp 1679235063
transform 1 0 3588 0 1 43520
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_76_29
timestamp 1679235063
transform 1 0 3772 0 1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_76_41
timestamp 1679235063
transform 1 0 4876 0 1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_76_53
timestamp 1679235063
transform 1 0 5980 0 1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_76_65
timestamp 1679235063
transform 1 0 7084 0 1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_76_77
timestamp 1679235063
transform 1 0 8188 0 1 43520
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_76_83
timestamp 1679235063
transform 1 0 8740 0 1 43520
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_76_85
timestamp 1679235063
transform 1 0 8924 0 1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_76_97
timestamp 1679235063
transform 1 0 10028 0 1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_76_109
timestamp 1679235063
transform 1 0 11132 0 1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_76_121
timestamp 1679235063
transform 1 0 12236 0 1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_76_133
timestamp 1679235063
transform 1 0 13340 0 1 43520
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_76_139
timestamp 1679235063
transform 1 0 13892 0 1 43520
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_76_141
timestamp 1679235063
transform 1 0 14076 0 1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_76_153
timestamp 1679235063
transform 1 0 15180 0 1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_76_165
timestamp 1679235063
transform 1 0 16284 0 1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_76_177
timestamp 1679235063
transform 1 0 17388 0 1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_76_189
timestamp 1679235063
transform 1 0 18492 0 1 43520
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_76_195
timestamp 1679235063
transform 1 0 19044 0 1 43520
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_76_197
timestamp 1679235063
transform 1 0 19228 0 1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_76_209
timestamp 1679235063
transform 1 0 20332 0 1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_76_221
timestamp 1679235063
transform 1 0 21436 0 1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_76_233
timestamp 1679235063
transform 1 0 22540 0 1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_76_245
timestamp 1679235063
transform 1 0 23644 0 1 43520
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_76_251
timestamp 1679235063
transform 1 0 24196 0 1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_76_253
timestamp 1679235063
transform 1 0 24380 0 1 43520
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_76_261
timestamp 1679235063
transform 1 0 25116 0 1 43520
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_77_3
timestamp 1679235063
transform 1 0 1380 0 -1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_77_15
timestamp 1679235063
transform 1 0 2484 0 -1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_77_27
timestamp 1679235063
transform 1 0 3588 0 -1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_77_39
timestamp 1679235063
transform 1 0 4692 0 -1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_77_51
timestamp 1679235063
transform 1 0 5796 0 -1 44608
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_77_55
timestamp 1679235063
transform 1 0 6164 0 -1 44608
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_77_57
timestamp 1679235063
transform 1 0 6348 0 -1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_77_69
timestamp 1679235063
transform 1 0 7452 0 -1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_77_81
timestamp 1679235063
transform 1 0 8556 0 -1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_77_93
timestamp 1679235063
transform 1 0 9660 0 -1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_77_105
timestamp 1679235063
transform 1 0 10764 0 -1 44608
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_77_111
timestamp 1679235063
transform 1 0 11316 0 -1 44608
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_77_113
timestamp 1679235063
transform 1 0 11500 0 -1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_77_125
timestamp 1679235063
transform 1 0 12604 0 -1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_77_137
timestamp 1679235063
transform 1 0 13708 0 -1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_77_149
timestamp 1679235063
transform 1 0 14812 0 -1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_77_161
timestamp 1679235063
transform 1 0 15916 0 -1 44608
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_77_167
timestamp 1679235063
transform 1 0 16468 0 -1 44608
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_77_169
timestamp 1679235063
transform 1 0 16652 0 -1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_77_181
timestamp 1679235063
transform 1 0 17756 0 -1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_77_193
timestamp 1679235063
transform 1 0 18860 0 -1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_77_205
timestamp 1679235063
transform 1 0 19964 0 -1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_77_217
timestamp 1679235063
transform 1 0 21068 0 -1 44608
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_77_223
timestamp 1679235063
transform 1 0 21620 0 -1 44608
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_77_225
timestamp 1679235063
transform 1 0 21804 0 -1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_77_237
timestamp 1679235063
transform 1 0 22908 0 -1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_77_249
timestamp 1679235063
transform 1 0 24012 0 -1 44608
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_77_255
timestamp 1679235063
transform 1 0 24564 0 -1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_77_258
timestamp 1679235063
transform 1 0 24840 0 -1 44608
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_77_264
timestamp 1679235063
transform 1 0 25392 0 -1 44608
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_78_3
timestamp 1679235063
transform 1 0 1380 0 1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_78_15
timestamp 1679235063
transform 1 0 2484 0 1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_78_27
timestamp 1679235063
transform 1 0 3588 0 1 44608
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_78_29
timestamp 1679235063
transform 1 0 3772 0 1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_78_41
timestamp 1679235063
transform 1 0 4876 0 1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_78_53
timestamp 1679235063
transform 1 0 5980 0 1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_78_65
timestamp 1679235063
transform 1 0 7084 0 1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_78_77
timestamp 1679235063
transform 1 0 8188 0 1 44608
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_78_83
timestamp 1679235063
transform 1 0 8740 0 1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_78_85
timestamp 1679235063
transform 1 0 8924 0 1 44608
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_78_93
timestamp 1679235063
transform 1 0 9660 0 1 44608
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_78_104
timestamp 1679235063
transform 1 0 10672 0 1 44608
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_78_115
timestamp 1679235063
transform 1 0 11684 0 1 44608
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_78_119
timestamp 1679235063
transform 1 0 12052 0 1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_78_131
timestamp 1679235063
transform 1 0 13156 0 1 44608
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_78_139
timestamp 1679235063
transform 1 0 13892 0 1 44608
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_78_141
timestamp 1679235063
transform 1 0 14076 0 1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_78_153
timestamp 1679235063
transform 1 0 15180 0 1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_78_165
timestamp 1679235063
transform 1 0 16284 0 1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_78_177
timestamp 1679235063
transform 1 0 17388 0 1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_78_189
timestamp 1679235063
transform 1 0 18492 0 1 44608
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_78_195
timestamp 1679235063
transform 1 0 19044 0 1 44608
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_78_197
timestamp 1679235063
transform 1 0 19228 0 1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_78_209
timestamp 1679235063
transform 1 0 20332 0 1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_78_230
timestamp 1679235063
transform 1 0 22264 0 1 44608
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_78_234
timestamp 1679235063
transform 1 0 22632 0 1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_78_246
timestamp 1679235063
transform 1 0 23736 0 1 44608
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_78_253
timestamp 1679235063
transform 1 0 24380 0 1 44608
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_78_264
timestamp 1679235063
transform 1 0 25392 0 1 44608
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_79_3
timestamp 1679235063
transform 1 0 1380 0 -1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_79_15
timestamp 1679235063
transform 1 0 2484 0 -1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_79_27
timestamp 1679235063
transform 1 0 3588 0 -1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_79_39
timestamp 1679235063
transform 1 0 4692 0 -1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_79_51
timestamp 1679235063
transform 1 0 5796 0 -1 45696
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_79_55
timestamp 1679235063
transform 1 0 6164 0 -1 45696
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_79_57
timestamp 1679235063
transform 1 0 6348 0 -1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_79_69
timestamp 1679235063
transform 1 0 7452 0 -1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_79_81
timestamp 1679235063
transform 1 0 8556 0 -1 45696
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_79_110
timestamp 1679235063
transform 1 0 11224 0 -1 45696
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_79_113
timestamp 1679235063
transform 1 0 11500 0 -1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_79_125
timestamp 1679235063
transform 1 0 12604 0 -1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_79_137
timestamp 1679235063
transform 1 0 13708 0 -1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_79_149
timestamp 1679235063
transform 1 0 14812 0 -1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_79_161
timestamp 1679235063
transform 1 0 15916 0 -1 45696
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_79_167
timestamp 1679235063
transform 1 0 16468 0 -1 45696
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_79_169
timestamp 1679235063
transform 1 0 16652 0 -1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_79_181
timestamp 1679235063
transform 1 0 17756 0 -1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_79_193
timestamp 1679235063
transform 1 0 18860 0 -1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_79_205
timestamp 1679235063
transform 1 0 19964 0 -1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_79_217
timestamp 1679235063
transform 1 0 21068 0 -1 45696
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_79_223
timestamp 1679235063
transform 1 0 21620 0 -1 45696
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_79_225
timestamp 1679235063
transform 1 0 21804 0 -1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_79_237
timestamp 1679235063
transform 1 0 22908 0 -1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_79_249
timestamp 1679235063
transform 1 0 24012 0 -1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_79_261
timestamp 1679235063
transform 1 0 25116 0 -1 45696
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_80_3
timestamp 1679235063
transform 1 0 1380 0 1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_80_15
timestamp 1679235063
transform 1 0 2484 0 1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_80_27
timestamp 1679235063
transform 1 0 3588 0 1 45696
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_80_29
timestamp 1679235063
transform 1 0 3772 0 1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_80_41
timestamp 1679235063
transform 1 0 4876 0 1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_80_53
timestamp 1679235063
transform 1 0 5980 0 1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_80_65
timestamp 1679235063
transform 1 0 7084 0 1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_80_77
timestamp 1679235063
transform 1 0 8188 0 1 45696
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_80_83
timestamp 1679235063
transform 1 0 8740 0 1 45696
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_80_85
timestamp 1679235063
transform 1 0 8924 0 1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_80_97
timestamp 1679235063
transform 1 0 10028 0 1 45696
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_80_122
timestamp 1679235063
transform 1 0 12328 0 1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_80_134
timestamp 1679235063
transform 1 0 13432 0 1 45696
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_80_141
timestamp 1679235063
transform 1 0 14076 0 1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_80_153
timestamp 1679235063
transform 1 0 15180 0 1 45696
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_80_157
timestamp 1679235063
transform 1 0 15548 0 1 45696
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_80_179
timestamp 1679235063
transform 1 0 17572 0 1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_80_191
timestamp 1679235063
transform 1 0 18676 0 1 45696
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_80_195
timestamp 1679235063
transform 1 0 19044 0 1 45696
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_80_197
timestamp 1679235063
transform 1 0 19228 0 1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_80_209
timestamp 1679235063
transform 1 0 20332 0 1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_80_221
timestamp 1679235063
transform 1 0 21436 0 1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_80_233
timestamp 1679235063
transform 1 0 22540 0 1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_80_245
timestamp 1679235063
transform 1 0 23644 0 1 45696
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_80_251
timestamp 1679235063
transform 1 0 24196 0 1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_80_253
timestamp 1679235063
transform 1 0 24380 0 1 45696
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_80_259
timestamp 1679235063
transform 1 0 24932 0 1 45696
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_80_264
timestamp 1679235063
transform 1 0 25392 0 1 45696
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_81_3
timestamp 1679235063
transform 1 0 1380 0 -1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_81_15
timestamp 1679235063
transform 1 0 2484 0 -1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_81_27
timestamp 1679235063
transform 1 0 3588 0 -1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_81_39
timestamp 1679235063
transform 1 0 4692 0 -1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_81_51
timestamp 1679235063
transform 1 0 5796 0 -1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_81_55
timestamp 1679235063
transform 1 0 6164 0 -1 46784
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_81_57
timestamp 1679235063
transform 1 0 6348 0 -1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_81_69
timestamp 1679235063
transform 1 0 7452 0 -1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_81_81
timestamp 1679235063
transform 1 0 8556 0 -1 46784
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_81_104
timestamp 1679235063
transform 1 0 10672 0 -1 46784
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_81_110
timestamp 1679235063
transform 1 0 11224 0 -1 46784
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_81_113
timestamp 1679235063
transform 1 0 11500 0 -1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_81_125
timestamp 1679235063
transform 1 0 12604 0 -1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_81_137
timestamp 1679235063
transform 1 0 13708 0 -1 46784
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_81_166
timestamp 1679235063
transform 1 0 16376 0 -1 46784
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_81_169
timestamp 1679235063
transform 1 0 16652 0 -1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_81_181
timestamp 1679235063
transform 1 0 17756 0 -1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_81_193
timestamp 1679235063
transform 1 0 18860 0 -1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_81_205
timestamp 1679235063
transform 1 0 19964 0 -1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_81_217
timestamp 1679235063
transform 1 0 21068 0 -1 46784
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_81_223
timestamp 1679235063
transform 1 0 21620 0 -1 46784
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_81_225
timestamp 1679235063
transform 1 0 21804 0 -1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_81_237
timestamp 1679235063
transform 1 0 22908 0 -1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_81_249
timestamp 1679235063
transform 1 0 24012 0 -1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_81_264
timestamp 1679235063
transform 1 0 25392 0 -1 46784
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_82_3
timestamp 1679235063
transform 1 0 1380 0 1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_82_15
timestamp 1679235063
transform 1 0 2484 0 1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_82_27
timestamp 1679235063
transform 1 0 3588 0 1 46784
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_82_29
timestamp 1679235063
transform 1 0 3772 0 1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_82_41
timestamp 1679235063
transform 1 0 4876 0 1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_82_53
timestamp 1679235063
transform 1 0 5980 0 1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_82_65
timestamp 1679235063
transform 1 0 7084 0 1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_82_77
timestamp 1679235063
transform 1 0 8188 0 1 46784
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_82_83
timestamp 1679235063
transform 1 0 8740 0 1 46784
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_82_85
timestamp 1679235063
transform 1 0 8924 0 1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_82_97
timestamp 1679235063
transform 1 0 10028 0 1 46784
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_82_107
timestamp 1679235063
transform 1 0 10948 0 1 46784
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_82_111
timestamp 1679235063
transform 1 0 11316 0 1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_82_123
timestamp 1679235063
transform 1 0 12420 0 1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_82_127
timestamp 1679235063
transform 1 0 12788 0 1 46784
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_82_136
timestamp 1679235063
transform 1 0 13616 0 1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_82_141
timestamp 1679235063
transform 1 0 14076 0 1 46784
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_82_164
timestamp 1679235063
transform 1 0 16192 0 1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_82_176
timestamp 1679235063
transform 1 0 17296 0 1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_82_188
timestamp 1679235063
transform 1 0 18400 0 1 46784
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_82_197
timestamp 1679235063
transform 1 0 19228 0 1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_82_209
timestamp 1679235063
transform 1 0 20332 0 1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_82_221
timestamp 1679235063
transform 1 0 21436 0 1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_82_233
timestamp 1679235063
transform 1 0 22540 0 1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_82_245
timestamp 1679235063
transform 1 0 23644 0 1 46784
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_82_251
timestamp 1679235063
transform 1 0 24196 0 1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_82_253
timestamp 1679235063
transform 1 0 24380 0 1 46784
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_82_261
timestamp 1679235063
transform 1 0 25116 0 1 46784
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_83_3
timestamp 1679235063
transform 1 0 1380 0 -1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_83_15
timestamp 1679235063
transform 1 0 2484 0 -1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_83_27
timestamp 1679235063
transform 1 0 3588 0 -1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_83_39
timestamp 1679235063
transform 1 0 4692 0 -1 47872
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_83_51
timestamp 1679235063
transform 1 0 5796 0 -1 47872
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_83_55
timestamp 1679235063
transform 1 0 6164 0 -1 47872
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_83_57
timestamp 1679235063
transform 1 0 6348 0 -1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_83_69
timestamp 1679235063
transform 1 0 7452 0 -1 47872
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_83_81
timestamp 1679235063
transform 1 0 8556 0 -1 47872
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_83_103
timestamp 1679235063
transform 1 0 10580 0 -1 47872
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_83_111
timestamp 1679235063
transform 1 0 11316 0 -1 47872
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_83_113
timestamp 1679235063
transform 1 0 11500 0 -1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_83_146
timestamp 1679235063
transform 1 0 14536 0 -1 47872
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_83_158
timestamp 1679235063
transform 1 0 15640 0 -1 47872
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_83_166
timestamp 1679235063
transform 1 0 16376 0 -1 47872
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_83_169
timestamp 1679235063
transform 1 0 16652 0 -1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_83_181
timestamp 1679235063
transform 1 0 17756 0 -1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_83_193
timestamp 1679235063
transform 1 0 18860 0 -1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_83_205
timestamp 1679235063
transform 1 0 19964 0 -1 47872
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_83_217
timestamp 1679235063
transform 1 0 21068 0 -1 47872
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_83_223
timestamp 1679235063
transform 1 0 21620 0 -1 47872
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_83_225
timestamp 1679235063
transform 1 0 21804 0 -1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_83_237
timestamp 1679235063
transform 1 0 22908 0 -1 47872
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_83_249
timestamp 1679235063
transform 1 0 24012 0 -1 47872
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_83_259
timestamp 1679235063
transform 1 0 24932 0 -1 47872
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_83_264
timestamp 1679235063
transform 1 0 25392 0 -1 47872
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_84_3
timestamp 1679235063
transform 1 0 1380 0 1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_84_15
timestamp 1679235063
transform 1 0 2484 0 1 47872
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_84_27
timestamp 1679235063
transform 1 0 3588 0 1 47872
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_84_29
timestamp 1679235063
transform 1 0 3772 0 1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_84_41
timestamp 1679235063
transform 1 0 4876 0 1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_84_53
timestamp 1679235063
transform 1 0 5980 0 1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_84_65
timestamp 1679235063
transform 1 0 7084 0 1 47872
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_84_77
timestamp 1679235063
transform 1 0 8188 0 1 47872
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_84_83
timestamp 1679235063
transform 1 0 8740 0 1 47872
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_84_85
timestamp 1679235063
transform 1 0 8924 0 1 47872
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_84_95
timestamp 1679235063
transform 1 0 9844 0 1 47872
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_84_107
timestamp 1679235063
transform 1 0 10948 0 1 47872
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_84_116
timestamp 1679235063
transform 1 0 11776 0 1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_84_128
timestamp 1679235063
transform 1 0 12880 0 1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_84_141
timestamp 1679235063
transform 1 0 14076 0 1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_84_153
timestamp 1679235063
transform 1 0 15180 0 1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_84_165
timestamp 1679235063
transform 1 0 16284 0 1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_84_177
timestamp 1679235063
transform 1 0 17388 0 1 47872
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_84_189
timestamp 1679235063
transform 1 0 18492 0 1 47872
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_84_195
timestamp 1679235063
transform 1 0 19044 0 1 47872
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_84_197
timestamp 1679235063
transform 1 0 19228 0 1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_84_209
timestamp 1679235063
transform 1 0 20332 0 1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_84_221
timestamp 1679235063
transform 1 0 21436 0 1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_84_233
timestamp 1679235063
transform 1 0 22540 0 1 47872
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_84_245
timestamp 1679235063
transform 1 0 23644 0 1 47872
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_84_251
timestamp 1679235063
transform 1 0 24196 0 1 47872
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_84_253
timestamp 1679235063
transform 1 0 24380 0 1 47872
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_84_259
timestamp 1679235063
transform 1 0 24932 0 1 47872
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_84_264
timestamp 1679235063
transform 1 0 25392 0 1 47872
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_85_3
timestamp 1679235063
transform 1 0 1380 0 -1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_85_15
timestamp 1679235063
transform 1 0 2484 0 -1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_85_27
timestamp 1679235063
transform 1 0 3588 0 -1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_85_39
timestamp 1679235063
transform 1 0 4692 0 -1 48960
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_85_51
timestamp 1679235063
transform 1 0 5796 0 -1 48960
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_85_55
timestamp 1679235063
transform 1 0 6164 0 -1 48960
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_85_57
timestamp 1679235063
transform 1 0 6348 0 -1 48960
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_85_69
timestamp 1679235063
transform 1 0 7452 0 -1 48960
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_85_93
timestamp 1679235063
transform 1 0 9660 0 -1 48960
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_85_102
timestamp 1679235063
transform 1 0 10488 0 -1 48960
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_85_110
timestamp 1679235063
transform 1 0 11224 0 -1 48960
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_85_113
timestamp 1679235063
transform 1 0 11500 0 -1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_85_125
timestamp 1679235063
transform 1 0 12604 0 -1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_85_137
timestamp 1679235063
transform 1 0 13708 0 -1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_85_149
timestamp 1679235063
transform 1 0 14812 0 -1 48960
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_85_161
timestamp 1679235063
transform 1 0 15916 0 -1 48960
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_85_167
timestamp 1679235063
transform 1 0 16468 0 -1 48960
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_85_169
timestamp 1679235063
transform 1 0 16652 0 -1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_85_181
timestamp 1679235063
transform 1 0 17756 0 -1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_85_193
timestamp 1679235063
transform 1 0 18860 0 -1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_85_205
timestamp 1679235063
transform 1 0 19964 0 -1 48960
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_85_217
timestamp 1679235063
transform 1 0 21068 0 -1 48960
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_85_223
timestamp 1679235063
transform 1 0 21620 0 -1 48960
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_85_225
timestamp 1679235063
transform 1 0 21804 0 -1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_85_237
timestamp 1679235063
transform 1 0 22908 0 -1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_85_249
timestamp 1679235063
transform 1 0 24012 0 -1 48960
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_85_261
timestamp 1679235063
transform 1 0 25116 0 -1 48960
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_86_3
timestamp 1679235063
transform 1 0 1380 0 1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_86_15
timestamp 1679235063
transform 1 0 2484 0 1 48960
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_86_27
timestamp 1679235063
transform 1 0 3588 0 1 48960
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_86_29
timestamp 1679235063
transform 1 0 3772 0 1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_86_41
timestamp 1679235063
transform 1 0 4876 0 1 48960
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_86_53
timestamp 1679235063
transform 1 0 5980 0 1 48960
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_86_59
timestamp 1679235063
transform 1 0 6532 0 1 48960
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_86_80
timestamp 1679235063
transform 1 0 8464 0 1 48960
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_86_87
timestamp 1679235063
transform 1 0 9108 0 1 48960
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_86_96
timestamp 1679235063
transform 1 0 9936 0 1 48960
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_86_100
timestamp 1679235063
transform 1 0 10304 0 1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_86_112
timestamp 1679235063
transform 1 0 11408 0 1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_86_124
timestamp 1679235063
transform 1 0 12512 0 1 48960
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_86_136
timestamp 1679235063
transform 1 0 13616 0 1 48960
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_86_141
timestamp 1679235063
transform 1 0 14076 0 1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_86_153
timestamp 1679235063
transform 1 0 15180 0 1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_86_165
timestamp 1679235063
transform 1 0 16284 0 1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_86_177
timestamp 1679235063
transform 1 0 17388 0 1 48960
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_86_189
timestamp 1679235063
transform 1 0 18492 0 1 48960
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_86_195
timestamp 1679235063
transform 1 0 19044 0 1 48960
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_86_197
timestamp 1679235063
transform 1 0 19228 0 1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_86_209
timestamp 1679235063
transform 1 0 20332 0 1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_86_221
timestamp 1679235063
transform 1 0 21436 0 1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_86_233
timestamp 1679235063
transform 1 0 22540 0 1 48960
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_86_245
timestamp 1679235063
transform 1 0 23644 0 1 48960
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_86_251
timestamp 1679235063
transform 1 0 24196 0 1 48960
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_86_253
timestamp 1679235063
transform 1 0 24380 0 1 48960
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_86_258
timestamp 1679235063
transform 1 0 24840 0 1 48960
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_86_264
timestamp 1679235063
transform 1 0 25392 0 1 48960
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_87_3
timestamp 1679235063
transform 1 0 1380 0 -1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_87_15
timestamp 1679235063
transform 1 0 2484 0 -1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_87_27
timestamp 1679235063
transform 1 0 3588 0 -1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_87_39
timestamp 1679235063
transform 1 0 4692 0 -1 50048
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_87_51
timestamp 1679235063
transform 1 0 5796 0 -1 50048
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_87_55
timestamp 1679235063
transform 1 0 6164 0 -1 50048
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_87_57
timestamp 1679235063
transform 1 0 6348 0 -1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_87_69
timestamp 1679235063
transform 1 0 7452 0 -1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_87_81
timestamp 1679235063
transform 1 0 8556 0 -1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_87_93
timestamp 1679235063
transform 1 0 9660 0 -1 50048
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_87_105
timestamp 1679235063
transform 1 0 10764 0 -1 50048
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_87_111
timestamp 1679235063
transform 1 0 11316 0 -1 50048
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_87_113
timestamp 1679235063
transform 1 0 11500 0 -1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_87_125
timestamp 1679235063
transform 1 0 12604 0 -1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_87_137
timestamp 1679235063
transform 1 0 13708 0 -1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_87_149
timestamp 1679235063
transform 1 0 14812 0 -1 50048
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_87_161
timestamp 1679235063
transform 1 0 15916 0 -1 50048
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_87_167
timestamp 1679235063
transform 1 0 16468 0 -1 50048
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_87_169
timestamp 1679235063
transform 1 0 16652 0 -1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_87_181
timestamp 1679235063
transform 1 0 17756 0 -1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_87_193
timestamp 1679235063
transform 1 0 18860 0 -1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_87_205
timestamp 1679235063
transform 1 0 19964 0 -1 50048
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_87_217
timestamp 1679235063
transform 1 0 21068 0 -1 50048
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_87_223
timestamp 1679235063
transform 1 0 21620 0 -1 50048
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_87_225
timestamp 1679235063
transform 1 0 21804 0 -1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_87_237
timestamp 1679235063
transform 1 0 22908 0 -1 50048
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_87_249
timestamp 1679235063
transform 1 0 24012 0 -1 50048
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_87_253
timestamp 1679235063
transform 1 0 24380 0 -1 50048
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_87_264
timestamp 1679235063
transform 1 0 25392 0 -1 50048
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_88_3
timestamp 1679235063
transform 1 0 1380 0 1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_88_15
timestamp 1679235063
transform 1 0 2484 0 1 50048
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_88_27
timestamp 1679235063
transform 1 0 3588 0 1 50048
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_88_29
timestamp 1679235063
transform 1 0 3772 0 1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_88_41
timestamp 1679235063
transform 1 0 4876 0 1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_88_53
timestamp 1679235063
transform 1 0 5980 0 1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_88_65
timestamp 1679235063
transform 1 0 7084 0 1 50048
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_88_77
timestamp 1679235063
transform 1 0 8188 0 1 50048
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_88_83
timestamp 1679235063
transform 1 0 8740 0 1 50048
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_88_85
timestamp 1679235063
transform 1 0 8924 0 1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_88_97
timestamp 1679235063
transform 1 0 10028 0 1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_88_109
timestamp 1679235063
transform 1 0 11132 0 1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_88_121
timestamp 1679235063
transform 1 0 12236 0 1 50048
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_88_133
timestamp 1679235063
transform 1 0 13340 0 1 50048
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_88_139
timestamp 1679235063
transform 1 0 13892 0 1 50048
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_88_141
timestamp 1679235063
transform 1 0 14076 0 1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_88_153
timestamp 1679235063
transform 1 0 15180 0 1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_88_165
timestamp 1679235063
transform 1 0 16284 0 1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_88_177
timestamp 1679235063
transform 1 0 17388 0 1 50048
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_88_189
timestamp 1679235063
transform 1 0 18492 0 1 50048
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_88_195
timestamp 1679235063
transform 1 0 19044 0 1 50048
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_88_197
timestamp 1679235063
transform 1 0 19228 0 1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_88_209
timestamp 1679235063
transform 1 0 20332 0 1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_88_221
timestamp 1679235063
transform 1 0 21436 0 1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_88_233
timestamp 1679235063
transform 1 0 22540 0 1 50048
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_88_245
timestamp 1679235063
transform 1 0 23644 0 1 50048
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_88_251
timestamp 1679235063
transform 1 0 24196 0 1 50048
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_88_253
timestamp 1679235063
transform 1 0 24380 0 1 50048
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_88_261
timestamp 1679235063
transform 1 0 25116 0 1 50048
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_89_3
timestamp 1679235063
transform 1 0 1380 0 -1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_89_15
timestamp 1679235063
transform 1 0 2484 0 -1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_89_27
timestamp 1679235063
transform 1 0 3588 0 -1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_89_39
timestamp 1679235063
transform 1 0 4692 0 -1 51136
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_89_51
timestamp 1679235063
transform 1 0 5796 0 -1 51136
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_89_55
timestamp 1679235063
transform 1 0 6164 0 -1 51136
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_89_57
timestamp 1679235063
transform 1 0 6348 0 -1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_89_69
timestamp 1679235063
transform 1 0 7452 0 -1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_89_81
timestamp 1679235063
transform 1 0 8556 0 -1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_89_93
timestamp 1679235063
transform 1 0 9660 0 -1 51136
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_89_105
timestamp 1679235063
transform 1 0 10764 0 -1 51136
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_89_111
timestamp 1679235063
transform 1 0 11316 0 -1 51136
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_89_113
timestamp 1679235063
transform 1 0 11500 0 -1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_89_125
timestamp 1679235063
transform 1 0 12604 0 -1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_89_137
timestamp 1679235063
transform 1 0 13708 0 -1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_89_149
timestamp 1679235063
transform 1 0 14812 0 -1 51136
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_89_161
timestamp 1679235063
transform 1 0 15916 0 -1 51136
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_89_167
timestamp 1679235063
transform 1 0 16468 0 -1 51136
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_89_169
timestamp 1679235063
transform 1 0 16652 0 -1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_89_181
timestamp 1679235063
transform 1 0 17756 0 -1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_89_193
timestamp 1679235063
transform 1 0 18860 0 -1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_89_205
timestamp 1679235063
transform 1 0 19964 0 -1 51136
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_89_217
timestamp 1679235063
transform 1 0 21068 0 -1 51136
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_89_223
timestamp 1679235063
transform 1 0 21620 0 -1 51136
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_89_225
timestamp 1679235063
transform 1 0 21804 0 -1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_89_237
timestamp 1679235063
transform 1 0 22908 0 -1 51136
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_89_249
timestamp 1679235063
transform 1 0 24012 0 -1 51136
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_89_253
timestamp 1679235063
transform 1 0 24380 0 -1 51136
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_89_256
timestamp 1679235063
transform 1 0 24656 0 -1 51136
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_89_264
timestamp 1679235063
transform 1 0 25392 0 -1 51136
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_90_3
timestamp 1679235063
transform 1 0 1380 0 1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_90_15
timestamp 1679235063
transform 1 0 2484 0 1 51136
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_90_27
timestamp 1679235063
transform 1 0 3588 0 1 51136
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_90_29
timestamp 1679235063
transform 1 0 3772 0 1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_90_41
timestamp 1679235063
transform 1 0 4876 0 1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_90_53
timestamp 1679235063
transform 1 0 5980 0 1 51136
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_90_65
timestamp 1679235063
transform 1 0 7084 0 1 51136
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_90_69
timestamp 1679235063
transform 1 0 7452 0 1 51136
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_90_77
timestamp 1679235063
transform 1 0 8188 0 1 51136
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_90_81
timestamp 1679235063
transform 1 0 8556 0 1 51136
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_90_85
timestamp 1679235063
transform 1 0 8924 0 1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_90_97
timestamp 1679235063
transform 1 0 10028 0 1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_90_109
timestamp 1679235063
transform 1 0 11132 0 1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_90_121
timestamp 1679235063
transform 1 0 12236 0 1 51136
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_90_133
timestamp 1679235063
transform 1 0 13340 0 1 51136
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_90_139
timestamp 1679235063
transform 1 0 13892 0 1 51136
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_90_141
timestamp 1679235063
transform 1 0 14076 0 1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_90_153
timestamp 1679235063
transform 1 0 15180 0 1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_90_165
timestamp 1679235063
transform 1 0 16284 0 1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_90_177
timestamp 1679235063
transform 1 0 17388 0 1 51136
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_90_189
timestamp 1679235063
transform 1 0 18492 0 1 51136
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_90_195
timestamp 1679235063
transform 1 0 19044 0 1 51136
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_90_197
timestamp 1679235063
transform 1 0 19228 0 1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_90_209
timestamp 1679235063
transform 1 0 20332 0 1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_90_221
timestamp 1679235063
transform 1 0 21436 0 1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_90_233
timestamp 1679235063
transform 1 0 22540 0 1 51136
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_90_245
timestamp 1679235063
transform 1 0 23644 0 1 51136
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_90_251
timestamp 1679235063
transform 1 0 24196 0 1 51136
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_90_253
timestamp 1679235063
transform 1 0 24380 0 1 51136
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_90_257
timestamp 1679235063
transform 1 0 24748 0 1 51136
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_90_264
timestamp 1679235063
transform 1 0 25392 0 1 51136
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_91_3
timestamp 1679235063
transform 1 0 1380 0 -1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_91_15
timestamp 1679235063
transform 1 0 2484 0 -1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_91_27
timestamp 1679235063
transform 1 0 3588 0 -1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_91_39
timestamp 1679235063
transform 1 0 4692 0 -1 52224
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_91_51
timestamp 1679235063
transform 1 0 5796 0 -1 52224
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_91_55
timestamp 1679235063
transform 1 0 6164 0 -1 52224
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_91_57
timestamp 1679235063
transform 1 0 6348 0 -1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_91_69
timestamp 1679235063
transform 1 0 7452 0 -1 52224
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_91_81
timestamp 1679235063
transform 1 0 8556 0 -1 52224
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_91_86
timestamp 1679235063
transform 1 0 9016 0 -1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_91_98
timestamp 1679235063
transform 1 0 10120 0 -1 52224
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_91_110
timestamp 1679235063
transform 1 0 11224 0 -1 52224
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_91_113
timestamp 1679235063
transform 1 0 11500 0 -1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_91_125
timestamp 1679235063
transform 1 0 12604 0 -1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_91_137
timestamp 1679235063
transform 1 0 13708 0 -1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_91_149
timestamp 1679235063
transform 1 0 14812 0 -1 52224
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_91_161
timestamp 1679235063
transform 1 0 15916 0 -1 52224
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_91_167
timestamp 1679235063
transform 1 0 16468 0 -1 52224
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_91_169
timestamp 1679235063
transform 1 0 16652 0 -1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_91_181
timestamp 1679235063
transform 1 0 17756 0 -1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_91_193
timestamp 1679235063
transform 1 0 18860 0 -1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_91_205
timestamp 1679235063
transform 1 0 19964 0 -1 52224
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_91_217
timestamp 1679235063
transform 1 0 21068 0 -1 52224
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_91_223
timestamp 1679235063
transform 1 0 21620 0 -1 52224
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_91_225
timestamp 1679235063
transform 1 0 21804 0 -1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_91_237
timestamp 1679235063
transform 1 0 22908 0 -1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_91_249
timestamp 1679235063
transform 1 0 24012 0 -1 52224
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_91_261
timestamp 1679235063
transform 1 0 25116 0 -1 52224
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_92_3
timestamp 1679235063
transform 1 0 1380 0 1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_92_15
timestamp 1679235063
transform 1 0 2484 0 1 52224
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_92_27
timestamp 1679235063
transform 1 0 3588 0 1 52224
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_92_29
timestamp 1679235063
transform 1 0 3772 0 1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_92_41
timestamp 1679235063
transform 1 0 4876 0 1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_92_53
timestamp 1679235063
transform 1 0 5980 0 1 52224
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_92_65
timestamp 1679235063
transform 1 0 7084 0 1 52224
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_92_74
timestamp 1679235063
transform 1 0 7912 0 1 52224
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_92_82
timestamp 1679235063
transform 1 0 8648 0 1 52224
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_92_85
timestamp 1679235063
transform 1 0 8924 0 1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_92_97
timestamp 1679235063
transform 1 0 10028 0 1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_92_109
timestamp 1679235063
transform 1 0 11132 0 1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_92_121
timestamp 1679235063
transform 1 0 12236 0 1 52224
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_92_133
timestamp 1679235063
transform 1 0 13340 0 1 52224
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_92_139
timestamp 1679235063
transform 1 0 13892 0 1 52224
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_92_141
timestamp 1679235063
transform 1 0 14076 0 1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_92_153
timestamp 1679235063
transform 1 0 15180 0 1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_92_165
timestamp 1679235063
transform 1 0 16284 0 1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_92_177
timestamp 1679235063
transform 1 0 17388 0 1 52224
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_92_189
timestamp 1679235063
transform 1 0 18492 0 1 52224
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_92_195
timestamp 1679235063
transform 1 0 19044 0 1 52224
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_92_197
timestamp 1679235063
transform 1 0 19228 0 1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_92_209
timestamp 1679235063
transform 1 0 20332 0 1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_92_221
timestamp 1679235063
transform 1 0 21436 0 1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_92_233
timestamp 1679235063
transform 1 0 22540 0 1 52224
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_92_245
timestamp 1679235063
transform 1 0 23644 0 1 52224
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_92_251
timestamp 1679235063
transform 1 0 24196 0 1 52224
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_92_253
timestamp 1679235063
transform 1 0 24380 0 1 52224
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_92_256
timestamp 1679235063
transform 1 0 24656 0 1 52224
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_92_264
timestamp 1679235063
transform 1 0 25392 0 1 52224
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_93_3
timestamp 1679235063
transform 1 0 1380 0 -1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_93_15
timestamp 1679235063
transform 1 0 2484 0 -1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_93_27
timestamp 1679235063
transform 1 0 3588 0 -1 53312
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_93_39
timestamp 1679235063
transform 1 0 4692 0 -1 53312
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_93_45
timestamp 1679235063
transform 1 0 5244 0 -1 53312
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_93_53
timestamp 1679235063
transform 1 0 5980 0 -1 53312
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_93_57
timestamp 1679235063
transform 1 0 6348 0 -1 53312
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_93_62
timestamp 1679235063
transform 1 0 6808 0 -1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_93_74
timestamp 1679235063
transform 1 0 7912 0 -1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_93_86
timestamp 1679235063
transform 1 0 9016 0 -1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_93_98
timestamp 1679235063
transform 1 0 10120 0 -1 53312
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_93_110
timestamp 1679235063
transform 1 0 11224 0 -1 53312
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_93_113
timestamp 1679235063
transform 1 0 11500 0 -1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_93_125
timestamp 1679235063
transform 1 0 12604 0 -1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_93_137
timestamp 1679235063
transform 1 0 13708 0 -1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_93_149
timestamp 1679235063
transform 1 0 14812 0 -1 53312
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_93_161
timestamp 1679235063
transform 1 0 15916 0 -1 53312
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_93_167
timestamp 1679235063
transform 1 0 16468 0 -1 53312
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_93_169
timestamp 1679235063
transform 1 0 16652 0 -1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_93_181
timestamp 1679235063
transform 1 0 17756 0 -1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_93_193
timestamp 1679235063
transform 1 0 18860 0 -1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_93_205
timestamp 1679235063
transform 1 0 19964 0 -1 53312
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_93_217
timestamp 1679235063
transform 1 0 21068 0 -1 53312
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_93_223
timestamp 1679235063
transform 1 0 21620 0 -1 53312
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_93_225
timestamp 1679235063
transform 1 0 21804 0 -1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_93_237
timestamp 1679235063
transform 1 0 22908 0 -1 53312
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_93_249
timestamp 1679235063
transform 1 0 24012 0 -1 53312
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_93_255
timestamp 1679235063
transform 1 0 24564 0 -1 53312
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_93_258
timestamp 1679235063
transform 1 0 24840 0 -1 53312
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_93_264
timestamp 1679235063
transform 1 0 25392 0 -1 53312
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_94_3
timestamp 1679235063
transform 1 0 1380 0 1 53312
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_94_21
timestamp 1679235063
transform 1 0 3036 0 1 53312
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_94_27
timestamp 1679235063
transform 1 0 3588 0 1 53312
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_94_29
timestamp 1679235063
transform 1 0 3772 0 1 53312
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_94_41
timestamp 1679235063
transform 1 0 4876 0 1 53312
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_94_61
timestamp 1679235063
transform 1 0 6716 0 1 53312
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_94_73
timestamp 1679235063
transform 1 0 7820 0 1 53312
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_94_81
timestamp 1679235063
transform 1 0 8556 0 1 53312
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_94_85
timestamp 1679235063
transform 1 0 8924 0 1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_94_97
timestamp 1679235063
transform 1 0 10028 0 1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_94_109
timestamp 1679235063
transform 1 0 11132 0 1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_94_121
timestamp 1679235063
transform 1 0 12236 0 1 53312
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_94_133
timestamp 1679235063
transform 1 0 13340 0 1 53312
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_94_139
timestamp 1679235063
transform 1 0 13892 0 1 53312
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_94_141
timestamp 1679235063
transform 1 0 14076 0 1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_94_153
timestamp 1679235063
transform 1 0 15180 0 1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_94_165
timestamp 1679235063
transform 1 0 16284 0 1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_94_177
timestamp 1679235063
transform 1 0 17388 0 1 53312
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_94_189
timestamp 1679235063
transform 1 0 18492 0 1 53312
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_94_195
timestamp 1679235063
transform 1 0 19044 0 1 53312
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_94_197
timestamp 1679235063
transform 1 0 19228 0 1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_94_209
timestamp 1679235063
transform 1 0 20332 0 1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_94_221
timestamp 1679235063
transform 1 0 21436 0 1 53312
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_94_233
timestamp 1679235063
transform 1 0 22540 0 1 53312
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_94_241
timestamp 1679235063
transform 1 0 23276 0 1 53312
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_94_244
timestamp 1679235063
transform 1 0 23552 0 1 53312
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_94_250
timestamp 1679235063
transform 1 0 24104 0 1 53312
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_94_255
timestamp 1679235063
transform 1 0 24564 0 1 53312
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_94_258
timestamp 1679235063
transform 1 0 24840 0 1 53312
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_94_264
timestamp 1679235063
transform 1 0 25392 0 1 53312
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_95_3
timestamp 1679235063
transform 1 0 1380 0 -1 54400
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_95_9
timestamp 1679235063
transform 1 0 1932 0 -1 54400
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_95_26
timestamp 1679235063
transform 1 0 3496 0 -1 54400
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_95_29
timestamp 1679235063
transform 1 0 3772 0 -1 54400
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_95_47
timestamp 1679235063
transform 1 0 5428 0 -1 54400
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_95_55
timestamp 1679235063
transform 1 0 6164 0 -1 54400
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_95_57
timestamp 1679235063
transform 1 0 6348 0 -1 54400
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_95_76
timestamp 1679235063
transform 1 0 8096 0 -1 54400
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_95_85
timestamp 1679235063
transform 1 0 8924 0 -1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_95_97
timestamp 1679235063
transform 1 0 10028 0 -1 54400
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_95_109
timestamp 1679235063
transform 1 0 11132 0 -1 54400
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_95_113
timestamp 1679235063
transform 1 0 11500 0 -1 54400
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_95_125
timestamp 1679235063
transform 1 0 12604 0 -1 54400
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_95_133
timestamp 1679235063
transform 1 0 13340 0 -1 54400
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_95_138
timestamp 1679235063
transform 1 0 13800 0 -1 54400
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_95_143
timestamp 1679235063
transform 1 0 14260 0 -1 54400
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_95_149
timestamp 1679235063
transform 1 0 14812 0 -1 54400
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_95_153
timestamp 1679235063
transform 1 0 15180 0 -1 54400
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_95_157
timestamp 1679235063
transform 1 0 15548 0 -1 54400
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_95_165
timestamp 1679235063
transform 1 0 16284 0 -1 54400
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_95_169
timestamp 1679235063
transform 1 0 16652 0 -1 54400
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_95_174
timestamp 1679235063
transform 1 0 17112 0 -1 54400
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_95_178
timestamp 1679235063
transform 1 0 17480 0 -1 54400
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_95_183
timestamp 1679235063
transform 1 0 17940 0 -1 54400
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_95_187
timestamp 1679235063
transform 1 0 18308 0 -1 54400
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_95_193
timestamp 1679235063
transform 1 0 18860 0 -1 54400
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_95_197
timestamp 1679235063
transform 1 0 19228 0 -1 54400
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_95_209
timestamp 1679235063
transform 1 0 20332 0 -1 54400
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_95_221
timestamp 1679235063
transform 1 0 21436 0 -1 54400
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_95_225
timestamp 1679235063
transform 1 0 21804 0 -1 54400
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_95_237
timestamp 1679235063
transform 1 0 22908 0 -1 54400
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_95_242
timestamp 1679235063
transform 1 0 23368 0 -1 54400
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_95_250
timestamp 1679235063
transform 1 0 24104 0 -1 54400
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_95_255
timestamp 1679235063
transform 1 0 24564 0 -1 54400
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_95_258
timestamp 1679235063
transform 1 0 24840 0 -1 54400
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_95_264
timestamp 1679235063
transform 1 0 25392 0 -1 54400
box -38 -48 222 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold1 pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1679235063
transform 1 0 24564 0 1 30464
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold2
timestamp 1679235063
transform 1 0 18124 0 -1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold3
timestamp 1679235063
transform 1 0 18676 0 -1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold4
timestamp 1679235063
transform 1 0 21988 0 -1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold5
timestamp 1679235063
transform 1 0 19044 0 -1 31552
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold6
timestamp 1679235063
transform 1 0 21528 0 1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold7
timestamp 1679235063
transform 1 0 14352 0 -1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold8
timestamp 1679235063
transform 1 0 21988 0 -1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold9
timestamp 1679235063
transform 1 0 20792 0 -1 34816
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold10
timestamp 1679235063
transform 1 0 9108 0 1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold11
timestamp 1679235063
transform 1 0 19412 0 -1 34816
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold12
timestamp 1679235063
transform 1 0 24656 0 1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold13
timestamp 1679235063
transform 1 0 11868 0 -1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold14
timestamp 1679235063
transform 1 0 21988 0 -1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold15
timestamp 1679235063
transform 1 0 14260 0 1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold16
timestamp 1679235063
transform 1 0 21988 0 -1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold17
timestamp 1679235063
transform 1 0 19504 0 -1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold18
timestamp 1679235063
transform 1 0 13064 0 1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold19
timestamp 1679235063
transform 1 0 14996 0 -1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold20
timestamp 1679235063
transform 1 0 17020 0 -1 31552
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold21
timestamp 1679235063
transform 1 0 9384 0 -1 33728
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold22
timestamp 1679235063
transform 1 0 17296 0 -1 30464
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold23
timestamp 1679235063
transform 1 0 11684 0 -1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold24
timestamp 1679235063
transform 1 0 11684 0 -1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold25
timestamp 1679235063
transform 1 0 11684 0 -1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold26
timestamp 1679235063
transform 1 0 16836 0 -1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold27
timestamp 1679235063
transform 1 0 9108 0 1 47872
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold28
timestamp 1679235063
transform 1 0 10580 0 1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold29
timestamp 1679235063
transform 1 0 15640 0 -1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold30
timestamp 1679235063
transform 1 0 9936 0 1 44608
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold31
timestamp 1679235063
transform 1 0 24656 0 -1 31552
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold32
timestamp 1679235063
transform 1 0 19412 0 1 30464
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold33
timestamp 1679235063
transform 1 0 19596 0 1 34816
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold34
timestamp 1679235063
transform 1 0 14444 0 -1 30464
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold35
timestamp 1679235063
transform 1 0 20792 0 1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold36
timestamp 1679235063
transform 1 0 19688 0 1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold37
timestamp 1679235063
transform 1 0 17112 0 1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold38
timestamp 1679235063
transform 1 0 23092 0 -1 34816
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold39
timestamp 1679235063
transform 1 0 17940 0 1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold40
timestamp 1679235063
transform 1 0 18216 0 1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold41
timestamp 1679235063
transform 1 0 14352 0 1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold42
timestamp 1679235063
transform 1 0 21528 0 1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold43
timestamp 1679235063
transform 1 0 14536 0 -1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold44
timestamp 1679235063
transform 1 0 24564 0 1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold45
timestamp 1679235063
transform 1 0 24564 0 1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold46
timestamp 1679235063
transform 1 0 21988 0 -1 34816
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold47
timestamp 1679235063
transform 1 0 12420 0 1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold48
timestamp 1679235063
transform 1 0 9292 0 1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold49
timestamp 1679235063
transform 1 0 11684 0 -1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold50
timestamp 1679235063
transform 1 0 24564 0 1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold51
timestamp 1679235063
transform 1 0 22816 0 1 31552
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold52
timestamp 1679235063
transform 1 0 24564 0 -1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold53
timestamp 1679235063
transform 1 0 22908 0 1 30464
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold54
timestamp 1679235063
transform 1 0 11684 0 -1 40256
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold55
timestamp 1679235063
transform 1 0 24564 0 1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold56
timestamp 1679235063
transform 1 0 24472 0 -1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold57
timestamp 1679235063
transform 1 0 22448 0 -1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold58
timestamp 1679235063
transform 1 0 12880 0 -1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold59
timestamp 1679235063
transform 1 0 18584 0 -1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold60
timestamp 1679235063
transform 1 0 18124 0 1 32640
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold61
timestamp 1679235063
transform 1 0 24564 0 1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold62
timestamp 1679235063
transform 1 0 7912 0 1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold63
timestamp 1679235063
transform 1 0 24564 0 1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold64
timestamp 1679235063
transform 1 0 20792 0 -1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold65
timestamp 1679235063
transform 1 0 13064 0 1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold66
timestamp 1679235063
transform 1 0 24564 0 1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold67
timestamp 1679235063
transform 1 0 20700 0 1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold68
timestamp 1679235063
transform 1 0 10488 0 -1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold69
timestamp 1679235063
transform 1 0 24564 0 1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold70
timestamp 1679235063
transform 1 0 24564 0 1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold71
timestamp 1679235063
transform 1 0 7912 0 1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold72
timestamp 1679235063
transform 1 0 12788 0 1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold73
timestamp 1679235063
transform 1 0 19228 0 -1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold74
timestamp 1679235063
transform 1 0 12788 0 1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold75
timestamp 1679235063
transform 1 0 24564 0 1 33728
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold76
timestamp 1679235063
transform 1 0 7820 0 -1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold77
timestamp 1679235063
transform 1 0 9476 0 1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold78
timestamp 1679235063
transform 1 0 16836 0 -1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold79
timestamp 1679235063
transform 1 0 23092 0 1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold80
timestamp 1679235063
transform 1 0 19412 0 1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold81
timestamp 1679235063
transform 1 0 15548 0 -1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold82
timestamp 1679235063
transform 1 0 24564 0 1 31552
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold83
timestamp 1679235063
transform 1 0 6716 0 -1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold84
timestamp 1679235063
transform 1 0 6624 0 -1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold85
timestamp 1679235063
transform 1 0 24656 0 1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold86
timestamp 1679235063
transform 1 0 24564 0 1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold87
timestamp 1679235063
transform 1 0 24564 0 1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold88
timestamp 1679235063
transform 1 0 11684 0 -1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold89
timestamp 1679235063
transform 1 0 14352 0 -1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold90
timestamp 1679235063
transform 1 0 6900 0 -1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold91
timestamp 1679235063
transform 1 0 9476 0 1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold92
timestamp 1679235063
transform 1 0 10488 0 -1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold93
timestamp 1679235063
transform 1 0 22448 0 -1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold94
timestamp 1679235063
transform 1 0 10488 0 -1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold95
timestamp 1679235063
transform 1 0 21988 0 -1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold96
timestamp 1679235063
transform 1 0 7912 0 1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold97
timestamp 1679235063
transform 1 0 10488 0 -1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold98
timestamp 1679235063
transform 1 0 19412 0 1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold99
timestamp 1679235063
transform 1 0 11868 0 -1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold100
timestamp 1679235063
transform 1 0 15456 0 -1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold101
timestamp 1679235063
transform 1 0 17572 0 1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s50_1  hold102 pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1679235063
transform 1 0 17664 0 1 38080
box -38 -48 774 592
use sky130_fd_sc_hd__clkbuf_1  input1
timestamp 1679235063
transform 1 0 23092 0 -1 54400
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input2
timestamp 1679235063
transform 1 0 1564 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input3
timestamp 1679235063
transform 1 0 22540 0 1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input4
timestamp 1679235063
transform 1 0 25116 0 -1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input5
timestamp 1679235063
transform 1 0 25116 0 1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input6
timestamp 1679235063
transform 1 0 25116 0 1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  input7
timestamp 1679235063
transform 1 0 25024 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input8
timestamp 1679235063
transform 1 0 25024 0 -1 38080
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  input9
timestamp 1679235063
transform 1 0 25116 0 1 38080
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input10
timestamp 1679235063
transform 1 0 25116 0 1 39168
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input11
timestamp 1679235063
transform 1 0 25116 0 -1 40256
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input12
timestamp 1679235063
transform 1 0 25116 0 -1 41344
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  input13
timestamp 1679235063
transform 1 0 25024 0 1 41344
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  input14
timestamp 1679235063
transform 1 0 16836 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  input15
timestamp 1679235063
transform 1 0 25024 0 1 42432
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input16
timestamp 1679235063
transform 1 0 25024 0 -1 43520
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input17
timestamp 1679235063
transform 1 0 25024 0 -1 44608
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  input18
timestamp 1679235063
transform 1 0 25116 0 1 44608
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input19
timestamp 1679235063
transform 1 0 25116 0 1 45696
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input20
timestamp 1679235063
transform 1 0 25116 0 -1 46784
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input21
timestamp 1679235063
transform 1 0 25116 0 -1 47872
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  input22
timestamp 1679235063
transform 1 0 25024 0 1 47872
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input23
timestamp 1679235063
transform 1 0 25024 0 1 48960
box -38 -48 406 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input24
timestamp 1679235063
transform 1 0 24472 0 -1 50048
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_1  input25
timestamp 1679235063
transform 1 0 17480 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input26
timestamp 1679235063
transform 1 0 18676 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input27
timestamp 1679235063
transform 1 0 23828 0 1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input28
timestamp 1679235063
transform 1 0 25116 0 -1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input29
timestamp 1679235063
transform 1 0 25116 0 1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input30
timestamp 1679235063
transform 1 0 25116 0 -1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input31
timestamp 1679235063
transform 1 0 25116 0 1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input32
timestamp 1679235063
transform 1 0 24472 0 -1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input33
timestamp 1679235063
transform 1 0 2208 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input34
timestamp 1679235063
transform 1 0 5152 0 1 2176
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_1  input35
timestamp 1679235063
transform 1 0 4508 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input36
timestamp 1679235063
transform 1 0 6348 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input37
timestamp 1679235063
transform 1 0 6532 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input38
timestamp 1679235063
transform 1 0 7084 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input39
timestamp 1679235063
transform 1 0 7176 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input40
timestamp 1679235063
transform 1 0 7820 0 -1 3264
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_1  input41
timestamp 1679235063
transform 1 0 7084 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input42
timestamp 1679235063
transform 1 0 8372 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input43
timestamp 1679235063
transform 1 0 6532 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input44
timestamp 1679235063
transform 1 0 2852 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input45
timestamp 1679235063
transform 1 0 9292 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input46
timestamp 1679235063
transform 1 0 9108 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input47
timestamp 1679235063
transform 1 0 9660 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input48
timestamp 1679235063
transform 1 0 7728 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input49
timestamp 1679235063
transform 1 0 9660 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input50
timestamp 1679235063
transform 1 0 8372 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input51
timestamp 1679235063
transform 1 0 11684 0 -1 3264
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_1  input52
timestamp 1679235063
transform 1 0 10948 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input53
timestamp 1679235063
transform 1 0 10304 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input54
timestamp 1679235063
transform 1 0 10304 0 1 2176
box -38 -48 958 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input55
timestamp 1679235063
transform 1 0 2116 0 -1 3264
box -38 -48 958 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input56
timestamp 1679235063
transform 1 0 2576 0 1 2176
box -38 -48 958 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input57
timestamp 1679235063
transform 1 0 3404 0 -1 3264
box -38 -48 958 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input58
timestamp 1679235063
transform 1 0 1564 0 1 3264
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_1  input59
timestamp 1679235063
transform 1 0 4140 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input60
timestamp 1679235063
transform 1 0 4232 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input61
timestamp 1679235063
transform 1 0 4876 0 1 3264
box -38 -48 958 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input62
timestamp 1679235063
transform 1 0 5152 0 -1 3264
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_1  input63
timestamp 1679235063
transform 1 0 13524 0 -1 54400
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input64
timestamp 1679235063
transform 1 0 14904 0 -1 54400
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input65
timestamp 1679235063
transform 1 0 16836 0 -1 54400
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input66
timestamp 1679235063
transform 1 0 17664 0 -1 54400
box -38 -48 314 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input67
timestamp 1679235063
transform 1 0 19412 0 -1 54400
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_16  input68
timestamp 1679235063
transform 1 0 23552 0 -1 3264
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_4  input69 pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1679235063
transform 1 0 24840 0 -1 51136
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  input70
timestamp 1679235063
transform 1 0 24840 0 1 51136
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  input71
timestamp 1679235063
transform 1 0 24840 0 1 52224
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  input72 pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1679235063
transform 1 0 25024 0 -1 53312
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  input73
timestamp 1679235063
transform 1 0 25024 0 -1 54400
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  input74
timestamp 1679235063
transform 1 0 25024 0 1 53312
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  input75
timestamp 1679235063
transform 1 0 23736 0 -1 54400
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input76
timestamp 1679235063
transform 1 0 23736 0 1 53312
box -38 -48 406 592
use sky130_fd_sc_hd__buf_12  output77 pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1679235063
transform 1 0 12328 0 1 3264
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output78
timestamp 1679235063
transform 1 0 1564 0 1 53312
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output79
timestamp 1679235063
transform 1 0 20792 0 1 8704
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output80
timestamp 1679235063
transform 1 0 22080 0 -1 9792
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output81
timestamp 1679235063
transform 1 0 23920 0 -1 9792
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output82
timestamp 1679235063
transform 1 0 23920 0 -1 10880
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output83
timestamp 1679235063
transform 1 0 22632 0 1 11968
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output84
timestamp 1679235063
transform 1 0 22632 0 1 13056
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output85
timestamp 1679235063
transform 1 0 22080 0 -1 14144
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output86
timestamp 1679235063
transform 1 0 23920 0 -1 14144
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output87
timestamp 1679235063
transform 1 0 23920 0 -1 15232
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output88
timestamp 1679235063
transform 1 0 22632 0 1 16320
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output89
timestamp 1679235063
transform 1 0 22080 0 -1 17408
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output90
timestamp 1679235063
transform 1 0 15640 0 1 5440
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output91
timestamp 1679235063
transform 1 0 22632 0 1 17408
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output92
timestamp 1679235063
transform 1 0 23920 0 -1 17408
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output93
timestamp 1679235063
transform 1 0 22632 0 1 18496
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output94
timestamp 1679235063
transform 1 0 20056 0 -1 20672
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output95
timestamp 1679235063
transform 1 0 20056 0 -1 21760
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output96
timestamp 1679235063
transform 1 0 22632 0 1 20672
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output97
timestamp 1679235063
transform 1 0 22080 0 -1 22848
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output98
timestamp 1679235063
transform 1 0 22632 0 1 22848
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output99
timestamp 1679235063
transform 1 0 23920 0 -1 22848
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output100
timestamp 1679235063
transform 1 0 22632 0 1 25024
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output101
timestamp 1679235063
transform 1 0 17480 0 1 6528
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output102
timestamp 1679235063
transform 1 0 18216 0 -1 7616
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output103
timestamp 1679235063
transform 1 0 20056 0 -1 7616
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output104
timestamp 1679235063
transform 1 0 22080 0 -1 7616
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output105
timestamp 1679235063
transform 1 0 23920 0 -1 5440
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output106
timestamp 1679235063
transform 1 0 23920 0 -1 6528
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output107
timestamp 1679235063
transform 1 0 23920 0 -1 7616
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output108
timestamp 1679235063
transform 1 0 22632 0 1 8704
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output109
timestamp 1679235063
transform 1 0 12972 0 -1 4352
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output110
timestamp 1679235063
transform 1 0 18676 0 -1 3264
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output111
timestamp 1679235063
transform 1 0 19412 0 1 2176
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output112
timestamp 1679235063
transform 1 0 17388 0 1 4352
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output113
timestamp 1679235063
transform 1 0 19412 0 1 3264
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output114
timestamp 1679235063
transform 1 0 18676 0 -1 4352
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output115
timestamp 1679235063
transform 1 0 21988 0 1 2176
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output116
timestamp 1679235063
transform 1 0 19412 0 1 4352
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output117
timestamp 1679235063
transform 1 0 21252 0 1 3264
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output118
timestamp 1679235063
transform 1 0 21252 0 1 4352
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output119
timestamp 1679235063
transform 1 0 21988 0 -1 4352
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output120
timestamp 1679235063
transform 1 0 12328 0 1 2176
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output121
timestamp 1679235063
transform 1 0 20332 0 1 5440
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output122
timestamp 1679235063
transform 1 0 21988 0 -1 5440
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output123
timestamp 1679235063
transform 1 0 23828 0 -1 4352
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output124
timestamp 1679235063
transform 1 0 22172 0 1 5440
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output125
timestamp 1679235063
transform 1 0 21988 0 -1 6528
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output126
timestamp 1679235063
transform 1 0 22172 0 1 7616
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output127
timestamp 1679235063
transform 1 0 20056 0 -1 6528
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output128
timestamp 1679235063
transform 1 0 17480 0 1 5440
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output129
timestamp 1679235063
transform 1 0 14904 0 -1 4352
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output130
timestamp 1679235063
transform 1 0 20332 0 1 7616
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output131
timestamp 1679235063
transform 1 0 12972 0 -1 3264
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output132
timestamp 1679235063
transform 1 0 14260 0 1 3264
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output133
timestamp 1679235063
transform 1 0 14444 0 1 2176
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output134
timestamp 1679235063
transform 1 0 14812 0 -1 3264
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output135
timestamp 1679235063
transform 1 0 16836 0 1 2176
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output136
timestamp 1679235063
transform 1 0 16100 0 1 3264
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output137
timestamp 1679235063
transform 1 0 16836 0 -1 3264
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output138
timestamp 1679235063
transform 1 0 16836 0 -1 4352
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output139
timestamp 1679235063
transform 1 0 2024 0 -1 54400
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output140
timestamp 1679235063
transform 1 0 3956 0 -1 54400
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output141
timestamp 1679235063
transform 1 0 5244 0 1 53312
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output142
timestamp 1679235063
transform 1 0 6624 0 -1 54400
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_3  PHY_0
timestamp 1679235063
transform 1 0 1104 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_1
timestamp 1679235063
transform -1 0 25852 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_2
timestamp 1679235063
transform 1 0 1104 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_3
timestamp 1679235063
transform -1 0 25852 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_4
timestamp 1679235063
transform 1 0 1104 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_5
timestamp 1679235063
transform -1 0 25852 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_6
timestamp 1679235063
transform 1 0 1104 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_7
timestamp 1679235063
transform -1 0 25852 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_8
timestamp 1679235063
transform 1 0 1104 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_9
timestamp 1679235063
transform -1 0 25852 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_10
timestamp 1679235063
transform 1 0 1104 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_11
timestamp 1679235063
transform -1 0 25852 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_12
timestamp 1679235063
transform 1 0 1104 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_13
timestamp 1679235063
transform -1 0 25852 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_14
timestamp 1679235063
transform 1 0 1104 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_15
timestamp 1679235063
transform -1 0 25852 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_16
timestamp 1679235063
transform 1 0 1104 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_17
timestamp 1679235063
transform -1 0 25852 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_18
timestamp 1679235063
transform 1 0 1104 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_19
timestamp 1679235063
transform -1 0 25852 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_20
timestamp 1679235063
transform 1 0 1104 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_21
timestamp 1679235063
transform -1 0 25852 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_22
timestamp 1679235063
transform 1 0 1104 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_23
timestamp 1679235063
transform -1 0 25852 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_24
timestamp 1679235063
transform 1 0 1104 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_25
timestamp 1679235063
transform -1 0 25852 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_26
timestamp 1679235063
transform 1 0 1104 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_27
timestamp 1679235063
transform -1 0 25852 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_28
timestamp 1679235063
transform 1 0 1104 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_29
timestamp 1679235063
transform -1 0 25852 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_30
timestamp 1679235063
transform 1 0 1104 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_31
timestamp 1679235063
transform -1 0 25852 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_32
timestamp 1679235063
transform 1 0 1104 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_33
timestamp 1679235063
transform -1 0 25852 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_34
timestamp 1679235063
transform 1 0 1104 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_35
timestamp 1679235063
transform -1 0 25852 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_36
timestamp 1679235063
transform 1 0 1104 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_37
timestamp 1679235063
transform -1 0 25852 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_38
timestamp 1679235063
transform 1 0 1104 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_39
timestamp 1679235063
transform -1 0 25852 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_40
timestamp 1679235063
transform 1 0 1104 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_41
timestamp 1679235063
transform -1 0 25852 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_42
timestamp 1679235063
transform 1 0 1104 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_43
timestamp 1679235063
transform -1 0 25852 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_44
timestamp 1679235063
transform 1 0 1104 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_45
timestamp 1679235063
transform -1 0 25852 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_46
timestamp 1679235063
transform 1 0 1104 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_47
timestamp 1679235063
transform -1 0 25852 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_48
timestamp 1679235063
transform 1 0 1104 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_49
timestamp 1679235063
transform -1 0 25852 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_50
timestamp 1679235063
transform 1 0 1104 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_51
timestamp 1679235063
transform -1 0 25852 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_52
timestamp 1679235063
transform 1 0 1104 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_53
timestamp 1679235063
transform -1 0 25852 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_54
timestamp 1679235063
transform 1 0 1104 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_55
timestamp 1679235063
transform -1 0 25852 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_56
timestamp 1679235063
transform 1 0 1104 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_57
timestamp 1679235063
transform -1 0 25852 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_58
timestamp 1679235063
transform 1 0 1104 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_59
timestamp 1679235063
transform -1 0 25852 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_60
timestamp 1679235063
transform 1 0 1104 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_61
timestamp 1679235063
transform -1 0 25852 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_62
timestamp 1679235063
transform 1 0 1104 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_63
timestamp 1679235063
transform -1 0 25852 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_64
timestamp 1679235063
transform 1 0 1104 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_65
timestamp 1679235063
transform -1 0 25852 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_66
timestamp 1679235063
transform 1 0 1104 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_67
timestamp 1679235063
transform -1 0 25852 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_68
timestamp 1679235063
transform 1 0 1104 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_69
timestamp 1679235063
transform -1 0 25852 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_70
timestamp 1679235063
transform 1 0 1104 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_71
timestamp 1679235063
transform -1 0 25852 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_72
timestamp 1679235063
transform 1 0 1104 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_73
timestamp 1679235063
transform -1 0 25852 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_74
timestamp 1679235063
transform 1 0 1104 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_75
timestamp 1679235063
transform -1 0 25852 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_76
timestamp 1679235063
transform 1 0 1104 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_77
timestamp 1679235063
transform -1 0 25852 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_78
timestamp 1679235063
transform 1 0 1104 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_79
timestamp 1679235063
transform -1 0 25852 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_80
timestamp 1679235063
transform 1 0 1104 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_81
timestamp 1679235063
transform -1 0 25852 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_82
timestamp 1679235063
transform 1 0 1104 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_83
timestamp 1679235063
transform -1 0 25852 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_84
timestamp 1679235063
transform 1 0 1104 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_85
timestamp 1679235063
transform -1 0 25852 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_86
timestamp 1679235063
transform 1 0 1104 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_87
timestamp 1679235063
transform -1 0 25852 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_88
timestamp 1679235063
transform 1 0 1104 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_89
timestamp 1679235063
transform -1 0 25852 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_90
timestamp 1679235063
transform 1 0 1104 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_91
timestamp 1679235063
transform -1 0 25852 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_92
timestamp 1679235063
transform 1 0 1104 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_93
timestamp 1679235063
transform -1 0 25852 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_94
timestamp 1679235063
transform 1 0 1104 0 -1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_95
timestamp 1679235063
transform -1 0 25852 0 -1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_96
timestamp 1679235063
transform 1 0 1104 0 1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_97
timestamp 1679235063
transform -1 0 25852 0 1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_98
timestamp 1679235063
transform 1 0 1104 0 -1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_99
timestamp 1679235063
transform -1 0 25852 0 -1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_100
timestamp 1679235063
transform 1 0 1104 0 1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_101
timestamp 1679235063
transform -1 0 25852 0 1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_102
timestamp 1679235063
transform 1 0 1104 0 -1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_103
timestamp 1679235063
transform -1 0 25852 0 -1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_104
timestamp 1679235063
transform 1 0 1104 0 1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_105
timestamp 1679235063
transform -1 0 25852 0 1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_106
timestamp 1679235063
transform 1 0 1104 0 -1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_107
timestamp 1679235063
transform -1 0 25852 0 -1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_108
timestamp 1679235063
transform 1 0 1104 0 1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_109
timestamp 1679235063
transform -1 0 25852 0 1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_110
timestamp 1679235063
transform 1 0 1104 0 -1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_111
timestamp 1679235063
transform -1 0 25852 0 -1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_112
timestamp 1679235063
transform 1 0 1104 0 1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_113
timestamp 1679235063
transform -1 0 25852 0 1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_114
timestamp 1679235063
transform 1 0 1104 0 -1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_115
timestamp 1679235063
transform -1 0 25852 0 -1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_116
timestamp 1679235063
transform 1 0 1104 0 1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_117
timestamp 1679235063
transform -1 0 25852 0 1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_118
timestamp 1679235063
transform 1 0 1104 0 -1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_119
timestamp 1679235063
transform -1 0 25852 0 -1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_120
timestamp 1679235063
transform 1 0 1104 0 1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_121
timestamp 1679235063
transform -1 0 25852 0 1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_122
timestamp 1679235063
transform 1 0 1104 0 -1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_123
timestamp 1679235063
transform -1 0 25852 0 -1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_124
timestamp 1679235063
transform 1 0 1104 0 1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_125
timestamp 1679235063
transform -1 0 25852 0 1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_126
timestamp 1679235063
transform 1 0 1104 0 -1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_127
timestamp 1679235063
transform -1 0 25852 0 -1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_128
timestamp 1679235063
transform 1 0 1104 0 1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_129
timestamp 1679235063
transform -1 0 25852 0 1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_130
timestamp 1679235063
transform 1 0 1104 0 -1 38080
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_131
timestamp 1679235063
transform -1 0 25852 0 -1 38080
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_132
timestamp 1679235063
transform 1 0 1104 0 1 38080
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_133
timestamp 1679235063
transform -1 0 25852 0 1 38080
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_134
timestamp 1679235063
transform 1 0 1104 0 -1 39168
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_135
timestamp 1679235063
transform -1 0 25852 0 -1 39168
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_136
timestamp 1679235063
transform 1 0 1104 0 1 39168
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_137
timestamp 1679235063
transform -1 0 25852 0 1 39168
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_138
timestamp 1679235063
transform 1 0 1104 0 -1 40256
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_139
timestamp 1679235063
transform -1 0 25852 0 -1 40256
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_140
timestamp 1679235063
transform 1 0 1104 0 1 40256
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_141
timestamp 1679235063
transform -1 0 25852 0 1 40256
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_142
timestamp 1679235063
transform 1 0 1104 0 -1 41344
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_143
timestamp 1679235063
transform -1 0 25852 0 -1 41344
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_144
timestamp 1679235063
transform 1 0 1104 0 1 41344
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_145
timestamp 1679235063
transform -1 0 25852 0 1 41344
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_146
timestamp 1679235063
transform 1 0 1104 0 -1 42432
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_147
timestamp 1679235063
transform -1 0 25852 0 -1 42432
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_148
timestamp 1679235063
transform 1 0 1104 0 1 42432
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_149
timestamp 1679235063
transform -1 0 25852 0 1 42432
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_150
timestamp 1679235063
transform 1 0 1104 0 -1 43520
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_151
timestamp 1679235063
transform -1 0 25852 0 -1 43520
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_152
timestamp 1679235063
transform 1 0 1104 0 1 43520
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_153
timestamp 1679235063
transform -1 0 25852 0 1 43520
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_154
timestamp 1679235063
transform 1 0 1104 0 -1 44608
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_155
timestamp 1679235063
transform -1 0 25852 0 -1 44608
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_156
timestamp 1679235063
transform 1 0 1104 0 1 44608
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_157
timestamp 1679235063
transform -1 0 25852 0 1 44608
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_158
timestamp 1679235063
transform 1 0 1104 0 -1 45696
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_159
timestamp 1679235063
transform -1 0 25852 0 -1 45696
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_160
timestamp 1679235063
transform 1 0 1104 0 1 45696
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_161
timestamp 1679235063
transform -1 0 25852 0 1 45696
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_162
timestamp 1679235063
transform 1 0 1104 0 -1 46784
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_163
timestamp 1679235063
transform -1 0 25852 0 -1 46784
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_164
timestamp 1679235063
transform 1 0 1104 0 1 46784
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_165
timestamp 1679235063
transform -1 0 25852 0 1 46784
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_166
timestamp 1679235063
transform 1 0 1104 0 -1 47872
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_167
timestamp 1679235063
transform -1 0 25852 0 -1 47872
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_168
timestamp 1679235063
transform 1 0 1104 0 1 47872
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_169
timestamp 1679235063
transform -1 0 25852 0 1 47872
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_170
timestamp 1679235063
transform 1 0 1104 0 -1 48960
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_171
timestamp 1679235063
transform -1 0 25852 0 -1 48960
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_172
timestamp 1679235063
transform 1 0 1104 0 1 48960
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_173
timestamp 1679235063
transform -1 0 25852 0 1 48960
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_174
timestamp 1679235063
transform 1 0 1104 0 -1 50048
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_175
timestamp 1679235063
transform -1 0 25852 0 -1 50048
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_176
timestamp 1679235063
transform 1 0 1104 0 1 50048
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_177
timestamp 1679235063
transform -1 0 25852 0 1 50048
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_178
timestamp 1679235063
transform 1 0 1104 0 -1 51136
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_179
timestamp 1679235063
transform -1 0 25852 0 -1 51136
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_180
timestamp 1679235063
transform 1 0 1104 0 1 51136
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_181
timestamp 1679235063
transform -1 0 25852 0 1 51136
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_182
timestamp 1679235063
transform 1 0 1104 0 -1 52224
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_183
timestamp 1679235063
transform -1 0 25852 0 -1 52224
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_184
timestamp 1679235063
transform 1 0 1104 0 1 52224
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_185
timestamp 1679235063
transform -1 0 25852 0 1 52224
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_186
timestamp 1679235063
transform 1 0 1104 0 -1 53312
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_187
timestamp 1679235063
transform -1 0 25852 0 -1 53312
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_188
timestamp 1679235063
transform 1 0 1104 0 1 53312
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_189
timestamp 1679235063
transform -1 0 25852 0 1 53312
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_190
timestamp 1679235063
transform 1 0 1104 0 -1 54400
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_191
timestamp 1679235063
transform -1 0 25852 0 -1 54400
box -38 -48 314 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__8_.mem_bottom_track_1.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1679235063
transform 1 0 19412 0 1 17408
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__8_.mem_bottom_track_1.sky130_fd_sc_hd__dfrtp_1_1_
timestamp 1679235063
transform 1 0 19872 0 1 19584
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__8_.mem_bottom_track_3.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1679235063
transform 1 0 22080 0 1 19584
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__8_.mem_bottom_track_3.sky130_fd_sc_hd__dfrtp_1_1_
timestamp 1679235063
transform 1 0 23368 0 -1 19584
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__8_.mem_bottom_track_5.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1679235063
transform 1 0 23552 0 -1 20672
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__8_.mem_bottom_track_5.sky130_fd_sc_hd__dfrtp_1_1_
timestamp 1679235063
transform 1 0 23276 0 -1 21760
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__8_.mem_bottom_track_7.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1679235063
transform 1 0 21528 0 1 21760
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__8_.mem_bottom_track_7.sky130_fd_sc_hd__dfrtp_1_1_
timestamp 1679235063
transform 1 0 19412 0 1 23936
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__8_.mem_bottom_track_9.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1679235063
transform 1 0 19688 0 -1 25024
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__8_.mem_bottom_track_9.sky130_fd_sc_hd__dfrtp_1_1_
timestamp 1679235063
transform 1 0 21896 0 1 23936
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__8_.mem_bottom_track_11.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1679235063
transform 1 0 23184 0 -1 23936
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__8_.mem_bottom_track_11.sky130_fd_sc_hd__dfrtp_1_1_
timestamp 1679235063
transform 1 0 23552 0 -1 25024
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__8_.mem_bottom_track_13.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1679235063
transform 1 0 23552 0 -1 26112
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__8_.mem_bottom_track_13.sky130_fd_sc_hd__dfrtp_1_1_
timestamp 1679235063
transform 1 0 23184 0 -1 27200
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__8_.mem_bottom_track_15.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1679235063
transform 1 0 21988 0 -1 28288
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__8_.mem_bottom_track_15.sky130_fd_sc_hd__dfrtp_1_1_
timestamp 1679235063
transform 1 0 19872 0 1 27200
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__8_.mem_bottom_track_17.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1679235063
transform 1 0 19412 0 1 26112
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__8_.mem_bottom_track_17.sky130_fd_sc_hd__dfrtp_1_1_
timestamp 1679235063
transform 1 0 17940 0 -1 27200
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__8_.mem_bottom_track_19.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1679235063
transform 1 0 17112 0 1 28288
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__8_.mem_bottom_track_19.sky130_fd_sc_hd__dfrtp_1_1_
timestamp 1679235063
transform 1 0 17112 0 1 29376
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__8_.mem_bottom_track_29.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1679235063
transform 1 0 16836 0 1 30464
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__8_.mem_bottom_track_29.sky130_fd_sc_hd__dfrtp_1_1_
timestamp 1679235063
transform 1 0 16836 0 1 31552
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__8_.mem_bottom_track_31.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1679235063
transform 1 0 17388 0 -1 32640
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__8_.mem_bottom_track_31.sky130_fd_sc_hd__dfrtp_1_1_
timestamp 1679235063
transform 1 0 19412 0 1 31552
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__8_.mem_bottom_track_33.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1679235063
transform 1 0 20700 0 1 30464
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__8_.mem_bottom_track_33.sky130_fd_sc_hd__dfrtp_1_1_
timestamp 1679235063
transform 1 0 22448 0 -1 31552
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__8_.mem_bottom_track_35.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1679235063
transform 1 0 23276 0 -1 30464
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__8_.mem_bottom_track_35.sky130_fd_sc_hd__dfrtp_1_1_
timestamp 1679235063
transform 1 0 23460 0 -1 32640
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__8_.mem_bottom_track_45.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1679235063
transform 1 0 22264 0 1 32640
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__8_.mem_bottom_track_45.sky130_fd_sc_hd__dfrtp_1_1_
timestamp 1679235063
transform 1 0 21988 0 -1 33728
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__8_.mem_bottom_track_47.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1679235063
transform 1 0 21620 0 1 33728
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__8_.mem_bottom_track_47.sky130_fd_sc_hd__dfrtp_1_1_
timestamp 1679235063
transform 1 0 19412 0 -1 33728
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__8_.mem_bottom_track_49.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1679235063
transform 1 0 19412 0 1 33728
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__8_.mem_bottom_track_49.sky130_fd_sc_hd__dfrtp_1_1_
timestamp 1679235063
transform 1 0 19412 0 1 32640
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__8_.mem_bottom_track_51.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1679235063
transform 1 0 20608 0 1 28288
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_4  sb_0__8_.mem_bottom_track_51.sky130_fd_sc_hd__dfrtp_1_1_
timestamp 1679235063
transform 1 0 23276 0 -1 18496
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__8_.mem_right_track_0.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1679235063
transform 1 0 20424 0 1 44608
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_2  sb_0__8_.mem_right_track_0.sky130_fd_sc_hd__dfrtp_1_1_
timestamp 1679235063
transform 1 0 13248 0 -1 31552
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__8_.mem_right_track_0.sky130_fd_sc_hd__dfrtp_1_2_
timestamp 1679235063
transform 1 0 9108 0 1 26112
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__8_.mem_right_track_2.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1679235063
transform 1 0 10212 0 1 27200
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__8_.mem_right_track_2.sky130_fd_sc_hd__dfrtp_1_1_
timestamp 1679235063
transform 1 0 9476 0 1 28288
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__8_.mem_right_track_2.sky130_fd_sc_hd__dfrtp_1_2_
timestamp 1679235063
transform 1 0 9384 0 -1 27200
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__8_.mem_right_track_4.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1679235063
transform 1 0 11500 0 1 29376
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__8_.mem_right_track_4.sky130_fd_sc_hd__dfrtp_1_1_
timestamp 1679235063
transform 1 0 12236 0 -1 30464
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__8_.mem_right_track_4.sky130_fd_sc_hd__dfrtp_1_2_
timestamp 1679235063
transform 1 0 11684 0 1 28288
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__8_.mem_right_track_6.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1679235063
transform 1 0 14260 0 1 29376
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__8_.mem_right_track_6.sky130_fd_sc_hd__dfrtp_1_1_
timestamp 1679235063
transform 1 0 12696 0 -1 27200
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__8_.mem_right_track_6.sky130_fd_sc_hd__dfrtp_1_2_
timestamp 1679235063
transform 1 0 11684 0 -1 25024
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__8_.mem_right_track_8.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1679235063
transform 1 0 12328 0 -1 26112
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__8_.mem_right_track_8.sky130_fd_sc_hd__dfrtp_1_1_
timestamp 1679235063
transform 1 0 10580 0 1 23936
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__8_.mem_right_track_8.sky130_fd_sc_hd__dfrtp_1_2_
timestamp 1679235063
transform 1 0 8556 0 -1 23936
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__8_.mem_right_track_10.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1679235063
transform 1 0 9200 0 -1 25024
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__8_.mem_right_track_10.sky130_fd_sc_hd__dfrtp_1_1_
timestamp 1679235063
transform 1 0 8188 0 -1 22848
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__8_.mem_right_track_10.sky130_fd_sc_hd__dfrtp_1_2_
timestamp 1679235063
transform 1 0 6348 0 1 19584
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__8_.mem_right_track_12.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1679235063
transform 1 0 6808 0 1 18496
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__8_.mem_right_track_12.sky130_fd_sc_hd__dfrtp_1_1_
timestamp 1679235063
transform 1 0 9108 0 1 19584
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__8_.mem_right_track_14.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1679235063
transform 1 0 11132 0 1 20672
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__8_.mem_right_track_14.sky130_fd_sc_hd__dfrtp_1_1_
timestamp 1679235063
transform 1 0 12788 0 -1 21760
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__8_.mem_right_track_16.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1679235063
transform 1 0 13432 0 -1 22848
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__8_.mem_right_track_16.sky130_fd_sc_hd__dfrtp_1_1_
timestamp 1679235063
transform 1 0 12788 0 -1 20672
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__8_.mem_right_track_18.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1679235063
transform 1 0 12328 0 -1 19584
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__8_.mem_right_track_18.sky130_fd_sc_hd__dfrtp_1_1_
timestamp 1679235063
transform 1 0 11684 0 -1 16320
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__8_.mem_right_track_20.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1679235063
transform 1 0 9752 0 1 13056
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__8_.mem_right_track_20.sky130_fd_sc_hd__dfrtp_1_1_
timestamp 1679235063
transform 1 0 9108 0 1 9792
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__8_.mem_right_track_22.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1679235063
transform 1 0 8556 0 -1 8704
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__8_.mem_right_track_22.sky130_fd_sc_hd__dfrtp_1_1_
timestamp 1679235063
transform 1 0 9016 0 -1 7616
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__8_.mem_right_track_24.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1679235063
transform 1 0 9936 0 1 5440
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__8_.mem_right_track_24.sky130_fd_sc_hd__dfrtp_1_1_
timestamp 1679235063
transform 1 0 10580 0 1 6528
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__8_.mem_right_track_26.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1679235063
transform 1 0 11684 0 -1 9792
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__8_.mem_right_track_26.sky130_fd_sc_hd__dfrtp_1_1_
timestamp 1679235063
transform 1 0 13524 0 -1 14144
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__8_.mem_right_track_28.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1679235063
transform 1 0 14444 0 -1 17408
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__8_.mem_right_track_28.sky130_fd_sc_hd__dfrtp_1_1_
timestamp 1679235063
transform 1 0 14260 0 1 19584
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__8_.mem_right_track_30.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1679235063
transform 1 0 15180 0 1 20672
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__8_.mem_right_track_30.sky130_fd_sc_hd__dfrtp_1_1_
timestamp 1679235063
transform 1 0 16100 0 1 21760
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__8_.mem_right_track_32.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1679235063
transform 1 0 16836 0 -1 20672
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__8_.mem_right_track_32.sky130_fd_sc_hd__dfrtp_1_1_
timestamp 1679235063
transform 1 0 16836 0 -1 18496
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__8_.mem_right_track_34.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1679235063
transform 1 0 16192 0 1 15232
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__8_.mem_right_track_34.sky130_fd_sc_hd__dfrtp_1_1_
timestamp 1679235063
transform 1 0 14628 0 1 10880
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__8_.mem_right_track_36.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1679235063
transform 1 0 14260 0 1 7616
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__8_.mem_right_track_36.sky130_fd_sc_hd__dfrtp_1_1_
timestamp 1679235063
transform 1 0 12972 0 -1 6528
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__8_.mem_right_track_38.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1679235063
transform 1 0 13708 0 -1 5440
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__8_.mem_right_track_38.sky130_fd_sc_hd__dfrtp_1_1_
timestamp 1679235063
transform 1 0 15088 0 1 4352
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__8_.mem_right_track_40.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1679235063
transform 1 0 16836 0 -1 5440
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__8_.mem_right_track_40.sky130_fd_sc_hd__dfrtp_1_1_
timestamp 1679235063
transform 1 0 16836 0 -1 6528
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__8_.mem_right_track_42.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1679235063
transform 1 0 17112 0 1 7616
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__8_.mem_right_track_42.sky130_fd_sc_hd__dfrtp_1_1_
timestamp 1679235063
transform 1 0 19688 0 -1 10880
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__8_.mem_right_track_44.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1679235063
transform 1 0 20332 0 1 11968
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__8_.mem_right_track_44.sky130_fd_sc_hd__dfrtp_1_1_
timestamp 1679235063
transform 1 0 19412 0 1 15232
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__8_.mem_right_track_46.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1679235063
transform 1 0 19688 0 -1 16320
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__8_.mem_right_track_46.sky130_fd_sc_hd__dfrtp_1_1_
timestamp 1679235063
transform 1 0 21988 0 -1 16320
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__8_.mem_right_track_48.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1679235063
transform 1 0 22264 0 1 15232
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__8_.mem_right_track_48.sky130_fd_sc_hd__dfrtp_1_1_
timestamp 1679235063
transform 1 0 22264 0 1 14144
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__8_.mem_right_track_50.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1679235063
transform 1 0 23000 0 -1 13056
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__8_.mem_right_track_50.sky130_fd_sc_hd__dfrtp_1_1_
timestamp 1679235063
transform 1 0 23092 0 -1 11968
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__8_.mem_right_track_52.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1679235063
transform 1 0 22264 0 1 9792
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__8_.mem_right_track_52.sky130_fd_sc_hd__dfrtp_1_1_
timestamp 1679235063
transform 1 0 22356 0 -1 8704
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__8_.mem_right_track_54.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1679235063
transform 1 0 21988 0 1 6528
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__8_.mem_right_track_54.sky130_fd_sc_hd__dfrtp_1_1_
timestamp 1679235063
transform 1 0 19688 0 -1 5440
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__8_.mem_right_track_56.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1679235063
transform 1 0 19780 0 1 6528
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__8_.mem_right_track_56.sky130_fd_sc_hd__dfrtp_1_1_
timestamp 1679235063
transform 1 0 19688 0 -1 8704
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__8_.mem_right_track_58.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1679235063
transform 1 0 17664 0 -1 9792
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__8_.mem_right_track_58.sky130_fd_sc_hd__dfrtp_1_1_
timestamp 1679235063
transform 1 0 16836 0 -1 14144
box -38 -48 1878 592
use sky130_fd_sc_hd__mux2_1  sb_0__8_.mux_bottom_track_1.mux_l1_in_0_
timestamp 1679235063
transform 1 0 20700 0 -1 22848
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  sb_0__8_.mux_bottom_track_1.mux_l1_in_1__190
timestamp 1679235063
transform 1 0 19964 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_0__8_.mux_bottom_track_1.mux_l1_in_1_
timestamp 1679235063
transform 1 0 18860 0 -1 21760
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_0__8_.mux_bottom_track_1.mux_l2_in_0_
timestamp 1679235063
transform 1 0 20056 0 -1 19584
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_2  sb_0__8_.mux_bottom_track_1.sky130_fd_sc_hd__buf_4_0_
timestamp 1679235063
transform 1 0 18492 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  sb_0__8_.mux_bottom_track_3.mux_l1_in_0_
timestamp 1679235063
transform 1 0 24564 0 1 20672
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_0__8_.mux_bottom_track_3.mux_l2_in_0_
timestamp 1679235063
transform 1 0 24564 0 1 17408
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  sb_0__8_.mux_bottom_track_3.mux_l2_in_0__145
timestamp 1679235063
transform 1 0 17940 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  sb_0__8_.mux_bottom_track_3.sky130_fd_sc_hd__buf_4_0_
timestamp 1679235063
transform 1 0 15456 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_0__8_.mux_bottom_track_5.mux_l1_in_0_
timestamp 1679235063
transform 1 0 24564 0 1 22848
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_0__8_.mux_bottom_track_5.mux_l2_in_0_
timestamp 1679235063
transform 1 0 22172 0 -1 19584
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  sb_0__8_.mux_bottom_track_5.mux_l2_in_0__152
timestamp 1679235063
transform 1 0 21804 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  sb_0__8_.mux_bottom_track_5.sky130_fd_sc_hd__buf_4_0_
timestamp 1679235063
transform 1 0 20884 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_0__8_.mux_bottom_track_7.mux_l1_in_0_
timestamp 1679235063
transform 1 0 21988 0 -1 26112
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  sb_0__8_.mux_bottom_track_7.mux_l1_in_1__154
timestamp 1679235063
transform 1 0 23828 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_0__8_.mux_bottom_track_7.mux_l1_in_1_
timestamp 1679235063
transform 1 0 19228 0 -1 23936
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_0__8_.mux_bottom_track_7.mux_l2_in_0_
timestamp 1679235063
transform 1 0 19504 0 1 22848
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_2  sb_0__8_.mux_bottom_track_7.sky130_fd_sc_hd__buf_4_0_
timestamp 1679235063
transform 1 0 19780 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  sb_0__8_.mux_bottom_track_9.mux_l1_in_0_
timestamp 1679235063
transform 1 0 22632 0 1 26112
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_0__8_.mux_bottom_track_9.mux_l2_in_0_
timestamp 1679235063
transform 1 0 21988 0 -1 21760
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  sb_0__8_.mux_bottom_track_9.mux_l2_in_0__155
timestamp 1679235063
transform 1 0 21896 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  sb_0__8_.mux_bottom_track_9.sky130_fd_sc_hd__buf_4_0_
timestamp 1679235063
transform 1 0 20148 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_0__8_.mux_bottom_track_11.mux_l1_in_0_
timestamp 1679235063
transform 1 0 24564 0 1 26112
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  sb_0__8_.mux_bottom_track_11.mux_l2_in_0__191
timestamp 1679235063
transform 1 0 19320 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_0__8_.mux_bottom_track_11.mux_l2_in_0_
timestamp 1679235063
transform 1 0 24564 0 1 21760
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  sb_0__8_.mux_bottom_track_11.sky130_fd_sc_hd__buf_4_0_
timestamp 1679235063
transform 1 0 24564 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_0__8_.mux_bottom_track_13.mux_l1_in_0_
timestamp 1679235063
transform 1 0 24196 0 -1 28288
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_0__8_.mux_bottom_track_13.mux_l2_in_0_
timestamp 1679235063
transform 1 0 22080 0 -1 25024
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  sb_0__8_.mux_bottom_track_13.mux_l2_in_0__192
timestamp 1679235063
transform 1 0 18676 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  sb_0__8_.mux_bottom_track_13.sky130_fd_sc_hd__buf_4_0_
timestamp 1679235063
transform 1 0 20608 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_0__8_.mux_bottom_track_15.mux_l1_in_0_
timestamp 1679235063
transform 1 0 22080 0 1 27200
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_0__8_.mux_bottom_track_15.mux_l2_in_0_
timestamp 1679235063
transform 1 0 20424 0 -1 23936
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  sb_0__8_.mux_bottom_track_15.mux_l2_in_0__193
timestamp 1679235063
transform 1 0 20884 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  sb_0__8_.mux_bottom_track_15.sky130_fd_sc_hd__buf_4_0_
timestamp 1679235063
transform 1 0 18492 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_0__8_.mux_bottom_track_17.mux_l1_in_0_
timestamp 1679235063
transform 1 0 20700 0 -1 27200
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  sb_0__8_.mux_bottom_track_17.mux_l2_in_0__194
timestamp 1679235063
transform 1 0 18860 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_0__8_.mux_bottom_track_17.mux_l2_in_0_
timestamp 1679235063
transform 1 0 18124 0 1 23936
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  sb_0__8_.mux_bottom_track_17.sky130_fd_sc_hd__buf_4_0_
timestamp 1679235063
transform 1 0 17572 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_0__8_.mux_bottom_track_19.mux_l1_in_0_
timestamp 1679235063
transform 1 0 20608 0 1 29376
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_0__8_.mux_bottom_track_19.mux_l2_in_0_
timestamp 1679235063
transform 1 0 17848 0 1 26112
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  sb_0__8_.mux_bottom_track_19.mux_l2_in_0__143
timestamp 1679235063
transform 1 0 18216 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  sb_0__8_.mux_bottom_track_19.sky130_fd_sc_hd__buf_4_0_
timestamp 1679235063
transform 1 0 16652 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_0__8_.mux_bottom_track_29.mux_l1_in_0_
timestamp 1679235063
transform 1 0 20148 0 -1 31552
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_0__8_.mux_bottom_track_29.mux_l2_in_0_
timestamp 1679235063
transform 1 0 18032 0 -1 28288
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  sb_0__8_.mux_bottom_track_29.mux_l2_in_0__144
timestamp 1679235063
transform 1 0 18032 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  sb_0__8_.mux_bottom_track_29.sky130_fd_sc_hd__buf_4_0_
timestamp 1679235063
transform 1 0 16008 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_0__8_.mux_bottom_track_31.mux_l1_in_0_
timestamp 1679235063
transform 1 0 21620 0 1 31552
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  sb_0__8_.mux_bottom_track_31.mux_l2_in_0__146
timestamp 1679235063
transform 1 0 19872 0 -1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_0__8_.mux_bottom_track_31.mux_l2_in_0_
timestamp 1679235063
transform 1 0 19412 0 1 28288
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  sb_0__8_.mux_bottom_track_31.sky130_fd_sc_hd__buf_4_0_
timestamp 1679235063
transform 1 0 18676 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_0__8_.mux_bottom_track_33.mux_l1_in_0_
timestamp 1679235063
transform 1 0 24564 0 1 32640
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  sb_0__8_.mux_bottom_track_33.mux_l2_in_0__147
timestamp 1679235063
transform 1 0 23184 0 1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_0__8_.mux_bottom_track_33.mux_l2_in_0_
timestamp 1679235063
transform 1 0 23276 0 1 27200
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  sb_0__8_.mux_bottom_track_33.sky130_fd_sc_hd__buf_4_0_
timestamp 1679235063
transform 1 0 21252 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_0__8_.mux_bottom_track_35.mux_l1_in_0_
timestamp 1679235063
transform 1 0 24196 0 -1 33728
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  sb_0__8_.mux_bottom_track_35.mux_l2_in_0__148
timestamp 1679235063
transform 1 0 24288 0 -1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_0__8_.mux_bottom_track_35.mux_l2_in_0_
timestamp 1679235063
transform 1 0 24564 0 1 28288
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  sb_0__8_.mux_bottom_track_35.sky130_fd_sc_hd__buf_4_0_
timestamp 1679235063
transform 1 0 21252 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_0__8_.mux_bottom_track_45.mux_l1_in_0_
timestamp 1679235063
transform 1 0 22724 0 1 34816
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  sb_0__8_.mux_bottom_track_45.mux_l2_in_0__149
timestamp 1679235063
transform 1 0 21252 0 -1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_0__8_.mux_bottom_track_45.mux_l2_in_0_
timestamp 1679235063
transform 1 0 21988 0 -1 30464
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  sb_0__8_.mux_bottom_track_45.sky130_fd_sc_hd__buf_4_0_
timestamp 1679235063
transform 1 0 19412 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_0__8_.mux_bottom_track_47.mux_l1_in_0_
timestamp 1679235063
transform 1 0 21988 0 -1 35904
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  sb_0__8_.mux_bottom_track_47.mux_l2_in_0__150
timestamp 1679235063
transform 1 0 19228 0 -1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_0__8_.mux_bottom_track_47.mux_l2_in_0_
timestamp 1679235063
transform 1 0 19872 0 -1 30464
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  sb_0__8_.mux_bottom_track_47.sky130_fd_sc_hd__buf_4_0_
timestamp 1679235063
transform 1 0 19044 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_0__8_.mux_bottom_track_49.mux_l1_in_0_
timestamp 1679235063
transform 1 0 20700 0 -1 35904
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_0__8_.mux_bottom_track_49.mux_l2_in_0_
timestamp 1679235063
transform 1 0 19412 0 1 29376
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  sb_0__8_.mux_bottom_track_49.mux_l2_in_0__151
timestamp 1679235063
transform 1 0 19228 0 -1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  sb_0__8_.mux_bottom_track_49.sky130_fd_sc_hd__buf_4_0_
timestamp 1679235063
transform 1 0 15640 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  sb_0__8_.mux_bottom_track_51.mux_l1_in_0_
timestamp 1679235063
transform 1 0 23092 0 -1 29376
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  sb_0__8_.mux_bottom_track_51.mux_l2_in_0__153
timestamp 1679235063
transform 1 0 17296 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_0__8_.mux_bottom_track_51.mux_l2_in_0_
timestamp 1679235063
transform 1 0 20700 0 -1 17408
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  sb_0__8_.mux_bottom_track_51.sky130_fd_sc_hd__buf_4_0_
timestamp 1679235063
transform 1 0 21988 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_0__8_.mux_right_track_0.mux_l1_in_0_
timestamp 1679235063
transform 1 0 15548 0 -1 32640
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_0__8_.mux_right_track_0.mux_l1_in_1_
timestamp 1679235063
transform 1 0 15640 0 1 31552
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_0__8_.mux_right_track_0.mux_l2_in_0_
timestamp 1679235063
transform 1 0 12972 0 -1 29376
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_0__8_.mux_right_track_0.mux_l2_in_1_
timestamp 1679235063
transform 1 0 7636 0 1 17408
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  sb_0__8_.mux_right_track_0.mux_l2_in_1__156
timestamp 1679235063
transform 1 0 8004 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_0__8_.mux_right_track_0.mux_l3_in_0_
timestamp 1679235063
transform 1 0 11500 0 1 25024
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  sb_0__8_.mux_right_track_0.sky130_fd_sc_hd__buf_4_0_
timestamp 1679235063
transform 1 0 17848 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_0__8_.mux_right_track_2.mux_l1_in_0_
timestamp 1679235063
transform 1 0 14720 0 1 28288
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_0__8_.mux_right_track_2.mux_l1_in_1_
timestamp 1679235063
transform 1 0 15916 0 1 28288
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_0__8_.mux_right_track_2.mux_l2_in_0_
timestamp 1679235063
transform 1 0 13156 0 -1 28288
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  sb_0__8_.mux_right_track_2.mux_l2_in_1__162
timestamp 1679235063
transform 1 0 9476 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_0__8_.mux_right_track_2.mux_l2_in_1_
timestamp 1679235063
transform 1 0 9660 0 1 20672
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_0__8_.mux_right_track_2.mux_l3_in_0_
timestamp 1679235063
transform 1 0 11776 0 1 26112
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  sb_0__8_.mux_right_track_2.sky130_fd_sc_hd__buf_4_0_
timestamp 1679235063
transform 1 0 16928 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_0__8_.mux_right_track_4.mux_l1_in_0_
timestamp 1679235063
transform 1 0 15364 0 -1 29376
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_0__8_.mux_right_track_4.mux_l1_in_1_
timestamp 1679235063
transform 1 0 15548 0 -1 30464
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_0__8_.mux_right_track_4.mux_l2_in_0_
timestamp 1679235063
transform 1 0 14168 0 -1 29376
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_0__8_.mux_right_track_4.mux_l2_in_1_
timestamp 1679235063
transform 1 0 12512 0 1 21760
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  sb_0__8_.mux_right_track_4.mux_l2_in_1__173
timestamp 1679235063
transform 1 0 13340 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_0__8_.mux_right_track_4.mux_l3_in_0_
timestamp 1679235063
transform 1 0 12972 0 1 26112
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  sb_0__8_.mux_right_track_4.sky130_fd_sc_hd__buf_4_0_
timestamp 1679235063
transform 1 0 17572 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_0__8_.mux_right_track_6.mux_l1_in_0_
timestamp 1679235063
transform 1 0 16836 0 -1 29376
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_0__8_.mux_right_track_6.mux_l1_in_1_
timestamp 1679235063
transform 1 0 16836 0 -1 28288
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_0__8_.mux_right_track_6.mux_l2_in_0_
timestamp 1679235063
transform 1 0 14444 0 1 26112
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_0__8_.mux_right_track_6.mux_l2_in_1_
timestamp 1679235063
transform 1 0 10948 0 1 18496
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  sb_0__8_.mux_right_track_6.mux_l2_in_1__184
timestamp 1679235063
transform 1 0 11684 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_0__8_.mux_right_track_6.mux_l3_in_0_
timestamp 1679235063
transform 1 0 13432 0 -1 23936
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  sb_0__8_.mux_right_track_6.sky130_fd_sc_hd__buf_4_0_
timestamp 1679235063
transform 1 0 18032 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_0__8_.mux_right_track_8.mux_l1_in_0_
timestamp 1679235063
transform 1 0 14996 0 -1 27200
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_0__8_.mux_right_track_8.mux_l1_in_1_
timestamp 1679235063
transform 1 0 15456 0 1 27200
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_0__8_.mux_right_track_8.mux_l2_in_0_
timestamp 1679235063
transform 1 0 13892 0 -1 25024
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  sb_0__8_.mux_right_track_8.mux_l2_in_1__185
timestamp 1679235063
transform 1 0 9108 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_0__8_.mux_right_track_8.mux_l2_in_1_
timestamp 1679235063
transform 1 0 9108 0 -1 17408
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_0__8_.mux_right_track_8.mux_l3_in_0_
timestamp 1679235063
transform 1 0 11776 0 -1 22848
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  sb_0__8_.mux_right_track_8.sky130_fd_sc_hd__buf_4_0_
timestamp 1679235063
transform 1 0 16836 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_0__8_.mux_right_track_10.mux_l1_in_0_
timestamp 1679235063
transform 1 0 14260 0 1 25024
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_0__8_.mux_right_track_10.mux_l1_in_1_
timestamp 1679235063
transform 1 0 14536 0 -1 26112
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_0__8_.mux_right_track_10.mux_l2_in_0_
timestamp 1679235063
transform 1 0 11316 0 1 21760
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_0__8_.mux_right_track_10.mux_l2_in_1_
timestamp 1679235063
transform 1 0 6992 0 1 13056
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  sb_0__8_.mux_right_track_10.mux_l2_in_1__157
timestamp 1679235063
transform 1 0 6532 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_0__8_.mux_right_track_10.mux_l3_in_0_
timestamp 1679235063
transform 1 0 9752 0 1 18496
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  sb_0__8_.mux_right_track_10.sky130_fd_sc_hd__buf_4_0_
timestamp 1679235063
transform 1 0 15640 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_0__8_.mux_right_track_12.mux_l1_in_0_
timestamp 1679235063
transform 1 0 12972 0 1 22848
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  sb_0__8_.mux_right_track_12.mux_l1_in_1__158
timestamp 1679235063
transform 1 0 9108 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_0__8_.mux_right_track_12.mux_l1_in_1_
timestamp 1679235063
transform 1 0 7820 0 1 11968
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_0__8_.mux_right_track_12.mux_l2_in_0_
timestamp 1679235063
transform 1 0 11868 0 1 19584
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  sb_0__8_.mux_right_track_12.sky130_fd_sc_hd__buf_4_0_
timestamp 1679235063
transform 1 0 16652 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_0__8_.mux_right_track_14.mux_l1_in_0_
timestamp 1679235063
transform 1 0 15548 0 -1 25024
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_0__8_.mux_right_track_14.mux_l1_in_1_
timestamp 1679235063
transform 1 0 14260 0 1 18496
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  sb_0__8_.mux_right_track_14.mux_l1_in_1__159
timestamp 1679235063
transform 1 0 14352 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_0__8_.mux_right_track_14.mux_l2_in_0_
timestamp 1679235063
transform 1 0 14904 0 1 21760
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  sb_0__8_.mux_right_track_14.sky130_fd_sc_hd__buf_4_0_
timestamp 1679235063
transform 1 0 18216 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_0__8_.mux_right_track_16.mux_l1_in_0_
timestamp 1679235063
transform 1 0 16836 0 -1 25024
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  sb_0__8_.mux_right_track_16.mux_l1_in_1__160
timestamp 1679235063
transform 1 0 14996 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_0__8_.mux_right_track_16.mux_l1_in_1_
timestamp 1679235063
transform 1 0 12880 0 -1 17408
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_0__8_.mux_right_track_16.mux_l2_in_0_
timestamp 1679235063
transform 1 0 14996 0 -1 20672
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  sb_0__8_.mux_right_track_16.sky130_fd_sc_hd__buf_4_0_
timestamp 1679235063
transform 1 0 19228 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_0__8_.mux_right_track_18.mux_l1_in_0_
timestamp 1679235063
transform 1 0 12972 0 1 15232
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_0__8_.mux_right_track_18.mux_l2_in_0_
timestamp 1679235063
transform 1 0 14076 0 -1 16320
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  sb_0__8_.mux_right_track_18.mux_l2_in_0__161
timestamp 1679235063
transform 1 0 15272 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  sb_0__8_.mux_right_track_18.sky130_fd_sc_hd__buf_4_0_
timestamp 1679235063
transform 1 0 18400 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_0__8_.mux_right_track_20.mux_l1_in_0_
timestamp 1679235063
transform 1 0 11316 0 1 10880
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_0__8_.mux_right_track_20.mux_l2_in_0_
timestamp 1679235063
transform 1 0 11500 0 1 9792
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  sb_0__8_.mux_right_track_20.mux_l2_in_0__163
timestamp 1679235063
transform 1 0 11684 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  sb_0__8_.mux_right_track_20.sky130_fd_sc_hd__buf_4_0_
timestamp 1679235063
transform 1 0 16100 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_0__8_.mux_right_track_22.mux_l1_in_0_
timestamp 1679235063
transform 1 0 10396 0 1 7616
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  sb_0__8_.mux_right_track_22.mux_l2_in_0__164
timestamp 1679235063
transform 1 0 10948 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_0__8_.mux_right_track_22.mux_l2_in_0_
timestamp 1679235063
transform 1 0 11776 0 1 7616
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  sb_0__8_.mux_right_track_22.sky130_fd_sc_hd__buf_4_0_
timestamp 1679235063
transform 1 0 16836 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_0__8_.mux_right_track_24.mux_l1_in_0_
timestamp 1679235063
transform 1 0 11684 0 -1 7616
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  sb_0__8_.mux_right_track_24.mux_l2_in_0__165
timestamp 1679235063
transform 1 0 13892 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_0__8_.mux_right_track_24.mux_l2_in_0_
timestamp 1679235063
transform 1 0 12972 0 1 7616
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  sb_0__8_.mux_right_track_24.sky130_fd_sc_hd__buf_4_0_
timestamp 1679235063
transform 1 0 21528 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_0__8_.mux_right_track_26.mux_l1_in_0_
timestamp 1679235063
transform 1 0 14076 0 -1 13056
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  sb_0__8_.mux_right_track_26.mux_l2_in_0__166
timestamp 1679235063
transform 1 0 16560 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_0__8_.mux_right_track_26.mux_l2_in_0_
timestamp 1679235063
transform 1 0 16376 0 1 13056
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  sb_0__8_.mux_right_track_26.sky130_fd_sc_hd__buf_4_0_
timestamp 1679235063
transform 1 0 18676 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_0__8_.mux_right_track_28.mux_l1_in_0_
timestamp 1679235063
transform 1 0 16836 0 -1 23936
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  sb_0__8_.mux_right_track_28.mux_l1_in_1__167
timestamp 1679235063
transform 1 0 14260 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_0__8_.mux_right_track_28.mux_l1_in_1_
timestamp 1679235063
transform 1 0 13616 0 -1 15232
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_0__8_.mux_right_track_28.mux_l2_in_0_
timestamp 1679235063
transform 1 0 16836 0 -1 19584
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  sb_0__8_.mux_right_track_28.sky130_fd_sc_hd__buf_4_0_
timestamp 1679235063
transform 1 0 20056 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_0__8_.mux_right_track_30.mux_l1_in_0_
timestamp 1679235063
transform 1 0 18032 0 -1 25024
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  sb_0__8_.mux_right_track_30.mux_l1_in_1__168
timestamp 1679235063
transform 1 0 15640 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_0__8_.mux_right_track_30.mux_l1_in_1_
timestamp 1679235063
transform 1 0 15272 0 1 16320
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_0__8_.mux_right_track_30.mux_l2_in_0_
timestamp 1679235063
transform 1 0 17480 0 1 19584
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  sb_0__8_.mux_right_track_30.sky130_fd_sc_hd__buf_4_0_
timestamp 1679235063
transform 1 0 21620 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_0__8_.mux_right_track_32.mux_l1_in_0_
timestamp 1679235063
transform 1 0 17848 0 1 22848
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  sb_0__8_.mux_right_track_32.mux_l1_in_1__169
timestamp 1679235063
transform 1 0 14904 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_0__8_.mux_right_track_32.mux_l1_in_1_
timestamp 1679235063
transform 1 0 15548 0 -1 15232
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_0__8_.mux_right_track_32.mux_l2_in_0_
timestamp 1679235063
transform 1 0 17940 0 1 17408
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  sb_0__8_.mux_right_track_32.sky130_fd_sc_hd__buf_4_0_
timestamp 1679235063
transform 1 0 19504 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_0__8_.mux_right_track_34.mux_l1_in_0_
timestamp 1679235063
transform 1 0 16744 0 1 18496
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  sb_0__8_.mux_right_track_34.mux_l1_in_1__170
timestamp 1679235063
transform 1 0 14260 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_0__8_.mux_right_track_34.mux_l1_in_1_
timestamp 1679235063
transform 1 0 13064 0 -1 7616
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_0__8_.mux_right_track_34.mux_l2_in_0_
timestamp 1679235063
transform 1 0 16836 0 -1 11968
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  sb_0__8_.mux_right_track_34.sky130_fd_sc_hd__buf_4_0_
timestamp 1679235063
transform 1 0 19044 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_0__8_.mux_right_track_36.mux_l1_in_0_
timestamp 1679235063
transform 1 0 12972 0 1 6528
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  sb_0__8_.mux_right_track_36.mux_l2_in_0__171
timestamp 1679235063
transform 1 0 19044 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_0__8_.mux_right_track_36.mux_l2_in_0_
timestamp 1679235063
transform 1 0 15180 0 -1 6528
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  sb_0__8_.mux_right_track_36.sky130_fd_sc_hd__buf_4_0_
timestamp 1679235063
transform 1 0 12328 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_0__8_.mux_right_track_38.mux_l1_in_0_
timestamp 1679235063
transform 1 0 14996 0 -1 7616
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_0__8_.mux_right_track_38.mux_l2_in_0_
timestamp 1679235063
transform 1 0 16284 0 1 6528
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  sb_0__8_.mux_right_track_38.mux_l2_in_0__172
timestamp 1679235063
transform 1 0 9660 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  sb_0__8_.mux_right_track_38.sky130_fd_sc_hd__buf_4_0_
timestamp 1679235063
transform 1 0 10948 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_0__8_.mux_right_track_40.mux_l1_in_0_
timestamp 1679235063
transform 1 0 16836 0 -1 8704
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_0__8_.mux_right_track_40.mux_l2_in_0_
timestamp 1679235063
transform 1 0 17020 0 -1 7616
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  sb_0__8_.mux_right_track_40.mux_l2_in_0__174
timestamp 1679235063
transform 1 0 21252 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  sb_0__8_.mux_right_track_40.sky130_fd_sc_hd__buf_4_0_
timestamp 1679235063
transform 1 0 21252 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_0__8_.mux_right_track_42.mux_l1_in_0_
timestamp 1679235063
transform 1 0 17756 0 1 10880
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  sb_0__8_.mux_right_track_42.mux_l2_in_0__175
timestamp 1679235063
transform 1 0 14536 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_0__8_.mux_right_track_42.mux_l2_in_0_
timestamp 1679235063
transform 1 0 20792 0 1 9792
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  sb_0__8_.mux_right_track_42.sky130_fd_sc_hd__buf_4_0_
timestamp 1679235063
transform 1 0 7912 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_0__8_.mux_right_track_44.mux_l1_in_0_
timestamp 1679235063
transform 1 0 19412 0 1 20672
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_0__8_.mux_right_track_44.mux_l1_in_1_
timestamp 1679235063
transform 1 0 18032 0 -1 11968
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  sb_0__8_.mux_right_track_44.mux_l1_in_1__176
timestamp 1679235063
transform 1 0 10672 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_0__8_.mux_right_track_44.mux_l2_in_0_
timestamp 1679235063
transform 1 0 19504 0 -1 15232
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  sb_0__8_.mux_right_track_44.sky130_fd_sc_hd__buf_4_0_
timestamp 1679235063
transform 1 0 13524 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_0__8_.mux_right_track_46.mux_l1_in_0_
timestamp 1679235063
transform 1 0 19688 0 1 21760
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_0__8_.mux_right_track_46.mux_l1_in_1_
timestamp 1679235063
transform 1 0 18676 0 -1 13056
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  sb_0__8_.mux_right_track_46.mux_l1_in_1__177
timestamp 1679235063
transform 1 0 24564 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_0__8_.mux_right_track_46.mux_l2_in_0_
timestamp 1679235063
transform 1 0 20700 0 -1 15232
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  sb_0__8_.mux_right_track_46.sky130_fd_sc_hd__buf_4_0_
timestamp 1679235063
transform 1 0 11960 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_0__8_.mux_right_track_48.mux_l1_in_0_
timestamp 1679235063
transform 1 0 20608 0 1 20672
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  sb_0__8_.mux_right_track_48.mux_l1_in_1__178
timestamp 1679235063
transform 1 0 15548 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_0__8_.mux_right_track_48.mux_l1_in_1_
timestamp 1679235063
transform 1 0 19596 0 -1 11968
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_0__8_.mux_right_track_48.mux_l2_in_0_
timestamp 1679235063
transform 1 0 21436 0 1 13056
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  sb_0__8_.mux_right_track_48.sky130_fd_sc_hd__buf_4_0_
timestamp 1679235063
transform 1 0 8648 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_0__8_.mux_right_track_50.mux_l1_in_0_
timestamp 1679235063
transform 1 0 20148 0 1 13056
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_0__8_.mux_right_track_50.mux_l2_in_0_
timestamp 1679235063
transform 1 0 22724 0 1 10880
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  sb_0__8_.mux_right_track_50.mux_l2_in_0__179
timestamp 1679235063
transform 1 0 10304 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  sb_0__8_.mux_right_track_50.sky130_fd_sc_hd__buf_4_0_
timestamp 1679235063
transform 1 0 10948 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_0__8_.mux_right_track_52.mux_l1_in_0_
timestamp 1679235063
transform 1 0 19872 0 -1 9792
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_0__8_.mux_right_track_52.mux_l2_in_0_
timestamp 1679235063
transform 1 0 24564 0 1 6528
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  sb_0__8_.mux_right_track_52.mux_l2_in_0__180
timestamp 1679235063
transform 1 0 9752 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  sb_0__8_.mux_right_track_52.sky130_fd_sc_hd__buf_4_0_
timestamp 1679235063
transform 1 0 10304 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_0__8_.mux_right_track_54.mux_l1_in_0_
timestamp 1679235063
transform 1 0 18308 0 -1 8704
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_0__8_.mux_right_track_54.mux_l2_in_0_
timestamp 1679235063
transform 1 0 20516 0 -1 4352
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  sb_0__8_.mux_right_track_54.mux_l2_in_0__181
timestamp 1679235063
transform 1 0 11684 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  sb_0__8_.mux_right_track_54.sky130_fd_sc_hd__buf_4_0_
timestamp 1679235063
transform 1 0 12328 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_0__8_.mux_right_track_56.mux_l1_in_0_
timestamp 1679235063
transform 1 0 18124 0 1 9792
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  sb_0__8_.mux_right_track_56.mux_l2_in_0__182
timestamp 1679235063
transform 1 0 16100 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_0__8_.mux_right_track_56.mux_l2_in_0_
timestamp 1679235063
transform 1 0 19596 0 1 8704
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  sb_0__8_.mux_right_track_56.sky130_fd_sc_hd__buf_4_0_
timestamp 1679235063
transform 1 0 10396 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_0__8_.mux_right_track_58.mux_l1_in_0_
timestamp 1679235063
transform 1 0 17940 0 1 18496
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  sb_0__8_.mux_right_track_58.mux_l1_in_1__183
timestamp 1679235063
transform 1 0 10580 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_0__8_.mux_right_track_58.mux_l1_in_1_
timestamp 1679235063
transform 1 0 11684 0 -1 8704
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_0__8_.mux_right_track_58.mux_l2_in_0_
timestamp 1679235063
transform 1 0 16836 0 1 11968
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  sb_0__8_.mux_right_track_58.sky130_fd_sc_hd__buf_4_0_
timestamp 1679235063
transform 1 0 16192 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_192 pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1679235063
transform 1 0 3680 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_193
timestamp 1679235063
transform 1 0 6256 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_194
timestamp 1679235063
transform 1 0 8832 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_195
timestamp 1679235063
transform 1 0 11408 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_196
timestamp 1679235063
transform 1 0 13984 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_197
timestamp 1679235063
transform 1 0 16560 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_198
timestamp 1679235063
transform 1 0 19136 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_199
timestamp 1679235063
transform 1 0 21712 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_200
timestamp 1679235063
transform 1 0 24288 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_201
timestamp 1679235063
transform 1 0 6256 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_202
timestamp 1679235063
transform 1 0 11408 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_203
timestamp 1679235063
transform 1 0 16560 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_204
timestamp 1679235063
transform 1 0 21712 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_205
timestamp 1679235063
transform 1 0 3680 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_206
timestamp 1679235063
transform 1 0 8832 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_207
timestamp 1679235063
transform 1 0 13984 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_208
timestamp 1679235063
transform 1 0 19136 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_209
timestamp 1679235063
transform 1 0 24288 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_210
timestamp 1679235063
transform 1 0 6256 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_211
timestamp 1679235063
transform 1 0 11408 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_212
timestamp 1679235063
transform 1 0 16560 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_213
timestamp 1679235063
transform 1 0 21712 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_214
timestamp 1679235063
transform 1 0 3680 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_215
timestamp 1679235063
transform 1 0 8832 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_216
timestamp 1679235063
transform 1 0 13984 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_217
timestamp 1679235063
transform 1 0 19136 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_218
timestamp 1679235063
transform 1 0 24288 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_219
timestamp 1679235063
transform 1 0 6256 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_220
timestamp 1679235063
transform 1 0 11408 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_221
timestamp 1679235063
transform 1 0 16560 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_222
timestamp 1679235063
transform 1 0 21712 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_223
timestamp 1679235063
transform 1 0 3680 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_224
timestamp 1679235063
transform 1 0 8832 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_225
timestamp 1679235063
transform 1 0 13984 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_226
timestamp 1679235063
transform 1 0 19136 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_227
timestamp 1679235063
transform 1 0 24288 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_228
timestamp 1679235063
transform 1 0 6256 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_229
timestamp 1679235063
transform 1 0 11408 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_230
timestamp 1679235063
transform 1 0 16560 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_231
timestamp 1679235063
transform 1 0 21712 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_232
timestamp 1679235063
transform 1 0 3680 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_233
timestamp 1679235063
transform 1 0 8832 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_234
timestamp 1679235063
transform 1 0 13984 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_235
timestamp 1679235063
transform 1 0 19136 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_236
timestamp 1679235063
transform 1 0 24288 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_237
timestamp 1679235063
transform 1 0 6256 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_238
timestamp 1679235063
transform 1 0 11408 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_239
timestamp 1679235063
transform 1 0 16560 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_240
timestamp 1679235063
transform 1 0 21712 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_241
timestamp 1679235063
transform 1 0 3680 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_242
timestamp 1679235063
transform 1 0 8832 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_243
timestamp 1679235063
transform 1 0 13984 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_244
timestamp 1679235063
transform 1 0 19136 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_245
timestamp 1679235063
transform 1 0 24288 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_246
timestamp 1679235063
transform 1 0 6256 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_247
timestamp 1679235063
transform 1 0 11408 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_248
timestamp 1679235063
transform 1 0 16560 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_249
timestamp 1679235063
transform 1 0 21712 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_250
timestamp 1679235063
transform 1 0 3680 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_251
timestamp 1679235063
transform 1 0 8832 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_252
timestamp 1679235063
transform 1 0 13984 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_253
timestamp 1679235063
transform 1 0 19136 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_254
timestamp 1679235063
transform 1 0 24288 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_255
timestamp 1679235063
transform 1 0 6256 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_256
timestamp 1679235063
transform 1 0 11408 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_257
timestamp 1679235063
transform 1 0 16560 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_258
timestamp 1679235063
transform 1 0 21712 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_259
timestamp 1679235063
transform 1 0 3680 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_260
timestamp 1679235063
transform 1 0 8832 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_261
timestamp 1679235063
transform 1 0 13984 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_262
timestamp 1679235063
transform 1 0 19136 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_263
timestamp 1679235063
transform 1 0 24288 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_264
timestamp 1679235063
transform 1 0 6256 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_265
timestamp 1679235063
transform 1 0 11408 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_266
timestamp 1679235063
transform 1 0 16560 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_267
timestamp 1679235063
transform 1 0 21712 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_268
timestamp 1679235063
transform 1 0 3680 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_269
timestamp 1679235063
transform 1 0 8832 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_270
timestamp 1679235063
transform 1 0 13984 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_271
timestamp 1679235063
transform 1 0 19136 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_272
timestamp 1679235063
transform 1 0 24288 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_273
timestamp 1679235063
transform 1 0 6256 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_274
timestamp 1679235063
transform 1 0 11408 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_275
timestamp 1679235063
transform 1 0 16560 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_276
timestamp 1679235063
transform 1 0 21712 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_277
timestamp 1679235063
transform 1 0 3680 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_278
timestamp 1679235063
transform 1 0 8832 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_279
timestamp 1679235063
transform 1 0 13984 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_280
timestamp 1679235063
transform 1 0 19136 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_281
timestamp 1679235063
transform 1 0 24288 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_282
timestamp 1679235063
transform 1 0 6256 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_283
timestamp 1679235063
transform 1 0 11408 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_284
timestamp 1679235063
transform 1 0 16560 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_285
timestamp 1679235063
transform 1 0 21712 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_286
timestamp 1679235063
transform 1 0 3680 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_287
timestamp 1679235063
transform 1 0 8832 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_288
timestamp 1679235063
transform 1 0 13984 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_289
timestamp 1679235063
transform 1 0 19136 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_290
timestamp 1679235063
transform 1 0 24288 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_291
timestamp 1679235063
transform 1 0 6256 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_292
timestamp 1679235063
transform 1 0 11408 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_293
timestamp 1679235063
transform 1 0 16560 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_294
timestamp 1679235063
transform 1 0 21712 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_295
timestamp 1679235063
transform 1 0 3680 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_296
timestamp 1679235063
transform 1 0 8832 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_297
timestamp 1679235063
transform 1 0 13984 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_298
timestamp 1679235063
transform 1 0 19136 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_299
timestamp 1679235063
transform 1 0 24288 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_300
timestamp 1679235063
transform 1 0 6256 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_301
timestamp 1679235063
transform 1 0 11408 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_302
timestamp 1679235063
transform 1 0 16560 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_303
timestamp 1679235063
transform 1 0 21712 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_304
timestamp 1679235063
transform 1 0 3680 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_305
timestamp 1679235063
transform 1 0 8832 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_306
timestamp 1679235063
transform 1 0 13984 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_307
timestamp 1679235063
transform 1 0 19136 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_308
timestamp 1679235063
transform 1 0 24288 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_309
timestamp 1679235063
transform 1 0 6256 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_310
timestamp 1679235063
transform 1 0 11408 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_311
timestamp 1679235063
transform 1 0 16560 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_312
timestamp 1679235063
transform 1 0 21712 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_313
timestamp 1679235063
transform 1 0 3680 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_314
timestamp 1679235063
transform 1 0 8832 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_315
timestamp 1679235063
transform 1 0 13984 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_316
timestamp 1679235063
transform 1 0 19136 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_317
timestamp 1679235063
transform 1 0 24288 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_318
timestamp 1679235063
transform 1 0 6256 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_319
timestamp 1679235063
transform 1 0 11408 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_320
timestamp 1679235063
transform 1 0 16560 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_321
timestamp 1679235063
transform 1 0 21712 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_322
timestamp 1679235063
transform 1 0 3680 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_323
timestamp 1679235063
transform 1 0 8832 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_324
timestamp 1679235063
transform 1 0 13984 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_325
timestamp 1679235063
transform 1 0 19136 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_326
timestamp 1679235063
transform 1 0 24288 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_327
timestamp 1679235063
transform 1 0 6256 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_328
timestamp 1679235063
transform 1 0 11408 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_329
timestamp 1679235063
transform 1 0 16560 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_330
timestamp 1679235063
transform 1 0 21712 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_331
timestamp 1679235063
transform 1 0 3680 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_332
timestamp 1679235063
transform 1 0 8832 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_333
timestamp 1679235063
transform 1 0 13984 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_334
timestamp 1679235063
transform 1 0 19136 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_335
timestamp 1679235063
transform 1 0 24288 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_336
timestamp 1679235063
transform 1 0 6256 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_337
timestamp 1679235063
transform 1 0 11408 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_338
timestamp 1679235063
transform 1 0 16560 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_339
timestamp 1679235063
transform 1 0 21712 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_340
timestamp 1679235063
transform 1 0 3680 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_341
timestamp 1679235063
transform 1 0 8832 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_342
timestamp 1679235063
transform 1 0 13984 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_343
timestamp 1679235063
transform 1 0 19136 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_344
timestamp 1679235063
transform 1 0 24288 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_345
timestamp 1679235063
transform 1 0 6256 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_346
timestamp 1679235063
transform 1 0 11408 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_347
timestamp 1679235063
transform 1 0 16560 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_348
timestamp 1679235063
transform 1 0 21712 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_349
timestamp 1679235063
transform 1 0 3680 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_350
timestamp 1679235063
transform 1 0 8832 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_351
timestamp 1679235063
transform 1 0 13984 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_352
timestamp 1679235063
transform 1 0 19136 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_353
timestamp 1679235063
transform 1 0 24288 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_354
timestamp 1679235063
transform 1 0 6256 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_355
timestamp 1679235063
transform 1 0 11408 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_356
timestamp 1679235063
transform 1 0 16560 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_357
timestamp 1679235063
transform 1 0 21712 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_358
timestamp 1679235063
transform 1 0 3680 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_359
timestamp 1679235063
transform 1 0 8832 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_360
timestamp 1679235063
transform 1 0 13984 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_361
timestamp 1679235063
transform 1 0 19136 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_362
timestamp 1679235063
transform 1 0 24288 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_363
timestamp 1679235063
transform 1 0 6256 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_364
timestamp 1679235063
transform 1 0 11408 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_365
timestamp 1679235063
transform 1 0 16560 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_366
timestamp 1679235063
transform 1 0 21712 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_367
timestamp 1679235063
transform 1 0 3680 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_368
timestamp 1679235063
transform 1 0 8832 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_369
timestamp 1679235063
transform 1 0 13984 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_370
timestamp 1679235063
transform 1 0 19136 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_371
timestamp 1679235063
transform 1 0 24288 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_372
timestamp 1679235063
transform 1 0 6256 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_373
timestamp 1679235063
transform 1 0 11408 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_374
timestamp 1679235063
transform 1 0 16560 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_375
timestamp 1679235063
transform 1 0 21712 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_376
timestamp 1679235063
transform 1 0 3680 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_377
timestamp 1679235063
transform 1 0 8832 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_378
timestamp 1679235063
transform 1 0 13984 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_379
timestamp 1679235063
transform 1 0 19136 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_380
timestamp 1679235063
transform 1 0 24288 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_381
timestamp 1679235063
transform 1 0 6256 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_382
timestamp 1679235063
transform 1 0 11408 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_383
timestamp 1679235063
transform 1 0 16560 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_384
timestamp 1679235063
transform 1 0 21712 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_385
timestamp 1679235063
transform 1 0 3680 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_386
timestamp 1679235063
transform 1 0 8832 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_387
timestamp 1679235063
transform 1 0 13984 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_388
timestamp 1679235063
transform 1 0 19136 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_389
timestamp 1679235063
transform 1 0 24288 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_390
timestamp 1679235063
transform 1 0 6256 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_391
timestamp 1679235063
transform 1 0 11408 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_392
timestamp 1679235063
transform 1 0 16560 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_393
timestamp 1679235063
transform 1 0 21712 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_394
timestamp 1679235063
transform 1 0 3680 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_395
timestamp 1679235063
transform 1 0 8832 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_396
timestamp 1679235063
transform 1 0 13984 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_397
timestamp 1679235063
transform 1 0 19136 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_398
timestamp 1679235063
transform 1 0 24288 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_399
timestamp 1679235063
transform 1 0 6256 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_400
timestamp 1679235063
transform 1 0 11408 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_401
timestamp 1679235063
transform 1 0 16560 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_402
timestamp 1679235063
transform 1 0 21712 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_403
timestamp 1679235063
transform 1 0 3680 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_404
timestamp 1679235063
transform 1 0 8832 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_405
timestamp 1679235063
transform 1 0 13984 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_406
timestamp 1679235063
transform 1 0 19136 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_407
timestamp 1679235063
transform 1 0 24288 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_408
timestamp 1679235063
transform 1 0 6256 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_409
timestamp 1679235063
transform 1 0 11408 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_410
timestamp 1679235063
transform 1 0 16560 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_411
timestamp 1679235063
transform 1 0 21712 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_412
timestamp 1679235063
transform 1 0 3680 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_413
timestamp 1679235063
transform 1 0 8832 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_414
timestamp 1679235063
transform 1 0 13984 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_415
timestamp 1679235063
transform 1 0 19136 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_416
timestamp 1679235063
transform 1 0 24288 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_417
timestamp 1679235063
transform 1 0 6256 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_418
timestamp 1679235063
transform 1 0 11408 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_419
timestamp 1679235063
transform 1 0 16560 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_420
timestamp 1679235063
transform 1 0 21712 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_421
timestamp 1679235063
transform 1 0 3680 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_422
timestamp 1679235063
transform 1 0 8832 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_423
timestamp 1679235063
transform 1 0 13984 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_424
timestamp 1679235063
transform 1 0 19136 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_425
timestamp 1679235063
transform 1 0 24288 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_426
timestamp 1679235063
transform 1 0 6256 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_427
timestamp 1679235063
transform 1 0 11408 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_428
timestamp 1679235063
transform 1 0 16560 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_429
timestamp 1679235063
transform 1 0 21712 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_430
timestamp 1679235063
transform 1 0 3680 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_431
timestamp 1679235063
transform 1 0 8832 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_432
timestamp 1679235063
transform 1 0 13984 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_433
timestamp 1679235063
transform 1 0 19136 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_434
timestamp 1679235063
transform 1 0 24288 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_435
timestamp 1679235063
transform 1 0 6256 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_436
timestamp 1679235063
transform 1 0 11408 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_437
timestamp 1679235063
transform 1 0 16560 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_438
timestamp 1679235063
transform 1 0 21712 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_439
timestamp 1679235063
transform 1 0 3680 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_440
timestamp 1679235063
transform 1 0 8832 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_441
timestamp 1679235063
transform 1 0 13984 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_442
timestamp 1679235063
transform 1 0 19136 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_443
timestamp 1679235063
transform 1 0 24288 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_444
timestamp 1679235063
transform 1 0 6256 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_445
timestamp 1679235063
transform 1 0 11408 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_446
timestamp 1679235063
transform 1 0 16560 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_447
timestamp 1679235063
transform 1 0 21712 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_448
timestamp 1679235063
transform 1 0 3680 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_449
timestamp 1679235063
transform 1 0 8832 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_450
timestamp 1679235063
transform 1 0 13984 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_451
timestamp 1679235063
transform 1 0 19136 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_452
timestamp 1679235063
transform 1 0 24288 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_453
timestamp 1679235063
transform 1 0 6256 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_454
timestamp 1679235063
transform 1 0 11408 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_455
timestamp 1679235063
transform 1 0 16560 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_456
timestamp 1679235063
transform 1 0 21712 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_457
timestamp 1679235063
transform 1 0 3680 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_458
timestamp 1679235063
transform 1 0 8832 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_459
timestamp 1679235063
transform 1 0 13984 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_460
timestamp 1679235063
transform 1 0 19136 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_461
timestamp 1679235063
transform 1 0 24288 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_462
timestamp 1679235063
transform 1 0 6256 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_463
timestamp 1679235063
transform 1 0 11408 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_464
timestamp 1679235063
transform 1 0 16560 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_465
timestamp 1679235063
transform 1 0 21712 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_466
timestamp 1679235063
transform 1 0 3680 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_467
timestamp 1679235063
transform 1 0 8832 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_468
timestamp 1679235063
transform 1 0 13984 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_469
timestamp 1679235063
transform 1 0 19136 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_470
timestamp 1679235063
transform 1 0 24288 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_471
timestamp 1679235063
transform 1 0 6256 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_472
timestamp 1679235063
transform 1 0 11408 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_473
timestamp 1679235063
transform 1 0 16560 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_474
timestamp 1679235063
transform 1 0 21712 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_475
timestamp 1679235063
transform 1 0 3680 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_476
timestamp 1679235063
transform 1 0 8832 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_477
timestamp 1679235063
transform 1 0 13984 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_478
timestamp 1679235063
transform 1 0 19136 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_479
timestamp 1679235063
transform 1 0 24288 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_480
timestamp 1679235063
transform 1 0 6256 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_481
timestamp 1679235063
transform 1 0 11408 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_482
timestamp 1679235063
transform 1 0 16560 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_483
timestamp 1679235063
transform 1 0 21712 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_484
timestamp 1679235063
transform 1 0 3680 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_485
timestamp 1679235063
transform 1 0 8832 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_486
timestamp 1679235063
transform 1 0 13984 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_487
timestamp 1679235063
transform 1 0 19136 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_488
timestamp 1679235063
transform 1 0 24288 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_489
timestamp 1679235063
transform 1 0 6256 0 -1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_490
timestamp 1679235063
transform 1 0 11408 0 -1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_491
timestamp 1679235063
transform 1 0 16560 0 -1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_492
timestamp 1679235063
transform 1 0 21712 0 -1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_493
timestamp 1679235063
transform 1 0 3680 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_494
timestamp 1679235063
transform 1 0 8832 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_495
timestamp 1679235063
transform 1 0 13984 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_496
timestamp 1679235063
transform 1 0 19136 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_497
timestamp 1679235063
transform 1 0 24288 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_498
timestamp 1679235063
transform 1 0 6256 0 -1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_499
timestamp 1679235063
transform 1 0 11408 0 -1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_500
timestamp 1679235063
transform 1 0 16560 0 -1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_501
timestamp 1679235063
transform 1 0 21712 0 -1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_502
timestamp 1679235063
transform 1 0 3680 0 1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_503
timestamp 1679235063
transform 1 0 8832 0 1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_504
timestamp 1679235063
transform 1 0 13984 0 1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_505
timestamp 1679235063
transform 1 0 19136 0 1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_506
timestamp 1679235063
transform 1 0 24288 0 1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_507
timestamp 1679235063
transform 1 0 6256 0 -1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_508
timestamp 1679235063
transform 1 0 11408 0 -1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_509
timestamp 1679235063
transform 1 0 16560 0 -1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_510
timestamp 1679235063
transform 1 0 21712 0 -1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_511
timestamp 1679235063
transform 1 0 3680 0 1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_512
timestamp 1679235063
transform 1 0 8832 0 1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_513
timestamp 1679235063
transform 1 0 13984 0 1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_514
timestamp 1679235063
transform 1 0 19136 0 1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_515
timestamp 1679235063
transform 1 0 24288 0 1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_516
timestamp 1679235063
transform 1 0 6256 0 -1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_517
timestamp 1679235063
transform 1 0 11408 0 -1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_518
timestamp 1679235063
transform 1 0 16560 0 -1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_519
timestamp 1679235063
transform 1 0 21712 0 -1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_520
timestamp 1679235063
transform 1 0 3680 0 1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_521
timestamp 1679235063
transform 1 0 8832 0 1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_522
timestamp 1679235063
transform 1 0 13984 0 1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_523
timestamp 1679235063
transform 1 0 19136 0 1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_524
timestamp 1679235063
transform 1 0 24288 0 1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_525
timestamp 1679235063
transform 1 0 6256 0 -1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_526
timestamp 1679235063
transform 1 0 11408 0 -1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_527
timestamp 1679235063
transform 1 0 16560 0 -1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_528
timestamp 1679235063
transform 1 0 21712 0 -1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_529
timestamp 1679235063
transform 1 0 3680 0 1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_530
timestamp 1679235063
transform 1 0 8832 0 1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_531
timestamp 1679235063
transform 1 0 13984 0 1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_532
timestamp 1679235063
transform 1 0 19136 0 1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_533
timestamp 1679235063
transform 1 0 24288 0 1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_534
timestamp 1679235063
transform 1 0 6256 0 -1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_535
timestamp 1679235063
transform 1 0 11408 0 -1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_536
timestamp 1679235063
transform 1 0 16560 0 -1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_537
timestamp 1679235063
transform 1 0 21712 0 -1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_538
timestamp 1679235063
transform 1 0 3680 0 1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_539
timestamp 1679235063
transform 1 0 8832 0 1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_540
timestamp 1679235063
transform 1 0 13984 0 1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_541
timestamp 1679235063
transform 1 0 19136 0 1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_542
timestamp 1679235063
transform 1 0 24288 0 1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_543
timestamp 1679235063
transform 1 0 6256 0 -1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_544
timestamp 1679235063
transform 1 0 11408 0 -1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_545
timestamp 1679235063
transform 1 0 16560 0 -1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_546
timestamp 1679235063
transform 1 0 21712 0 -1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_547
timestamp 1679235063
transform 1 0 3680 0 1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_548
timestamp 1679235063
transform 1 0 8832 0 1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_549
timestamp 1679235063
transform 1 0 13984 0 1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_550
timestamp 1679235063
transform 1 0 19136 0 1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_551
timestamp 1679235063
transform 1 0 24288 0 1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_552
timestamp 1679235063
transform 1 0 6256 0 -1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_553
timestamp 1679235063
transform 1 0 11408 0 -1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_554
timestamp 1679235063
transform 1 0 16560 0 -1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_555
timestamp 1679235063
transform 1 0 21712 0 -1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_556
timestamp 1679235063
transform 1 0 3680 0 1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_557
timestamp 1679235063
transform 1 0 8832 0 1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_558
timestamp 1679235063
transform 1 0 13984 0 1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_559
timestamp 1679235063
transform 1 0 19136 0 1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_560
timestamp 1679235063
transform 1 0 24288 0 1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_561
timestamp 1679235063
transform 1 0 6256 0 -1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_562
timestamp 1679235063
transform 1 0 11408 0 -1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_563
timestamp 1679235063
transform 1 0 16560 0 -1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_564
timestamp 1679235063
transform 1 0 21712 0 -1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_565
timestamp 1679235063
transform 1 0 3680 0 1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_566
timestamp 1679235063
transform 1 0 8832 0 1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_567
timestamp 1679235063
transform 1 0 13984 0 1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_568
timestamp 1679235063
transform 1 0 19136 0 1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_569
timestamp 1679235063
transform 1 0 24288 0 1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_570
timestamp 1679235063
transform 1 0 6256 0 -1 47872
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_571
timestamp 1679235063
transform 1 0 11408 0 -1 47872
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_572
timestamp 1679235063
transform 1 0 16560 0 -1 47872
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_573
timestamp 1679235063
transform 1 0 21712 0 -1 47872
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_574
timestamp 1679235063
transform 1 0 3680 0 1 47872
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_575
timestamp 1679235063
transform 1 0 8832 0 1 47872
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_576
timestamp 1679235063
transform 1 0 13984 0 1 47872
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_577
timestamp 1679235063
transform 1 0 19136 0 1 47872
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_578
timestamp 1679235063
transform 1 0 24288 0 1 47872
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_579
timestamp 1679235063
transform 1 0 6256 0 -1 48960
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_580
timestamp 1679235063
transform 1 0 11408 0 -1 48960
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_581
timestamp 1679235063
transform 1 0 16560 0 -1 48960
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_582
timestamp 1679235063
transform 1 0 21712 0 -1 48960
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_583
timestamp 1679235063
transform 1 0 3680 0 1 48960
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_584
timestamp 1679235063
transform 1 0 8832 0 1 48960
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_585
timestamp 1679235063
transform 1 0 13984 0 1 48960
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_586
timestamp 1679235063
transform 1 0 19136 0 1 48960
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_587
timestamp 1679235063
transform 1 0 24288 0 1 48960
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_588
timestamp 1679235063
transform 1 0 6256 0 -1 50048
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_589
timestamp 1679235063
transform 1 0 11408 0 -1 50048
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_590
timestamp 1679235063
transform 1 0 16560 0 -1 50048
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_591
timestamp 1679235063
transform 1 0 21712 0 -1 50048
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_592
timestamp 1679235063
transform 1 0 3680 0 1 50048
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_593
timestamp 1679235063
transform 1 0 8832 0 1 50048
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_594
timestamp 1679235063
transform 1 0 13984 0 1 50048
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_595
timestamp 1679235063
transform 1 0 19136 0 1 50048
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_596
timestamp 1679235063
transform 1 0 24288 0 1 50048
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_597
timestamp 1679235063
transform 1 0 6256 0 -1 51136
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_598
timestamp 1679235063
transform 1 0 11408 0 -1 51136
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_599
timestamp 1679235063
transform 1 0 16560 0 -1 51136
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_600
timestamp 1679235063
transform 1 0 21712 0 -1 51136
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_601
timestamp 1679235063
transform 1 0 3680 0 1 51136
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_602
timestamp 1679235063
transform 1 0 8832 0 1 51136
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_603
timestamp 1679235063
transform 1 0 13984 0 1 51136
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_604
timestamp 1679235063
transform 1 0 19136 0 1 51136
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_605
timestamp 1679235063
transform 1 0 24288 0 1 51136
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_606
timestamp 1679235063
transform 1 0 6256 0 -1 52224
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_607
timestamp 1679235063
transform 1 0 11408 0 -1 52224
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_608
timestamp 1679235063
transform 1 0 16560 0 -1 52224
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_609
timestamp 1679235063
transform 1 0 21712 0 -1 52224
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_610
timestamp 1679235063
transform 1 0 3680 0 1 52224
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_611
timestamp 1679235063
transform 1 0 8832 0 1 52224
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_612
timestamp 1679235063
transform 1 0 13984 0 1 52224
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_613
timestamp 1679235063
transform 1 0 19136 0 1 52224
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_614
timestamp 1679235063
transform 1 0 24288 0 1 52224
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_615
timestamp 1679235063
transform 1 0 6256 0 -1 53312
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_616
timestamp 1679235063
transform 1 0 11408 0 -1 53312
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_617
timestamp 1679235063
transform 1 0 16560 0 -1 53312
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_618
timestamp 1679235063
transform 1 0 21712 0 -1 53312
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_619
timestamp 1679235063
transform 1 0 3680 0 1 53312
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_620
timestamp 1679235063
transform 1 0 8832 0 1 53312
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_621
timestamp 1679235063
transform 1 0 13984 0 1 53312
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_622
timestamp 1679235063
transform 1 0 19136 0 1 53312
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_623
timestamp 1679235063
transform 1 0 24288 0 1 53312
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_624
timestamp 1679235063
transform 1 0 3680 0 -1 54400
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_625
timestamp 1679235063
transform 1 0 6256 0 -1 54400
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_626
timestamp 1679235063
transform 1 0 8832 0 -1 54400
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_627
timestamp 1679235063
transform 1 0 11408 0 -1 54400
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_628
timestamp 1679235063
transform 1 0 13984 0 -1 54400
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_629
timestamp 1679235063
transform 1 0 16560 0 -1 54400
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_630
timestamp 1679235063
transform 1 0 19136 0 -1 54400
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_631
timestamp 1679235063
transform 1 0 21712 0 -1 54400
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_632
timestamp 1679235063
transform 1 0 24288 0 -1 54400
box -38 -48 130 592
<< labels >>
flabel metal4 s 7944 2128 8264 54448 0 FreeSans 1920 90 0 0 VGND
port 0 nsew ground bidirectional
flabel metal4 s 17944 2128 18264 54448 0 FreeSans 1920 90 0 0 VGND
port 0 nsew ground bidirectional
flabel metal4 s 2944 2128 3264 54448 0 FreeSans 1920 90 0 0 VPWR
port 1 nsew power bidirectional
flabel metal4 s 12944 2128 13264 54448 0 FreeSans 1920 90 0 0 VPWR
port 1 nsew power bidirectional
flabel metal4 s 22944 2128 23264 54448 0 FreeSans 1920 90 0 0 VPWR
port 1 nsew power bidirectional
flabel metal2 s 25870 56200 25926 57000 0 FreeSans 224 90 0 0 ccff_head
port 2 nsew signal input
flabel metal2 s 1490 0 1546 800 0 FreeSans 224 90 0 0 ccff_head_0
port 3 nsew signal input
flabel metal3 s 26200 688 27000 808 0 FreeSans 480 0 0 0 ccff_tail
port 4 nsew signal tristate
flabel metal2 s 1030 56200 1086 57000 0 FreeSans 224 90 0 0 ccff_tail_0
port 5 nsew signal tristate
flabel metal3 s 26200 25984 27000 26104 0 FreeSans 480 0 0 0 chanx_right_in[0]
port 6 nsew signal input
flabel metal3 s 26200 34144 27000 34264 0 FreeSans 480 0 0 0 chanx_right_in[10]
port 7 nsew signal input
flabel metal3 s 26200 34960 27000 35080 0 FreeSans 480 0 0 0 chanx_right_in[11]
port 8 nsew signal input
flabel metal3 s 26200 35776 27000 35896 0 FreeSans 480 0 0 0 chanx_right_in[12]
port 9 nsew signal input
flabel metal3 s 26200 36592 27000 36712 0 FreeSans 480 0 0 0 chanx_right_in[13]
port 10 nsew signal input
flabel metal3 s 26200 37408 27000 37528 0 FreeSans 480 0 0 0 chanx_right_in[14]
port 11 nsew signal input
flabel metal3 s 26200 38224 27000 38344 0 FreeSans 480 0 0 0 chanx_right_in[15]
port 12 nsew signal input
flabel metal3 s 26200 39040 27000 39160 0 FreeSans 480 0 0 0 chanx_right_in[16]
port 13 nsew signal input
flabel metal3 s 26200 39856 27000 39976 0 FreeSans 480 0 0 0 chanx_right_in[17]
port 14 nsew signal input
flabel metal3 s 26200 40672 27000 40792 0 FreeSans 480 0 0 0 chanx_right_in[18]
port 15 nsew signal input
flabel metal3 s 26200 41488 27000 41608 0 FreeSans 480 0 0 0 chanx_right_in[19]
port 16 nsew signal input
flabel metal3 s 26200 26800 27000 26920 0 FreeSans 480 0 0 0 chanx_right_in[1]
port 17 nsew signal input
flabel metal3 s 26200 42304 27000 42424 0 FreeSans 480 0 0 0 chanx_right_in[20]
port 18 nsew signal input
flabel metal3 s 26200 43120 27000 43240 0 FreeSans 480 0 0 0 chanx_right_in[21]
port 19 nsew signal input
flabel metal3 s 26200 43936 27000 44056 0 FreeSans 480 0 0 0 chanx_right_in[22]
port 20 nsew signal input
flabel metal3 s 26200 44752 27000 44872 0 FreeSans 480 0 0 0 chanx_right_in[23]
port 21 nsew signal input
flabel metal3 s 26200 45568 27000 45688 0 FreeSans 480 0 0 0 chanx_right_in[24]
port 22 nsew signal input
flabel metal3 s 26200 46384 27000 46504 0 FreeSans 480 0 0 0 chanx_right_in[25]
port 23 nsew signal input
flabel metal3 s 26200 47200 27000 47320 0 FreeSans 480 0 0 0 chanx_right_in[26]
port 24 nsew signal input
flabel metal3 s 26200 48016 27000 48136 0 FreeSans 480 0 0 0 chanx_right_in[27]
port 25 nsew signal input
flabel metal3 s 26200 48832 27000 48952 0 FreeSans 480 0 0 0 chanx_right_in[28]
port 26 nsew signal input
flabel metal3 s 26200 49648 27000 49768 0 FreeSans 480 0 0 0 chanx_right_in[29]
port 27 nsew signal input
flabel metal3 s 26200 27616 27000 27736 0 FreeSans 480 0 0 0 chanx_right_in[2]
port 28 nsew signal input
flabel metal3 s 26200 28432 27000 28552 0 FreeSans 480 0 0 0 chanx_right_in[3]
port 29 nsew signal input
flabel metal3 s 26200 29248 27000 29368 0 FreeSans 480 0 0 0 chanx_right_in[4]
port 30 nsew signal input
flabel metal3 s 26200 30064 27000 30184 0 FreeSans 480 0 0 0 chanx_right_in[5]
port 31 nsew signal input
flabel metal3 s 26200 30880 27000 31000 0 FreeSans 480 0 0 0 chanx_right_in[6]
port 32 nsew signal input
flabel metal3 s 26200 31696 27000 31816 0 FreeSans 480 0 0 0 chanx_right_in[7]
port 33 nsew signal input
flabel metal3 s 26200 32512 27000 32632 0 FreeSans 480 0 0 0 chanx_right_in[8]
port 34 nsew signal input
flabel metal3 s 26200 33328 27000 33448 0 FreeSans 480 0 0 0 chanx_right_in[9]
port 35 nsew signal input
flabel metal3 s 26200 1504 27000 1624 0 FreeSans 480 0 0 0 chanx_right_out[0]
port 36 nsew signal tristate
flabel metal3 s 26200 9664 27000 9784 0 FreeSans 480 0 0 0 chanx_right_out[10]
port 37 nsew signal tristate
flabel metal3 s 26200 10480 27000 10600 0 FreeSans 480 0 0 0 chanx_right_out[11]
port 38 nsew signal tristate
flabel metal3 s 26200 11296 27000 11416 0 FreeSans 480 0 0 0 chanx_right_out[12]
port 39 nsew signal tristate
flabel metal3 s 26200 12112 27000 12232 0 FreeSans 480 0 0 0 chanx_right_out[13]
port 40 nsew signal tristate
flabel metal3 s 26200 12928 27000 13048 0 FreeSans 480 0 0 0 chanx_right_out[14]
port 41 nsew signal tristate
flabel metal3 s 26200 13744 27000 13864 0 FreeSans 480 0 0 0 chanx_right_out[15]
port 42 nsew signal tristate
flabel metal3 s 26200 14560 27000 14680 0 FreeSans 480 0 0 0 chanx_right_out[16]
port 43 nsew signal tristate
flabel metal3 s 26200 15376 27000 15496 0 FreeSans 480 0 0 0 chanx_right_out[17]
port 44 nsew signal tristate
flabel metal3 s 26200 16192 27000 16312 0 FreeSans 480 0 0 0 chanx_right_out[18]
port 45 nsew signal tristate
flabel metal3 s 26200 17008 27000 17128 0 FreeSans 480 0 0 0 chanx_right_out[19]
port 46 nsew signal tristate
flabel metal3 s 26200 2320 27000 2440 0 FreeSans 480 0 0 0 chanx_right_out[1]
port 47 nsew signal tristate
flabel metal3 s 26200 17824 27000 17944 0 FreeSans 480 0 0 0 chanx_right_out[20]
port 48 nsew signal tristate
flabel metal3 s 26200 18640 27000 18760 0 FreeSans 480 0 0 0 chanx_right_out[21]
port 49 nsew signal tristate
flabel metal3 s 26200 19456 27000 19576 0 FreeSans 480 0 0 0 chanx_right_out[22]
port 50 nsew signal tristate
flabel metal3 s 26200 20272 27000 20392 0 FreeSans 480 0 0 0 chanx_right_out[23]
port 51 nsew signal tristate
flabel metal3 s 26200 21088 27000 21208 0 FreeSans 480 0 0 0 chanx_right_out[24]
port 52 nsew signal tristate
flabel metal3 s 26200 21904 27000 22024 0 FreeSans 480 0 0 0 chanx_right_out[25]
port 53 nsew signal tristate
flabel metal3 s 26200 22720 27000 22840 0 FreeSans 480 0 0 0 chanx_right_out[26]
port 54 nsew signal tristate
flabel metal3 s 26200 23536 27000 23656 0 FreeSans 480 0 0 0 chanx_right_out[27]
port 55 nsew signal tristate
flabel metal3 s 26200 24352 27000 24472 0 FreeSans 480 0 0 0 chanx_right_out[28]
port 56 nsew signal tristate
flabel metal3 s 26200 25168 27000 25288 0 FreeSans 480 0 0 0 chanx_right_out[29]
port 57 nsew signal tristate
flabel metal3 s 26200 3136 27000 3256 0 FreeSans 480 0 0 0 chanx_right_out[2]
port 58 nsew signal tristate
flabel metal3 s 26200 3952 27000 4072 0 FreeSans 480 0 0 0 chanx_right_out[3]
port 59 nsew signal tristate
flabel metal3 s 26200 4768 27000 4888 0 FreeSans 480 0 0 0 chanx_right_out[4]
port 60 nsew signal tristate
flabel metal3 s 26200 5584 27000 5704 0 FreeSans 480 0 0 0 chanx_right_out[5]
port 61 nsew signal tristate
flabel metal3 s 26200 6400 27000 6520 0 FreeSans 480 0 0 0 chanx_right_out[6]
port 62 nsew signal tristate
flabel metal3 s 26200 7216 27000 7336 0 FreeSans 480 0 0 0 chanx_right_out[7]
port 63 nsew signal tristate
flabel metal3 s 26200 8032 27000 8152 0 FreeSans 480 0 0 0 chanx_right_out[8]
port 64 nsew signal tristate
flabel metal3 s 26200 8848 27000 8968 0 FreeSans 480 0 0 0 chanx_right_out[9]
port 65 nsew signal tristate
flabel metal2 s 1858 0 1914 800 0 FreeSans 224 90 0 0 chany_bottom_in_0[0]
port 66 nsew signal input
flabel metal2 s 5538 0 5594 800 0 FreeSans 224 90 0 0 chany_bottom_in_0[10]
port 67 nsew signal input
flabel metal2 s 5906 0 5962 800 0 FreeSans 224 90 0 0 chany_bottom_in_0[11]
port 68 nsew signal input
flabel metal2 s 6274 0 6330 800 0 FreeSans 224 90 0 0 chany_bottom_in_0[12]
port 69 nsew signal input
flabel metal2 s 6642 0 6698 800 0 FreeSans 224 90 0 0 chany_bottom_in_0[13]
port 70 nsew signal input
flabel metal2 s 7010 0 7066 800 0 FreeSans 224 90 0 0 chany_bottom_in_0[14]
port 71 nsew signal input
flabel metal2 s 7378 0 7434 800 0 FreeSans 224 90 0 0 chany_bottom_in_0[15]
port 72 nsew signal input
flabel metal2 s 7746 0 7802 800 0 FreeSans 224 90 0 0 chany_bottom_in_0[16]
port 73 nsew signal input
flabel metal2 s 8114 0 8170 800 0 FreeSans 224 90 0 0 chany_bottom_in_0[17]
port 74 nsew signal input
flabel metal2 s 8482 0 8538 800 0 FreeSans 224 90 0 0 chany_bottom_in_0[18]
port 75 nsew signal input
flabel metal2 s 8850 0 8906 800 0 FreeSans 224 90 0 0 chany_bottom_in_0[19]
port 76 nsew signal input
flabel metal2 s 2226 0 2282 800 0 FreeSans 224 90 0 0 chany_bottom_in_0[1]
port 77 nsew signal input
flabel metal2 s 9218 0 9274 800 0 FreeSans 224 90 0 0 chany_bottom_in_0[20]
port 78 nsew signal input
flabel metal2 s 9586 0 9642 800 0 FreeSans 224 90 0 0 chany_bottom_in_0[21]
port 79 nsew signal input
flabel metal2 s 9954 0 10010 800 0 FreeSans 224 90 0 0 chany_bottom_in_0[22]
port 80 nsew signal input
flabel metal2 s 10322 0 10378 800 0 FreeSans 224 90 0 0 chany_bottom_in_0[23]
port 81 nsew signal input
flabel metal2 s 10690 0 10746 800 0 FreeSans 224 90 0 0 chany_bottom_in_0[24]
port 82 nsew signal input
flabel metal2 s 11058 0 11114 800 0 FreeSans 224 90 0 0 chany_bottom_in_0[25]
port 83 nsew signal input
flabel metal2 s 11426 0 11482 800 0 FreeSans 224 90 0 0 chany_bottom_in_0[26]
port 84 nsew signal input
flabel metal2 s 11794 0 11850 800 0 FreeSans 224 90 0 0 chany_bottom_in_0[27]
port 85 nsew signal input
flabel metal2 s 12162 0 12218 800 0 FreeSans 224 90 0 0 chany_bottom_in_0[28]
port 86 nsew signal input
flabel metal2 s 12530 0 12586 800 0 FreeSans 224 90 0 0 chany_bottom_in_0[29]
port 87 nsew signal input
flabel metal2 s 2594 0 2650 800 0 FreeSans 224 90 0 0 chany_bottom_in_0[2]
port 88 nsew signal input
flabel metal2 s 2962 0 3018 800 0 FreeSans 224 90 0 0 chany_bottom_in_0[3]
port 89 nsew signal input
flabel metal2 s 3330 0 3386 800 0 FreeSans 224 90 0 0 chany_bottom_in_0[4]
port 90 nsew signal input
flabel metal2 s 3698 0 3754 800 0 FreeSans 224 90 0 0 chany_bottom_in_0[5]
port 91 nsew signal input
flabel metal2 s 4066 0 4122 800 0 FreeSans 224 90 0 0 chany_bottom_in_0[6]
port 92 nsew signal input
flabel metal2 s 4434 0 4490 800 0 FreeSans 224 90 0 0 chany_bottom_in_0[7]
port 93 nsew signal input
flabel metal2 s 4802 0 4858 800 0 FreeSans 224 90 0 0 chany_bottom_in_0[8]
port 94 nsew signal input
flabel metal2 s 5170 0 5226 800 0 FreeSans 224 90 0 0 chany_bottom_in_0[9]
port 95 nsew signal input
flabel metal2 s 12898 0 12954 800 0 FreeSans 224 90 0 0 chany_bottom_out_0[0]
port 96 nsew signal tristate
flabel metal2 s 16578 0 16634 800 0 FreeSans 224 90 0 0 chany_bottom_out_0[10]
port 97 nsew signal tristate
flabel metal2 s 16946 0 17002 800 0 FreeSans 224 90 0 0 chany_bottom_out_0[11]
port 98 nsew signal tristate
flabel metal2 s 17314 0 17370 800 0 FreeSans 224 90 0 0 chany_bottom_out_0[12]
port 99 nsew signal tristate
flabel metal2 s 17682 0 17738 800 0 FreeSans 224 90 0 0 chany_bottom_out_0[13]
port 100 nsew signal tristate
flabel metal2 s 18050 0 18106 800 0 FreeSans 224 90 0 0 chany_bottom_out_0[14]
port 101 nsew signal tristate
flabel metal2 s 18418 0 18474 800 0 FreeSans 224 90 0 0 chany_bottom_out_0[15]
port 102 nsew signal tristate
flabel metal2 s 18786 0 18842 800 0 FreeSans 224 90 0 0 chany_bottom_out_0[16]
port 103 nsew signal tristate
flabel metal2 s 19154 0 19210 800 0 FreeSans 224 90 0 0 chany_bottom_out_0[17]
port 104 nsew signal tristate
flabel metal2 s 19522 0 19578 800 0 FreeSans 224 90 0 0 chany_bottom_out_0[18]
port 105 nsew signal tristate
flabel metal2 s 19890 0 19946 800 0 FreeSans 224 90 0 0 chany_bottom_out_0[19]
port 106 nsew signal tristate
flabel metal2 s 13266 0 13322 800 0 FreeSans 224 90 0 0 chany_bottom_out_0[1]
port 107 nsew signal tristate
flabel metal2 s 20258 0 20314 800 0 FreeSans 224 90 0 0 chany_bottom_out_0[20]
port 108 nsew signal tristate
flabel metal2 s 20626 0 20682 800 0 FreeSans 224 90 0 0 chany_bottom_out_0[21]
port 109 nsew signal tristate
flabel metal2 s 20994 0 21050 800 0 FreeSans 224 90 0 0 chany_bottom_out_0[22]
port 110 nsew signal tristate
flabel metal2 s 21362 0 21418 800 0 FreeSans 224 90 0 0 chany_bottom_out_0[23]
port 111 nsew signal tristate
flabel metal2 s 21730 0 21786 800 0 FreeSans 224 90 0 0 chany_bottom_out_0[24]
port 112 nsew signal tristate
flabel metal2 s 22098 0 22154 800 0 FreeSans 224 90 0 0 chany_bottom_out_0[25]
port 113 nsew signal tristate
flabel metal2 s 22466 0 22522 800 0 FreeSans 224 90 0 0 chany_bottom_out_0[26]
port 114 nsew signal tristate
flabel metal2 s 22834 0 22890 800 0 FreeSans 224 90 0 0 chany_bottom_out_0[27]
port 115 nsew signal tristate
flabel metal2 s 23202 0 23258 800 0 FreeSans 224 90 0 0 chany_bottom_out_0[28]
port 116 nsew signal tristate
flabel metal2 s 23570 0 23626 800 0 FreeSans 224 90 0 0 chany_bottom_out_0[29]
port 117 nsew signal tristate
flabel metal2 s 13634 0 13690 800 0 FreeSans 224 90 0 0 chany_bottom_out_0[2]
port 118 nsew signal tristate
flabel metal2 s 14002 0 14058 800 0 FreeSans 224 90 0 0 chany_bottom_out_0[3]
port 119 nsew signal tristate
flabel metal2 s 14370 0 14426 800 0 FreeSans 224 90 0 0 chany_bottom_out_0[4]
port 120 nsew signal tristate
flabel metal2 s 14738 0 14794 800 0 FreeSans 224 90 0 0 chany_bottom_out_0[5]
port 121 nsew signal tristate
flabel metal2 s 15106 0 15162 800 0 FreeSans 224 90 0 0 chany_bottom_out_0[6]
port 122 nsew signal tristate
flabel metal2 s 15474 0 15530 800 0 FreeSans 224 90 0 0 chany_bottom_out_0[7]
port 123 nsew signal tristate
flabel metal2 s 15842 0 15898 800 0 FreeSans 224 90 0 0 chany_bottom_out_0[8]
port 124 nsew signal tristate
flabel metal2 s 16210 0 16266 800 0 FreeSans 224 90 0 0 chany_bottom_out_0[9]
port 125 nsew signal tristate
flabel metal2 s 2410 56200 2466 57000 0 FreeSans 224 90 0 0 gfpga_pad_io_soc_dir[0]
port 126 nsew signal tristate
flabel metal2 s 3790 56200 3846 57000 0 FreeSans 224 90 0 0 gfpga_pad_io_soc_dir[1]
port 127 nsew signal tristate
flabel metal2 s 5170 56200 5226 57000 0 FreeSans 224 90 0 0 gfpga_pad_io_soc_dir[2]
port 128 nsew signal tristate
flabel metal2 s 6550 56200 6606 57000 0 FreeSans 224 90 0 0 gfpga_pad_io_soc_dir[3]
port 129 nsew signal tristate
flabel metal2 s 13450 56200 13506 57000 0 FreeSans 224 90 0 0 gfpga_pad_io_soc_in[0]
port 130 nsew signal input
flabel metal2 s 14830 56200 14886 57000 0 FreeSans 224 90 0 0 gfpga_pad_io_soc_in[1]
port 131 nsew signal input
flabel metal2 s 16210 56200 16266 57000 0 FreeSans 224 90 0 0 gfpga_pad_io_soc_in[2]
port 132 nsew signal input
flabel metal2 s 17590 56200 17646 57000 0 FreeSans 224 90 0 0 gfpga_pad_io_soc_in[3]
port 133 nsew signal input
flabel metal2 s 7930 56200 7986 57000 0 FreeSans 224 90 0 0 gfpga_pad_io_soc_out[0]
port 134 nsew signal tristate
flabel metal2 s 9310 56200 9366 57000 0 FreeSans 224 90 0 0 gfpga_pad_io_soc_out[1]
port 135 nsew signal tristate
flabel metal2 s 10690 56200 10746 57000 0 FreeSans 224 90 0 0 gfpga_pad_io_soc_out[2]
port 136 nsew signal tristate
flabel metal2 s 12070 56200 12126 57000 0 FreeSans 224 90 0 0 gfpga_pad_io_soc_out[3]
port 137 nsew signal tristate
flabel metal2 s 18970 56200 19026 57000 0 FreeSans 224 90 0 0 isol_n
port 138 nsew signal input
flabel metal2 s 23938 0 23994 800 0 FreeSans 224 90 0 0 prog_clk
port 139 nsew signal input
flabel metal2 s 24306 0 24362 800 0 FreeSans 224 90 0 0 prog_reset
port 140 nsew signal input
flabel metal2 s 24674 0 24730 800 0 FreeSans 224 90 0 0 reset
port 141 nsew signal input
flabel metal3 s 26200 50464 27000 50584 0 FreeSans 480 0 0 0 right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_
port 142 nsew signal input
flabel metal3 s 26200 51280 27000 51400 0 FreeSans 480 0 0 0 right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_
port 143 nsew signal input
flabel metal3 s 26200 52096 27000 52216 0 FreeSans 480 0 0 0 right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_
port 144 nsew signal input
flabel metal3 s 26200 52912 27000 53032 0 FreeSans 480 0 0 0 right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_
port 145 nsew signal input
flabel metal3 s 26200 53728 27000 53848 0 FreeSans 480 0 0 0 right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_4_
port 146 nsew signal input
flabel metal3 s 26200 54544 27000 54664 0 FreeSans 480 0 0 0 right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_5_
port 147 nsew signal input
flabel metal3 s 26200 55360 27000 55480 0 FreeSans 480 0 0 0 right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_6_
port 148 nsew signal input
flabel metal3 s 26200 56176 27000 56296 0 FreeSans 480 0 0 0 right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_7_
port 149 nsew signal input
flabel metal2 s 20350 56200 20406 57000 0 FreeSans 224 90 0 0 right_top_grid_bottom_width_0_height_0_subtile_0__pin_inpad_0_
port 150 nsew signal input
flabel metal2 s 21730 56200 21786 57000 0 FreeSans 224 90 0 0 right_top_grid_bottom_width_0_height_0_subtile_1__pin_inpad_0_
port 151 nsew signal input
flabel metal2 s 23110 56200 23166 57000 0 FreeSans 224 90 0 0 right_top_grid_bottom_width_0_height_0_subtile_2__pin_inpad_0_
port 152 nsew signal input
flabel metal2 s 24490 56200 24546 57000 0 FreeSans 224 90 0 0 right_top_grid_bottom_width_0_height_0_subtile_3__pin_inpad_0_
port 153 nsew signal input
flabel metal3 s 0 1776 800 1896 0 FreeSans 480 0 0 0 right_width_0_height_0_subtile_0__pin_inpad_0_
port 154 nsew signal tristate
flabel metal3 s 0 4088 800 4208 0 FreeSans 480 0 0 0 right_width_0_height_0_subtile_1__pin_inpad_0_
port 155 nsew signal tristate
flabel metal3 s 0 6400 800 6520 0 FreeSans 480 0 0 0 right_width_0_height_0_subtile_2__pin_inpad_0_
port 156 nsew signal tristate
flabel metal3 s 0 8712 800 8832 0 FreeSans 480 0 0 0 right_width_0_height_0_subtile_3__pin_inpad_0_
port 157 nsew signal tristate
flabel metal2 s 25042 0 25098 800 0 FreeSans 224 90 0 0 test_enable
port 158 nsew signal input
rlabel metal1 13478 54400 13478 54400 0 VGND
rlabel metal1 13478 53856 13478 53856 0 VPWR
rlabel metal1 9844 33490 9844 33490 0 cby_0__8_.cby_0__1_.ccff_tail
rlabel metal1 9798 33082 9798 33082 0 cby_0__8_.cby_0__1_.left_grid_right_width_0_height_0_subtile_0__pin_outpad_0_
rlabel metal1 9154 45390 9154 45390 0 cby_0__8_.cby_0__1_.left_grid_right_width_0_height_0_subtile_1__pin_outpad_0_
rlabel metal1 9108 36346 9108 36346 0 cby_0__8_.cby_0__1_.left_grid_right_width_0_height_0_subtile_2__pin_outpad_0_
rlabel metal1 8464 39610 8464 39610 0 cby_0__8_.cby_0__1_.left_grid_right_width_0_height_0_subtile_3__pin_outpad_0_
rlabel metal2 7682 18530 7682 18530 0 cby_0__8_.cby_0__1_.mem_right_ipin_0.ccff_tail
rlabel metal1 15640 9418 15640 9418 0 cby_0__8_.cby_0__1_.mem_right_ipin_0.mem_out\[0\]
rlabel metal1 9568 11662 9568 11662 0 cby_0__8_.cby_0__1_.mem_right_ipin_0.mem_out\[1\]
rlabel metal1 7958 13838 7958 13838 0 cby_0__8_.cby_0__1_.mem_right_ipin_0.mem_out\[2\]
rlabel metal1 7958 15674 7958 15674 0 cby_0__8_.cby_0__1_.mem_right_ipin_1.ccff_tail
rlabel metal1 15778 13328 15778 13328 0 cby_0__8_.cby_0__1_.mem_right_ipin_1.mem_out\[0\]
rlabel metal1 13386 11186 13386 11186 0 cby_0__8_.cby_0__1_.mem_right_ipin_1.mem_out\[1\]
rlabel metal1 9568 13838 9568 13838 0 cby_0__8_.cby_0__1_.mem_right_ipin_1.mem_out\[2\]
rlabel metal1 8556 21862 8556 21862 0 cby_0__8_.cby_0__1_.mem_right_ipin_2.ccff_tail
rlabel metal1 16790 10574 16790 10574 0 cby_0__8_.cby_0__1_.mem_right_ipin_2.mem_out\[0\]
rlabel metal1 12926 13804 12926 13804 0 cby_0__8_.cby_0__1_.mem_right_ipin_2.mem_out\[1\]
rlabel metal1 9292 19482 9292 19482 0 cby_0__8_.cby_0__1_.mem_right_ipin_2.mem_out\[2\]
rlabel metal1 9522 18326 9522 18326 0 cby_0__8_.cby_0__1_.mem_right_ipin_3.mem_out\[0\]
rlabel metal1 16238 26384 16238 26384 0 cby_0__8_.cby_0__1_.mem_right_ipin_3.mem_out\[1\]
rlabel metal1 10258 25330 10258 25330 0 cby_0__8_.cby_0__1_.mem_right_ipin_3.mem_out\[2\]
rlabel metal2 15686 11288 15686 11288 0 cby_0__8_.cby_0__1_.mux_right_ipin_0.sky130_fd_sc_hd__mux2_1_0_X
rlabel metal1 9108 14586 9108 14586 0 cby_0__8_.cby_0__1_.mux_right_ipin_0.sky130_fd_sc_hd__mux2_1_10_X
rlabel metal1 8694 20570 8694 20570 0 cby_0__8_.cby_0__1_.mux_right_ipin_0.sky130_fd_sc_hd__mux2_1_11_X
rlabel metal1 13846 10778 13846 10778 0 cby_0__8_.cby_0__1_.mux_right_ipin_0.sky130_fd_sc_hd__mux2_1_1_X
rlabel metal1 13478 10166 13478 10166 0 cby_0__8_.cby_0__1_.mux_right_ipin_0.sky130_fd_sc_hd__mux2_1_2_X
rlabel metal2 12328 13532 12328 13532 0 cby_0__8_.cby_0__1_.mux_right_ipin_0.sky130_fd_sc_hd__mux2_1_3_X
rlabel metal1 11178 12682 11178 12682 0 cby_0__8_.cby_0__1_.mux_right_ipin_0.sky130_fd_sc_hd__mux2_1_4_X
rlabel metal1 11086 14858 11086 14858 0 cby_0__8_.cby_0__1_.mux_right_ipin_0.sky130_fd_sc_hd__mux2_1_5_X
rlabel metal1 11408 15062 11408 15062 0 cby_0__8_.cby_0__1_.mux_right_ipin_0.sky130_fd_sc_hd__mux2_1_6_X
rlabel metal1 8970 11832 8970 11832 0 cby_0__8_.cby_0__1_.mux_right_ipin_0.sky130_fd_sc_hd__mux2_1_7_X
rlabel metal1 9982 14042 9982 14042 0 cby_0__8_.cby_0__1_.mux_right_ipin_0.sky130_fd_sc_hd__mux2_1_8_X
rlabel metal1 10212 14858 10212 14858 0 cby_0__8_.cby_0__1_.mux_right_ipin_0.sky130_fd_sc_hd__mux2_1_9_X
rlabel metal1 14536 8602 14536 8602 0 cby_0__8_.cby_0__1_.mux_right_ipin_1.sky130_fd_sc_hd__mux2_1_0_X
rlabel metal1 8740 14042 8740 14042 0 cby_0__8_.cby_0__1_.mux_right_ipin_1.sky130_fd_sc_hd__mux2_1_10_X
rlabel metal1 8924 32402 8924 32402 0 cby_0__8_.cby_0__1_.mux_right_ipin_1.sky130_fd_sc_hd__mux2_1_11_X
rlabel metal1 14490 8942 14490 8942 0 cby_0__8_.cby_0__1_.mux_right_ipin_1.sky130_fd_sc_hd__mux2_1_1_X
rlabel metal1 14490 9418 14490 9418 0 cby_0__8_.cby_0__1_.mux_right_ipin_1.sky130_fd_sc_hd__mux2_1_2_X
rlabel metal1 15318 13158 15318 13158 0 cby_0__8_.cby_0__1_.mux_right_ipin_1.sky130_fd_sc_hd__mux2_1_3_X
rlabel metal1 12926 14246 12926 14246 0 cby_0__8_.cby_0__1_.mux_right_ipin_1.sky130_fd_sc_hd__mux2_1_4_X
rlabel metal1 11408 12818 11408 12818 0 cby_0__8_.cby_0__1_.mux_right_ipin_1.sky130_fd_sc_hd__mux2_1_5_X
rlabel metal2 12650 12104 12650 12104 0 cby_0__8_.cby_0__1_.mux_right_ipin_1.sky130_fd_sc_hd__mux2_1_6_X
rlabel metal1 9706 13906 9706 13906 0 cby_0__8_.cby_0__1_.mux_right_ipin_1.sky130_fd_sc_hd__mux2_1_7_X
rlabel metal1 9844 13974 9844 13974 0 cby_0__8_.cby_0__1_.mux_right_ipin_1.sky130_fd_sc_hd__mux2_1_8_X
rlabel metal1 9384 12954 9384 12954 0 cby_0__8_.cby_0__1_.mux_right_ipin_1.sky130_fd_sc_hd__mux2_1_9_X
rlabel metal1 16744 10234 16744 10234 0 cby_0__8_.cby_0__1_.mux_right_ipin_2.sky130_fd_sc_hd__mux2_1_0_X
rlabel metal1 10074 21658 10074 21658 0 cby_0__8_.cby_0__1_.mux_right_ipin_2.sky130_fd_sc_hd__mux2_1_10_X
rlabel metal1 9292 36142 9292 36142 0 cby_0__8_.cby_0__1_.mux_right_ipin_2.sky130_fd_sc_hd__mux2_1_11_X
rlabel metal1 15548 10506 15548 10506 0 cby_0__8_.cby_0__1_.mux_right_ipin_2.sky130_fd_sc_hd__mux2_1_1_X
rlabel metal2 12742 12240 12742 12240 0 cby_0__8_.cby_0__1_.mux_right_ipin_2.sky130_fd_sc_hd__mux2_1_2_X
rlabel metal2 12558 12546 12558 12546 0 cby_0__8_.cby_0__1_.mux_right_ipin_2.sky130_fd_sc_hd__mux2_1_3_X
rlabel metal1 10718 16660 10718 16660 0 cby_0__8_.cby_0__1_.mux_right_ipin_2.sky130_fd_sc_hd__mux2_1_4_X
rlabel metal1 12328 14042 12328 14042 0 cby_0__8_.cby_0__1_.mux_right_ipin_2.sky130_fd_sc_hd__mux2_1_5_X
rlabel metal2 11730 15878 11730 15878 0 cby_0__8_.cby_0__1_.mux_right_ipin_2.sky130_fd_sc_hd__mux2_1_6_X
rlabel metal1 10350 16422 10350 16422 0 cby_0__8_.cby_0__1_.mux_right_ipin_2.sky130_fd_sc_hd__mux2_1_7_X
rlabel metal2 14674 22576 14674 22576 0 cby_0__8_.cby_0__1_.mux_right_ipin_2.sky130_fd_sc_hd__mux2_1_8_X
rlabel metal1 10350 17272 10350 17272 0 cby_0__8_.cby_0__1_.mux_right_ipin_2.sky130_fd_sc_hd__mux2_1_9_X
rlabel metal2 12466 16592 12466 16592 0 cby_0__8_.cby_0__1_.mux_right_ipin_3.sky130_fd_sc_hd__mux2_1_0_X
rlabel metal2 10350 27846 10350 27846 0 cby_0__8_.cby_0__1_.mux_right_ipin_3.sky130_fd_sc_hd__mux2_1_10_X
rlabel metal1 9568 39406 9568 39406 0 cby_0__8_.cby_0__1_.mux_right_ipin_3.sky130_fd_sc_hd__mux2_1_11_X
rlabel metal1 14030 12410 14030 12410 0 cby_0__8_.cby_0__1_.mux_right_ipin_3.sky130_fd_sc_hd__mux2_1_1_X
rlabel metal2 12190 14484 12190 14484 0 cby_0__8_.cby_0__1_.mux_right_ipin_3.sky130_fd_sc_hd__mux2_1_2_X
rlabel metal2 12098 14790 12098 14790 0 cby_0__8_.cby_0__1_.mux_right_ipin_3.sky130_fd_sc_hd__mux2_1_3_X
rlabel metal1 12972 18394 12972 18394 0 cby_0__8_.cby_0__1_.mux_right_ipin_3.sky130_fd_sc_hd__mux2_1_4_X
rlabel metal1 11822 16456 11822 16456 0 cby_0__8_.cby_0__1_.mux_right_ipin_3.sky130_fd_sc_hd__mux2_1_5_X
rlabel metal1 11684 17306 11684 17306 0 cby_0__8_.cby_0__1_.mux_right_ipin_3.sky130_fd_sc_hd__mux2_1_6_X
rlabel metal1 10258 19482 10258 19482 0 cby_0__8_.cby_0__1_.mux_right_ipin_3.sky130_fd_sc_hd__mux2_1_7_X
rlabel metal2 12742 25568 12742 25568 0 cby_0__8_.cby_0__1_.mux_right_ipin_3.sky130_fd_sc_hd__mux2_1_8_X
rlabel metal1 10120 21862 10120 21862 0 cby_0__8_.cby_0__1_.mux_right_ipin_3.sky130_fd_sc_hd__mux2_1_9_X
rlabel metal1 11546 40018 11546 40018 0 cby_0__8_.grid_io_left_left_0__1_.logical_tile_io_mode_io__0.ccff_tail
rlabel metal1 10488 46002 10488 46002 0 cby_0__8_.grid_io_left_left_0__1_.logical_tile_io_mode_io__0.gfpga_pad_io_soc_dir
rlabel metal1 15042 46002 15042 46002 0 cby_0__8_.grid_io_left_left_0__1_.logical_tile_io_mode_io__0.logical_tile_io_mode_physical__iopad_0.io_0_.SOC_DIR_N
rlabel metal2 9982 44132 9982 44132 0 cby_0__8_.grid_io_left_left_0__1_.logical_tile_io_mode_io__1.ccff_tail
rlabel metal1 10166 47158 10166 47158 0 cby_0__8_.grid_io_left_left_0__1_.logical_tile_io_mode_io__1.gfpga_pad_io_soc_dir
rlabel metal1 14490 46614 14490 46614 0 cby_0__8_.grid_io_left_left_0__1_.logical_tile_io_mode_io__1.logical_tile_io_mode_physical__iopad_0.io_0_.SOC_DIR_N
rlabel metal2 9154 47396 9154 47396 0 cby_0__8_.grid_io_left_left_0__1_.logical_tile_io_mode_io__2.ccff_tail
rlabel metal1 9706 49402 9706 49402 0 cby_0__8_.grid_io_left_left_0__1_.logical_tile_io_mode_io__2.gfpga_pad_io_soc_dir
rlabel metal2 14490 47464 14490 47464 0 cby_0__8_.grid_io_left_left_0__1_.logical_tile_io_mode_io__2.logical_tile_io_mode_physical__iopad_0.io_0_.SOC_DIR_N
rlabel metal1 5198 53040 5198 53040 0 cby_0__8_.grid_io_left_left_0__1_.logical_tile_io_mode_io__3.gfpga_pad_io_soc_dir
rlabel metal1 12604 47702 12604 47702 0 cby_0__8_.grid_io_left_left_0__1_.logical_tile_io_mode_io__3.logical_tile_io_mode_physical__iopad_0.io_0_.SOC_DIR_N
rlabel metal1 24702 53754 24702 53754 0 ccff_head
rlabel metal1 1656 4114 1656 4114 0 ccff_head_0
rlabel metal3 25630 748 25630 748 0 ccff_tail
rlabel metal1 1564 53618 1564 53618 0 ccff_tail_0
rlabel metal1 22632 29614 22632 29614 0 chanx_right_in[0]
rlabel metal1 24840 35462 24840 35462 0 chanx_right_in[10]
rlabel metal1 24840 36006 24840 36006 0 chanx_right_in[11]
rlabel metal1 25116 37230 25116 37230 0 chanx_right_in[12]
rlabel metal2 25162 36703 25162 36703 0 chanx_right_in[13]
rlabel metal2 25162 37655 25162 37655 0 chanx_right_in[14]
rlabel via2 25346 38301 25346 38301 0 chanx_right_in[15]
rlabel metal2 25346 39253 25346 39253 0 chanx_right_in[16]
rlabel metal1 25346 40052 25346 40052 0 chanx_right_in[17]
rlabel metal2 25346 40919 25346 40919 0 chanx_right_in[18]
rlabel via2 25162 41565 25162 41565 0 chanx_right_in[19]
rlabel metal2 17066 24412 17066 24412 0 chanx_right_in[1]
rlabel metal2 25162 42483 25162 42483 0 chanx_right_in[20]
rlabel metal2 25530 43401 25530 43401 0 chanx_right_in[21]
rlabel metal2 24794 44183 24794 44183 0 chanx_right_in[22]
rlabel via2 25346 44829 25346 44829 0 chanx_right_in[23]
rlabel metal2 25346 45781 25346 45781 0 chanx_right_in[24]
rlabel metal2 25346 46495 25346 46495 0 chanx_right_in[25]
rlabel metal2 25346 47447 25346 47447 0 chanx_right_in[26]
rlabel via2 25162 48093 25162 48093 0 chanx_right_in[27]
rlabel metal2 25162 49011 25162 49011 0 chanx_right_in[28]
rlabel metal2 25530 49929 25530 49929 0 chanx_right_in[29]
rlabel metal1 19044 23290 19044 23290 0 chanx_right_in[2]
rlabel metal1 19780 27506 19780 27506 0 chanx_right_in[3]
rlabel metal1 24702 29546 24702 29546 0 chanx_right_in[4]
rlabel metal1 25392 29138 25392 29138 0 chanx_right_in[5]
rlabel metal2 25346 30277 25346 30277 0 chanx_right_in[6]
rlabel metal1 25346 34544 25346 34544 0 chanx_right_in[7]
rlabel metal2 24610 33745 24610 33745 0 chanx_right_in[8]
rlabel metal2 24702 33983 24702 33983 0 chanx_right_in[9]
rlabel metal3 24112 1564 24112 1564 0 chanx_right_out[0]
rlabel metal2 23322 9673 23322 9673 0 chanx_right_out[10]
rlabel metal2 24702 10013 24702 10013 0 chanx_right_out[11]
rlabel metal2 24794 10965 24794 10965 0 chanx_right_out[12]
rlabel metal3 25676 12172 25676 12172 0 chanx_right_out[13]
rlabel metal3 25676 12988 25676 12988 0 chanx_right_out[14]
rlabel metal1 24104 13974 24104 13974 0 chanx_right_out[15]
rlabel metal2 25162 14297 25162 14297 0 chanx_right_out[16]
rlabel metal2 24794 15181 24794 15181 0 chanx_right_out[17]
rlabel metal3 25676 16252 25676 16252 0 chanx_right_out[18]
rlabel metal1 24104 17238 24104 17238 0 chanx_right_out[19]
rlabel metal1 17342 2414 17342 2414 0 chanx_right_out[1]
rlabel metal1 24380 17714 24380 17714 0 chanx_right_out[20]
rlabel metal2 24794 17901 24794 17901 0 chanx_right_out[21]
rlabel metal1 23460 18802 23460 18802 0 chanx_right_out[22]
rlabel via2 23230 20349 23230 20349 0 chanx_right_out[23]
rlabel metal1 21689 21454 21689 21454 0 chanx_right_out[24]
rlabel metal1 24380 20978 24380 20978 0 chanx_right_out[25]
rlabel metal1 24104 22678 24104 22678 0 chanx_right_out[26]
rlabel metal2 23782 23375 23782 23375 0 chanx_right_out[27]
rlabel metal2 24794 23477 24794 23477 0 chanx_right_out[28]
rlabel metal3 25676 25228 25676 25228 0 chanx_right_out[29]
rlabel metal2 18998 5032 18998 5032 0 chanx_right_out[2]
rlabel metal2 22034 7055 22034 7055 0 chanx_right_out[3]
rlabel metal2 21942 6205 21942 6205 0 chanx_right_out[4]
rlabel metal2 23322 6477 23322 6477 0 chanx_right_out[5]
rlabel metal2 24794 5797 24794 5797 0 chanx_right_out[6]
rlabel metal2 24702 6749 24702 6749 0 chanx_right_out[7]
rlabel metal2 25162 7769 25162 7769 0 chanx_right_out[8]
rlabel metal3 25676 8908 25676 8908 0 chanx_right_out[9]
rlabel metal1 2162 4114 2162 4114 0 chany_bottom_in_0[0]
rlabel metal1 5842 1734 5842 1734 0 chany_bottom_in_0[10]
rlabel metal1 4738 2380 4738 2380 0 chany_bottom_in_0[11]
rlabel metal1 6348 3502 6348 3502 0 chany_bottom_in_0[12]
rlabel metal1 6716 4114 6716 4114 0 chany_bottom_in_0[13]
rlabel metal1 7176 3502 7176 3502 0 chany_bottom_in_0[14]
rlabel metal2 7406 3468 7406 3468 0 chany_bottom_in_0[15]
rlabel metal1 7820 3026 7820 3026 0 chany_bottom_in_0[16]
rlabel metal1 7590 2414 7590 2414 0 chany_bottom_in_0[17]
rlabel metal1 8280 3502 8280 3502 0 chany_bottom_in_0[18]
rlabel metal1 6716 2618 6716 2618 0 chany_bottom_in_0[19]
rlabel metal2 2254 2132 2254 2132 0 chany_bottom_in_0[1]
rlabel metal1 9384 4114 9384 4114 0 chany_bottom_in_0[20]
rlabel metal1 9338 3536 9338 3536 0 chany_bottom_in_0[21]
rlabel metal1 9936 4590 9936 4590 0 chany_bottom_in_0[22]
rlabel metal1 9798 2278 9798 2278 0 chany_bottom_in_0[23]
rlabel metal1 9476 3026 9476 3026 0 chany_bottom_in_0[24]
rlabel metal1 10028 2346 10028 2346 0 chany_bottom_in_0[25]
rlabel metal2 11454 1761 11454 1761 0 chany_bottom_in_0[26]
rlabel via1 11178 3028 11178 3028 0 chany_bottom_in_0[27]
rlabel metal1 10672 3026 10672 3026 0 chany_bottom_in_0[28]
rlabel metal2 12558 1588 12558 1588 0 chany_bottom_in_0[29]
rlabel metal1 2392 3026 2392 3026 0 chany_bottom_in_0[2]
rlabel metal1 2691 2414 2691 2414 0 chany_bottom_in_0[3]
rlabel metal1 3404 3026 3404 3026 0 chany_bottom_in_0[4]
rlabel metal1 1886 3502 1886 3502 0 chany_bottom_in_0[5]
rlabel metal1 4232 4114 4232 4114 0 chany_bottom_in_0[6]
rlabel metal1 4508 3162 4508 3162 0 chany_bottom_in_0[7]
rlabel metal2 4830 1761 4830 1761 0 chany_bottom_in_0[8]
rlabel metal1 5796 2278 5796 2278 0 chany_bottom_in_0[9]
rlabel metal2 12926 1418 12926 1418 0 chany_bottom_out_0[0]
rlabel metal1 17066 3094 17066 3094 0 chany_bottom_out_0[10]
rlabel metal1 18446 2822 18446 2822 0 chany_bottom_out_0[11]
rlabel metal2 17342 1503 17342 1503 0 chany_bottom_out_0[12]
rlabel metal1 18814 3570 18814 3570 0 chany_bottom_out_0[13]
rlabel metal2 18078 823 18078 823 0 chany_bottom_out_0[14]
rlabel metal2 18446 891 18446 891 0 chany_bottom_out_0[15]
rlabel metal1 19366 4658 19366 4658 0 chany_bottom_out_0[16]
rlabel metal1 20470 3434 20470 3434 0 chany_bottom_out_0[17]
rlabel metal1 20654 3706 20654 3706 0 chany_bottom_out_0[18]
rlabel metal2 19918 1418 19918 1418 0 chany_bottom_out_0[19]
rlabel metal2 13294 1554 13294 1554 0 chany_bottom_out_0[1]
rlabel metal1 20562 5746 20562 5746 0 chany_bottom_out_0[20]
rlabel metal2 20654 1761 20654 1761 0 chany_bottom_out_0[21]
rlabel metal2 21022 1418 21022 1418 0 chany_bottom_out_0[22]
rlabel metal2 21390 1792 21390 1792 0 chany_bottom_out_0[23]
rlabel metal2 21758 1860 21758 1860 0 chany_bottom_out_0[24]
rlabel metal2 22126 823 22126 823 0 chany_bottom_out_0[25]
rlabel metal2 22494 840 22494 840 0 chany_bottom_out_0[26]
rlabel metal1 21850 3604 21850 3604 0 chany_bottom_out_0[27]
rlabel metal2 23230 1163 23230 1163 0 chany_bottom_out_0[28]
rlabel metal1 22954 7752 22954 7752 0 chany_bottom_out_0[29]
rlabel metal2 13662 1860 13662 1860 0 chany_bottom_out_0[2]
rlabel metal1 14398 3570 14398 3570 0 chany_bottom_out_0[3]
rlabel metal2 14398 1554 14398 1554 0 chany_bottom_out_0[4]
rlabel metal1 15042 2958 15042 2958 0 chany_bottom_out_0[5]
rlabel metal1 16238 2890 16238 2890 0 chany_bottom_out_0[6]
rlabel metal1 16054 3570 16054 3570 0 chany_bottom_out_0[7]
rlabel metal1 16652 2958 16652 2958 0 chany_bottom_out_0[8]
rlabel metal1 16790 4046 16790 4046 0 chany_bottom_out_0[9]
rlabel metal2 22126 32300 22126 32300 0 clknet_0_prog_clk
rlabel metal2 9982 14960 9982 14960 0 clknet_4_0_0_prog_clk
rlabel metal1 9430 36618 9430 36618 0 clknet_4_10_0_prog_clk
rlabel metal1 18768 33966 18768 33966 0 clknet_4_11_0_prog_clk
rlabel metal2 19918 20094 19918 20094 0 clknet_4_12_0_prog_clk
rlabel metal2 20470 27132 20470 27132 0 clknet_4_13_0_prog_clk
rlabel metal2 19458 32674 19458 32674 0 clknet_4_14_0_prog_clk
rlabel metal1 19964 44846 19964 44846 0 clknet_4_15_0_prog_clk
rlabel metal1 13202 13362 13202 13362 0 clknet_4_1_0_prog_clk
rlabel metal1 9292 18190 9292 18190 0 clknet_4_2_0_prog_clk
rlabel metal1 12742 20366 12742 20366 0 clknet_4_3_0_prog_clk
rlabel metal2 19734 10948 19734 10948 0 clknet_4_4_0_prog_clk
rlabel metal1 20102 13838 20102 13838 0 clknet_4_5_0_prog_clk
rlabel metal1 15686 21114 15686 21114 0 clknet_4_6_0_prog_clk
rlabel metal1 17848 15538 17848 15538 0 clknet_4_7_0_prog_clk
rlabel metal1 13294 31790 13294 31790 0 clknet_4_8_0_prog_clk
rlabel metal2 12558 28798 12558 28798 0 clknet_4_9_0_prog_clk
rlabel metal1 2484 54094 2484 54094 0 gfpga_pad_io_soc_dir[0]
rlabel metal2 4002 56236 4002 56236 0 gfpga_pad_io_soc_dir[1]
rlabel metal1 5474 53618 5474 53618 0 gfpga_pad_io_soc_dir[2]
rlabel metal2 6762 56236 6762 56236 0 gfpga_pad_io_soc_dir[3]
rlabel metal1 13616 54162 13616 54162 0 gfpga_pad_io_soc_in[0]
rlabel metal1 14996 54162 14996 54162 0 gfpga_pad_io_soc_in[1]
rlabel metal1 16836 54162 16836 54162 0 gfpga_pad_io_soc_in[2]
rlabel metal1 17756 54162 17756 54162 0 gfpga_pad_io_soc_in[3]
rlabel metal2 7958 55711 7958 55711 0 gfpga_pad_io_soc_out[0]
rlabel metal2 9338 51894 9338 51894 0 gfpga_pad_io_soc_out[1]
rlabel metal2 10902 56236 10902 56236 0 gfpga_pad_io_soc_out[2]
rlabel metal2 12098 51112 12098 51112 0 gfpga_pad_io_soc_out[3]
rlabel metal1 19228 54094 19228 54094 0 isol_n
rlabel metal1 21942 53958 21942 53958 0 net1
rlabel metal2 22034 35564 22034 35564 0 net10
rlabel metal1 20493 25330 20493 25330 0 net100
rlabel metal2 15042 4964 15042 4964 0 net101
rlabel metal1 13340 4658 13340 4658 0 net102
rlabel metal1 19458 7378 19458 7378 0 net103
rlabel metal2 15134 7922 15134 7922 0 net104
rlabel metal1 23828 5202 23828 5202 0 net105
rlabel metal2 23966 6086 23966 6086 0 net106
rlabel metal2 11914 5491 11914 5491 0 net107
rlabel metal2 10626 5151 10626 5151 0 net108
rlabel via3 20125 12580 20125 12580 0 net109
rlabel metal1 25116 40154 25116 40154 0 net11
rlabel metal1 19090 3026 19090 3026 0 net110
rlabel metal1 20056 12138 20056 12138 0 net111
rlabel metal1 18400 4590 18400 4590 0 net112
rlabel metal1 20240 3502 20240 3502 0 net113
rlabel metal1 18630 4114 18630 4114 0 net114
rlabel metal2 22034 2176 22034 2176 0 net115
rlabel metal1 20102 4590 20102 4590 0 net116
rlabel metal1 21160 3502 21160 3502 0 net117
rlabel via3 21413 18020 21413 18020 0 net118
rlabel via3 22149 17068 22149 17068 0 net119
rlabel metal1 25208 40902 25208 40902 0 net12
rlabel metal1 15226 2278 15226 2278 0 net120
rlabel metal2 20930 4114 20930 4114 0 net121
rlabel metal1 22034 5168 22034 5168 0 net122
rlabel metal1 20838 7752 20838 7752 0 net123
rlabel metal1 21114 3026 21114 3026 0 net124
rlabel metal1 22218 6324 22218 6324 0 net125
rlabel metal2 22218 5508 22218 5508 0 net126
rlabel metal1 17204 4998 17204 4998 0 net127
rlabel metal2 20378 4641 20378 4641 0 net128
rlabel metal1 20838 2074 20838 2074 0 net129
rlabel metal1 25622 41514 25622 41514 0 net13
rlabel metal1 21206 7854 21206 7854 0 net130
rlabel metal3 15111 16660 15111 16660 0 net131
rlabel via3 17365 15300 17365 15300 0 net132
rlabel metal2 14490 3434 14490 3434 0 net133
rlabel metal1 14720 3026 14720 3026 0 net134
rlabel metal2 17066 5882 17066 5882 0 net135
rlabel metal1 18262 10438 18262 10438 0 net136
rlabel metal1 19504 13158 19504 13158 0 net137
rlabel metal1 17756 4114 17756 4114 0 net138
rlabel metal1 4462 53210 4462 53210 0 net139
rlabel metal1 20286 22678 20286 22678 0 net14
rlabel metal2 6578 53686 6578 53686 0 net140
rlabel metal2 7682 53108 7682 53108 0 net141
rlabel metal2 6762 53142 6762 53142 0 net142
rlabel metal1 18308 26010 18308 26010 0 net143
rlabel metal1 18262 27506 18262 27506 0 net144
rlabel metal1 18952 16150 18952 16150 0 net145
rlabel metal2 19826 28798 19826 28798 0 net146
rlabel metal2 23690 28458 23690 28458 0 net147
rlabel metal1 24932 28458 24932 28458 0 net148
rlabel metal1 21850 30226 21850 30226 0 net149
rlabel metal1 25760 42602 25760 42602 0 net15
rlabel metal1 19780 30226 19780 30226 0 net150
rlabel metal1 19550 29274 19550 29274 0 net151
rlabel metal2 22586 19074 22586 19074 0 net152
rlabel metal1 20194 17306 20194 17306 0 net153
rlabel metal1 19642 23630 19642 23630 0 net154
rlabel metal2 22586 17153 22586 17153 0 net155
rlabel metal1 7958 17306 7958 17306 0 net156
rlabel metal1 6992 12954 6992 12954 0 net157
rlabel metal1 8694 12206 8694 12206 0 net158
rlabel metal1 14536 17714 14536 17714 0 net159
rlabel metal1 25484 43146 25484 43146 0 net16
rlabel metal1 13616 17306 13616 17306 0 net160
rlabel metal2 15318 15810 15318 15810 0 net161
rlabel metal1 9798 20910 9798 20910 0 net162
rlabel metal1 11822 8942 11822 8942 0 net163
rlabel metal1 12098 7854 12098 7854 0 net164
rlabel metal2 13386 8670 13386 8670 0 net165
rlabel metal1 16698 13294 16698 13294 0 net166
rlabel metal1 14168 15130 14168 15130 0 net167
rlabel metal2 15686 17034 15686 17034 0 net168
rlabel metal1 15456 14994 15456 14994 0 net169
rlabel metal1 25576 44234 25576 44234 0 net17
rlabel metal1 13892 7378 13892 7378 0 net170
rlabel metal1 17342 6426 17342 6426 0 net171
rlabel metal1 16330 2482 16330 2482 0 net172
rlabel metal2 13386 21454 13386 21454 0 net173
rlabel metal2 21298 5168 21298 5168 0 net174
rlabel metal1 16054 13226 16054 13226 0 net175
rlabel metal1 10994 10982 10994 10982 0 net176
rlabel metal2 19090 12619 19090 12619 0 net177
rlabel metal1 18078 11798 18078 11798 0 net178
rlabel metal2 13570 4794 13570 4794 0 net179
rlabel metal1 24334 44710 24334 44710 0 net18
rlabel metal1 24610 5882 24610 5882 0 net180
rlabel metal1 16238 2380 16238 2380 0 net181
rlabel metal1 16652 13974 16652 13974 0 net182
rlabel metal1 11362 8602 11362 8602 0 net183
rlabel metal2 11730 18496 11730 18496 0 net184
rlabel metal2 9522 17952 9522 17952 0 net185
rlabel metal1 11270 13906 11270 13906 0 net186
rlabel metal1 11592 10778 11592 10778 0 net187
rlabel metal1 15456 23698 15456 23698 0 net188
rlabel metal1 15916 26010 15916 26010 0 net189
rlabel metal1 23368 38522 23368 38522 0 net19
rlabel metal1 19642 22610 19642 22610 0 net190
rlabel metal1 20010 22542 20010 22542 0 net191
rlabel metal1 20010 21998 20010 21998 0 net192
rlabel metal1 20884 22066 20884 22066 0 net193
rlabel metal1 18722 24174 18722 24174 0 net194
rlabel metal2 23598 30464 23598 30464 0 net195
rlabel metal2 18814 19924 18814 19924 0 net196
rlabel metal1 16560 15402 16560 15402 0 net197
rlabel metal2 20654 12002 20654 12002 0 net198
rlabel metal1 20516 28594 20516 28594 0 net199
rlabel metal2 5382 4250 5382 4250 0 net2
rlabel metal1 24242 46342 24242 46342 0 net20
rlabel metal2 22218 24616 22218 24616 0 net200
rlabel metal1 14950 28186 14950 28186 0 net201
rlabel metal1 22540 18394 22540 18394 0 net202
rlabel metal1 20010 32946 20010 32946 0 net203
rlabel metal2 8878 8670 8878 8670 0 net204
rlabel metal1 19918 31858 19918 31858 0 net205
rlabel metal1 25392 18938 25392 18938 0 net206
rlabel metal1 13984 3978 13984 3978 0 net207
rlabel metal2 22678 26656 22678 26656 0 net208
rlabel metal1 13432 6358 13432 6358 0 net209
rlabel metal1 25576 47430 25576 47430 0 net21
rlabel metal2 21206 28322 21206 28322 0 net210
rlabel metal1 20148 26010 20148 26010 0 net211
rlabel metal1 13202 25466 13202 25466 0 net212
rlabel metal1 14720 22202 14720 22202 0 net213
rlabel metal1 17434 31450 17434 31450 0 net214
rlabel metal1 9890 33626 9890 33626 0 net215
rlabel metal2 17434 29852 17434 29852 0 net216
rlabel metal1 11776 6426 11776 6426 0 net217
rlabel metal1 10212 13226 10212 13226 0 net218
rlabel metal1 11914 20570 11914 20570 0 net219
rlabel metal1 21436 47974 21436 47974 0 net22
rlabel metal2 15502 21148 15502 21148 0 net220
rlabel metal1 9062 48246 9062 48246 0 net221
rlabel metal1 11132 23290 11132 23290 0 net222
rlabel metal1 15916 16218 15916 16218 0 net223
rlabel metal1 9890 46478 9890 46478 0 net224
rlabel metal1 24564 32334 24564 32334 0 net225
rlabel metal1 19320 30634 19320 30634 0 net226
rlabel metal2 19734 34408 19734 34408 0 net227
rlabel metal1 13846 30158 13846 30158 0 net228
rlabel metal2 20010 16286 20010 16286 0 net229
rlabel metal1 22126 47226 22126 47226 0 net23
rlabel metal2 20010 24990 20010 24990 0 net230
rlabel metal2 17434 8364 17434 8364 0 net231
rlabel metal1 23046 33422 23046 33422 0 net232
rlabel metal2 18630 4420 18630 4420 0 net233
rlabel metal1 18446 9146 18446 9146 0 net234
rlabel metal2 14030 5406 14030 5406 0 net235
rlabel metal1 22908 22950 22908 22950 0 net236
rlabel metal1 13662 19278 13662 19278 0 net237
rlabel metal1 23920 10098 23920 10098 0 net238
rlabel metal2 25254 17918 25254 17918 0 net239
rlabel metal1 22862 49742 22862 49742 0 net24
rlabel metal2 21574 33966 21574 33966 0 net240
rlabel metal1 11822 27506 11822 27506 0 net241
rlabel metal2 9338 7582 9338 7582 0 net242
rlabel metal1 12098 28186 12098 28186 0 net243
rlabel metal2 25254 26180 25254 26180 0 net244
rlabel metal1 23414 31790 23414 31790 0 net245
rlabel metal1 23775 6970 23775 6970 0 net246
rlabel metal1 23184 30906 23184 30906 0 net247
rlabel metal2 12374 41684 12374 41684 0 net248
rlabel metal1 23920 15538 23920 15538 0 net249
rlabel metal2 21114 23834 21114 23834 0 net25
rlabel metal1 25116 16218 25116 16218 0 net250
rlabel metal2 21850 21250 21850 21250 0 net251
rlabel metal2 13570 8840 13570 8840 0 net252
rlabel metal1 19320 16218 19320 16218 0 net253
rlabel metal2 17710 32606 17710 32606 0 net254
rlabel metal1 25300 20026 25300 20026 0 net255
rlabel metal2 8602 14756 8602 14756 0 net256
rlabel metal1 23506 23800 23506 23800 0 net257
rlabel metal1 22678 25942 22678 25942 0 net258
rlabel metal1 15456 5882 15456 5882 0 net259
rlabel metal2 21022 26826 21022 26826 0 net26
rlabel metal2 23322 13022 23322 13022 0 net260
rlabel metal1 20792 18870 20792 18870 0 net261
rlabel metal2 10258 5916 10258 5916 0 net262
rlabel metal2 22678 8670 22678 8670 0 net263
rlabel metal2 25254 27744 25254 27744 0 net264
rlabel metal2 8602 21284 8602 21284 0 net265
rlabel metal2 13478 16762 13478 16762 0 net266
rlabel metal1 18676 28186 18676 28186 0 net267
rlabel metal1 12949 24106 12949 24106 0 net268
rlabel metal1 24288 33898 24288 33898 0 net269
rlabel metal1 23138 26010 23138 26010 0 net27
rlabel metal2 9430 10846 9430 10846 0 net270
rlabel metal2 8510 22814 8510 22814 0 net271
rlabel metal1 15633 8058 15633 8058 0 net272
rlabel metal2 23782 5984 23782 5984 0 net273
rlabel metal2 20102 10404 20102 10404 0 net274
rlabel metal1 14529 13702 14529 13702 0 net275
rlabel metal1 23920 31994 23920 31994 0 net276
rlabel metal1 7176 18802 7176 18802 0 net277
rlabel metal1 6762 15130 6762 15130 0 net278
rlabel metal2 23414 11934 23414 11934 0 net279
rlabel metal1 24242 26350 24242 26350 0 net28
rlabel metal1 24334 7786 24334 7786 0 net280
rlabel metal1 20010 5304 20010 5304 0 net281
rlabel metal2 12742 20910 12742 20910 0 net282
rlabel metal1 14812 18394 14812 18394 0 net283
rlabel metal2 7866 16558 7866 16558 0 net284
rlabel metal1 8878 23800 8878 23800 0 net285
rlabel metal1 11592 24854 11592 24854 0 net286
rlabel metal2 22586 14620 22586 14620 0 net287
rlabel metal1 10488 28186 10488 28186 0 net288
rlabel metal2 19734 23970 19734 23970 0 net289
rlabel metal2 25070 27948 25070 27948 0 net29
rlabel metal1 8602 12716 8602 12716 0 net290
rlabel metal1 9476 26418 9476 26418 0 net291
rlabel metal1 17158 18360 17158 18360 0 net292
rlabel metal2 12466 28764 12466 28764 0 net293
rlabel metal1 13524 26894 13524 26894 0 net294
rlabel metal1 18308 13158 18308 13158 0 net295
rlabel metal1 17572 38182 17572 38182 0 net296
rlabel via2 20930 12971 20930 12971 0 net3
rlabel metal1 24932 28186 24932 28186 0 net30
rlabel metal1 24656 35190 24656 35190 0 net31
rlabel metal1 24104 34714 24104 34714 0 net32
rlabel metal2 2254 5032 2254 5032 0 net33
rlabel metal1 13202 14858 13202 14858 0 net34
rlabel metal1 13248 12818 13248 12818 0 net35
rlabel metal2 6394 3774 6394 3774 0 net36
rlabel metal1 6900 3978 6900 3978 0 net37
rlabel metal1 14398 12818 14398 12818 0 net38
rlabel metal1 14352 14994 14352 14994 0 net39
rlabel metal1 24012 35802 24012 35802 0 net4
rlabel metal1 14628 12682 14628 12682 0 net40
rlabel via2 16054 14229 16054 14229 0 net41
rlabel metal1 8510 3366 8510 3366 0 net42
rlabel metal2 13386 4998 13386 4998 0 net43
rlabel metal1 5566 17510 5566 17510 0 net44
rlabel metal1 14076 7514 14076 7514 0 net45
rlabel metal1 12926 10030 12926 10030 0 net46
rlabel metal1 15686 9622 15686 9622 0 net47
rlabel via2 8234 2533 8234 2533 0 net48
rlabel metal1 15640 9554 15640 9554 0 net49
rlabel metal1 25346 36006 25346 36006 0 net5
rlabel metal2 19090 11526 19090 11526 0 net50
rlabel metal2 20562 13328 20562 13328 0 net51
rlabel metal1 16974 9894 16974 9894 0 net52
rlabel metal1 14720 8534 14720 8534 0 net53
rlabel metal1 14030 2346 14030 2346 0 net54
rlabel metal1 10442 19346 10442 19346 0 net55
rlabel metal1 12742 22066 12742 22066 0 net56
rlabel metal1 11408 18666 11408 18666 0 net57
rlabel metal2 8878 15725 8878 15725 0 net58
rlabel metal1 6854 13226 6854 13226 0 net59
rlabel metal1 25438 37094 25438 37094 0 net6
rlabel metal1 5612 3706 5612 3706 0 net60
rlabel metal2 5198 10812 5198 10812 0 net61
rlabel metal1 12972 16626 12972 16626 0 net62
rlabel metal2 12650 50796 12650 50796 0 net63
rlabel metal1 14628 47090 14628 47090 0 net64
rlabel metal2 15502 50218 15502 50218 0 net65
rlabel metal2 17158 49912 17158 49912 0 net66
rlabel metal1 18170 54128 18170 54128 0 net67
rlabel metal1 21896 44914 21896 44914 0 net68
rlabel metal2 25070 50592 25070 50592 0 net69
rlabel metal1 26036 36618 26036 36618 0 net7
rlabel metal1 23230 51238 23230 51238 0 net70
rlabel metal1 25944 52462 25944 52462 0 net71
rlabel metal1 26174 32946 26174 32946 0 net72
rlabel metal1 26036 53958 26036 53958 0 net73
rlabel metal1 22218 32334 22218 32334 0 net74
rlabel metal1 21390 54026 21390 54026 0 net75
rlabel metal1 20424 41446 20424 41446 0 net76
rlabel metal1 14030 2618 14030 2618 0 net77
rlabel metal1 1794 53516 1794 53516 0 net78
rlabel metal1 21551 8942 21551 8942 0 net79
rlabel metal1 25990 37706 25990 37706 0 net8
rlabel metal2 21942 7463 21942 7463 0 net80
rlabel metal2 8418 9945 8418 9945 0 net81
rlabel metal2 10902 10897 10902 10897 0 net82
rlabel metal2 19826 14688 19826 14688 0 net83
rlabel metal1 23322 13294 23322 13294 0 net84
rlabel metal2 19458 14110 19458 14110 0 net85
rlabel metal2 19826 14178 19826 14178 0 net86
rlabel metal2 21482 13974 21482 13974 0 net87
rlabel metal1 23046 10778 23046 10778 0 net88
rlabel metal2 22310 14569 22310 14569 0 net89
rlabel metal1 22862 38182 22862 38182 0 net9
rlabel metal1 14122 4998 14122 4998 0 net90
rlabel metal2 22678 16116 22678 16116 0 net91
rlabel metal2 20838 17952 20838 17952 0 net92
rlabel metal2 14398 16864 14398 16864 0 net93
rlabel metal1 19734 20434 19734 20434 0 net94
rlabel metal2 22034 21318 22034 21318 0 net95
rlabel metal1 21758 23222 21758 23222 0 net96
rlabel metal1 18837 21114 18837 21114 0 net97
rlabel metal2 23874 22644 23874 22644 0 net98
rlabel metal1 23184 22610 23184 22610 0 net99
rlabel via2 19366 25109 19366 25109 0 prog_clk
rlabel metal1 25116 2618 25116 2618 0 prog_reset
rlabel metal2 24978 50711 24978 50711 0 right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_
rlabel metal2 25530 51561 25530 51561 0 right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_
rlabel metal2 24978 52275 24978 52275 0 right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_
rlabel metal2 25070 53023 25070 53023 0 right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_
rlabel metal2 24794 53975 24794 53975 0 right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_4_
rlabel metal2 24702 54077 24702 54077 0 right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_5_
rlabel metal3 25446 55420 25446 55420 0 right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_6_
rlabel via2 23437 56100 23437 56100 0 right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_7_
rlabel metal1 18676 52462 18676 52462 0 right_top_grid_bottom_width_0_height_0_subtile_0__pin_inpad_0_
rlabel metal2 21758 43981 21758 43981 0 right_top_grid_bottom_width_0_height_0_subtile_1__pin_inpad_0_
rlabel metal2 22908 56236 22908 56236 0 right_top_grid_bottom_width_0_height_0_subtile_2__pin_inpad_0_
rlabel metal2 24472 55692 24472 55692 0 right_top_grid_bottom_width_0_height_0_subtile_3__pin_inpad_0_
rlabel metal1 22770 35054 22770 35054 0 right_width_0_height_0_subtile_0__pin_inpad_0_
rlabel metal1 16330 15640 16330 15640 0 right_width_0_height_0_subtile_1__pin_inpad_0_
rlabel metal1 24932 35258 24932 35258 0 right_width_0_height_0_subtile_2__pin_inpad_0_
rlabel metal1 24518 33626 24518 33626 0 right_width_0_height_0_subtile_3__pin_inpad_0_
rlabel metal2 18630 15062 18630 15062 0 sb_0__8_.mem_bottom_track_1.ccff_head
rlabel metal1 21850 19686 21850 19686 0 sb_0__8_.mem_bottom_track_1.ccff_tail
rlabel metal1 20976 18734 20976 18734 0 sb_0__8_.mem_bottom_track_1.mem_out\[0\]
rlabel metal1 22816 21454 22816 21454 0 sb_0__8_.mem_bottom_track_11.ccff_head
rlabel metal2 20838 25398 20838 25398 0 sb_0__8_.mem_bottom_track_11.ccff_tail
rlabel metal1 24886 19822 24886 19822 0 sb_0__8_.mem_bottom_track_11.mem_out\[0\]
rlabel metal1 24334 26758 24334 26758 0 sb_0__8_.mem_bottom_track_13.ccff_tail
rlabel metal1 25070 26010 25070 26010 0 sb_0__8_.mem_bottom_track_13.mem_out\[0\]
rlabel metal1 21436 27302 21436 27302 0 sb_0__8_.mem_bottom_track_15.ccff_tail
rlabel metal2 22678 28322 22678 28322 0 sb_0__8_.mem_bottom_track_15.mem_out\[0\]
rlabel metal1 19504 26826 19504 26826 0 sb_0__8_.mem_bottom_track_17.ccff_tail
rlabel metal1 20976 26418 20976 26418 0 sb_0__8_.mem_bottom_track_17.mem_out\[0\]
rlabel metal2 18906 27948 18906 27948 0 sb_0__8_.mem_bottom_track_19.ccff_tail
rlabel metal1 18860 28730 18860 28730 0 sb_0__8_.mem_bottom_track_19.mem_out\[0\]
rlabel metal2 18630 32436 18630 32436 0 sb_0__8_.mem_bottom_track_29.ccff_tail
rlabel metal1 18676 30906 18676 30906 0 sb_0__8_.mem_bottom_track_29.mem_out\[0\]
rlabel metal2 25162 18428 25162 18428 0 sb_0__8_.mem_bottom_track_3.ccff_tail
rlabel metal1 23920 19686 23920 19686 0 sb_0__8_.mem_bottom_track_3.mem_out\[0\]
rlabel metal1 20102 28662 20102 28662 0 sb_0__8_.mem_bottom_track_31.ccff_tail
rlabel metal1 22218 31892 22218 31892 0 sb_0__8_.mem_bottom_track_31.mem_out\[0\]
rlabel metal1 24288 30702 24288 30702 0 sb_0__8_.mem_bottom_track_33.ccff_tail
rlabel metal1 24564 32878 24564 32878 0 sb_0__8_.mem_bottom_track_33.mem_out\[0\]
rlabel metal1 24932 31790 24932 31790 0 sb_0__8_.mem_bottom_track_35.ccff_tail
rlabel metal1 24748 31314 24748 31314 0 sb_0__8_.mem_bottom_track_35.mem_out\[0\]
rlabel metal1 23644 33286 23644 33286 0 sb_0__8_.mem_bottom_track_45.ccff_tail
rlabel metal1 23230 34578 23230 34578 0 sb_0__8_.mem_bottom_track_45.mem_out\[0\]
rlabel metal1 20424 33626 20424 33626 0 sb_0__8_.mem_bottom_track_47.ccff_tail
rlabel metal2 22126 34374 22126 34374 0 sb_0__8_.mem_bottom_track_47.mem_out\[0\]
rlabel metal1 20378 32742 20378 32742 0 sb_0__8_.mem_bottom_track_49.ccff_tail
rlabel metal1 21068 34578 21068 34578 0 sb_0__8_.mem_bottom_track_49.mem_out\[0\]
rlabel metal1 22632 20434 22632 20434 0 sb_0__8_.mem_bottom_track_5.ccff_tail
rlabel metal1 25300 20570 25300 20570 0 sb_0__8_.mem_bottom_track_5.mem_out\[0\]
rlabel metal1 22494 28390 22494 28390 0 sb_0__8_.mem_bottom_track_51.mem_out\[0\]
rlabel metal1 20470 24378 20470 24378 0 sb_0__8_.mem_bottom_track_7.ccff_tail
rlabel metal1 21482 23698 21482 23698 0 sb_0__8_.mem_bottom_track_7.mem_out\[0\]
rlabel metal2 21574 25840 21574 25840 0 sb_0__8_.mem_bottom_track_9.mem_out\[0\]
rlabel metal2 12098 26384 12098 26384 0 sb_0__8_.mem_right_track_0.ccff_tail
rlabel metal2 22218 41514 22218 41514 0 sb_0__8_.mem_right_track_0.mem_out\[0\]
rlabel metal1 13754 29070 13754 29070 0 sb_0__8_.mem_right_track_0.mem_out\[1\]
rlabel metal2 10626 22882 10626 22882 0 sb_0__8_.mem_right_track_10.ccff_head
rlabel metal1 8234 19686 8234 19686 0 sb_0__8_.mem_right_track_10.ccff_tail
rlabel metal1 13938 25330 13938 25330 0 sb_0__8_.mem_right_track_10.mem_out\[0\]
rlabel metal1 6854 19754 6854 19754 0 sb_0__8_.mem_right_track_10.mem_out\[1\]
rlabel metal2 11730 20162 11730 20162 0 sb_0__8_.mem_right_track_12.ccff_tail
rlabel metal1 8556 18598 8556 18598 0 sb_0__8_.mem_right_track_12.mem_out\[0\]
rlabel metal1 15272 21522 15272 21522 0 sb_0__8_.mem_right_track_14.ccff_tail
rlabel metal1 13846 20774 13846 20774 0 sb_0__8_.mem_right_track_14.mem_out\[0\]
rlabel metal1 15088 20366 15088 20366 0 sb_0__8_.mem_right_track_16.ccff_tail
rlabel metal2 12788 21522 12788 21522 0 sb_0__8_.mem_right_track_16.mem_out\[0\]
rlabel metal2 13478 15436 13478 15436 0 sb_0__8_.mem_right_track_18.ccff_tail
rlabel metal2 12834 18564 12834 18564 0 sb_0__8_.mem_right_track_18.mem_out\[0\]
rlabel metal2 11178 26588 11178 26588 0 sb_0__8_.mem_right_track_2.ccff_tail
rlabel metal1 14352 28594 14352 28594 0 sb_0__8_.mem_right_track_2.mem_out\[0\]
rlabel metal1 13754 27948 13754 27948 0 sb_0__8_.mem_right_track_2.mem_out\[1\]
rlabel metal1 10672 9894 10672 9894 0 sb_0__8_.mem_right_track_20.ccff_tail
rlabel metal1 11316 13158 11316 13158 0 sb_0__8_.mem_right_track_20.mem_out\[0\]
rlabel metal1 10856 7514 10856 7514 0 sb_0__8_.mem_right_track_22.ccff_tail
rlabel via1 10350 8058 10350 8058 0 sb_0__8_.mem_right_track_22.mem_out\[0\]
rlabel metal1 12880 8466 12880 8466 0 sb_0__8_.mem_right_track_24.ccff_tail
rlabel metal1 12006 6290 12006 6290 0 sb_0__8_.mem_right_track_24.mem_out\[0\]
rlabel metal1 15594 13838 15594 13838 0 sb_0__8_.mem_right_track_26.ccff_tail
rlabel metal1 14950 12750 14950 12750 0 sb_0__8_.mem_right_track_26.mem_out\[0\]
rlabel metal1 16330 19890 16330 19890 0 sb_0__8_.mem_right_track_28.ccff_tail
rlabel metal1 14398 18292 14398 18292 0 sb_0__8_.mem_right_track_28.mem_out\[0\]
rlabel metal1 18078 19924 18078 19924 0 sb_0__8_.mem_right_track_30.ccff_tail
rlabel metal1 16238 16626 16238 16626 0 sb_0__8_.mem_right_track_30.mem_out\[0\]
rlabel metal2 18630 17884 18630 17884 0 sb_0__8_.mem_right_track_32.ccff_tail
rlabel metal1 19090 18734 19090 18734 0 sb_0__8_.mem_right_track_32.mem_out\[0\]
rlabel metal1 16928 11322 16928 11322 0 sb_0__8_.mem_right_track_34.ccff_tail
rlabel metal1 17894 15674 17894 15674 0 sb_0__8_.mem_right_track_34.mem_out\[0\]
rlabel metal1 15272 6154 15272 6154 0 sb_0__8_.mem_right_track_36.ccff_tail
rlabel metal1 14306 6800 14306 6800 0 sb_0__8_.mem_right_track_36.mem_out\[0\]
rlabel metal1 16928 4794 16928 4794 0 sb_0__8_.mem_right_track_38.ccff_tail
rlabel metal2 15502 4522 15502 4522 0 sb_0__8_.mem_right_track_38.mem_out\[0\]
rlabel metal1 13938 28050 13938 28050 0 sb_0__8_.mem_right_track_4.ccff_tail
rlabel metal1 14444 30226 14444 30226 0 sb_0__8_.mem_right_track_4.mem_out\[0\]
rlabel metal2 12650 28322 12650 28322 0 sb_0__8_.mem_right_track_4.mem_out\[1\]
rlabel metal2 17710 6766 17710 6766 0 sb_0__8_.mem_right_track_40.ccff_tail
rlabel metal1 18446 4998 18446 4998 0 sb_0__8_.mem_right_track_40.mem_out\[0\]
rlabel metal2 21482 11254 21482 11254 0 sb_0__8_.mem_right_track_42.ccff_tail
rlabel metal2 18906 10098 18906 10098 0 sb_0__8_.mem_right_track_42.mem_out\[0\]
rlabel metal1 21114 15334 21114 15334 0 sb_0__8_.mem_right_track_44.ccff_tail
rlabel metal1 19826 15402 19826 15402 0 sb_0__8_.mem_right_track_44.mem_out\[0\]
rlabel metal2 23782 15402 23782 15402 0 sb_0__8_.mem_right_track_46.ccff_tail
rlabel metal1 21482 15912 21482 15912 0 sb_0__8_.mem_right_track_46.mem_out\[0\]
rlabel metal1 24610 13328 24610 13328 0 sb_0__8_.mem_right_track_48.ccff_tail
rlabel metal3 22609 19652 22609 19652 0 sb_0__8_.mem_right_track_48.mem_out\[0\]
rlabel metal2 24610 11322 24610 11322 0 sb_0__8_.mem_right_track_50.ccff_tail
rlabel metal2 24794 13192 24794 13192 0 sb_0__8_.mem_right_track_50.mem_out\[0\]
rlabel metal1 24748 8466 24748 8466 0 sb_0__8_.mem_right_track_52.ccff_tail
rlabel metal2 24058 9690 24058 9690 0 sb_0__8_.mem_right_track_52.mem_out\[0\]
rlabel metal2 21482 4522 21482 4522 0 sb_0__8_.mem_right_track_54.ccff_tail
rlabel metal1 19412 8398 19412 8398 0 sb_0__8_.mem_right_track_54.mem_out\[0\]
rlabel metal1 20884 9010 20884 9010 0 sb_0__8_.mem_right_track_56.ccff_tail
rlabel metal2 21114 9044 21114 9044 0 sb_0__8_.mem_right_track_56.mem_out\[0\]
rlabel metal1 19274 9350 19274 9350 0 sb_0__8_.mem_right_track_58.mem_out\[0\]
rlabel metal2 13478 24106 13478 24106 0 sb_0__8_.mem_right_track_6.ccff_tail
rlabel metal1 15778 28050 15778 28050 0 sb_0__8_.mem_right_track_6.mem_out\[0\]
rlabel metal2 15042 26758 15042 26758 0 sb_0__8_.mem_right_track_6.mem_out\[1\]
rlabel metal2 14122 24922 14122 24922 0 sb_0__8_.mem_right_track_8.mem_out\[0\]
rlabel metal1 13478 24684 13478 24684 0 sb_0__8_.mem_right_track_8.mem_out\[1\]
rlabel metal1 16790 8942 16790 8942 0 sb_0__8_.mux_bottom_track_1.out
rlabel metal1 20654 19482 20654 19482 0 sb_0__8_.mux_bottom_track_1.sky130_fd_sc_hd__mux2_1_0_X
rlabel metal2 20470 20400 20470 20400 0 sb_0__8_.mux_bottom_track_1.sky130_fd_sc_hd__mux2_1_1_X
rlabel metal1 18814 15062 18814 15062 0 sb_0__8_.mux_bottom_track_1.sky130_fd_sc_hd__mux2_1_2_X
rlabel metal2 20194 10336 20194 10336 0 sb_0__8_.mux_bottom_track_11.out
rlabel metal1 24886 22066 24886 22066 0 sb_0__8_.mux_bottom_track_11.sky130_fd_sc_hd__mux2_1_0_X
rlabel metal2 24610 19992 24610 19992 0 sb_0__8_.mux_bottom_track_11.sky130_fd_sc_hd__mux2_1_1_X
rlabel metal2 20654 13061 20654 13061 0 sb_0__8_.mux_bottom_track_13.out
rlabel metal1 23046 24786 23046 24786 0 sb_0__8_.mux_bottom_track_13.sky130_fd_sc_hd__mux2_1_0_X
rlabel metal2 21390 14076 21390 14076 0 sb_0__8_.mux_bottom_track_13.sky130_fd_sc_hd__mux2_1_1_X
rlabel metal3 18262 12444 18262 12444 0 sb_0__8_.mux_bottom_track_15.out
rlabel metal2 22310 25534 22310 25534 0 sb_0__8_.mux_bottom_track_15.sky130_fd_sc_hd__mux2_1_0_X
rlabel metal1 20378 21658 20378 21658 0 sb_0__8_.mux_bottom_track_15.sky130_fd_sc_hd__mux2_1_1_X
rlabel metal1 17526 16422 17526 16422 0 sb_0__8_.mux_bottom_track_17.out
rlabel metal1 18630 24276 18630 24276 0 sb_0__8_.mux_bottom_track_17.sky130_fd_sc_hd__mux2_1_0_X
rlabel metal1 17756 16558 17756 16558 0 sb_0__8_.mux_bottom_track_17.sky130_fd_sc_hd__mux2_1_1_X
rlabel metal2 17020 9452 17020 9452 0 sb_0__8_.mux_bottom_track_19.out
rlabel metal1 18354 26248 18354 26248 0 sb_0__8_.mux_bottom_track_19.sky130_fd_sc_hd__mux2_1_0_X
rlabel metal1 16836 17646 16836 17646 0 sb_0__8_.mux_bottom_track_19.sky130_fd_sc_hd__mux2_1_1_X
rlabel metal1 16100 18598 16100 18598 0 sb_0__8_.mux_bottom_track_29.out
rlabel metal1 18998 28118 18998 28118 0 sb_0__8_.mux_bottom_track_29.sky130_fd_sc_hd__mux2_1_0_X
rlabel metal1 16882 18734 16882 18734 0 sb_0__8_.mux_bottom_track_29.sky130_fd_sc_hd__mux2_1_1_X
rlabel metal1 24702 2312 24702 2312 0 sb_0__8_.mux_bottom_track_3.out
rlabel metal1 25024 17714 25024 17714 0 sb_0__8_.mux_bottom_track_3.sky130_fd_sc_hd__mux2_1_0_X
rlabel metal1 19458 17068 19458 17068 0 sb_0__8_.mux_bottom_track_3.sky130_fd_sc_hd__mux2_1_1_X
rlabel metal1 16468 19958 16468 19958 0 sb_0__8_.mux_bottom_track_31.out
rlabel metal1 20102 28390 20102 28390 0 sb_0__8_.mux_bottom_track_31.sky130_fd_sc_hd__mux2_1_0_X
rlabel metal1 19044 19822 19044 19822 0 sb_0__8_.mux_bottom_track_31.sky130_fd_sc_hd__mux2_1_1_X
rlabel metal1 21252 9622 21252 9622 0 sb_0__8_.mux_bottom_track_33.out
rlabel metal1 24334 32742 24334 32742 0 sb_0__8_.mux_bottom_track_33.sky130_fd_sc_hd__mux2_1_0_X
rlabel metal1 21482 13872 21482 13872 0 sb_0__8_.mux_bottom_track_33.sky130_fd_sc_hd__mux2_1_1_X
rlabel metal2 21252 15844 21252 15844 0 sb_0__8_.mux_bottom_track_35.out
rlabel metal1 24610 33286 24610 33286 0 sb_0__8_.mux_bottom_track_35.sky130_fd_sc_hd__mux2_1_0_X
rlabel metal1 21988 19346 21988 19346 0 sb_0__8_.mux_bottom_track_35.sky130_fd_sc_hd__mux2_1_1_X
rlabel metal1 19550 18054 19550 18054 0 sb_0__8_.mux_bottom_track_45.out
rlabel metal1 22632 34918 22632 34918 0 sb_0__8_.mux_bottom_track_45.sky130_fd_sc_hd__mux2_1_0_X
rlabel metal1 20332 18326 20332 18326 0 sb_0__8_.mux_bottom_track_45.sky130_fd_sc_hd__mux2_1_1_X
rlabel metal3 19159 19380 19159 19380 0 sb_0__8_.mux_bottom_track_47.out
rlabel metal1 21344 35462 21344 35462 0 sb_0__8_.mux_bottom_track_47.sky130_fd_sc_hd__mux2_1_0_X
rlabel metal1 19458 20502 19458 20502 0 sb_0__8_.mux_bottom_track_47.sky130_fd_sc_hd__mux2_1_1_X
rlabel metal1 13570 15062 13570 15062 0 sb_0__8_.mux_bottom_track_49.out
rlabel metal1 20332 35530 20332 35530 0 sb_0__8_.mux_bottom_track_49.sky130_fd_sc_hd__mux2_1_0_X
rlabel metal1 16054 22678 16054 22678 0 sb_0__8_.mux_bottom_track_49.sky130_fd_sc_hd__mux2_1_1_X
rlabel metal2 20930 10472 20930 10472 0 sb_0__8_.mux_bottom_track_5.out
rlabel metal1 23598 19482 23598 19482 0 sb_0__8_.mux_bottom_track_5.sky130_fd_sc_hd__mux2_1_0_X
rlabel metal2 21344 13804 21344 13804 0 sb_0__8_.mux_bottom_track_5.sky130_fd_sc_hd__mux2_1_1_X
rlabel metal1 19366 12716 19366 12716 0 sb_0__8_.mux_bottom_track_51.out
rlabel via2 21206 17323 21206 17323 0 sb_0__8_.mux_bottom_track_51.sky130_fd_sc_hd__mux2_1_0_X
rlabel metal2 22402 14926 22402 14926 0 sb_0__8_.mux_bottom_track_51.sky130_fd_sc_hd__mux2_1_1_X
rlabel metal1 15778 5270 15778 5270 0 sb_0__8_.mux_bottom_track_7.out
rlabel metal1 21022 22950 21022 22950 0 sb_0__8_.mux_bottom_track_7.sky130_fd_sc_hd__mux2_1_0_X
rlabel metal2 19918 23290 19918 23290 0 sb_0__8_.mux_bottom_track_7.sky130_fd_sc_hd__mux2_1_1_X
rlabel metal1 19734 17238 19734 17238 0 sb_0__8_.mux_bottom_track_7.sky130_fd_sc_hd__mux2_1_2_X
rlabel metal1 20056 14246 20056 14246 0 sb_0__8_.mux_bottom_track_9.out
rlabel metal1 22540 21658 22540 21658 0 sb_0__8_.mux_bottom_track_9.sky130_fd_sc_hd__mux2_1_0_X
rlabel metal1 20378 14348 20378 14348 0 sb_0__8_.mux_bottom_track_9.sky130_fd_sc_hd__mux2_1_1_X
rlabel metal1 18722 25160 18722 25160 0 sb_0__8_.mux_right_track_0.out
rlabel metal1 14536 32198 14536 32198 0 sb_0__8_.mux_right_track_0.sky130_fd_sc_hd__mux2_1_0_X
rlabel metal1 14536 31926 14536 31926 0 sb_0__8_.mux_right_track_0.sky130_fd_sc_hd__mux2_1_1_X
rlabel metal1 12098 25194 12098 25194 0 sb_0__8_.mux_right_track_0.sky130_fd_sc_hd__mux2_1_2_X
rlabel metal1 7958 17782 7958 17782 0 sb_0__8_.mux_right_track_0.sky130_fd_sc_hd__mux2_1_3_X
rlabel metal1 18078 25330 18078 25330 0 sb_0__8_.mux_right_track_0.sky130_fd_sc_hd__mux2_1_4_X
rlabel metal1 15870 19482 15870 19482 0 sb_0__8_.mux_right_track_10.out
rlabel metal1 13386 25160 13386 25160 0 sb_0__8_.mux_right_track_10.sky130_fd_sc_hd__mux2_1_0_X
rlabel metal1 13662 25704 13662 25704 0 sb_0__8_.mux_right_track_10.sky130_fd_sc_hd__mux2_1_1_X
rlabel metal1 11316 21862 11316 21862 0 sb_0__8_.mux_right_track_10.sky130_fd_sc_hd__mux2_1_2_X
rlabel metal1 7222 13498 7222 13498 0 sb_0__8_.mux_right_track_10.sky130_fd_sc_hd__mux2_1_3_X
rlabel metal2 14122 19040 14122 19040 0 sb_0__8_.mux_right_track_10.sky130_fd_sc_hd__mux2_1_4_X
rlabel metal1 16698 19720 16698 19720 0 sb_0__8_.mux_right_track_12.out
rlabel metal2 12374 21386 12374 21386 0 sb_0__8_.mux_right_track_12.sky130_fd_sc_hd__mux2_1_0_X
rlabel metal1 8602 16626 8602 16626 0 sb_0__8_.mux_right_track_12.sky130_fd_sc_hd__mux2_1_1_X
rlabel metal1 15778 19924 15778 19924 0 sb_0__8_.mux_right_track_12.sky130_fd_sc_hd__mux2_1_2_X
rlabel metal1 14904 14382 14904 14382 0 sb_0__8_.mux_right_track_14.out
rlabel metal1 15502 24582 15502 24582 0 sb_0__8_.mux_right_track_14.sky130_fd_sc_hd__mux2_1_0_X
rlabel metal1 14306 18802 14306 18802 0 sb_0__8_.mux_right_track_14.sky130_fd_sc_hd__mux2_1_1_X
rlabel metal2 14950 21726 14950 21726 0 sb_0__8_.mux_right_track_14.sky130_fd_sc_hd__mux2_1_2_X
rlabel metal1 16146 18258 16146 18258 0 sb_0__8_.mux_right_track_16.out
rlabel metal1 15686 20570 15686 20570 0 sb_0__8_.mux_right_track_16.sky130_fd_sc_hd__mux2_1_0_X
rlabel metal1 12926 17272 12926 17272 0 sb_0__8_.mux_right_track_16.sky130_fd_sc_hd__mux2_1_1_X
rlabel metal1 19366 19346 19366 19346 0 sb_0__8_.mux_right_track_16.sky130_fd_sc_hd__mux2_1_2_X
rlabel metal1 20930 14382 20930 14382 0 sb_0__8_.mux_right_track_18.out
rlabel metal1 13800 15674 13800 15674 0 sb_0__8_.mux_right_track_18.sky130_fd_sc_hd__mux2_1_0_X
rlabel metal1 14122 16184 14122 16184 0 sb_0__8_.mux_right_track_18.sky130_fd_sc_hd__mux2_1_1_X
rlabel metal1 19458 25738 19458 25738 0 sb_0__8_.mux_right_track_2.out
rlabel metal1 14214 28186 14214 28186 0 sb_0__8_.mux_right_track_2.sky130_fd_sc_hd__mux2_1_0_X
rlabel metal1 14766 28118 14766 28118 0 sb_0__8_.mux_right_track_2.sky130_fd_sc_hd__mux2_1_1_X
rlabel metal2 12834 27098 12834 27098 0 sb_0__8_.mux_right_track_2.sky130_fd_sc_hd__mux2_1_2_X
rlabel metal1 10212 21114 10212 21114 0 sb_0__8_.mux_right_track_2.sky130_fd_sc_hd__mux2_1_3_X
rlabel metal2 12926 26248 12926 26248 0 sb_0__8_.mux_right_track_2.sky130_fd_sc_hd__mux2_1_4_X
rlabel metal1 17158 12954 17158 12954 0 sb_0__8_.mux_right_track_20.out
rlabel metal1 11684 10098 11684 10098 0 sb_0__8_.mux_right_track_20.sky130_fd_sc_hd__mux2_1_0_X
rlabel metal1 16054 12818 16054 12818 0 sb_0__8_.mux_right_track_20.sky130_fd_sc_hd__mux2_1_1_X
rlabel metal1 20378 11084 20378 11084 0 sb_0__8_.mux_right_track_22.out
rlabel metal1 11362 7786 11362 7786 0 sb_0__8_.mux_right_track_22.sky130_fd_sc_hd__mux2_1_0_X
rlabel metal2 11822 8211 11822 8211 0 sb_0__8_.mux_right_track_22.sky130_fd_sc_hd__mux2_1_1_X
rlabel metal1 21436 12818 21436 12818 0 sb_0__8_.mux_right_track_24.out
rlabel metal1 12052 7514 12052 7514 0 sb_0__8_.mux_right_track_24.sky130_fd_sc_hd__mux2_1_0_X
rlabel metal1 14306 7718 14306 7718 0 sb_0__8_.mux_right_track_24.sky130_fd_sc_hd__mux2_1_1_X
rlabel metal1 18722 13192 18722 13192 0 sb_0__8_.mux_right_track_26.out
rlabel metal1 14950 12954 14950 12954 0 sb_0__8_.mux_right_track_26.sky130_fd_sc_hd__mux2_1_0_X
rlabel metal1 18906 13362 18906 13362 0 sb_0__8_.mux_right_track_26.sky130_fd_sc_hd__mux2_1_1_X
rlabel metal1 19136 14382 19136 14382 0 sb_0__8_.mux_right_track_28.out
rlabel metal1 17158 19482 17158 19482 0 sb_0__8_.mux_right_track_28.sky130_fd_sc_hd__mux2_1_0_X
rlabel metal1 13708 15130 13708 15130 0 sb_0__8_.mux_right_track_28.sky130_fd_sc_hd__mux2_1_1_X
rlabel metal2 20286 18836 20286 18836 0 sb_0__8_.mux_right_track_28.sky130_fd_sc_hd__mux2_1_2_X
rlabel metal1 22862 2550 22862 2550 0 sb_0__8_.mux_right_track_30.out
rlabel metal1 17940 19890 17940 19890 0 sb_0__8_.mux_right_track_30.sky130_fd_sc_hd__mux2_1_0_X
rlabel metal1 15870 16422 15870 16422 0 sb_0__8_.mux_right_track_30.sky130_fd_sc_hd__mux2_1_1_X
rlabel metal1 21850 15504 21850 15504 0 sb_0__8_.mux_right_track_30.sky130_fd_sc_hd__mux2_1_2_X
rlabel metal1 19504 14586 19504 14586 0 sb_0__8_.mux_right_track_32.out
rlabel metal1 18492 17714 18492 17714 0 sb_0__8_.mux_right_track_32.sky130_fd_sc_hd__mux2_1_0_X
rlabel metal2 15594 16218 15594 16218 0 sb_0__8_.mux_right_track_32.sky130_fd_sc_hd__mux2_1_1_X
rlabel metal1 19734 14416 19734 14416 0 sb_0__8_.mux_right_track_32.sky130_fd_sc_hd__mux2_1_2_X
rlabel metal2 9522 8126 9522 8126 0 sb_0__8_.mux_right_track_34.out
rlabel metal1 16928 18598 16928 18598 0 sb_0__8_.mux_right_track_34.sky130_fd_sc_hd__mux2_1_0_X
rlabel metal1 13570 7174 13570 7174 0 sb_0__8_.mux_right_track_34.sky130_fd_sc_hd__mux2_1_1_X
rlabel metal1 19274 5236 19274 5236 0 sb_0__8_.mux_right_track_34.sky130_fd_sc_hd__mux2_1_2_X
rlabel metal1 11040 9146 11040 9146 0 sb_0__8_.mux_right_track_36.out
rlabel metal1 15134 6358 15134 6358 0 sb_0__8_.mux_right_track_36.sky130_fd_sc_hd__mux2_1_0_X
rlabel metal1 14766 6086 14766 6086 0 sb_0__8_.mux_right_track_36.sky130_fd_sc_hd__mux2_1_1_X
rlabel metal2 10994 4794 10994 4794 0 sb_0__8_.mux_right_track_38.out
rlabel metal1 16790 6664 16790 6664 0 sb_0__8_.mux_right_track_38.sky130_fd_sc_hd__mux2_1_0_X
rlabel metal2 15318 5576 15318 5576 0 sb_0__8_.mux_right_track_38.sky130_fd_sc_hd__mux2_1_1_X
rlabel metal1 19228 21522 19228 21522 0 sb_0__8_.mux_right_track_4.out
rlabel metal1 15042 29274 15042 29274 0 sb_0__8_.mux_right_track_4.sky130_fd_sc_hd__mux2_1_0_X
rlabel metal2 14582 29648 14582 29648 0 sb_0__8_.mux_right_track_4.sky130_fd_sc_hd__mux2_1_1_X
rlabel metal1 13570 26282 13570 26282 0 sb_0__8_.mux_right_track_4.sky130_fd_sc_hd__mux2_1_2_X
rlabel metal1 12972 26282 12972 26282 0 sb_0__8_.mux_right_track_4.sky130_fd_sc_hd__mux2_1_3_X
rlabel metal1 17802 25908 17802 25908 0 sb_0__8_.mux_right_track_4.sky130_fd_sc_hd__mux2_1_4_X
rlabel metal2 21298 2244 21298 2244 0 sb_0__8_.mux_right_track_40.out
rlabel metal2 17526 7888 17526 7888 0 sb_0__8_.mux_right_track_40.sky130_fd_sc_hd__mux2_1_0_X
rlabel metal1 21482 2482 21482 2482 0 sb_0__8_.mux_right_track_40.sky130_fd_sc_hd__mux2_1_1_X
rlabel metal1 10074 4658 10074 4658 0 sb_0__8_.mux_right_track_42.out
rlabel metal1 20608 10098 20608 10098 0 sb_0__8_.mux_right_track_42.sky130_fd_sc_hd__mux2_1_0_X
rlabel metal2 20746 8976 20746 8976 0 sb_0__8_.mux_right_track_42.sky130_fd_sc_hd__mux2_1_1_X
rlabel metal1 13110 9044 13110 9044 0 sb_0__8_.mux_right_track_44.out
rlabel metal1 19918 15130 19918 15130 0 sb_0__8_.mux_right_track_44.sky130_fd_sc_hd__mux2_1_0_X
rlabel metal1 19412 14994 19412 14994 0 sb_0__8_.mux_right_track_44.sky130_fd_sc_hd__mux2_1_1_X
rlabel metal1 14536 13294 14536 13294 0 sb_0__8_.mux_right_track_44.sky130_fd_sc_hd__mux2_1_2_X
rlabel metal2 22034 10353 22034 10353 0 sb_0__8_.mux_right_track_46.out
rlabel metal1 19734 21896 19734 21896 0 sb_0__8_.mux_right_track_46.sky130_fd_sc_hd__mux2_1_0_X
rlabel metal1 19320 12614 19320 12614 0 sb_0__8_.mux_right_track_46.sky130_fd_sc_hd__mux2_1_1_X
rlabel metal1 12926 12852 12926 12852 0 sb_0__8_.mux_right_track_46.sky130_fd_sc_hd__mux2_1_2_X
rlabel metal2 14306 6052 14306 6052 0 sb_0__8_.mux_right_track_48.out
rlabel metal1 21942 13260 21942 13260 0 sb_0__8_.mux_right_track_48.sky130_fd_sc_hd__mux2_1_0_X
rlabel metal1 20102 11866 20102 11866 0 sb_0__8_.mux_right_track_48.sky130_fd_sc_hd__mux2_1_1_X
rlabel metal1 21620 13158 21620 13158 0 sb_0__8_.mux_right_track_48.sky130_fd_sc_hd__mux2_1_2_X
rlabel metal2 12834 4896 12834 4896 0 sb_0__8_.mux_right_track_50.out
rlabel metal2 20194 12172 20194 12172 0 sb_0__8_.mux_right_track_50.sky130_fd_sc_hd__mux2_1_0_X
rlabel metal1 13478 4216 13478 4216 0 sb_0__8_.mux_right_track_50.sky130_fd_sc_hd__mux2_1_1_X
rlabel metal1 12673 4658 12673 4658 0 sb_0__8_.mux_right_track_52.out
rlabel metal2 19918 9248 19918 9248 0 sb_0__8_.mux_right_track_52.sky130_fd_sc_hd__mux2_1_0_X
rlabel metal1 10488 4590 10488 4590 0 sb_0__8_.mux_right_track_52.sky130_fd_sc_hd__mux2_1_1_X
rlabel metal1 11730 3502 11730 3502 0 sb_0__8_.mux_right_track_54.out
rlabel metal1 20148 4046 20148 4046 0 sb_0__8_.mux_right_track_54.sky130_fd_sc_hd__mux2_1_0_X
rlabel metal1 16652 3910 16652 3910 0 sb_0__8_.mux_right_track_54.sky130_fd_sc_hd__mux2_1_1_X
rlabel metal1 12811 5202 12811 5202 0 sb_0__8_.mux_right_track_56.out
rlabel metal1 19274 9010 19274 9010 0 sb_0__8_.mux_right_track_56.sky130_fd_sc_hd__mux2_1_0_X
rlabel metal3 17572 3536 17572 3536 0 sb_0__8_.mux_right_track_56.sky130_fd_sc_hd__mux2_1_1_X
rlabel metal2 16330 3944 16330 3944 0 sb_0__8_.mux_right_track_58.out
rlabel metal2 19044 14892 19044 14892 0 sb_0__8_.mux_right_track_58.sky130_fd_sc_hd__mux2_1_0_X
rlabel metal2 16790 10200 16790 10200 0 sb_0__8_.mux_right_track_58.sky130_fd_sc_hd__mux2_1_1_X
rlabel metal1 16652 12206 16652 12206 0 sb_0__8_.mux_right_track_58.sky130_fd_sc_hd__mux2_1_2_X
rlabel metal1 17894 20978 17894 20978 0 sb_0__8_.mux_right_track_6.out
rlabel metal1 15778 26282 15778 26282 0 sb_0__8_.mux_right_track_6.sky130_fd_sc_hd__mux2_1_0_X
rlabel metal2 14858 27098 14858 27098 0 sb_0__8_.mux_right_track_6.sky130_fd_sc_hd__mux2_1_1_X
rlabel metal1 14214 23834 14214 23834 0 sb_0__8_.mux_right_track_6.sky130_fd_sc_hd__mux2_1_2_X
rlabel metal2 12558 20145 12558 20145 0 sb_0__8_.mux_right_track_6.sky130_fd_sc_hd__mux2_1_3_X
rlabel metal1 18262 23732 18262 23732 0 sb_0__8_.mux_right_track_6.sky130_fd_sc_hd__mux2_1_4_X
rlabel metal1 18446 22474 18446 22474 0 sb_0__8_.mux_right_track_8.out
rlabel metal2 14398 25772 14398 25772 0 sb_0__8_.mux_right_track_8.sky130_fd_sc_hd__mux2_1_0_X
rlabel metal1 14904 24922 14904 24922 0 sb_0__8_.mux_right_track_8.sky130_fd_sc_hd__mux2_1_1_X
rlabel via1 13386 22491 13386 22491 0 sb_0__8_.mux_right_track_8.sky130_fd_sc_hd__mux2_1_2_X
rlabel metal1 10580 16966 10580 16966 0 sb_0__8_.mux_right_track_8.sky130_fd_sc_hd__mux2_1_3_X
rlabel metal1 17066 22678 17066 22678 0 sb_0__8_.mux_right_track_8.sky130_fd_sc_hd__mux2_1_4_X
<< properties >>
string FIXED_BBOX 0 0 27000 57000
<< end >>
