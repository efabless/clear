magic
tech sky130A
magscale 1 2
timestamp 1682506515
<< viali >>
rect 14565 54281 14599 54315
rect 16405 54281 16439 54315
rect 24501 54281 24535 54315
rect 24685 54281 24719 54315
rect 5825 54213 5859 54247
rect 8401 54213 8435 54247
rect 10977 54213 11011 54247
rect 14105 54213 14139 54247
rect 18429 54213 18463 54247
rect 21465 54213 21499 54247
rect 23305 54213 23339 54247
rect 2237 54145 2271 54179
rect 4629 54145 4663 54179
rect 7389 54145 7423 54179
rect 9965 54145 9999 54179
rect 11897 54145 11931 54179
rect 12357 54145 12391 54179
rect 14841 54145 14875 54179
rect 15577 54145 15611 54179
rect 16129 54145 16163 54179
rect 16865 54145 16899 54179
rect 17601 54145 17635 54179
rect 18981 54145 19015 54179
rect 19441 54145 19475 54179
rect 20177 54145 20211 54179
rect 20913 54145 20947 54179
rect 22017 54145 22051 54179
rect 22753 54145 22787 54179
rect 23765 54145 23799 54179
rect 25053 54145 25087 54179
rect 3249 54077 3283 54111
rect 12817 54077 12851 54111
rect 15025 54009 15059 54043
rect 17785 54009 17819 54043
rect 20361 54009 20395 54043
rect 25237 54009 25271 54043
rect 11713 53941 11747 53975
rect 15761 53941 15795 53975
rect 17049 53941 17083 53975
rect 18521 53941 18555 53975
rect 19625 53941 19659 53975
rect 21097 53941 21131 53975
rect 22201 53941 22235 53975
rect 22937 53941 22971 53975
rect 23949 53941 23983 53975
rect 16405 53737 16439 53771
rect 18889 53737 18923 53771
rect 21281 53669 21315 53703
rect 23121 53669 23155 53703
rect 3249 53601 3283 53635
rect 6561 53601 6595 53635
rect 8401 53601 8435 53635
rect 11069 53601 11103 53635
rect 12725 53601 12759 53635
rect 24409 53601 24443 53635
rect 2237 53533 2271 53567
rect 5549 53533 5583 53567
rect 7297 53533 7331 53567
rect 10425 53533 10459 53567
rect 12449 53533 12483 53567
rect 14289 53533 14323 53567
rect 14841 53533 14875 53567
rect 15669 53533 15703 53567
rect 16129 53533 16163 53567
rect 16681 53533 16715 53567
rect 17601 53533 17635 53567
rect 18245 53533 18279 53567
rect 18705 53533 18739 53567
rect 19441 53533 19475 53567
rect 20269 53533 20303 53567
rect 20729 53533 20763 53567
rect 21097 53533 21131 53567
rect 22017 53533 22051 53567
rect 22661 53533 22695 53567
rect 23305 53533 23339 53567
rect 23857 53533 23891 53567
rect 24961 53533 24995 53567
rect 18429 53465 18463 53499
rect 20453 53465 20487 53499
rect 14473 53397 14507 53431
rect 15761 53397 15795 53431
rect 16865 53397 16899 53431
rect 17417 53397 17451 53431
rect 19625 53397 19659 53431
rect 21833 53397 21867 53431
rect 22477 53397 22511 53431
rect 23949 53397 23983 53431
rect 25053 53397 25087 53431
rect 2145 53193 2179 53227
rect 17325 53193 17359 53227
rect 19533 53193 19567 53227
rect 19717 53193 19751 53227
rect 21005 53193 21039 53227
rect 21833 53193 21867 53227
rect 22293 53193 22327 53227
rect 22569 53193 22603 53227
rect 23029 53193 23063 53227
rect 3985 53125 4019 53159
rect 5825 53125 5859 53159
rect 9137 53125 9171 53159
rect 13829 53125 13863 53159
rect 21189 53125 21223 53159
rect 1777 53057 1811 53091
rect 2973 53057 3007 53091
rect 4813 53057 4847 53091
rect 8125 53057 8159 53091
rect 9781 53057 9815 53091
rect 11897 53057 11931 53091
rect 14657 53057 14691 53091
rect 14933 53057 14967 53091
rect 16129 53057 16163 53091
rect 16405 53057 16439 53091
rect 19073 53057 19107 53091
rect 19349 53057 19383 53091
rect 20545 53057 20579 53091
rect 20821 53057 20855 53091
rect 23489 53057 23523 53091
rect 24133 53057 24167 53091
rect 24409 53057 24443 53091
rect 24777 53057 24811 53091
rect 25053 53057 25087 53091
rect 10425 52989 10459 53023
rect 12357 52989 12391 53023
rect 14013 52921 14047 52955
rect 1593 52853 1627 52887
rect 14473 52853 14507 52887
rect 15945 52853 15979 52887
rect 18889 52853 18923 52887
rect 20361 52853 20395 52887
rect 23305 52853 23339 52887
rect 23949 52853 23983 52887
rect 25237 52853 25271 52887
rect 12633 52649 12667 52683
rect 14105 52649 14139 52683
rect 24593 52649 24627 52683
rect 25237 52581 25271 52615
rect 3249 52513 3283 52547
rect 6561 52513 6595 52547
rect 7757 52513 7791 52547
rect 11253 52513 11287 52547
rect 13645 52513 13679 52547
rect 2237 52445 2271 52479
rect 5457 52445 5491 52479
rect 7205 52445 7239 52479
rect 10793 52445 10827 52479
rect 12817 52445 12851 52479
rect 24777 52445 24811 52479
rect 25053 52445 25087 52479
rect 13461 52377 13495 52411
rect 7021 52105 7055 52139
rect 11713 52105 11747 52139
rect 12357 52105 12391 52139
rect 13277 52105 13311 52139
rect 25329 52105 25363 52139
rect 6929 52037 6963 52071
rect 2973 51969 3007 52003
rect 4813 51969 4847 52003
rect 7849 51969 7883 52003
rect 9873 51969 9907 52003
rect 11897 51969 11931 52003
rect 12541 51969 12575 52003
rect 3341 51901 3375 51935
rect 5089 51901 5123 51935
rect 8493 51901 8527 51935
rect 10149 51901 10183 51935
rect 25513 51765 25547 51799
rect 10241 51561 10275 51595
rect 2881 51425 2915 51459
rect 5733 51425 5767 51459
rect 7573 51425 7607 51459
rect 2237 51357 2271 51391
rect 5457 51357 5491 51391
rect 7113 51357 7147 51391
rect 10425 51357 10459 51391
rect 25053 51357 25087 51391
rect 25237 51221 25271 51255
rect 6929 51017 6963 51051
rect 9597 50949 9631 50983
rect 2513 50881 2547 50915
rect 4353 50881 4387 50915
rect 6837 50881 6871 50915
rect 7757 50881 7791 50915
rect 9413 50881 9447 50915
rect 24777 50881 24811 50915
rect 25053 50881 25087 50915
rect 2789 50813 2823 50847
rect 4629 50813 4663 50847
rect 7481 50813 7515 50847
rect 25237 50677 25271 50711
rect 6837 50473 6871 50507
rect 9229 50473 9263 50507
rect 25145 50405 25179 50439
rect 3249 50337 3283 50371
rect 2237 50269 2271 50303
rect 7021 50269 7055 50303
rect 9413 50269 9447 50303
rect 24685 50269 24719 50303
rect 25329 50269 25363 50303
rect 24777 50133 24811 50167
rect 6377 49929 6411 49963
rect 3157 49861 3191 49895
rect 6561 49861 6595 49895
rect 9413 49861 9447 49895
rect 2145 49793 2179 49827
rect 3985 49793 4019 49827
rect 9229 49793 9263 49827
rect 24777 49793 24811 49827
rect 6009 49725 6043 49759
rect 24501 49725 24535 49759
rect 4242 49589 4276 49623
rect 11621 49385 11655 49419
rect 12725 49385 12759 49419
rect 2053 49249 2087 49283
rect 1777 49181 1811 49215
rect 11805 49181 11839 49215
rect 12909 49181 12943 49215
rect 24869 49181 24903 49215
rect 25329 49181 25363 49215
rect 3341 49045 3375 49079
rect 25145 49045 25179 49079
rect 24501 48637 24535 48671
rect 24777 48637 24811 48671
rect 18153 48229 18187 48263
rect 17141 48093 17175 48127
rect 17785 47957 17819 47991
rect 25237 47957 25271 47991
rect 25513 47957 25547 47991
rect 9229 47753 9263 47787
rect 17233 47753 17267 47787
rect 18429 47753 18463 47787
rect 18521 47753 18555 47787
rect 19257 47753 19291 47787
rect 19165 47685 19199 47719
rect 9413 47617 9447 47651
rect 17325 47617 17359 47651
rect 24501 47617 24535 47651
rect 17417 47549 17451 47583
rect 18705 47549 18739 47583
rect 24777 47549 24811 47583
rect 11989 47413 12023 47447
rect 16865 47413 16899 47447
rect 18061 47413 18095 47447
rect 18153 47141 18187 47175
rect 10149 47073 10183 47107
rect 15761 47073 15795 47107
rect 17509 47073 17543 47107
rect 18613 47073 18647 47107
rect 18797 47073 18831 47107
rect 12357 47005 12391 47039
rect 18521 47005 18555 47039
rect 19441 47005 19475 47039
rect 20545 47005 20579 47039
rect 23213 47005 23247 47039
rect 23489 47005 23523 47039
rect 10425 46937 10459 46971
rect 16037 46937 16071 46971
rect 20085 46937 20119 46971
rect 24409 46937 24443 46971
rect 25237 46937 25271 46971
rect 11897 46869 11931 46903
rect 13001 46869 13035 46903
rect 14289 46869 14323 46903
rect 17785 46869 17819 46903
rect 21189 46869 21223 46903
rect 25421 46869 25455 46903
rect 7297 46665 7331 46699
rect 11161 46665 11195 46699
rect 11713 46665 11747 46699
rect 16313 46665 16347 46699
rect 18613 46665 18647 46699
rect 19441 46665 19475 46699
rect 20085 46665 20119 46699
rect 20177 46665 20211 46699
rect 21557 46665 21591 46699
rect 22385 46665 22419 46699
rect 22477 46665 22511 46699
rect 7481 46529 7515 46563
rect 10517 46529 10551 46563
rect 11897 46529 11931 46563
rect 16865 46529 16899 46563
rect 12357 46461 12391 46495
rect 12633 46461 12667 46495
rect 14565 46461 14599 46495
rect 14841 46461 14875 46495
rect 17141 46461 17175 46495
rect 20361 46461 20395 46495
rect 22569 46461 22603 46495
rect 24501 46461 24535 46495
rect 24777 46461 24811 46495
rect 14105 46325 14139 46359
rect 18981 46325 19015 46359
rect 19165 46325 19199 46359
rect 19717 46325 19751 46359
rect 22017 46325 22051 46359
rect 24225 46325 24259 46359
rect 8125 46121 8159 46155
rect 9137 46121 9171 46155
rect 10701 46121 10735 46155
rect 14197 46121 14231 46155
rect 16497 46121 16531 46155
rect 22017 46121 22051 46155
rect 10057 46053 10091 46087
rect 16865 46053 16899 46087
rect 11345 45985 11379 46019
rect 11897 45985 11931 46019
rect 17141 45985 17175 46019
rect 17417 45985 17451 46019
rect 19809 45985 19843 46019
rect 22845 45985 22879 46019
rect 9321 45917 9355 45951
rect 10241 45917 10275 45951
rect 11069 45917 11103 45951
rect 15853 45917 15887 45951
rect 19533 45917 19567 45951
rect 22661 45917 22695 45951
rect 22753 45917 22787 45951
rect 24593 45917 24627 45951
rect 8033 45849 8067 45883
rect 12173 45849 12207 45883
rect 8585 45781 8619 45815
rect 11161 45781 11195 45815
rect 13645 45781 13679 45815
rect 18889 45781 18923 45815
rect 21281 45781 21315 45815
rect 21649 45781 21683 45815
rect 22293 45781 22327 45815
rect 23857 45781 23891 45815
rect 23949 45781 23983 45815
rect 24225 45781 24259 45815
rect 25237 45781 25271 45815
rect 11897 45577 11931 45611
rect 19993 45577 20027 45611
rect 8769 45509 8803 45543
rect 9413 45509 9447 45543
rect 20913 45509 20947 45543
rect 9137 45441 9171 45475
rect 11805 45441 11839 45475
rect 12265 45441 12299 45475
rect 13553 45441 13587 45475
rect 16865 45441 16899 45475
rect 20821 45441 20855 45475
rect 22109 45441 22143 45475
rect 13645 45373 13679 45407
rect 13737 45373 13771 45407
rect 14381 45373 14415 45407
rect 14657 45373 14691 45407
rect 17509 45373 17543 45407
rect 18245 45373 18279 45407
rect 18521 45373 18555 45407
rect 21097 45373 21131 45407
rect 22385 45373 22419 45407
rect 24133 45373 24167 45407
rect 24501 45373 24535 45407
rect 24777 45373 24811 45407
rect 11161 45305 11195 45339
rect 13185 45305 13219 45339
rect 10885 45237 10919 45271
rect 16129 45237 16163 45271
rect 16497 45237 16531 45271
rect 20453 45237 20487 45271
rect 21557 45237 21591 45271
rect 23857 45237 23891 45271
rect 7849 45033 7883 45067
rect 8401 45033 8435 45067
rect 11253 45033 11287 45067
rect 18889 45033 18923 45067
rect 21465 45033 21499 45067
rect 21833 45033 21867 45067
rect 12449 44965 12483 44999
rect 9413 44897 9447 44931
rect 11897 44897 11931 44931
rect 15117 44897 15151 44931
rect 19993 44897 20027 44931
rect 22569 44897 22603 44931
rect 25237 44897 25271 44931
rect 8585 44829 8619 44863
rect 13093 44829 13127 44863
rect 18245 44829 18279 44863
rect 19717 44829 19751 44863
rect 22293 44829 22327 44863
rect 24593 44829 24627 44863
rect 7757 44761 7791 44795
rect 9229 44761 9263 44795
rect 11161 44761 11195 44795
rect 12265 44761 12299 44795
rect 12725 44761 12759 44795
rect 15393 44761 15427 44795
rect 6469 44693 6503 44727
rect 7297 44693 7331 44727
rect 9781 44693 9815 44727
rect 11621 44693 11655 44727
rect 13737 44693 13771 44727
rect 16865 44693 16899 44727
rect 17233 44693 17267 44727
rect 19349 44693 19383 44727
rect 24041 44693 24075 44727
rect 5825 44489 5859 44523
rect 6745 44489 6779 44523
rect 9045 44489 9079 44523
rect 11069 44489 11103 44523
rect 11897 44489 11931 44523
rect 15209 44489 15243 44523
rect 20821 44489 20855 44523
rect 7573 44421 7607 44455
rect 13369 44421 13403 44455
rect 6009 44353 6043 44387
rect 6653 44353 6687 44387
rect 7389 44353 7423 44387
rect 8953 44353 8987 44387
rect 9873 44353 9907 44387
rect 10241 44353 10275 44387
rect 10977 44353 11011 44387
rect 12265 44353 12299 44387
rect 13093 44353 13127 44387
rect 16865 44353 16899 44387
rect 19073 44353 19107 44387
rect 20177 44353 20211 44387
rect 24777 44353 24811 44387
rect 12357 44285 12391 44319
rect 12449 44285 12483 44319
rect 17141 44285 17175 44319
rect 22293 44285 22327 44319
rect 22569 44285 22603 44319
rect 24501 44285 24535 44319
rect 11621 44217 11655 44251
rect 7849 44149 7883 44183
rect 9413 44149 9447 44183
rect 10333 44149 10367 44183
rect 14841 44149 14875 44183
rect 18613 44149 18647 44183
rect 19717 44149 19751 44183
rect 21925 44149 21959 44183
rect 24041 44149 24075 44183
rect 6745 43945 6779 43979
rect 8401 43945 8435 43979
rect 10885 43945 10919 43979
rect 11345 43945 11379 43979
rect 21557 43945 21591 43979
rect 7205 43877 7239 43911
rect 18153 43877 18187 43911
rect 9137 43809 9171 43843
rect 17509 43809 17543 43843
rect 17601 43809 17635 43843
rect 18337 43809 18371 43843
rect 22569 43809 22603 43843
rect 22753 43809 22787 43843
rect 6653 43741 6687 43775
rect 8585 43741 8619 43775
rect 14289 43741 14323 43775
rect 15393 43741 15427 43775
rect 17417 43741 17451 43775
rect 19441 43741 19475 43775
rect 20913 43741 20947 43775
rect 23305 43741 23339 43775
rect 25329 43741 25363 43775
rect 9413 43673 9447 43707
rect 20453 43673 20487 43707
rect 22477 43673 22511 43707
rect 14933 43605 14967 43639
rect 16037 43605 16071 43639
rect 17049 43605 17083 43639
rect 18797 43605 18831 43639
rect 20085 43605 20119 43639
rect 20545 43605 20579 43639
rect 22109 43605 22143 43639
rect 23949 43605 23983 43639
rect 24501 43605 24535 43639
rect 24685 43605 24719 43639
rect 25145 43605 25179 43639
rect 7757 43401 7791 43435
rect 9137 43401 9171 43435
rect 15209 43401 15243 43435
rect 17325 43401 17359 43435
rect 22477 43401 22511 43435
rect 23305 43401 23339 43435
rect 8677 43333 8711 43367
rect 9505 43333 9539 43367
rect 12817 43333 12851 43367
rect 21373 43333 21407 43367
rect 1685 43265 1719 43299
rect 2145 43265 2179 43299
rect 7941 43265 7975 43299
rect 8493 43265 8527 43299
rect 10149 43265 10183 43299
rect 15301 43265 15335 43299
rect 18245 43265 18279 43299
rect 20545 43265 20579 43299
rect 22385 43265 22419 43299
rect 23029 43265 23063 43299
rect 9597 43197 9631 43231
rect 9689 43197 9723 43231
rect 12541 43197 12575 43231
rect 15393 43197 15427 43231
rect 17417 43197 17451 43231
rect 17601 43197 17635 43231
rect 18521 43197 18555 43231
rect 22569 43197 22603 43231
rect 23581 43197 23615 43231
rect 23857 43197 23891 43231
rect 1869 43129 1903 43163
rect 14289 43129 14323 43163
rect 15853 43129 15887 43163
rect 7481 43061 7515 43095
rect 14841 43061 14875 43095
rect 16037 43061 16071 43095
rect 16405 43061 16439 43095
rect 16957 43061 16991 43095
rect 19993 43061 20027 43095
rect 22017 43061 22051 43095
rect 25329 43061 25363 43095
rect 8953 42857 8987 42891
rect 9229 42857 9263 42891
rect 16865 42857 16899 42891
rect 19888 42857 19922 42891
rect 13001 42789 13035 42823
rect 16497 42789 16531 42823
rect 4997 42721 5031 42755
rect 9413 42721 9447 42755
rect 10885 42721 10919 42755
rect 12633 42721 12667 42755
rect 14749 42721 14783 42755
rect 22477 42721 22511 42755
rect 23489 42721 23523 42755
rect 7849 42653 7883 42687
rect 9781 42653 9815 42687
rect 18705 42653 18739 42687
rect 19625 42653 19659 42687
rect 22937 42653 22971 42687
rect 23213 42653 23247 42687
rect 24685 42653 24719 42687
rect 4813 42585 4847 42619
rect 10425 42585 10459 42619
rect 11161 42585 11195 42619
rect 15025 42585 15059 42619
rect 17693 42585 17727 42619
rect 17969 42585 18003 42619
rect 22293 42585 22327 42619
rect 5365 42517 5399 42551
rect 8493 42517 8527 42551
rect 21373 42517 21407 42551
rect 21833 42517 21867 42551
rect 22201 42517 22235 42551
rect 25329 42517 25363 42551
rect 5825 42313 5859 42347
rect 9781 42313 9815 42347
rect 11069 42313 11103 42347
rect 11713 42313 11747 42347
rect 12909 42313 12943 42347
rect 15301 42313 15335 42347
rect 15761 42313 15795 42347
rect 17141 42313 17175 42347
rect 17601 42313 17635 42347
rect 18245 42313 18279 42347
rect 23029 42313 23063 42347
rect 25237 42313 25271 42347
rect 7849 42245 7883 42279
rect 10241 42245 10275 42279
rect 13369 42245 13403 42279
rect 19073 42245 19107 42279
rect 23765 42245 23799 42279
rect 5365 42177 5399 42211
rect 5733 42177 5767 42211
rect 7573 42177 7607 42211
rect 10149 42177 10183 42211
rect 12081 42177 12115 42211
rect 13277 42177 13311 42211
rect 14105 42177 14139 42211
rect 15669 42177 15703 42211
rect 17509 42177 17543 42211
rect 18797 42177 18831 42211
rect 21465 42177 21499 42211
rect 22385 42177 22419 42211
rect 9321 42109 9355 42143
rect 10333 42109 10367 42143
rect 12173 42109 12207 42143
rect 12357 42109 12391 42143
rect 13553 42109 13587 42143
rect 15853 42109 15887 42143
rect 17693 42109 17727 42143
rect 22017 42109 22051 42143
rect 23489 42109 23523 42143
rect 16865 42041 16899 42075
rect 20545 42041 20579 42075
rect 21281 42041 21315 42075
rect 21925 42041 21959 42075
rect 10793 41973 10827 42007
rect 20913 41973 20947 42007
rect 4169 41769 4203 41803
rect 4905 41769 4939 41803
rect 8033 41769 8067 41803
rect 8769 41769 8803 41803
rect 11529 41769 11563 41803
rect 22661 41769 22695 41803
rect 25237 41769 25271 41803
rect 7757 41701 7791 41735
rect 21373 41701 21407 41735
rect 6009 41633 6043 41667
rect 6285 41633 6319 41667
rect 9597 41633 9631 41667
rect 9781 41633 9815 41667
rect 10885 41633 10919 41667
rect 12081 41633 12115 41667
rect 14841 41633 14875 41667
rect 15669 41633 15703 41667
rect 15761 41633 15795 41667
rect 16957 41633 16991 41667
rect 18613 41633 18647 41667
rect 18705 41633 18739 41667
rect 20177 41633 20211 41667
rect 22017 41633 22051 41667
rect 23121 41633 23155 41667
rect 23305 41633 23339 41667
rect 8309 41565 8343 41599
rect 12725 41565 12759 41599
rect 16865 41565 16899 41599
rect 17509 41565 17543 41599
rect 20085 41565 20119 41599
rect 24041 41565 24075 41599
rect 24593 41565 24627 41599
rect 3617 41497 3651 41531
rect 4077 41497 4111 41531
rect 4813 41497 4847 41531
rect 5273 41497 5307 41531
rect 11897 41497 11931 41531
rect 11989 41497 12023 41531
rect 15577 41497 15611 41531
rect 19349 41497 19383 41531
rect 21833 41497 21867 41531
rect 8493 41429 8527 41463
rect 9137 41429 9171 41463
rect 9505 41429 9539 41463
rect 10333 41429 10367 41463
rect 10701 41429 10735 41463
rect 10793 41429 10827 41463
rect 13369 41429 13403 41463
rect 14657 41429 14691 41463
rect 15209 41429 15243 41463
rect 16405 41429 16439 41463
rect 16773 41429 16807 41463
rect 18153 41429 18187 41463
rect 18521 41429 18555 41463
rect 19625 41429 19659 41463
rect 19993 41429 20027 41463
rect 21741 41429 21775 41463
rect 23029 41429 23063 41463
rect 23857 41429 23891 41463
rect 3617 41225 3651 41259
rect 4721 41225 4755 41259
rect 10793 41225 10827 41259
rect 11069 41225 11103 41259
rect 13185 41225 13219 41259
rect 19809 41225 19843 41259
rect 22017 41225 22051 41259
rect 24593 41225 24627 41259
rect 11713 41157 11747 41191
rect 16129 41157 16163 41191
rect 19717 41157 19751 41191
rect 20453 41157 20487 41191
rect 1777 41089 1811 41123
rect 2053 41089 2087 41123
rect 3525 41089 3559 41123
rect 3985 41089 4019 41123
rect 4629 41089 4663 41123
rect 7941 41089 7975 41123
rect 12541 41089 12575 41123
rect 13829 41089 13863 41123
rect 15945 41089 15979 41123
rect 16957 41089 16991 41123
rect 21097 41089 21131 41123
rect 22845 41089 22879 41123
rect 25329 41089 25363 41123
rect 9045 41021 9079 41055
rect 9321 41021 9355 41055
rect 14105 41021 14139 41055
rect 17233 41021 17267 41055
rect 19901 41021 19935 41055
rect 21189 41021 21223 41055
rect 21373 41021 21407 41055
rect 23121 41021 23155 41055
rect 15577 40953 15611 40987
rect 1593 40885 1627 40919
rect 5089 40885 5123 40919
rect 8585 40885 8619 40919
rect 11345 40885 11379 40919
rect 13001 40885 13035 40919
rect 18705 40885 18739 40919
rect 18981 40885 19015 40919
rect 19349 40885 19383 40919
rect 20729 40885 20763 40919
rect 22569 40885 22603 40919
rect 25145 40885 25179 40919
rect 8677 40681 8711 40715
rect 10425 40681 10459 40715
rect 14289 40681 14323 40715
rect 16129 40681 16163 40715
rect 18613 40681 18647 40715
rect 20913 40681 20947 40715
rect 23857 40681 23891 40715
rect 8217 40613 8251 40647
rect 10885 40613 10919 40647
rect 11437 40613 11471 40647
rect 13737 40613 13771 40647
rect 16773 40613 16807 40647
rect 6745 40545 6779 40579
rect 11989 40545 12023 40579
rect 13093 40545 13127 40579
rect 13277 40545 13311 40579
rect 14841 40545 14875 40579
rect 17233 40545 17267 40579
rect 17325 40545 17359 40579
rect 21465 40545 21499 40579
rect 22937 40545 22971 40579
rect 23121 40545 23155 40579
rect 6469 40477 6503 40511
rect 9873 40477 9907 40511
rect 11805 40477 11839 40511
rect 13001 40477 13035 40511
rect 14749 40477 14783 40511
rect 15485 40477 15519 40511
rect 17969 40477 18003 40511
rect 21373 40477 21407 40511
rect 22845 40477 22879 40511
rect 23581 40477 23615 40511
rect 24041 40477 24075 40511
rect 24593 40477 24627 40511
rect 9137 40409 9171 40443
rect 21925 40409 21959 40443
rect 8493 40341 8527 40375
rect 10609 40341 10643 40375
rect 11069 40341 11103 40375
rect 11897 40341 11931 40375
rect 12633 40341 12667 40375
rect 14657 40341 14691 40375
rect 17141 40341 17175 40375
rect 21281 40341 21315 40375
rect 22201 40341 22235 40375
rect 22477 40341 22511 40375
rect 25237 40341 25271 40375
rect 7481 40137 7515 40171
rect 7849 40137 7883 40171
rect 11713 40137 11747 40171
rect 12081 40137 12115 40171
rect 14749 40137 14783 40171
rect 15577 40137 15611 40171
rect 18245 40137 18279 40171
rect 19901 40137 19935 40171
rect 20637 40137 20671 40171
rect 21005 40137 21039 40171
rect 22109 40137 22143 40171
rect 22385 40137 22419 40171
rect 25145 40137 25179 40171
rect 6837 40069 6871 40103
rect 8953 40069 8987 40103
rect 10701 40069 10735 40103
rect 15945 40069 15979 40103
rect 18613 40069 18647 40103
rect 7941 40001 7975 40035
rect 11161 40001 11195 40035
rect 15117 40001 15151 40035
rect 16037 40001 16071 40035
rect 16865 40001 16899 40035
rect 19809 40001 19843 40035
rect 22293 40001 22327 40035
rect 8033 39933 8067 39967
rect 8677 39933 8711 39967
rect 12173 39933 12207 39967
rect 12265 39933 12299 39967
rect 13001 39933 13035 39967
rect 13277 39933 13311 39967
rect 16129 39933 16163 39967
rect 18705 39933 18739 39967
rect 18889 39933 18923 39967
rect 20085 39933 20119 39967
rect 21097 39933 21131 39967
rect 21281 39933 21315 39967
rect 23397 39933 23431 39967
rect 23673 39933 23707 39967
rect 17509 39865 17543 39899
rect 19441 39865 19475 39899
rect 11345 39797 11379 39831
rect 21925 39797 21959 39831
rect 22845 39797 22879 39831
rect 23121 39797 23155 39831
rect 8125 39593 8159 39627
rect 8493 39593 8527 39627
rect 9781 39593 9815 39627
rect 11240 39593 11274 39627
rect 12725 39593 12759 39627
rect 14473 39593 14507 39627
rect 21373 39593 21407 39627
rect 15669 39525 15703 39559
rect 20453 39525 20487 39559
rect 6929 39457 6963 39491
rect 10241 39457 10275 39491
rect 10333 39457 10367 39491
rect 10977 39457 11011 39491
rect 15117 39457 15151 39491
rect 16313 39457 16347 39491
rect 19993 39457 20027 39491
rect 21833 39457 21867 39491
rect 21925 39457 21959 39491
rect 23213 39457 23247 39491
rect 25053 39457 25087 39491
rect 25145 39457 25179 39491
rect 5181 39389 5215 39423
rect 7481 39389 7515 39423
rect 13369 39389 13403 39423
rect 17693 39389 17727 39423
rect 19901 39389 19935 39423
rect 23029 39389 23063 39423
rect 5457 39321 5491 39355
rect 8677 39321 8711 39355
rect 10149 39321 10183 39355
rect 14933 39321 14967 39355
rect 16129 39321 16163 39355
rect 21741 39321 21775 39355
rect 22937 39321 22971 39355
rect 23765 39321 23799 39355
rect 24961 39321 24995 39355
rect 9137 39253 9171 39287
rect 13093 39253 13127 39287
rect 13553 39253 13587 39287
rect 14105 39253 14139 39287
rect 14841 39253 14875 39287
rect 16037 39253 16071 39287
rect 18337 39253 18371 39287
rect 19441 39253 19475 39287
rect 19809 39253 19843 39287
rect 22569 39253 22603 39287
rect 24593 39253 24627 39287
rect 6009 39049 6043 39083
rect 6561 39049 6595 39083
rect 9505 39049 9539 39083
rect 10425 39049 10459 39083
rect 12265 39049 12299 39083
rect 12725 39049 12759 39083
rect 18613 39049 18647 39083
rect 19441 39049 19475 39083
rect 21005 39049 21039 39083
rect 21097 39049 21131 39083
rect 21925 39049 21959 39083
rect 22109 39049 22143 39083
rect 25237 39049 25271 39083
rect 17141 38981 17175 39015
rect 18889 38981 18923 39015
rect 19809 38981 19843 39015
rect 5365 38913 5399 38947
rect 6929 38913 6963 38947
rect 7757 38913 7791 38947
rect 10793 38913 10827 38947
rect 12633 38913 12667 38947
rect 13461 38913 13495 38947
rect 15301 38913 15335 38947
rect 16865 38913 16899 38947
rect 24593 38913 24627 38947
rect 7021 38845 7055 38879
rect 7113 38845 7147 38879
rect 9597 38845 9631 38879
rect 9781 38845 9815 38879
rect 10885 38845 10919 38879
rect 10977 38845 11011 38879
rect 12817 38845 12851 38879
rect 15393 38845 15427 38879
rect 15577 38845 15611 38879
rect 19901 38845 19935 38879
rect 19993 38845 20027 38879
rect 21281 38845 21315 38879
rect 22385 38845 22419 38879
rect 22661 38845 22695 38879
rect 9137 38777 9171 38811
rect 8401 38709 8435 38743
rect 8861 38709 8895 38743
rect 14105 38709 14139 38743
rect 14933 38709 14967 38743
rect 15945 38709 15979 38743
rect 20637 38709 20671 38743
rect 24133 38709 24167 38743
rect 7665 38505 7699 38539
rect 10425 38505 10459 38539
rect 12252 38505 12286 38539
rect 16221 38505 16255 38539
rect 17417 38505 17451 38539
rect 18797 38505 18831 38539
rect 13737 38437 13771 38471
rect 15853 38437 15887 38471
rect 24133 38437 24167 38471
rect 24593 38437 24627 38471
rect 5457 38369 5491 38403
rect 8217 38369 8251 38403
rect 9689 38369 9723 38403
rect 9781 38369 9815 38403
rect 10977 38369 11011 38403
rect 11989 38369 12023 38403
rect 14289 38369 14323 38403
rect 16681 38369 16715 38403
rect 16865 38369 16899 38403
rect 17969 38369 18003 38403
rect 18429 38369 18463 38403
rect 23213 38369 23247 38403
rect 23305 38369 23339 38403
rect 25145 38369 25179 38403
rect 1777 38301 1811 38335
rect 2053 38301 2087 38335
rect 8677 38301 8711 38335
rect 10793 38301 10827 38335
rect 18613 38301 18647 38335
rect 19441 38301 19475 38335
rect 21005 38301 21039 38335
rect 21373 38301 21407 38335
rect 23121 38301 23155 38335
rect 24961 38301 24995 38335
rect 25053 38301 25087 38335
rect 5733 38233 5767 38267
rect 9597 38233 9631 38267
rect 17785 38233 17819 38267
rect 20177 38233 20211 38267
rect 22201 38233 22235 38267
rect 24041 38233 24075 38267
rect 1593 38165 1627 38199
rect 7205 38165 7239 38199
rect 8033 38165 8067 38199
rect 8125 38165 8159 38199
rect 9229 38165 9263 38199
rect 10885 38165 10919 38199
rect 15393 38165 15427 38199
rect 16589 38165 16623 38199
rect 17877 38165 17911 38199
rect 18981 38165 19015 38199
rect 22753 38165 22787 38199
rect 23857 38165 23891 38199
rect 6009 37961 6043 37995
rect 9413 37961 9447 37995
rect 11345 37961 11379 37995
rect 11713 37961 11747 37995
rect 13921 37961 13955 37995
rect 15393 37961 15427 37995
rect 16865 37961 16899 37995
rect 17509 37961 17543 37995
rect 18337 37961 18371 37995
rect 21097 37961 21131 37995
rect 22017 37961 22051 37995
rect 22385 37961 22419 37995
rect 23029 37961 23063 37995
rect 6837 37893 6871 37927
rect 8861 37893 8895 37927
rect 10425 37893 10459 37927
rect 10701 37893 10735 37927
rect 21005 37893 21039 37927
rect 22477 37893 22511 37927
rect 23305 37893 23339 37927
rect 5365 37825 5399 37859
rect 9045 37825 9079 37859
rect 9781 37825 9815 37859
rect 9873 37825 9907 37859
rect 12909 37825 12943 37859
rect 13829 37825 13863 37859
rect 18429 37825 18463 37859
rect 19533 37825 19567 37859
rect 19625 37825 19659 37859
rect 20269 37825 20303 37859
rect 6561 37757 6595 37791
rect 8585 37757 8619 37791
rect 9965 37757 9999 37791
rect 13001 37757 13035 37791
rect 13185 37757 13219 37791
rect 15485 37757 15519 37791
rect 15669 37757 15703 37791
rect 18521 37757 18555 37791
rect 19809 37757 19843 37791
rect 21189 37757 21223 37791
rect 22661 37757 22695 37791
rect 23581 37757 23615 37791
rect 23857 37757 23891 37791
rect 15025 37689 15059 37723
rect 17969 37689 18003 37723
rect 19165 37689 19199 37723
rect 12265 37621 12299 37655
rect 12541 37621 12575 37655
rect 13553 37621 13587 37655
rect 14657 37621 14691 37655
rect 17417 37621 17451 37655
rect 20637 37621 20671 37655
rect 25329 37621 25363 37655
rect 6193 37417 6227 37451
rect 8585 37417 8619 37451
rect 9689 37417 9723 37451
rect 11069 37417 11103 37451
rect 19349 37417 19383 37451
rect 21281 37417 21315 37451
rect 22753 37417 22787 37451
rect 24041 37417 24075 37451
rect 9965 37349 9999 37383
rect 4353 37281 4387 37315
rect 6837 37281 6871 37315
rect 7113 37281 7147 37315
rect 10609 37281 10643 37315
rect 11897 37281 11931 37315
rect 13139 37281 13173 37315
rect 13921 37281 13955 37315
rect 15485 37281 15519 37315
rect 16589 37281 16623 37315
rect 16681 37281 16715 37315
rect 17785 37281 17819 37315
rect 17877 37281 17911 37315
rect 20729 37281 20763 37315
rect 22201 37281 22235 37315
rect 4077 37213 4111 37247
rect 11713 37213 11747 37247
rect 11805 37213 11839 37247
rect 15301 37213 15335 37247
rect 17693 37213 17727 37247
rect 20545 37213 20579 37247
rect 20637 37213 20671 37247
rect 21925 37213 21959 37247
rect 22937 37213 22971 37247
rect 23397 37213 23431 37247
rect 24593 37213 24627 37247
rect 25237 37213 25271 37247
rect 9137 37145 9171 37179
rect 10333 37145 10367 37179
rect 10425 37145 10459 37179
rect 13001 37145 13035 37179
rect 16497 37145 16531 37179
rect 18981 37145 19015 37179
rect 5825 37077 5859 37111
rect 11345 37077 11379 37111
rect 12541 37077 12575 37111
rect 12909 37077 12943 37111
rect 13553 37077 13587 37111
rect 14289 37077 14323 37111
rect 14933 37077 14967 37111
rect 15393 37077 15427 37111
rect 16129 37077 16163 37111
rect 17325 37077 17359 37111
rect 18521 37077 18555 37111
rect 20177 37077 20211 37111
rect 21557 37077 21591 37111
rect 22017 37077 22051 37111
rect 7297 36873 7331 36907
rect 10425 36873 10459 36907
rect 13001 36873 13035 36907
rect 13369 36873 13403 36907
rect 14933 36873 14967 36907
rect 17049 36873 17083 36907
rect 17417 36873 17451 36907
rect 19993 36873 20027 36907
rect 22201 36873 22235 36907
rect 24593 36873 24627 36907
rect 9137 36805 9171 36839
rect 11529 36805 11563 36839
rect 13461 36805 13495 36839
rect 21925 36805 21959 36839
rect 11897 36737 11931 36771
rect 14841 36737 14875 36771
rect 16681 36737 16715 36771
rect 17509 36737 17543 36771
rect 18245 36737 18279 36771
rect 20361 36737 20395 36771
rect 20453 36737 20487 36771
rect 22385 36737 22419 36771
rect 25329 36737 25363 36771
rect 9873 36669 9907 36703
rect 13645 36669 13679 36703
rect 15117 36669 15151 36703
rect 17693 36669 17727 36703
rect 20637 36669 20671 36703
rect 22845 36669 22879 36703
rect 23121 36669 23155 36703
rect 25145 36601 25179 36635
rect 7205 36533 7239 36567
rect 8677 36533 8711 36567
rect 12541 36533 12575 36567
rect 14197 36533 14231 36567
rect 14473 36533 14507 36567
rect 15485 36533 15519 36567
rect 18889 36533 18923 36567
rect 19625 36533 19659 36567
rect 21097 36533 21131 36567
rect 7021 36329 7055 36363
rect 7297 36329 7331 36363
rect 7757 36329 7791 36363
rect 9137 36329 9171 36363
rect 10793 36329 10827 36363
rect 11069 36329 11103 36363
rect 11253 36329 11287 36363
rect 12909 36329 12943 36363
rect 14289 36329 14323 36363
rect 16221 36329 16255 36363
rect 19441 36261 19475 36295
rect 23305 36261 23339 36295
rect 5273 36193 5307 36227
rect 8309 36193 8343 36227
rect 9689 36193 9723 36227
rect 13461 36193 13495 36227
rect 14933 36193 14967 36227
rect 16865 36193 16899 36227
rect 19901 36193 19935 36227
rect 19993 36193 20027 36227
rect 21373 36193 21407 36227
rect 21465 36193 21499 36227
rect 23949 36193 23983 36227
rect 1777 36125 1811 36159
rect 2053 36125 2087 36159
rect 9597 36125 9631 36159
rect 11529 36125 11563 36159
rect 19073 36125 19107 36159
rect 23765 36125 23799 36159
rect 25329 36125 25363 36159
rect 5549 36057 5583 36091
rect 8217 36057 8251 36091
rect 9505 36057 9539 36091
rect 12265 36057 12299 36091
rect 14657 36057 14691 36091
rect 15485 36057 15519 36091
rect 16589 36057 16623 36091
rect 17417 36057 17451 36091
rect 19809 36057 19843 36091
rect 1593 35989 1627 36023
rect 8125 35989 8159 36023
rect 13277 35989 13311 36023
rect 13369 35989 13403 36023
rect 14749 35989 14783 36023
rect 16681 35989 16715 36023
rect 20913 35989 20947 36023
rect 21281 35989 21315 36023
rect 22661 35989 22695 36023
rect 23673 35989 23707 36023
rect 24409 35989 24443 36023
rect 24685 35989 24719 36023
rect 24869 35989 24903 36023
rect 25145 35989 25179 36023
rect 6009 35785 6043 35819
rect 6469 35785 6503 35819
rect 9873 35785 9907 35819
rect 14105 35785 14139 35819
rect 14933 35785 14967 35819
rect 20361 35785 20395 35819
rect 22385 35785 22419 35819
rect 24961 35785 24995 35819
rect 13829 35717 13863 35751
rect 20269 35717 20303 35751
rect 4261 35649 4295 35683
rect 7021 35649 7055 35683
rect 11713 35649 11747 35683
rect 14841 35649 14875 35683
rect 17693 35649 17727 35683
rect 23213 35649 23247 35683
rect 4537 35581 4571 35615
rect 8125 35581 8159 35615
rect 8401 35581 8435 35615
rect 11989 35581 12023 35615
rect 15025 35581 15059 35615
rect 17969 35581 18003 35615
rect 19441 35581 19475 35615
rect 20453 35581 20487 35615
rect 22477 35581 22511 35615
rect 22661 35581 22695 35615
rect 23489 35581 23523 35615
rect 13461 35513 13495 35547
rect 15577 35513 15611 35547
rect 7665 35445 7699 35479
rect 10149 35445 10183 35479
rect 14473 35445 14507 35479
rect 16037 35445 16071 35479
rect 19901 35445 19935 35479
rect 21005 35445 21039 35479
rect 21281 35445 21315 35479
rect 22017 35445 22051 35479
rect 25421 35445 25455 35479
rect 8033 35241 8067 35275
rect 9137 35241 9171 35275
rect 10596 35241 10630 35275
rect 12817 35241 12851 35275
rect 14933 35241 14967 35275
rect 17233 35241 17267 35275
rect 25237 35241 25271 35275
rect 8309 35173 8343 35207
rect 6561 35105 6595 35139
rect 9689 35105 9723 35139
rect 10333 35105 10367 35139
rect 13277 35105 13311 35139
rect 13369 35105 13403 35139
rect 15485 35105 15519 35139
rect 19441 35105 19475 35139
rect 22293 35105 22327 35139
rect 5181 35037 5215 35071
rect 6285 35037 6319 35071
rect 14289 35037 14323 35071
rect 18245 35037 18279 35071
rect 24593 35037 24627 35071
rect 9505 34969 9539 35003
rect 12449 34969 12483 35003
rect 15761 34969 15795 35003
rect 18889 34969 18923 35003
rect 19717 34969 19751 35003
rect 22569 34969 22603 35003
rect 5825 34901 5859 34935
rect 9597 34901 9631 34935
rect 12081 34901 12115 34935
rect 13185 34901 13219 34935
rect 17509 34901 17543 34935
rect 21189 34901 21223 34935
rect 21649 34901 21683 34935
rect 24041 34901 24075 34935
rect 7481 34697 7515 34731
rect 9505 34697 9539 34731
rect 9873 34697 9907 34731
rect 12449 34697 12483 34731
rect 13093 34697 13127 34731
rect 13553 34697 13587 34731
rect 15577 34697 15611 34731
rect 17969 34697 18003 34731
rect 18797 34697 18831 34731
rect 18889 34697 18923 34731
rect 19441 34697 19475 34731
rect 22477 34697 22511 34731
rect 23029 34697 23063 34731
rect 15945 34629 15979 34663
rect 21097 34629 21131 34663
rect 24317 34629 24351 34663
rect 7757 34561 7791 34595
rect 11805 34561 11839 34595
rect 13461 34561 13495 34595
rect 14197 34561 14231 34595
rect 17325 34561 17359 34595
rect 21005 34561 21039 34595
rect 22385 34561 22419 34595
rect 23949 34561 23983 34595
rect 25329 34561 25363 34595
rect 13645 34493 13679 34527
rect 16037 34493 16071 34527
rect 16129 34493 16163 34527
rect 18981 34493 19015 34527
rect 19993 34493 20027 34527
rect 21189 34493 21223 34527
rect 22569 34493 22603 34527
rect 23765 34425 23799 34459
rect 8020 34357 8054 34391
rect 18429 34357 18463 34391
rect 20637 34357 20671 34391
rect 22017 34357 22051 34391
rect 25145 34357 25179 34391
rect 7849 34153 7883 34187
rect 9781 34153 9815 34187
rect 10241 34153 10275 34187
rect 17417 34153 17451 34187
rect 21833 34153 21867 34187
rect 25329 34153 25363 34187
rect 25421 34153 25455 34187
rect 13185 34085 13219 34119
rect 5825 34017 5859 34051
rect 8401 34017 8435 34051
rect 10701 34017 10735 34051
rect 10793 34017 10827 34051
rect 11437 34017 11471 34051
rect 17693 34017 17727 34051
rect 22845 34017 22879 34051
rect 23029 34017 23063 34051
rect 5549 33949 5583 33983
rect 9137 33949 9171 33983
rect 10609 33949 10643 33983
rect 13461 33949 13495 33983
rect 15669 33949 15703 33983
rect 19809 33949 19843 33983
rect 20913 33949 20947 33983
rect 22753 33949 22787 33983
rect 24777 33949 24811 33983
rect 11713 33881 11747 33915
rect 15945 33881 15979 33915
rect 21557 33881 21591 33915
rect 7297 33813 7331 33847
rect 8217 33813 8251 33847
rect 8309 33813 8343 33847
rect 19533 33813 19567 33847
rect 20453 33813 20487 33847
rect 22385 33813 22419 33847
rect 24593 33813 24627 33847
rect 7297 33609 7331 33643
rect 10517 33609 10551 33643
rect 12817 33609 12851 33643
rect 13277 33609 13311 33643
rect 20545 33609 20579 33643
rect 20913 33609 20947 33643
rect 22385 33609 22419 33643
rect 25237 33609 25271 33643
rect 12725 33541 12759 33575
rect 18613 33541 18647 33575
rect 21005 33541 21039 33575
rect 22477 33541 22511 33575
rect 1777 33473 1811 33507
rect 2053 33473 2087 33507
rect 7573 33473 7607 33507
rect 13185 33473 13219 33507
rect 14013 33473 14047 33507
rect 18337 33473 18371 33507
rect 5641 33405 5675 33439
rect 9781 33405 9815 33439
rect 13369 33405 13403 33439
rect 14289 33405 14323 33439
rect 20085 33405 20119 33439
rect 21189 33405 21223 33439
rect 22569 33405 22603 33439
rect 23489 33405 23523 33439
rect 23765 33405 23799 33439
rect 21557 33337 21591 33371
rect 1593 33269 1627 33303
rect 8217 33269 8251 33303
rect 12541 33269 12575 33303
rect 15761 33269 15795 33303
rect 16037 33269 16071 33303
rect 22017 33269 22051 33303
rect 7573 33065 7607 33099
rect 9413 33065 9447 33099
rect 10885 33065 10919 33099
rect 11897 33065 11931 33099
rect 16129 33065 16163 33099
rect 16589 33065 16623 33099
rect 17693 33065 17727 33099
rect 19533 33065 19567 33099
rect 25145 33065 25179 33099
rect 7113 32997 7147 33031
rect 14289 32997 14323 33031
rect 23029 32997 23063 33031
rect 23673 32997 23707 33031
rect 5365 32929 5399 32963
rect 8217 32929 8251 32963
rect 10057 32929 10091 32963
rect 10609 32929 10643 32963
rect 11345 32929 11379 32963
rect 11529 32929 11563 32963
rect 14749 32929 14783 32963
rect 14841 32929 14875 32963
rect 17049 32929 17083 32963
rect 17233 32929 17267 32963
rect 20177 32929 20211 32963
rect 21373 32929 21407 32963
rect 22569 32929 22603 32963
rect 23397 32929 23431 32963
rect 9781 32861 9815 32895
rect 15485 32861 15519 32895
rect 18797 32861 18831 32895
rect 21281 32861 21315 32895
rect 22385 32861 22419 32895
rect 24869 32861 24903 32895
rect 25329 32861 25363 32895
rect 5641 32793 5675 32827
rect 8033 32793 8067 32827
rect 19993 32793 20027 32827
rect 21189 32793 21223 32827
rect 7941 32725 7975 32759
rect 9873 32725 9907 32759
rect 11253 32725 11287 32759
rect 14657 32725 14691 32759
rect 16957 32725 16991 32759
rect 19073 32725 19107 32759
rect 19901 32725 19935 32759
rect 20821 32725 20855 32759
rect 22017 32725 22051 32759
rect 22477 32725 22511 32759
rect 23213 32725 23247 32759
rect 4813 32521 4847 32555
rect 5181 32521 5215 32555
rect 5549 32521 5583 32555
rect 7021 32521 7055 32555
rect 13737 32521 13771 32555
rect 14197 32521 14231 32555
rect 16129 32521 16163 32555
rect 17785 32521 17819 32555
rect 19073 32521 19107 32555
rect 5641 32453 5675 32487
rect 7941 32453 7975 32487
rect 13369 32453 13403 32487
rect 16773 32453 16807 32487
rect 20177 32453 20211 32487
rect 7665 32385 7699 32419
rect 9781 32385 9815 32419
rect 10241 32385 10275 32419
rect 14105 32385 14139 32419
rect 15485 32385 15519 32419
rect 18981 32385 19015 32419
rect 21189 32385 21223 32419
rect 22201 32385 22235 32419
rect 22845 32385 22879 32419
rect 23489 32385 23523 32419
rect 24869 32385 24903 32419
rect 25329 32385 25363 32419
rect 5825 32317 5859 32351
rect 11713 32317 11747 32351
rect 12541 32317 12575 32351
rect 14289 32317 14323 32351
rect 17877 32317 17911 32351
rect 17969 32317 18003 32351
rect 19257 32317 19291 32351
rect 20269 32317 20303 32351
rect 20453 32317 20487 32351
rect 9413 32249 9447 32283
rect 21465 32249 21499 32283
rect 25145 32249 25179 32283
rect 10885 32181 10919 32215
rect 13277 32181 13311 32215
rect 16405 32181 16439 32215
rect 17417 32181 17451 32215
rect 18613 32181 18647 32215
rect 19809 32181 19843 32215
rect 21005 32181 21039 32215
rect 22017 32181 22051 32215
rect 22661 32181 22695 32215
rect 23305 32181 23339 32215
rect 8033 31977 8067 32011
rect 8585 31977 8619 32011
rect 11253 31977 11287 32011
rect 12081 31977 12115 32011
rect 17049 31977 17083 32011
rect 19441 31977 19475 32011
rect 21005 31977 21039 32011
rect 24041 31977 24075 32011
rect 11713 31909 11747 31943
rect 17509 31909 17543 31943
rect 18705 31909 18739 31943
rect 19809 31909 19843 31943
rect 20821 31909 20855 31943
rect 22017 31909 22051 31943
rect 25145 31909 25179 31943
rect 6285 31841 6319 31875
rect 6561 31841 6595 31875
rect 8309 31841 8343 31875
rect 9505 31841 9539 31875
rect 9781 31841 9815 31875
rect 12725 31841 12759 31875
rect 18061 31841 18095 31875
rect 18889 31841 18923 31875
rect 19349 31841 19383 31875
rect 20269 31841 20303 31875
rect 20361 31841 20395 31875
rect 22477 31841 22511 31875
rect 22569 31841 22603 31875
rect 12449 31773 12483 31807
rect 15301 31773 15335 31807
rect 17969 31773 18003 31807
rect 20177 31773 20211 31807
rect 23397 31773 23431 31807
rect 24869 31773 24903 31807
rect 25329 31773 25363 31807
rect 15577 31705 15611 31739
rect 22385 31705 22419 31739
rect 11621 31637 11655 31671
rect 12541 31637 12575 31671
rect 17877 31637 17911 31671
rect 18521 31637 18555 31671
rect 7297 31433 7331 31467
rect 16313 31433 16347 31467
rect 16865 31433 16899 31467
rect 17325 31433 17359 31467
rect 19993 31433 20027 31467
rect 25145 31433 25179 31467
rect 12909 31365 12943 31399
rect 18613 31365 18647 31399
rect 19901 31365 19935 31399
rect 22385 31365 22419 31399
rect 3617 31297 3651 31331
rect 7665 31297 7699 31331
rect 8493 31297 8527 31331
rect 9413 31297 9447 31331
rect 15669 31297 15703 31331
rect 17233 31297 17267 31331
rect 18521 31297 18555 31331
rect 24501 31297 24535 31331
rect 25329 31297 25363 31331
rect 3801 31229 3835 31263
rect 4997 31229 5031 31263
rect 6837 31229 6871 31263
rect 7757 31229 7791 31263
rect 7941 31229 7975 31263
rect 9689 31229 9723 31263
rect 12633 31229 12667 31263
rect 14749 31229 14783 31263
rect 17417 31229 17451 31263
rect 18705 31229 18739 31263
rect 20085 31229 20119 31263
rect 22109 31229 22143 31263
rect 7021 31161 7055 31195
rect 11161 31161 11195 31195
rect 18153 31161 18187 31195
rect 11621 31093 11655 31127
rect 14381 31093 14415 31127
rect 19533 31093 19567 31127
rect 23857 31093 23891 31127
rect 24317 31093 24351 31127
rect 24869 31093 24903 31127
rect 7757 30889 7791 30923
rect 8953 30889 8987 30923
rect 12541 30889 12575 30923
rect 15577 30889 15611 30923
rect 22845 30889 22879 30923
rect 24869 30889 24903 30923
rect 19441 30821 19475 30855
rect 21833 30821 21867 30855
rect 8401 30753 8435 30787
rect 11989 30753 12023 30787
rect 13093 30753 13127 30787
rect 14841 30753 14875 30787
rect 17141 30753 17175 30787
rect 18889 30753 18923 30787
rect 20085 30753 20119 30787
rect 22293 30753 22327 30787
rect 22477 30753 22511 30787
rect 9689 30685 9723 30719
rect 14657 30685 14691 30719
rect 16037 30685 16071 30719
rect 22201 30685 22235 30719
rect 23949 30685 23983 30719
rect 25329 30685 25363 30719
rect 8125 30617 8159 30651
rect 12265 30617 12299 30651
rect 17417 30617 17451 30651
rect 19809 30617 19843 30651
rect 7481 30549 7515 30583
rect 8217 30549 8251 30583
rect 10333 30549 10367 30583
rect 12909 30549 12943 30583
rect 13001 30549 13035 30583
rect 14289 30549 14323 30583
rect 14749 30549 14783 30583
rect 15393 30549 15427 30583
rect 16681 30549 16715 30583
rect 19901 30549 19935 30583
rect 20453 30549 20487 30583
rect 23765 30549 23799 30583
rect 25145 30549 25179 30583
rect 25421 30345 25455 30379
rect 16773 30277 16807 30311
rect 18981 30277 19015 30311
rect 23673 30277 23707 30311
rect 8861 30209 8895 30243
rect 10793 30209 10827 30243
rect 11713 30209 11747 30243
rect 12909 30209 12943 30243
rect 14565 30209 14599 30243
rect 17785 30209 17819 30243
rect 19809 30209 19843 30243
rect 23397 30209 23431 30243
rect 10149 30141 10183 30175
rect 10885 30141 10919 30175
rect 10977 30141 11011 30175
rect 13001 30141 13035 30175
rect 13093 30141 13127 30175
rect 14841 30141 14875 30175
rect 17877 30141 17911 30175
rect 18061 30141 18095 30175
rect 10425 30073 10459 30107
rect 17049 30073 17083 30107
rect 19349 30073 19383 30107
rect 9505 30005 9539 30039
rect 12541 30005 12575 30039
rect 16313 30005 16347 30039
rect 17417 30005 17451 30039
rect 18521 30005 18555 30039
rect 19625 30005 19659 30039
rect 25145 30005 25179 30039
rect 15945 29801 15979 29835
rect 25145 29733 25179 29767
rect 3985 29665 4019 29699
rect 9689 29665 9723 29699
rect 9965 29665 9999 29699
rect 12541 29665 12575 29699
rect 17693 29665 17727 29699
rect 19993 29665 20027 29699
rect 20177 29665 20211 29699
rect 23305 29665 23339 29699
rect 23397 29665 23431 29699
rect 11897 29597 11931 29631
rect 19901 29597 19935 29631
rect 23213 29597 23247 29631
rect 25329 29597 25363 29631
rect 4169 29529 4203 29563
rect 5825 29529 5859 29563
rect 14657 29529 14691 29563
rect 17417 29529 17451 29563
rect 18245 29529 18279 29563
rect 7481 29461 7515 29495
rect 11437 29461 11471 29495
rect 12909 29461 12943 29495
rect 16773 29461 16807 29495
rect 17049 29461 17083 29495
rect 17509 29461 17543 29495
rect 19533 29461 19567 29495
rect 22845 29461 22879 29495
rect 3387 29257 3421 29291
rect 9229 29257 9263 29291
rect 9781 29257 9815 29291
rect 11069 29257 11103 29291
rect 11529 29257 11563 29291
rect 13921 29257 13955 29291
rect 15945 29257 15979 29291
rect 17233 29257 17267 29291
rect 18061 29257 18095 29291
rect 18521 29257 18555 29291
rect 22385 29257 22419 29291
rect 23949 29257 23983 29291
rect 25329 29257 25363 29291
rect 25513 29257 25547 29291
rect 12449 29189 12483 29223
rect 13093 29189 13127 29223
rect 15853 29189 15887 29223
rect 22477 29189 22511 29223
rect 24685 29189 24719 29223
rect 3284 29121 3318 29155
rect 10149 29121 10183 29155
rect 12357 29121 12391 29155
rect 13829 29121 13863 29155
rect 17325 29121 17359 29155
rect 18429 29121 18463 29155
rect 19533 29121 19567 29155
rect 20177 29121 20211 29155
rect 20821 29121 20855 29155
rect 23673 29121 23707 29155
rect 24133 29121 24167 29155
rect 7021 29053 7055 29087
rect 10241 29053 10275 29087
rect 10425 29053 10459 29087
rect 12541 29053 12575 29087
rect 14105 29053 14139 29087
rect 16037 29053 16071 29087
rect 17417 29053 17451 29087
rect 18613 29053 18647 29087
rect 20269 29053 20303 29087
rect 20453 29053 20487 29087
rect 21281 29053 21315 29087
rect 22661 29053 22695 29087
rect 8769 28985 8803 29019
rect 9505 28985 9539 29019
rect 11989 28985 12023 29019
rect 13461 28985 13495 29019
rect 15485 28985 15519 29019
rect 16865 28985 16899 29019
rect 19809 28985 19843 29019
rect 22017 28985 22051 29019
rect 24869 28985 24903 29019
rect 7284 28917 7318 28951
rect 9137 28917 9171 28951
rect 6377 28713 6411 28747
rect 7849 28713 7883 28747
rect 10885 28713 10919 28747
rect 11437 28713 11471 28747
rect 17969 28713 18003 28747
rect 21097 28713 21131 28747
rect 12633 28645 12667 28679
rect 13737 28645 13771 28679
rect 23857 28645 23891 28679
rect 3985 28577 4019 28611
rect 8401 28577 8435 28611
rect 12081 28577 12115 28611
rect 13185 28577 13219 28611
rect 14841 28577 14875 28611
rect 16773 28577 16807 28611
rect 21741 28577 21775 28611
rect 6745 28509 6779 28543
rect 9137 28509 9171 28543
rect 13001 28509 13035 28543
rect 14657 28509 14691 28543
rect 15485 28509 15519 28543
rect 16589 28509 16623 28543
rect 21465 28509 21499 28543
rect 24041 28509 24075 28543
rect 24777 28509 24811 28543
rect 4169 28441 4203 28475
rect 5825 28441 5859 28475
rect 8309 28441 8343 28475
rect 9413 28441 9447 28475
rect 11805 28441 11839 28475
rect 13093 28441 13127 28475
rect 16681 28441 16715 28475
rect 7389 28373 7423 28407
rect 8217 28373 8251 28407
rect 11897 28373 11931 28407
rect 13829 28373 13863 28407
rect 14289 28373 14323 28407
rect 14749 28373 14783 28407
rect 15301 28373 15335 28407
rect 16221 28373 16255 28407
rect 17325 28373 17359 28407
rect 17693 28373 17727 28407
rect 20729 28373 20763 28407
rect 21557 28373 21591 28407
rect 24593 28373 24627 28407
rect 8309 28169 8343 28203
rect 8677 28169 8711 28203
rect 12357 28169 12391 28203
rect 14749 28169 14783 28203
rect 17141 28169 17175 28203
rect 17785 28169 17819 28203
rect 23765 28169 23799 28203
rect 25237 28169 25271 28203
rect 6837 28101 6871 28135
rect 21189 28101 21223 28135
rect 24685 28101 24719 28135
rect 11713 28033 11747 28067
rect 15393 28033 15427 28067
rect 18613 28033 18647 28067
rect 2053 27965 2087 27999
rect 2237 27965 2271 27999
rect 2789 27965 2823 27999
rect 6561 27965 6595 27999
rect 9229 27965 9263 27999
rect 9505 27965 9539 27999
rect 10977 27965 11011 27999
rect 13001 27965 13035 27999
rect 13277 27965 13311 27999
rect 17877 27965 17911 27999
rect 18061 27965 18095 27999
rect 19165 27965 19199 27999
rect 19441 27965 19475 27999
rect 20913 27965 20947 27999
rect 22017 27965 22051 27999
rect 22293 27965 22327 27999
rect 18521 27897 18555 27931
rect 24869 27897 24903 27931
rect 11253 27829 11287 27863
rect 15117 27829 15151 27863
rect 16037 27829 16071 27863
rect 17417 27829 17451 27863
rect 24133 27829 24167 27863
rect 7757 27625 7791 27659
rect 11069 27625 11103 27659
rect 15656 27625 15690 27659
rect 13001 27557 13035 27591
rect 18981 27557 19015 27591
rect 20637 27557 20671 27591
rect 11989 27489 12023 27523
rect 13553 27489 13587 27523
rect 15393 27489 15427 27523
rect 18245 27489 18279 27523
rect 20085 27489 20119 27523
rect 21097 27489 21131 27523
rect 21281 27489 21315 27523
rect 24041 27489 24075 27523
rect 4020 27421 4054 27455
rect 6653 27421 6687 27455
rect 11897 27421 11931 27455
rect 14289 27421 14323 27455
rect 18153 27421 18187 27455
rect 19809 27421 19843 27455
rect 22293 27421 22327 27455
rect 4123 27353 4157 27387
rect 11805 27353 11839 27387
rect 13461 27353 13495 27387
rect 18061 27353 18095 27387
rect 22569 27353 22603 27387
rect 24685 27353 24719 27387
rect 24869 27353 24903 27387
rect 7297 27285 7331 27319
rect 9597 27285 9631 27319
rect 11437 27285 11471 27319
rect 12633 27285 12667 27319
rect 13369 27285 13403 27319
rect 14933 27285 14967 27319
rect 17141 27285 17175 27319
rect 17693 27285 17727 27319
rect 18705 27285 18739 27319
rect 19441 27285 19475 27319
rect 19901 27285 19935 27319
rect 21005 27285 21039 27319
rect 8677 27081 8711 27115
rect 9137 27081 9171 27115
rect 9505 27081 9539 27115
rect 15025 27081 15059 27115
rect 18521 27081 18555 27115
rect 20453 27081 20487 27115
rect 23765 27081 23799 27115
rect 6837 27013 6871 27047
rect 10701 27013 10735 27047
rect 13553 27013 13587 27047
rect 24685 27013 24719 27047
rect 3433 26945 3467 26979
rect 11713 26945 11747 26979
rect 13277 26945 13311 26979
rect 17233 26945 17267 26979
rect 18429 26945 18463 26979
rect 19441 26945 19475 26979
rect 20821 26945 20855 26979
rect 3617 26877 3651 26911
rect 5181 26877 5215 26911
rect 6561 26877 6595 26911
rect 8769 26877 8803 26911
rect 9597 26877 9631 26911
rect 9781 26877 9815 26911
rect 17325 26877 17359 26911
rect 17417 26877 17451 26911
rect 18705 26877 18739 26911
rect 19901 26877 19935 26911
rect 22017 26877 22051 26911
rect 22293 26877 22327 26911
rect 24133 26877 24167 26911
rect 25145 26877 25179 26911
rect 8309 26809 8343 26843
rect 19257 26809 19291 26843
rect 24869 26809 24903 26843
rect 10793 26741 10827 26775
rect 12357 26741 12391 26775
rect 15393 26741 15427 26775
rect 16405 26741 16439 26775
rect 16865 26741 16899 26775
rect 18061 26741 18095 26775
rect 21465 26741 21499 26775
rect 3617 26537 3651 26571
rect 4261 26537 4295 26571
rect 8217 26537 8251 26571
rect 8585 26537 8619 26571
rect 10425 26537 10459 26571
rect 13001 26537 13035 26571
rect 17693 26537 17727 26571
rect 17969 26537 18003 26571
rect 20545 26537 20579 26571
rect 20821 26537 20855 26571
rect 23949 26537 23983 26571
rect 25237 26537 25271 26571
rect 10793 26469 10827 26503
rect 14933 26469 14967 26503
rect 21005 26469 21039 26503
rect 21281 26469 21315 26503
rect 4445 26401 4479 26435
rect 6745 26401 6779 26435
rect 11253 26401 11287 26435
rect 11437 26401 11471 26435
rect 12357 26401 12391 26435
rect 13461 26401 13495 26435
rect 13645 26401 13679 26435
rect 14197 26401 14231 26435
rect 15577 26401 15611 26435
rect 19901 26401 19935 26435
rect 20085 26401 20119 26435
rect 21741 26401 21775 26435
rect 21833 26401 21867 26435
rect 22937 26401 22971 26435
rect 23121 26401 23155 26435
rect 3985 26333 4019 26367
rect 6469 26333 6503 26367
rect 9413 26333 9447 26367
rect 16129 26333 16163 26367
rect 19809 26333 19843 26367
rect 21649 26333 21683 26367
rect 23857 26333 23891 26367
rect 24593 26333 24627 26367
rect 14657 26265 14691 26299
rect 15301 26265 15335 26299
rect 15393 26265 15427 26299
rect 22845 26265 22879 26299
rect 10057 26197 10091 26231
rect 11161 26197 11195 26231
rect 13369 26197 13403 26231
rect 16773 26197 16807 26231
rect 19441 26197 19475 26231
rect 22477 26197 22511 26231
rect 3479 25993 3513 26027
rect 9505 25993 9539 26027
rect 10609 25993 10643 26027
rect 11713 25993 11747 26027
rect 13001 25993 13035 26027
rect 13093 25993 13127 26027
rect 18337 25993 18371 26027
rect 19625 25993 19659 26027
rect 19717 25993 19751 26027
rect 22569 25993 22603 26027
rect 7757 25925 7791 25959
rect 12173 25925 12207 25959
rect 14565 25925 14599 25959
rect 16313 25925 16347 25959
rect 18245 25925 18279 25959
rect 3376 25857 3410 25891
rect 3985 25857 4019 25891
rect 7481 25857 7515 25891
rect 10517 25857 10551 25891
rect 21005 25857 21039 25891
rect 21465 25857 21499 25891
rect 22477 25857 22511 25891
rect 23305 25857 23339 25891
rect 24133 25857 24167 25891
rect 3065 25789 3099 25823
rect 6837 25789 6871 25823
rect 10701 25789 10735 25823
rect 13185 25789 13219 25823
rect 14289 25789 14323 25823
rect 18521 25789 18555 25823
rect 19901 25789 19935 25823
rect 22753 25789 22787 25823
rect 25145 25789 25179 25823
rect 4445 25721 4479 25755
rect 21281 25721 21315 25755
rect 4261 25653 4295 25687
rect 9229 25653 9263 25687
rect 10149 25653 10183 25687
rect 11253 25653 11287 25687
rect 12633 25653 12667 25687
rect 16681 25653 16715 25687
rect 17877 25653 17911 25687
rect 19257 25653 19291 25687
rect 22109 25653 22143 25687
rect 4077 25449 4111 25483
rect 7481 25449 7515 25483
rect 10977 25449 11011 25483
rect 12173 25449 12207 25483
rect 23213 25449 23247 25483
rect 7113 25313 7147 25347
rect 7941 25313 7975 25347
rect 8033 25313 8067 25347
rect 9229 25313 9263 25347
rect 12633 25313 12667 25347
rect 12817 25313 12851 25347
rect 15117 25313 15151 25347
rect 17233 25313 17267 25347
rect 17417 25313 17451 25347
rect 20637 25313 20671 25347
rect 4261 25245 4295 25279
rect 4813 25245 4847 25279
rect 7849 25245 7883 25279
rect 14933 25245 14967 25279
rect 15025 25245 15059 25279
rect 20361 25245 20395 25279
rect 22569 25245 22603 25279
rect 23857 25245 23891 25279
rect 24869 25245 24903 25279
rect 9505 25177 9539 25211
rect 11529 25177 11563 25211
rect 12541 25177 12575 25211
rect 16497 25177 16531 25211
rect 17141 25177 17175 25211
rect 5457 25109 5491 25143
rect 14565 25109 14599 25143
rect 16773 25109 16807 25143
rect 22109 25109 22143 25143
rect 23949 25109 23983 25143
rect 24685 25109 24719 25143
rect 9965 24905 9999 24939
rect 11345 24905 11379 24939
rect 12265 24905 12299 24939
rect 19993 24905 20027 24939
rect 22017 24905 22051 24939
rect 25053 24905 25087 24939
rect 4261 24837 4295 24871
rect 12173 24837 12207 24871
rect 17601 24837 17635 24871
rect 23305 24837 23339 24871
rect 6561 24769 6595 24803
rect 8677 24769 8711 24803
rect 9873 24769 9907 24803
rect 10701 24769 10735 24803
rect 13369 24769 13403 24803
rect 15945 24769 15979 24803
rect 16037 24769 16071 24803
rect 17325 24769 17359 24803
rect 20085 24769 20119 24803
rect 21925 24769 21959 24803
rect 22569 24769 22603 24803
rect 1685 24701 1719 24735
rect 1869 24701 1903 24735
rect 2881 24701 2915 24735
rect 3985 24701 4019 24735
rect 5733 24701 5767 24735
rect 8033 24701 8067 24735
rect 8769 24701 8803 24735
rect 8861 24701 8895 24735
rect 10057 24701 10091 24735
rect 12357 24701 12391 24735
rect 13461 24701 13495 24735
rect 13553 24701 13587 24735
rect 14933 24701 14967 24735
rect 16221 24701 16255 24735
rect 19073 24701 19107 24735
rect 20269 24701 20303 24735
rect 23029 24701 23063 24735
rect 8309 24633 8343 24667
rect 19625 24633 19659 24667
rect 22385 24633 22419 24667
rect 6101 24565 6135 24599
rect 7205 24565 7239 24599
rect 9505 24565 9539 24599
rect 11805 24565 11839 24599
rect 13001 24565 13035 24599
rect 15577 24565 15611 24599
rect 24777 24565 24811 24599
rect 5733 24361 5767 24395
rect 6469 24361 6503 24395
rect 10333 24361 10367 24395
rect 17417 24361 17451 24395
rect 25145 24361 25179 24395
rect 6101 24293 6135 24327
rect 10517 24293 10551 24327
rect 12725 24293 12759 24327
rect 19993 24293 20027 24327
rect 7113 24225 7147 24259
rect 9137 24225 9171 24259
rect 10977 24225 11011 24259
rect 11253 24225 11287 24259
rect 14933 24225 14967 24259
rect 15669 24225 15703 24259
rect 20453 24225 20487 24259
rect 20545 24225 20579 24259
rect 21925 24225 21959 24259
rect 22017 24225 22051 24259
rect 23857 24225 23891 24259
rect 2237 24157 2271 24191
rect 3985 24157 4019 24191
rect 13185 24157 13219 24191
rect 14289 24157 14323 24191
rect 17877 24157 17911 24191
rect 19625 24157 19659 24191
rect 21833 24157 21867 24191
rect 22845 24157 22879 24191
rect 24685 24157 24719 24191
rect 4261 24089 4295 24123
rect 10149 24089 10183 24123
rect 13001 24089 13035 24123
rect 15945 24089 15979 24123
rect 18521 24089 18555 24123
rect 2053 24021 2087 24055
rect 6837 24021 6871 24055
rect 6929 24021 6963 24055
rect 13461 24021 13495 24055
rect 18797 24021 18831 24055
rect 19257 24021 19291 24055
rect 20361 24021 20395 24055
rect 21465 24021 21499 24055
rect 24777 24021 24811 24055
rect 3847 23817 3881 23851
rect 5549 23817 5583 23851
rect 8309 23817 8343 23851
rect 8585 23817 8619 23851
rect 9689 23817 9723 23851
rect 10885 23817 10919 23851
rect 12541 23817 12575 23851
rect 13737 23817 13771 23851
rect 14381 23817 14415 23851
rect 14657 23817 14691 23851
rect 15025 23817 15059 23851
rect 15393 23817 15427 23851
rect 15761 23817 15795 23851
rect 17233 23817 17267 23851
rect 17325 23817 17359 23851
rect 18061 23817 18095 23851
rect 21465 23817 21499 23851
rect 21833 23817 21867 23851
rect 24593 23817 24627 23851
rect 6837 23749 6871 23783
rect 13829 23749 13863 23783
rect 15853 23749 15887 23783
rect 19993 23749 20027 23783
rect 23121 23749 23155 23783
rect 25145 23749 25179 23783
rect 3744 23681 3778 23715
rect 4905 23681 4939 23715
rect 9597 23681 9631 23715
rect 10793 23681 10827 23715
rect 12633 23681 12667 23715
rect 18245 23681 18279 23715
rect 22845 23681 22879 23715
rect 6561 23613 6595 23647
rect 9873 23613 9907 23647
rect 10977 23613 11011 23647
rect 11805 23613 11839 23647
rect 12725 23613 12759 23647
rect 13921 23613 13955 23647
rect 16037 23613 16071 23647
rect 17417 23613 17451 23647
rect 18981 23613 19015 23647
rect 19717 23613 19751 23647
rect 25329 23613 25363 23647
rect 9229 23545 9263 23579
rect 10425 23545 10459 23579
rect 13369 23545 13403 23579
rect 11621 23477 11655 23511
rect 12173 23477 12207 23511
rect 16865 23477 16899 23511
rect 8033 23273 8067 23307
rect 8401 23273 8435 23307
rect 18889 23273 18923 23307
rect 21189 23273 21223 23307
rect 21557 23273 21591 23307
rect 11713 23205 11747 23239
rect 14289 23205 14323 23239
rect 1593 23137 1627 23171
rect 2973 23137 3007 23171
rect 6285 23137 6319 23171
rect 11069 23137 11103 23171
rect 11989 23137 12023 23171
rect 14749 23137 14783 23171
rect 14841 23137 14875 23171
rect 17141 23137 17175 23171
rect 17417 23137 17451 23171
rect 19441 23137 19475 23171
rect 22017 23137 22051 23171
rect 25053 23137 25087 23171
rect 25145 23137 25179 23171
rect 4261 23069 4295 23103
rect 9597 23069 9631 23103
rect 22845 23069 22879 23103
rect 23857 23069 23891 23103
rect 24961 23069 24995 23103
rect 1777 23001 1811 23035
rect 6561 23001 6595 23035
rect 10241 23001 10275 23035
rect 12265 23001 12299 23035
rect 14657 23001 14691 23035
rect 19717 23001 19751 23035
rect 4905 22933 4939 22967
rect 11437 22933 11471 22967
rect 13737 22933 13771 22967
rect 15393 22933 15427 22967
rect 24593 22933 24627 22967
rect 4813 22729 4847 22763
rect 10149 22729 10183 22763
rect 10793 22729 10827 22763
rect 12541 22729 12575 22763
rect 13829 22729 13863 22763
rect 13921 22729 13955 22763
rect 17693 22729 17727 22763
rect 24593 22729 24627 22763
rect 25145 22729 25179 22763
rect 3985 22661 4019 22695
rect 8217 22661 8251 22695
rect 9413 22661 9447 22695
rect 10885 22661 10919 22695
rect 11713 22661 11747 22695
rect 18797 22661 18831 22695
rect 4353 22593 4387 22627
rect 7113 22593 7147 22627
rect 8953 22593 8987 22627
rect 13001 22593 13035 22627
rect 14657 22593 14691 22627
rect 16313 22593 16347 22627
rect 18061 22593 18095 22627
rect 19441 22593 19475 22627
rect 20547 22593 20581 22627
rect 24777 22593 24811 22627
rect 10977 22525 11011 22559
rect 14105 22525 14139 22559
rect 21281 22525 21315 22559
rect 22109 22525 22143 22559
rect 22385 22525 22419 22559
rect 24133 22525 24167 22559
rect 13461 22457 13495 22491
rect 4629 22389 4663 22423
rect 7757 22389 7791 22423
rect 10425 22389 10459 22423
rect 12817 22389 12851 22423
rect 15301 22389 15335 22423
rect 16129 22389 16163 22423
rect 20085 22389 20119 22423
rect 4432 22185 4466 22219
rect 20821 22185 20855 22219
rect 25145 22185 25179 22219
rect 14749 22117 14783 22151
rect 4169 22049 4203 22083
rect 5917 22049 5951 22083
rect 8125 22049 8159 22083
rect 9689 22049 9723 22083
rect 10793 22049 10827 22083
rect 11621 22049 11655 22083
rect 11713 22049 11747 22083
rect 13093 22049 13127 22083
rect 13553 22049 13587 22083
rect 14197 22049 14231 22083
rect 15209 22049 15243 22083
rect 15301 22049 15335 22083
rect 16497 22049 16531 22083
rect 17877 22049 17911 22083
rect 18061 22049 18095 22083
rect 20085 22049 20119 22083
rect 22845 22049 22879 22083
rect 24041 22049 24075 22083
rect 2237 21981 2271 22015
rect 3341 21981 3375 22015
rect 7941 21981 7975 22015
rect 9505 21981 9539 22015
rect 12909 21981 12943 22015
rect 19441 21981 19475 22015
rect 21097 21981 21131 22015
rect 23397 21981 23431 22015
rect 8033 21913 8067 21947
rect 16313 21913 16347 21947
rect 20545 21913 20579 21947
rect 21373 21913 21407 21947
rect 24685 21913 24719 21947
rect 2053 21845 2087 21879
rect 3157 21845 3191 21879
rect 6193 21845 6227 21879
rect 7573 21845 7607 21879
rect 8677 21845 8711 21879
rect 9137 21845 9171 21879
rect 9597 21845 9631 21879
rect 11161 21845 11195 21879
rect 11529 21845 11563 21879
rect 12449 21845 12483 21879
rect 12817 21845 12851 21879
rect 14381 21845 14415 21879
rect 15117 21845 15151 21879
rect 15945 21845 15979 21879
rect 16405 21845 16439 21879
rect 17417 21845 17451 21879
rect 17785 21845 17819 21879
rect 18613 21845 18647 21879
rect 20453 21845 20487 21879
rect 24777 21845 24811 21879
rect 5181 21641 5215 21675
rect 5549 21641 5583 21675
rect 6653 21641 6687 21675
rect 7021 21641 7055 21675
rect 10793 21641 10827 21675
rect 12909 21641 12943 21675
rect 14289 21641 14323 21675
rect 14657 21641 14691 21675
rect 17141 21641 17175 21675
rect 17601 21641 17635 21675
rect 20085 21641 20119 21675
rect 21189 21641 21223 21675
rect 22477 21641 22511 21675
rect 24961 21641 24995 21675
rect 8125 21573 8159 21607
rect 9873 21573 9907 21607
rect 15393 21573 15427 21607
rect 25237 21573 25271 21607
rect 1869 21505 1903 21539
rect 5641 21505 5675 21539
rect 7849 21505 7883 21539
rect 10885 21505 10919 21539
rect 16129 21505 16163 21539
rect 17509 21505 17543 21539
rect 20545 21505 20579 21539
rect 22385 21505 22419 21539
rect 23213 21505 23247 21539
rect 2053 21437 2087 21471
rect 2881 21437 2915 21471
rect 5825 21437 5859 21471
rect 7113 21437 7147 21471
rect 7205 21437 7239 21471
rect 10977 21437 11011 21471
rect 12081 21437 12115 21471
rect 14749 21437 14783 21471
rect 14841 21437 14875 21471
rect 17785 21437 17819 21471
rect 18337 21437 18371 21471
rect 18613 21437 18647 21471
rect 22661 21437 22695 21471
rect 23489 21437 23523 21471
rect 12265 21369 12299 21403
rect 10425 21301 10459 21335
rect 13921 21301 13955 21335
rect 15669 21301 15703 21335
rect 16865 21301 16899 21335
rect 22017 21301 22051 21335
rect 7021 21097 7055 21131
rect 8585 21097 8619 21131
rect 9137 21097 9171 21131
rect 16037 21097 16071 21131
rect 21925 21097 21959 21131
rect 17325 21029 17359 21063
rect 2053 20961 2087 20995
rect 4169 20961 4203 20995
rect 4445 20961 4479 20995
rect 9689 20961 9723 20995
rect 11805 20961 11839 20995
rect 14565 20961 14599 20995
rect 16957 20961 16991 20995
rect 17785 20961 17819 20995
rect 17969 20961 18003 20995
rect 19901 20961 19935 20995
rect 23857 20961 23891 20995
rect 1777 20893 1811 20927
rect 6377 20893 6411 20927
rect 7941 20893 7975 20927
rect 9597 20893 9631 20927
rect 11621 20893 11655 20927
rect 14289 20893 14323 20927
rect 16681 20893 16715 20927
rect 17693 20893 17727 20927
rect 18705 20893 18739 20927
rect 22845 20893 22879 20927
rect 9505 20825 9539 20859
rect 20177 20825 20211 20859
rect 5917 20757 5951 20791
rect 10241 20757 10275 20791
rect 11253 20757 11287 20791
rect 11713 20757 11747 20791
rect 16497 20757 16531 20791
rect 18521 20757 18555 20791
rect 21649 20757 21683 20791
rect 3341 20553 3375 20587
rect 4169 20553 4203 20587
rect 8217 20553 8251 20587
rect 8585 20553 8619 20587
rect 9321 20553 9355 20587
rect 12173 20553 12207 20587
rect 12817 20553 12851 20587
rect 15025 20553 15059 20587
rect 18245 20553 18279 20587
rect 19349 20553 19383 20587
rect 21281 20553 21315 20587
rect 9413 20485 9447 20519
rect 17693 20485 17727 20519
rect 23305 20485 23339 20519
rect 3525 20417 3559 20451
rect 4353 20417 4387 20451
rect 7113 20417 7147 20451
rect 8677 20417 8711 20451
rect 10977 20417 11011 20451
rect 12081 20417 12115 20451
rect 13277 20417 13311 20451
rect 15485 20417 15519 20451
rect 17049 20417 17083 20451
rect 19257 20417 19291 20451
rect 20637 20417 20671 20451
rect 22293 20417 22327 20451
rect 24133 20417 24167 20451
rect 8861 20349 8895 20383
rect 12265 20349 12299 20383
rect 13553 20349 13587 20383
rect 16129 20349 16163 20383
rect 19533 20349 19567 20383
rect 24409 20349 24443 20383
rect 11713 20281 11747 20315
rect 16865 20281 16899 20315
rect 6101 20213 6135 20247
rect 7757 20213 7791 20247
rect 17785 20213 17819 20247
rect 18889 20213 18923 20247
rect 7849 20009 7883 20043
rect 10609 20009 10643 20043
rect 11253 20009 11287 20043
rect 18981 20009 19015 20043
rect 7389 19941 7423 19975
rect 9137 19941 9171 19975
rect 10425 19941 10459 19975
rect 15117 19941 15151 19975
rect 17969 19941 18003 19975
rect 5365 19873 5399 19907
rect 5641 19873 5675 19907
rect 8401 19873 8435 19907
rect 9689 19873 9723 19907
rect 11805 19873 11839 19907
rect 23857 19873 23891 19907
rect 8217 19805 8251 19839
rect 9505 19805 9539 19839
rect 9597 19805 9631 19839
rect 13001 19805 13035 19839
rect 15853 19805 15887 19839
rect 17049 19805 17083 19839
rect 17785 19805 17819 19839
rect 18613 19805 18647 19839
rect 20453 19805 20487 19839
rect 21557 19805 21591 19839
rect 22845 19805 22879 19839
rect 8309 19737 8343 19771
rect 11621 19737 11655 19771
rect 16037 19737 16071 19771
rect 20637 19737 20671 19771
rect 24685 19737 24719 19771
rect 7113 19669 7147 19703
rect 10241 19669 10275 19703
rect 11713 19669 11747 19703
rect 13645 19669 13679 19703
rect 16865 19669 16899 19703
rect 18429 19669 18463 19703
rect 22201 19669 22235 19703
rect 24777 19669 24811 19703
rect 10425 19465 10459 19499
rect 10885 19465 10919 19499
rect 12173 19465 12207 19499
rect 13277 19465 13311 19499
rect 23765 19465 23799 19499
rect 2145 19397 2179 19431
rect 10793 19397 10827 19431
rect 13645 19397 13679 19431
rect 8125 19329 8159 19363
rect 12081 19329 12115 19363
rect 17693 19329 17727 19363
rect 18337 19329 18371 19363
rect 18981 19329 19015 19363
rect 8401 19261 8435 19295
rect 10977 19261 11011 19295
rect 12265 19261 12299 19295
rect 13001 19261 13035 19295
rect 13737 19261 13771 19295
rect 13829 19261 13863 19295
rect 19257 19261 19291 19295
rect 21189 19261 21223 19295
rect 22017 19261 22051 19295
rect 22293 19261 22327 19295
rect 24041 19261 24075 19295
rect 24225 19261 24259 19295
rect 14473 19193 14507 19227
rect 2237 19125 2271 19159
rect 6837 19125 6871 19159
rect 7665 19125 7699 19159
rect 9873 19125 9907 19159
rect 11713 19125 11747 19159
rect 12725 19125 12759 19159
rect 14381 19125 14415 19159
rect 14749 19125 14783 19159
rect 17509 19125 17543 19159
rect 18153 19125 18187 19159
rect 20729 19125 20763 19159
rect 7205 18921 7239 18955
rect 10885 18921 10919 18955
rect 13001 18921 13035 18955
rect 14289 18921 14323 18955
rect 16497 18921 16531 18955
rect 16865 18921 16899 18955
rect 24041 18921 24075 18955
rect 7389 18853 7423 18887
rect 11805 18853 11839 18887
rect 21097 18853 21131 18887
rect 2053 18785 2087 18819
rect 9137 18785 9171 18819
rect 12357 18785 12391 18819
rect 13461 18785 13495 18819
rect 13645 18785 13679 18819
rect 14841 18785 14875 18819
rect 17417 18785 17451 18819
rect 21557 18785 21591 18819
rect 21649 18785 21683 18819
rect 22569 18785 22603 18819
rect 25237 18785 25271 18819
rect 1777 18717 1811 18751
rect 5825 18717 5859 18751
rect 6929 18717 6963 18751
rect 7941 18717 7975 18751
rect 11437 18717 11471 18751
rect 14657 18717 14691 18751
rect 17233 18717 17267 18751
rect 18705 18717 18739 18751
rect 19349 18717 19383 18751
rect 19809 18717 19843 18751
rect 22293 18717 22327 18751
rect 24593 18717 24627 18751
rect 9413 18649 9447 18683
rect 12173 18649 12207 18683
rect 17325 18649 17359 18683
rect 17877 18649 17911 18683
rect 18889 18649 18923 18683
rect 21465 18649 21499 18683
rect 6469 18581 6503 18615
rect 8585 18581 8619 18615
rect 11253 18581 11287 18615
rect 12265 18581 12299 18615
rect 13369 18581 13403 18615
rect 14749 18581 14783 18615
rect 20453 18581 20487 18615
rect 5273 18377 5307 18411
rect 5641 18377 5675 18411
rect 9505 18377 9539 18411
rect 10057 18377 10091 18411
rect 10425 18377 10459 18411
rect 10793 18377 10827 18411
rect 12817 18377 12851 18411
rect 13185 18377 13219 18411
rect 13277 18377 13311 18411
rect 14013 18377 14047 18411
rect 14381 18377 14415 18411
rect 15117 18377 15151 18411
rect 19993 18377 20027 18411
rect 6837 18309 6871 18343
rect 8585 18309 8619 18343
rect 12357 18309 12391 18343
rect 12541 18309 12575 18343
rect 20177 18309 20211 18343
rect 20453 18309 20487 18343
rect 9413 18241 9447 18275
rect 10885 18241 10919 18275
rect 22293 18241 22327 18275
rect 24133 18241 24167 18275
rect 5733 18173 5767 18207
rect 5917 18173 5951 18207
rect 6561 18173 6595 18207
rect 9597 18173 9631 18207
rect 10977 18173 11011 18207
rect 13461 18173 13495 18207
rect 14473 18173 14507 18207
rect 14657 18173 14691 18207
rect 17877 18173 17911 18207
rect 18153 18173 18187 18207
rect 21281 18173 21315 18207
rect 23305 18173 23339 18207
rect 24777 18173 24811 18207
rect 19625 18105 19659 18139
rect 9045 18037 9079 18071
rect 6561 17833 6595 17867
rect 7113 17833 7147 17867
rect 10425 17833 10459 17867
rect 17509 17833 17543 17867
rect 19349 17833 19383 17867
rect 21465 17833 21499 17867
rect 23673 17833 23707 17867
rect 23949 17765 23983 17799
rect 7573 17697 7607 17731
rect 7757 17697 7791 17731
rect 8401 17697 8435 17731
rect 11069 17697 11103 17731
rect 11345 17697 11379 17731
rect 19717 17697 19751 17731
rect 22201 17697 22235 17731
rect 4813 17629 4847 17663
rect 7481 17629 7515 17663
rect 9137 17629 9171 17663
rect 15577 17629 15611 17663
rect 16221 17629 16255 17663
rect 16865 17629 16899 17663
rect 17969 17629 18003 17663
rect 21925 17629 21959 17663
rect 5089 17561 5123 17595
rect 9873 17561 9907 17595
rect 18705 17561 18739 17595
rect 19993 17561 20027 17595
rect 10517 17493 10551 17527
rect 12817 17493 12851 17527
rect 13185 17493 13219 17527
rect 13829 17493 13863 17527
rect 15393 17493 15427 17527
rect 16313 17493 16347 17527
rect 6009 17289 6043 17323
rect 6745 17289 6779 17323
rect 7481 17289 7515 17323
rect 7849 17289 7883 17323
rect 9873 17289 9907 17323
rect 10333 17289 10367 17323
rect 13093 17289 13127 17323
rect 16037 17289 16071 17323
rect 21281 17289 21315 17323
rect 2237 17221 2271 17255
rect 12449 17221 12483 17255
rect 13461 17221 13495 17255
rect 19533 17221 19567 17255
rect 20085 17221 20119 17255
rect 21557 17221 21591 17255
rect 23213 17221 23247 17255
rect 5365 17153 5399 17187
rect 9045 17153 9079 17187
rect 9137 17153 9171 17187
rect 10241 17153 10275 17187
rect 11713 17153 11747 17187
rect 15945 17153 15979 17187
rect 16865 17153 16899 17187
rect 19441 17153 19475 17187
rect 20637 17153 20671 17187
rect 22017 17153 22051 17187
rect 23949 17153 23983 17187
rect 7941 17085 7975 17119
rect 8033 17085 8067 17119
rect 9321 17085 9355 17119
rect 10425 17085 10459 17119
rect 13553 17085 13587 17119
rect 13645 17085 13679 17119
rect 16129 17085 16163 17119
rect 17141 17085 17175 17119
rect 19717 17085 19751 17119
rect 24685 17085 24719 17119
rect 8677 17017 8711 17051
rect 10977 17017 11011 17051
rect 23397 17017 23431 17051
rect 2329 16949 2363 16983
rect 15209 16949 15243 16983
rect 15577 16949 15611 16983
rect 18613 16949 18647 16983
rect 19073 16949 19107 16983
rect 22661 16949 22695 16983
rect 6272 16745 6306 16779
rect 8493 16745 8527 16779
rect 12725 16745 12759 16779
rect 12909 16745 12943 16779
rect 16405 16745 16439 16779
rect 19349 16745 19383 16779
rect 21189 16745 21223 16779
rect 6009 16609 6043 16643
rect 7757 16609 7791 16643
rect 9781 16609 9815 16643
rect 10885 16609 10919 16643
rect 14841 16609 14875 16643
rect 15577 16609 15611 16643
rect 15669 16609 15703 16643
rect 18889 16609 18923 16643
rect 20545 16609 20579 16643
rect 21741 16609 21775 16643
rect 22017 16609 22051 16643
rect 23765 16609 23799 16643
rect 1777 16541 1811 16575
rect 9505 16541 9539 16575
rect 10701 16541 10735 16575
rect 11529 16541 11563 16575
rect 17969 16541 18003 16575
rect 18613 16541 18647 16575
rect 20361 16541 20395 16575
rect 2513 16473 2547 16507
rect 12173 16473 12207 16507
rect 21097 16473 21131 16507
rect 8125 16405 8159 16439
rect 8677 16405 8711 16439
rect 9137 16405 9171 16439
rect 9597 16405 9631 16439
rect 10333 16405 10367 16439
rect 10793 16405 10827 16439
rect 15117 16405 15151 16439
rect 15485 16405 15519 16439
rect 16221 16405 16255 16439
rect 19625 16405 19659 16439
rect 23489 16405 23523 16439
rect 7021 16201 7055 16235
rect 7389 16201 7423 16235
rect 9597 16201 9631 16235
rect 10057 16201 10091 16235
rect 16221 16201 16255 16235
rect 17233 16201 17267 16235
rect 18797 16201 18831 16235
rect 19165 16201 19199 16235
rect 19533 16201 19567 16235
rect 20821 16201 20855 16235
rect 7481 16133 7515 16167
rect 12081 16133 12115 16167
rect 15669 16133 15703 16167
rect 19625 16133 19659 16167
rect 8217 16065 8251 16099
rect 9965 16065 9999 16099
rect 20729 16065 20763 16099
rect 22385 16065 22419 16099
rect 23213 16065 23247 16099
rect 24133 16065 24167 16099
rect 7665 15997 7699 16031
rect 10241 15997 10275 16031
rect 11805 15997 11839 16031
rect 19809 15997 19843 16031
rect 21005 15997 21039 16031
rect 22477 15997 22511 16031
rect 22661 15997 22695 16031
rect 24777 15997 24811 16031
rect 9229 15929 9263 15963
rect 15853 15929 15887 15963
rect 18613 15929 18647 15963
rect 8861 15861 8895 15895
rect 13553 15861 13587 15895
rect 14013 15861 14047 15895
rect 17509 15861 17543 15895
rect 17877 15861 17911 15895
rect 20361 15861 20395 15895
rect 22017 15861 22051 15895
rect 8493 15657 8527 15691
rect 13001 15657 13035 15691
rect 15025 15657 15059 15691
rect 17417 15657 17451 15691
rect 14105 15589 14139 15623
rect 18981 15589 19015 15623
rect 19441 15589 19475 15623
rect 7021 15521 7055 15555
rect 10241 15521 10275 15555
rect 12725 15521 12759 15555
rect 13553 15521 13587 15555
rect 18429 15521 18463 15555
rect 18613 15521 18647 15555
rect 19901 15521 19935 15555
rect 20085 15521 20119 15555
rect 21281 15521 21315 15555
rect 6745 15453 6779 15487
rect 9137 15453 9171 15487
rect 12541 15453 12575 15487
rect 13461 15453 13495 15487
rect 14565 15453 14599 15487
rect 15669 15453 15703 15487
rect 19809 15453 19843 15487
rect 20821 15453 20855 15487
rect 22109 15453 22143 15487
rect 22753 15453 22787 15487
rect 24593 15453 24627 15487
rect 10517 15385 10551 15419
rect 13369 15385 13403 15419
rect 15945 15385 15979 15419
rect 23857 15385 23891 15419
rect 9781 15317 9815 15351
rect 11989 15317 12023 15351
rect 14657 15317 14691 15351
rect 17969 15317 18003 15351
rect 18337 15317 18371 15351
rect 20637 15317 20671 15351
rect 21925 15317 21959 15351
rect 25237 15317 25271 15351
rect 11805 15113 11839 15147
rect 13001 15113 13035 15147
rect 13369 15113 13403 15147
rect 14565 15113 14599 15147
rect 14657 15113 14691 15147
rect 15301 15113 15335 15147
rect 16313 15113 16347 15147
rect 18061 15113 18095 15147
rect 20545 15113 20579 15147
rect 21465 15113 21499 15147
rect 7757 15045 7791 15079
rect 8401 15045 8435 15079
rect 10149 15045 10183 15079
rect 16957 15045 16991 15079
rect 23305 15045 23339 15079
rect 10517 14977 10551 15011
rect 12173 14977 12207 15011
rect 15669 14977 15703 15011
rect 17969 14977 18003 15011
rect 21189 14977 21223 15011
rect 22569 14977 22603 15011
rect 24133 14977 24167 15011
rect 8125 14909 8159 14943
rect 12265 14909 12299 14943
rect 12357 14909 12391 14943
rect 13461 14909 13495 14943
rect 13553 14909 13587 14943
rect 14749 14909 14783 14943
rect 18245 14909 18279 14943
rect 18797 14909 18831 14943
rect 19073 14909 19107 14943
rect 24685 14909 24719 14943
rect 14197 14841 14231 14875
rect 22753 14841 22787 14875
rect 23489 14841 23523 14875
rect 17049 14773 17083 14807
rect 17601 14773 17635 14807
rect 21005 14773 21039 14807
rect 8585 14569 8619 14603
rect 13001 14569 13035 14603
rect 14841 14569 14875 14603
rect 17049 14569 17083 14603
rect 20269 14501 20303 14535
rect 10057 14433 10091 14467
rect 12173 14433 12207 14467
rect 12357 14433 12391 14467
rect 13553 14433 13587 14467
rect 19441 14433 19475 14467
rect 21281 14433 21315 14467
rect 7941 14365 7975 14399
rect 13369 14365 13403 14399
rect 15301 14365 15335 14399
rect 17601 14365 17635 14399
rect 18429 14365 18463 14399
rect 18889 14365 18923 14399
rect 21005 14365 21039 14399
rect 10333 14297 10367 14331
rect 12725 14297 12759 14331
rect 14381 14297 14415 14331
rect 15577 14297 15611 14331
rect 18613 14297 18647 14331
rect 23029 14297 23063 14331
rect 11805 14229 11839 14263
rect 13461 14229 13495 14263
rect 14473 14229 14507 14263
rect 17693 14229 17727 14263
rect 22753 14229 22787 14263
rect 9873 14025 9907 14059
rect 10241 14025 10275 14059
rect 12081 14025 12115 14059
rect 12449 14025 12483 14059
rect 12909 14025 12943 14059
rect 13829 14025 13863 14059
rect 14933 14025 14967 14059
rect 17509 14025 17543 14059
rect 19165 14025 19199 14059
rect 20085 14025 20119 14059
rect 23029 14025 23063 14059
rect 17969 13957 18003 13991
rect 20545 13957 20579 13991
rect 25145 13957 25179 13991
rect 1777 13889 1811 13923
rect 12817 13889 12851 13923
rect 13461 13889 13495 13923
rect 14381 13889 14415 13923
rect 16313 13889 16347 13923
rect 16865 13889 16899 13923
rect 18521 13889 18555 13923
rect 20453 13889 20487 13923
rect 21281 13889 21315 13923
rect 23213 13889 23247 13923
rect 23949 13889 23983 13923
rect 2053 13821 2087 13855
rect 8125 13821 8159 13855
rect 8401 13821 8435 13855
rect 13001 13821 13035 13855
rect 14565 13821 14599 13855
rect 20637 13821 20671 13855
rect 16129 13753 16163 13787
rect 17785 13685 17819 13719
rect 12265 13481 12299 13515
rect 17693 13481 17727 13515
rect 16497 13413 16531 13447
rect 18797 13413 18831 13447
rect 10793 13345 10827 13379
rect 10977 13345 11011 13379
rect 16957 13345 16991 13379
rect 17049 13345 17083 13379
rect 18153 13345 18187 13379
rect 18337 13345 18371 13379
rect 11621 13277 11655 13311
rect 14289 13277 14323 13311
rect 15485 13277 15519 13311
rect 15945 13277 15979 13311
rect 19533 13277 19567 13311
rect 20269 13277 20303 13311
rect 20729 13277 20763 13311
rect 21097 13277 21131 13311
rect 22661 13277 22695 13311
rect 10701 13209 10735 13243
rect 13553 13209 13587 13243
rect 15669 13209 15703 13243
rect 18061 13209 18095 13243
rect 19717 13209 19751 13243
rect 20453 13209 20487 13243
rect 23857 13209 23891 13243
rect 10333 13141 10367 13175
rect 13645 13141 13679 13175
rect 14933 13141 14967 13175
rect 16865 13141 16899 13175
rect 21741 13141 21775 13175
rect 10609 12937 10643 12971
rect 13369 12937 13403 12971
rect 13829 12937 13863 12971
rect 19625 12937 19659 12971
rect 19901 12937 19935 12971
rect 21189 12937 21223 12971
rect 9137 12869 9171 12903
rect 13093 12869 13127 12903
rect 16957 12869 16991 12903
rect 21097 12869 21131 12903
rect 22753 12869 22787 12903
rect 11713 12801 11747 12835
rect 13737 12801 13771 12835
rect 14565 12801 14599 12835
rect 17877 12801 17911 12835
rect 22109 12801 22143 12835
rect 23213 12801 23247 12835
rect 23949 12801 23983 12835
rect 8861 12733 8895 12767
rect 10885 12733 10919 12767
rect 13921 12733 13955 12767
rect 14841 12733 14875 12767
rect 16313 12733 16347 12767
rect 18153 12733 18187 12767
rect 21373 12733 21407 12767
rect 24777 12733 24811 12767
rect 12357 12597 12391 12631
rect 17509 12597 17543 12631
rect 20177 12597 20211 12631
rect 20729 12597 20763 12631
rect 22201 12597 22235 12631
rect 11345 12393 11379 12427
rect 15209 12393 15243 12427
rect 16405 12393 16439 12427
rect 21373 12393 21407 12427
rect 22661 12325 22695 12359
rect 9597 12257 9631 12291
rect 12081 12257 12115 12291
rect 13553 12257 13587 12291
rect 15853 12257 15887 12291
rect 16957 12257 16991 12291
rect 19625 12257 19659 12291
rect 11805 12189 11839 12223
rect 14381 12189 14415 12223
rect 14841 12189 14875 12223
rect 18245 12189 18279 12223
rect 22017 12189 22051 12223
rect 22845 12189 22879 12223
rect 23489 12189 23523 12223
rect 9873 12121 9907 12155
rect 16773 12121 16807 12155
rect 19901 12121 19935 12155
rect 13829 12053 13863 12087
rect 14473 12053 14507 12087
rect 15577 12053 15611 12087
rect 15669 12053 15703 12087
rect 16865 12053 16899 12087
rect 17601 12053 17635 12087
rect 18889 12053 18923 12087
rect 21833 12053 21867 12087
rect 22385 12053 22419 12087
rect 23305 12053 23339 12087
rect 10885 11849 10919 11883
rect 14749 11849 14783 11883
rect 15577 11849 15611 11883
rect 20821 11849 20855 11883
rect 21189 11849 21223 11883
rect 15669 11781 15703 11815
rect 16221 11781 16255 11815
rect 25145 11781 25179 11815
rect 10241 11713 10275 11747
rect 13001 11713 13035 11747
rect 17969 11713 18003 11747
rect 20177 11713 20211 11747
rect 23949 11713 23983 11747
rect 11529 11645 11563 11679
rect 13277 11645 13311 11679
rect 15761 11645 15795 11679
rect 18245 11645 18279 11679
rect 15209 11577 15243 11611
rect 16405 11509 16439 11543
rect 19717 11509 19751 11543
rect 15485 11305 15519 11339
rect 16681 11305 16715 11339
rect 17141 11237 17175 11271
rect 20177 11237 20211 11271
rect 21189 11237 21223 11271
rect 23213 11237 23247 11271
rect 18889 11169 18923 11203
rect 14841 11101 14875 11135
rect 16037 11101 16071 11135
rect 16865 11101 16899 11135
rect 18429 11101 18463 11135
rect 20361 11101 20395 11135
rect 21741 11101 21775 11135
rect 23397 11101 23431 11135
rect 16221 11033 16255 11067
rect 18613 11033 18647 11067
rect 21005 11033 21039 11067
rect 21925 11033 21959 11067
rect 19533 10965 19567 10999
rect 19533 10761 19567 10795
rect 19625 10761 19659 10795
rect 21281 10761 21315 10795
rect 11989 10693 12023 10727
rect 12449 10693 12483 10727
rect 18521 10625 18555 10659
rect 22937 10625 22971 10659
rect 23949 10625 23983 10659
rect 19717 10557 19751 10591
rect 24777 10557 24811 10591
rect 12173 10489 12207 10523
rect 18337 10489 18371 10523
rect 19165 10421 19199 10455
rect 22753 10421 22787 10455
rect 14565 10013 14599 10047
rect 16865 10013 16899 10047
rect 22201 10013 22235 10047
rect 22661 10013 22695 10047
rect 24869 10013 24903 10047
rect 14749 9945 14783 9979
rect 23857 9945 23891 9979
rect 16957 9877 16991 9911
rect 22017 9877 22051 9911
rect 24685 9877 24719 9911
rect 22477 9673 22511 9707
rect 16957 9605 16991 9639
rect 18889 9605 18923 9639
rect 22661 9537 22695 9571
rect 23397 9537 23431 9571
rect 23949 9537 23983 9571
rect 7573 9469 7607 9503
rect 24685 9469 24719 9503
rect 17141 9401 17175 9435
rect 19073 9401 19107 9435
rect 23213 9333 23247 9367
rect 7113 9129 7147 9163
rect 7757 8993 7791 9027
rect 7481 8925 7515 8959
rect 23857 8925 23891 8959
rect 24869 8925 24903 8959
rect 7573 8857 7607 8891
rect 23949 8789 23983 8823
rect 24685 8789 24719 8823
rect 6377 8517 6411 8551
rect 18889 8517 18923 8551
rect 20821 8517 20855 8551
rect 25145 8517 25179 8551
rect 3985 8449 4019 8483
rect 6009 8449 6043 8483
rect 22293 8449 22327 8483
rect 23949 8449 23983 8483
rect 4261 8381 4295 8415
rect 22753 8381 22787 8415
rect 19073 8313 19107 8347
rect 21005 8313 21039 8347
rect 23305 7905 23339 7939
rect 20637 7837 20671 7871
rect 21649 7837 21683 7871
rect 22845 7837 22879 7871
rect 20453 7701 20487 7735
rect 21465 7701 21499 7735
rect 18521 7429 18555 7463
rect 19441 7429 19475 7463
rect 25145 7429 25179 7463
rect 20269 7361 20303 7395
rect 22109 7361 22143 7395
rect 23949 7361 23983 7395
rect 21281 7293 21315 7327
rect 22569 7293 22603 7327
rect 19625 7225 19659 7259
rect 18613 7157 18647 7191
rect 20269 6749 20303 6783
rect 20821 6749 20855 6783
rect 22845 6749 22879 6783
rect 22017 6681 22051 6715
rect 23857 6681 23891 6715
rect 20085 6613 20119 6647
rect 17969 6409 18003 6443
rect 18245 6273 18279 6307
rect 20269 6273 20303 6307
rect 22201 6273 22235 6307
rect 23949 6273 23983 6307
rect 19257 6205 19291 6239
rect 21281 6205 21315 6239
rect 22477 6205 22511 6239
rect 24777 6205 24811 6239
rect 24777 5865 24811 5899
rect 21005 5729 21039 5763
rect 22845 5729 22879 5763
rect 20545 5661 20579 5695
rect 22385 5661 22419 5695
rect 24685 5593 24719 5627
rect 18797 5253 18831 5287
rect 17785 5185 17819 5219
rect 19441 5185 19475 5219
rect 22109 5185 22143 5219
rect 23949 5185 23983 5219
rect 19901 5117 19935 5151
rect 22477 5117 22511 5151
rect 24777 5117 24811 5151
rect 24777 4777 24811 4811
rect 19901 4641 19935 4675
rect 21741 4641 21775 4675
rect 23213 4641 23247 4675
rect 23489 4641 23523 4675
rect 17693 4573 17727 4607
rect 19441 4573 19475 4607
rect 21281 4573 21315 4607
rect 24685 4573 24719 4607
rect 18613 4505 18647 4539
rect 1777 4097 1811 4131
rect 11989 4097 12023 4131
rect 13553 4097 13587 4131
rect 16129 4097 16163 4131
rect 16313 4097 16347 4131
rect 16865 4097 16899 4131
rect 18889 4097 18923 4131
rect 22017 4097 22051 4131
rect 23857 4097 23891 4131
rect 11345 4029 11379 4063
rect 11713 4029 11747 4063
rect 14013 4029 14047 4063
rect 17325 4029 17359 4063
rect 19165 4029 19199 4063
rect 22477 4029 22511 4063
rect 24317 4029 24351 4063
rect 1593 3961 1627 3995
rect 9965 3961 9999 3995
rect 2053 3893 2087 3927
rect 6377 3893 6411 3927
rect 9505 3893 9539 3927
rect 9781 3893 9815 3927
rect 11069 3893 11103 3927
rect 5273 3689 5307 3723
rect 6745 3689 6779 3723
rect 8217 3689 8251 3723
rect 9321 3689 9355 3723
rect 10057 3689 10091 3723
rect 1777 3621 1811 3655
rect 5917 3621 5951 3655
rect 7573 3553 7607 3587
rect 12817 3553 12851 3587
rect 15485 3553 15519 3587
rect 17325 3553 17359 3587
rect 19901 3553 19935 3587
rect 21741 3553 21775 3587
rect 1961 3485 1995 3519
rect 2421 3485 2455 3519
rect 5089 3485 5123 3519
rect 6101 3485 6135 3519
rect 6561 3485 6595 3519
rect 8033 3485 8067 3519
rect 9137 3485 9171 3519
rect 9873 3485 9907 3519
rect 10517 3485 10551 3519
rect 10977 3485 11011 3519
rect 11253 3485 11287 3519
rect 12541 3485 12575 3519
rect 15117 3485 15151 3519
rect 16865 3485 16899 3519
rect 19441 3485 19475 3519
rect 21281 3485 21315 3519
rect 3157 3417 3191 3451
rect 2237 3349 2271 3383
rect 2881 3349 2915 3383
rect 3249 3349 3283 3383
rect 3617 3349 3651 3383
rect 4813 3349 4847 3383
rect 7205 3349 7239 3383
rect 7757 3349 7791 3383
rect 8677 3349 8711 3383
rect 10701 3349 10735 3383
rect 25421 3349 25455 3383
rect 2697 3145 2731 3179
rect 5181 3145 5215 3179
rect 5917 3145 5951 3179
rect 7021 3145 7055 3179
rect 7757 3145 7791 3179
rect 8493 3145 8527 3179
rect 11897 3145 11931 3179
rect 24869 3145 24903 3179
rect 23581 3077 23615 3111
rect 1869 3009 1903 3043
rect 2513 3009 2547 3043
rect 4721 3009 4755 3043
rect 4997 3009 5031 3043
rect 5733 3009 5767 3043
rect 6837 3009 6871 3043
rect 7573 3009 7607 3043
rect 8309 3009 8343 3043
rect 9321 3009 9355 3043
rect 10609 3009 10643 3043
rect 11713 3009 11747 3043
rect 12633 3009 12667 3043
rect 14289 3009 14323 3043
rect 16865 3009 16899 3043
rect 18705 3009 18739 3043
rect 3249 2941 3283 2975
rect 3525 2941 3559 2975
rect 9045 2941 9079 2975
rect 10333 2941 10367 2975
rect 13369 2941 13403 2975
rect 14749 2941 14783 2975
rect 17325 2941 17359 2975
rect 19165 2941 19199 2975
rect 2053 2873 2087 2907
rect 1501 2805 1535 2839
rect 4353 2805 4387 2839
rect 6469 2805 6503 2839
rect 1869 2601 1903 2635
rect 2605 2601 2639 2635
rect 3341 2601 3375 2635
rect 7113 2601 7147 2635
rect 9781 2601 9815 2635
rect 11713 2601 11747 2635
rect 4169 2533 4203 2567
rect 4997 2465 5031 2499
rect 7941 2465 7975 2499
rect 10609 2465 10643 2499
rect 14105 2465 14139 2499
rect 15209 2465 15243 2499
rect 17325 2465 17359 2499
rect 18521 2465 18555 2499
rect 19901 2465 19935 2499
rect 22477 2465 22511 2499
rect 1685 2397 1719 2431
rect 2421 2397 2455 2431
rect 3985 2397 4019 2431
rect 4721 2397 4755 2431
rect 5825 2397 5859 2431
rect 6469 2397 6503 2431
rect 6929 2397 6963 2431
rect 7665 2397 7699 2431
rect 9137 2397 9171 2431
rect 9597 2397 9631 2431
rect 10333 2397 10367 2431
rect 11897 2397 11931 2431
rect 12541 2397 12575 2431
rect 14657 2397 14691 2431
rect 16957 2397 16991 2431
rect 19441 2397 19475 2431
rect 22017 2397 22051 2431
rect 25329 2397 25363 2431
rect 3249 2329 3283 2363
rect 6101 2329 6135 2363
rect 6653 2329 6687 2363
rect 9321 2329 9355 2363
rect 13553 2329 13587 2363
<< metal1 >>
rect 1104 54426 25852 54448
rect 1104 54374 7950 54426
rect 8002 54374 8014 54426
rect 8066 54374 8078 54426
rect 8130 54374 8142 54426
rect 8194 54374 8206 54426
rect 8258 54374 17950 54426
rect 18002 54374 18014 54426
rect 18066 54374 18078 54426
rect 18130 54374 18142 54426
rect 18194 54374 18206 54426
rect 18258 54374 25852 54426
rect 1104 54352 25852 54374
rect 9950 54272 9956 54324
rect 10008 54272 10014 54324
rect 14553 54315 14611 54321
rect 14553 54281 14565 54315
rect 14599 54312 14611 54315
rect 14734 54312 14740 54324
rect 14599 54284 14740 54312
rect 14599 54281 14611 54284
rect 14553 54275 14611 54281
rect 14734 54272 14740 54284
rect 14792 54272 14798 54324
rect 16206 54272 16212 54324
rect 16264 54312 16270 54324
rect 16393 54315 16451 54321
rect 16393 54312 16405 54315
rect 16264 54284 16405 54312
rect 16264 54272 16270 54284
rect 16393 54281 16405 54284
rect 16439 54312 16451 54315
rect 16439 54284 16574 54312
rect 16439 54281 16451 54284
rect 16393 54275 16451 54281
rect 5813 54247 5871 54253
rect 5813 54213 5825 54247
rect 5859 54244 5871 54247
rect 7834 54244 7840 54256
rect 5859 54216 7840 54244
rect 5859 54213 5871 54216
rect 5813 54207 5871 54213
rect 7834 54204 7840 54216
rect 7892 54204 7898 54256
rect 8389 54247 8447 54253
rect 8389 54213 8401 54247
rect 8435 54244 8447 54247
rect 9968 54244 9996 54272
rect 8435 54216 9996 54244
rect 10965 54247 11023 54253
rect 8435 54213 8447 54216
rect 8389 54207 8447 54213
rect 10965 54213 10977 54247
rect 11011 54244 11023 54247
rect 11422 54244 11428 54256
rect 11011 54216 11428 54244
rect 11011 54213 11023 54216
rect 10965 54207 11023 54213
rect 11422 54204 11428 54216
rect 11480 54204 11486 54256
rect 12894 54244 12900 54256
rect 11900 54216 12900 54244
rect 2225 54179 2283 54185
rect 2225 54145 2237 54179
rect 2271 54176 2283 54179
rect 4338 54176 4344 54188
rect 2271 54148 4344 54176
rect 2271 54145 2283 54148
rect 2225 54139 2283 54145
rect 4338 54136 4344 54148
rect 4396 54136 4402 54188
rect 4614 54136 4620 54188
rect 4672 54136 4678 54188
rect 7377 54179 7435 54185
rect 7377 54145 7389 54179
rect 7423 54145 7435 54179
rect 7377 54139 7435 54145
rect 3237 54111 3295 54117
rect 3237 54077 3249 54111
rect 3283 54108 3295 54111
rect 5902 54108 5908 54120
rect 3283 54080 5908 54108
rect 3283 54077 3295 54080
rect 3237 54071 3295 54077
rect 5902 54068 5908 54080
rect 5960 54068 5966 54120
rect 7392 54108 7420 54139
rect 9950 54136 9956 54188
rect 10008 54136 10014 54188
rect 11900 54185 11928 54216
rect 12894 54204 12900 54216
rect 12952 54244 12958 54256
rect 14093 54247 14151 54253
rect 14093 54244 14105 54247
rect 12952 54216 14105 54244
rect 12952 54204 12958 54216
rect 14093 54213 14105 54216
rect 14139 54213 14151 54247
rect 14093 54207 14151 54213
rect 11885 54179 11943 54185
rect 11885 54145 11897 54179
rect 11931 54145 11943 54179
rect 11885 54139 11943 54145
rect 12342 54136 12348 54188
rect 12400 54136 12406 54188
rect 14752 54176 14780 54272
rect 14829 54179 14887 54185
rect 14829 54176 14841 54179
rect 14752 54148 14841 54176
rect 14829 54145 14841 54148
rect 14875 54145 14887 54179
rect 14829 54139 14887 54145
rect 15194 54136 15200 54188
rect 15252 54176 15258 54188
rect 15565 54179 15623 54185
rect 15565 54176 15577 54179
rect 15252 54148 15577 54176
rect 15252 54136 15258 54148
rect 15565 54145 15577 54148
rect 15611 54176 15623 54179
rect 16117 54179 16175 54185
rect 16117 54176 16129 54179
rect 15611 54148 16129 54176
rect 15611 54145 15623 54148
rect 15565 54139 15623 54145
rect 16117 54145 16129 54148
rect 16163 54145 16175 54179
rect 16546 54176 16574 54284
rect 24486 54272 24492 54324
rect 24544 54272 24550 54324
rect 24670 54272 24676 54324
rect 24728 54272 24734 54324
rect 17678 54204 17684 54256
rect 17736 54244 17742 54256
rect 18417 54247 18475 54253
rect 18417 54244 18429 54247
rect 17736 54216 18429 54244
rect 17736 54204 17742 54216
rect 18417 54213 18429 54216
rect 18463 54244 18475 54247
rect 18874 54244 18880 54256
rect 18463 54216 18880 54244
rect 18463 54213 18475 54216
rect 18417 54207 18475 54213
rect 18874 54204 18880 54216
rect 18932 54204 18938 54256
rect 21453 54247 21511 54253
rect 21453 54244 21465 54247
rect 20180 54216 21465 54244
rect 16853 54179 16911 54185
rect 16853 54176 16865 54179
rect 16546 54148 16865 54176
rect 16117 54139 16175 54145
rect 16853 54145 16865 54148
rect 16899 54145 16911 54179
rect 16853 54139 16911 54145
rect 16942 54136 16948 54188
rect 17000 54176 17006 54188
rect 17589 54179 17647 54185
rect 17589 54176 17601 54179
rect 17000 54148 17601 54176
rect 17000 54136 17006 54148
rect 17589 54145 17601 54148
rect 17635 54176 17647 54179
rect 18969 54179 19027 54185
rect 18969 54176 18981 54179
rect 17635 54148 18981 54176
rect 17635 54145 17647 54148
rect 17589 54139 17647 54145
rect 18969 54145 18981 54148
rect 19015 54145 19027 54179
rect 18969 54139 19027 54145
rect 19429 54179 19487 54185
rect 19429 54145 19441 54179
rect 19475 54145 19487 54179
rect 19429 54139 19487 54145
rect 10226 54108 10232 54120
rect 7392 54080 10232 54108
rect 10226 54068 10232 54080
rect 10284 54068 10290 54120
rect 12526 54068 12532 54120
rect 12584 54108 12590 54120
rect 12805 54111 12863 54117
rect 12805 54108 12817 54111
rect 12584 54080 12817 54108
rect 12584 54068 12590 54080
rect 12805 54077 12817 54080
rect 12851 54077 12863 54111
rect 12805 54071 12863 54077
rect 18414 54068 18420 54120
rect 18472 54108 18478 54120
rect 19444 54108 19472 54139
rect 19518 54136 19524 54188
rect 19576 54176 19582 54188
rect 20180 54185 20208 54216
rect 21453 54213 21465 54216
rect 21499 54213 21511 54247
rect 23293 54247 23351 54253
rect 23293 54244 23305 54247
rect 21453 54207 21511 54213
rect 22020 54216 23305 54244
rect 20165 54179 20223 54185
rect 20165 54176 20177 54179
rect 19576 54148 20177 54176
rect 19576 54136 19582 54148
rect 20165 54145 20177 54148
rect 20211 54145 20223 54179
rect 20165 54139 20223 54145
rect 20714 54136 20720 54188
rect 20772 54176 20778 54188
rect 20901 54179 20959 54185
rect 20901 54176 20913 54179
rect 20772 54148 20913 54176
rect 20772 54136 20778 54148
rect 20901 54145 20913 54148
rect 20947 54145 20959 54179
rect 20901 54139 20959 54145
rect 21358 54136 21364 54188
rect 21416 54176 21422 54188
rect 22020 54185 22048 54216
rect 23293 54213 23305 54216
rect 23339 54213 23351 54247
rect 23293 54207 23351 54213
rect 22005 54179 22063 54185
rect 22005 54176 22017 54179
rect 21416 54148 22017 54176
rect 21416 54136 21422 54148
rect 22005 54145 22017 54148
rect 22051 54145 22063 54179
rect 22005 54139 22063 54145
rect 22462 54136 22468 54188
rect 22520 54176 22526 54188
rect 22741 54179 22799 54185
rect 22741 54176 22753 54179
rect 22520 54148 22753 54176
rect 22520 54136 22526 54148
rect 22741 54145 22753 54148
rect 22787 54145 22799 54179
rect 22741 54139 22799 54145
rect 23753 54179 23811 54185
rect 23753 54145 23765 54179
rect 23799 54176 23811 54179
rect 24688 54176 24716 54272
rect 23799 54148 24716 54176
rect 23799 54145 23811 54148
rect 23753 54139 23811 54145
rect 25038 54136 25044 54188
rect 25096 54136 25102 54188
rect 19702 54108 19708 54120
rect 18472 54080 19708 54108
rect 18472 54068 18478 54080
rect 19702 54068 19708 54080
rect 19760 54068 19766 54120
rect 15013 54043 15071 54049
rect 15013 54009 15025 54043
rect 15059 54040 15071 54043
rect 16206 54040 16212 54052
rect 15059 54012 16212 54040
rect 15059 54009 15071 54012
rect 15013 54003 15071 54009
rect 16206 54000 16212 54012
rect 16264 54000 16270 54052
rect 17773 54043 17831 54049
rect 17773 54040 17785 54043
rect 16546 54012 17785 54040
rect 11698 53932 11704 53984
rect 11756 53932 11762 53984
rect 15746 53932 15752 53984
rect 15804 53932 15810 53984
rect 16114 53932 16120 53984
rect 16172 53972 16178 53984
rect 16546 53972 16574 54012
rect 17773 54009 17785 54012
rect 17819 54009 17831 54043
rect 17773 54003 17831 54009
rect 19334 54000 19340 54052
rect 19392 54040 19398 54052
rect 20349 54043 20407 54049
rect 20349 54040 20361 54043
rect 19392 54012 20361 54040
rect 19392 54000 19398 54012
rect 20349 54009 20361 54012
rect 20395 54009 20407 54043
rect 20349 54003 20407 54009
rect 22278 54000 22284 54052
rect 22336 54040 22342 54052
rect 25225 54043 25283 54049
rect 25225 54040 25237 54043
rect 22336 54012 25237 54040
rect 22336 54000 22342 54012
rect 25225 54009 25237 54012
rect 25271 54009 25283 54043
rect 25225 54003 25283 54009
rect 16172 53944 16574 53972
rect 16172 53932 16178 53944
rect 17034 53932 17040 53984
rect 17092 53932 17098 53984
rect 18414 53932 18420 53984
rect 18472 53972 18478 53984
rect 18509 53975 18567 53981
rect 18509 53972 18521 53975
rect 18472 53944 18521 53972
rect 18472 53932 18478 53944
rect 18509 53941 18521 53944
rect 18555 53941 18567 53975
rect 18509 53935 18567 53941
rect 19426 53932 19432 53984
rect 19484 53972 19490 53984
rect 19613 53975 19671 53981
rect 19613 53972 19625 53975
rect 19484 53944 19625 53972
rect 19484 53932 19490 53944
rect 19613 53941 19625 53944
rect 19659 53941 19671 53975
rect 19613 53935 19671 53941
rect 21082 53932 21088 53984
rect 21140 53932 21146 53984
rect 22186 53932 22192 53984
rect 22244 53932 22250 53984
rect 22370 53932 22376 53984
rect 22428 53972 22434 53984
rect 22925 53975 22983 53981
rect 22925 53972 22937 53975
rect 22428 53944 22937 53972
rect 22428 53932 22434 53944
rect 22925 53941 22937 53944
rect 22971 53941 22983 53975
rect 22925 53935 22983 53941
rect 23566 53932 23572 53984
rect 23624 53972 23630 53984
rect 23937 53975 23995 53981
rect 23937 53972 23949 53975
rect 23624 53944 23949 53972
rect 23624 53932 23630 53944
rect 23937 53941 23949 53944
rect 23983 53941 23995 53975
rect 23937 53935 23995 53941
rect 1104 53882 25852 53904
rect 1104 53830 2950 53882
rect 3002 53830 3014 53882
rect 3066 53830 3078 53882
rect 3130 53830 3142 53882
rect 3194 53830 3206 53882
rect 3258 53830 12950 53882
rect 13002 53830 13014 53882
rect 13066 53830 13078 53882
rect 13130 53830 13142 53882
rect 13194 53830 13206 53882
rect 13258 53830 22950 53882
rect 23002 53830 23014 53882
rect 23066 53830 23078 53882
rect 23130 53830 23142 53882
rect 23194 53830 23206 53882
rect 23258 53830 25852 53882
rect 1104 53808 25852 53830
rect 16393 53771 16451 53777
rect 16393 53737 16405 53771
rect 16439 53768 16451 53771
rect 16574 53768 16580 53780
rect 16439 53740 16580 53768
rect 16439 53737 16451 53740
rect 16393 53731 16451 53737
rect 16574 53728 16580 53740
rect 16632 53728 16638 53780
rect 18874 53728 18880 53780
rect 18932 53728 18938 53780
rect 5534 53660 5540 53712
rect 5592 53660 5598 53712
rect 21269 53703 21327 53709
rect 21269 53669 21281 53703
rect 21315 53700 21327 53703
rect 21910 53700 21916 53712
rect 21315 53672 21916 53700
rect 21315 53669 21327 53672
rect 21269 53663 21327 53669
rect 21910 53660 21916 53672
rect 21968 53660 21974 53712
rect 22370 53660 22376 53712
rect 22428 53700 22434 53712
rect 23109 53703 23167 53709
rect 23109 53700 23121 53703
rect 22428 53672 23121 53700
rect 22428 53660 22434 53672
rect 23109 53669 23121 53672
rect 23155 53669 23167 53703
rect 23109 53663 23167 53669
rect 3237 53635 3295 53641
rect 3237 53601 3249 53635
rect 3283 53632 3295 53635
rect 5552 53632 5580 53660
rect 3283 53604 5580 53632
rect 6549 53635 6607 53641
rect 3283 53601 3295 53604
rect 3237 53595 3295 53601
rect 6549 53601 6561 53635
rect 6595 53632 6607 53635
rect 7374 53632 7380 53644
rect 6595 53604 7380 53632
rect 6595 53601 6607 53604
rect 6549 53595 6607 53601
rect 7374 53592 7380 53604
rect 7432 53592 7438 53644
rect 8389 53635 8447 53641
rect 8389 53601 8401 53635
rect 8435 53632 8447 53635
rect 8846 53632 8852 53644
rect 8435 53604 8852 53632
rect 8435 53601 8447 53604
rect 8389 53595 8447 53601
rect 8846 53592 8852 53604
rect 8904 53592 8910 53644
rect 11054 53592 11060 53644
rect 11112 53592 11118 53644
rect 12158 53592 12164 53644
rect 12216 53632 12222 53644
rect 12713 53635 12771 53641
rect 12713 53632 12725 53635
rect 12216 53604 12725 53632
rect 12216 53592 12222 53604
rect 12713 53601 12725 53604
rect 12759 53601 12771 53635
rect 24397 53635 24455 53641
rect 24397 53632 24409 53635
rect 12713 53595 12771 53601
rect 23308 53604 24409 53632
rect 2225 53567 2283 53573
rect 2225 53533 2237 53567
rect 2271 53564 2283 53567
rect 5537 53567 5595 53573
rect 2271 53536 4476 53564
rect 2271 53533 2283 53536
rect 2225 53527 2283 53533
rect 4448 53496 4476 53536
rect 5537 53533 5549 53567
rect 5583 53564 5595 53567
rect 6822 53564 6828 53576
rect 5583 53536 6828 53564
rect 5583 53533 5595 53536
rect 5537 53527 5595 53533
rect 6822 53524 6828 53536
rect 6880 53524 6886 53576
rect 7285 53567 7343 53573
rect 7285 53533 7297 53567
rect 7331 53564 7343 53567
rect 9122 53564 9128 53576
rect 7331 53536 9128 53564
rect 7331 53533 7343 53536
rect 7285 53527 7343 53533
rect 9122 53524 9128 53536
rect 9180 53524 9186 53576
rect 10318 53524 10324 53576
rect 10376 53564 10382 53576
rect 10413 53567 10471 53573
rect 10413 53564 10425 53567
rect 10376 53536 10425 53564
rect 10376 53524 10382 53536
rect 10413 53533 10425 53536
rect 10459 53533 10471 53567
rect 10413 53527 10471 53533
rect 12437 53567 12495 53573
rect 12437 53533 12449 53567
rect 12483 53564 12495 53567
rect 12618 53564 12624 53576
rect 12483 53536 12624 53564
rect 12483 53533 12495 53536
rect 12437 53527 12495 53533
rect 12618 53524 12624 53536
rect 12676 53524 12682 53576
rect 13998 53524 14004 53576
rect 14056 53564 14062 53576
rect 14277 53567 14335 53573
rect 14277 53564 14289 53567
rect 14056 53536 14289 53564
rect 14056 53524 14062 53536
rect 14277 53533 14289 53536
rect 14323 53564 14335 53567
rect 14829 53567 14887 53573
rect 14829 53564 14841 53567
rect 14323 53536 14841 53564
rect 14323 53533 14335 53536
rect 14277 53527 14335 53533
rect 14829 53533 14841 53536
rect 14875 53533 14887 53567
rect 14829 53527 14887 53533
rect 15470 53524 15476 53576
rect 15528 53564 15534 53576
rect 15657 53567 15715 53573
rect 15657 53564 15669 53567
rect 15528 53536 15669 53564
rect 15528 53524 15534 53536
rect 15657 53533 15669 53536
rect 15703 53564 15715 53567
rect 16117 53567 16175 53573
rect 16117 53564 16129 53567
rect 15703 53536 16129 53564
rect 15703 53533 15715 53536
rect 15657 53527 15715 53533
rect 16117 53533 16129 53536
rect 16163 53533 16175 53567
rect 16117 53527 16175 53533
rect 16574 53524 16580 53576
rect 16632 53564 16638 53576
rect 16669 53567 16727 53573
rect 16669 53564 16681 53567
rect 16632 53536 16681 53564
rect 16632 53524 16638 53536
rect 16669 53533 16681 53536
rect 16715 53533 16727 53567
rect 16669 53527 16727 53533
rect 17310 53524 17316 53576
rect 17368 53564 17374 53576
rect 17589 53567 17647 53573
rect 17589 53564 17601 53567
rect 17368 53536 17601 53564
rect 17368 53524 17374 53536
rect 17589 53533 17601 53536
rect 17635 53533 17647 53567
rect 17589 53527 17647 53533
rect 18233 53567 18291 53573
rect 18233 53533 18245 53567
rect 18279 53564 18291 53567
rect 18322 53564 18328 53576
rect 18279 53536 18328 53564
rect 18279 53533 18291 53536
rect 18233 53527 18291 53533
rect 18322 53524 18328 53536
rect 18380 53564 18386 53576
rect 18693 53567 18751 53573
rect 18693 53564 18705 53567
rect 18380 53536 18705 53564
rect 18380 53524 18386 53536
rect 18693 53533 18705 53536
rect 18739 53533 18751 53567
rect 18693 53527 18751 53533
rect 19150 53524 19156 53576
rect 19208 53564 19214 53576
rect 19429 53567 19487 53573
rect 19429 53564 19441 53567
rect 19208 53536 19441 53564
rect 19208 53524 19214 53536
rect 19429 53533 19441 53536
rect 19475 53533 19487 53567
rect 19429 53527 19487 53533
rect 19886 53524 19892 53576
rect 19944 53564 19950 53576
rect 20257 53567 20315 53573
rect 20257 53564 20269 53567
rect 19944 53536 20269 53564
rect 19944 53524 19950 53536
rect 20257 53533 20269 53536
rect 20303 53564 20315 53567
rect 20717 53567 20775 53573
rect 20717 53564 20729 53567
rect 20303 53536 20729 53564
rect 20303 53533 20315 53536
rect 20257 53527 20315 53533
rect 20717 53533 20729 53536
rect 20763 53533 20775 53567
rect 20717 53527 20775 53533
rect 20990 53524 20996 53576
rect 21048 53564 21054 53576
rect 21085 53567 21143 53573
rect 21085 53564 21097 53567
rect 21048 53536 21097 53564
rect 21048 53524 21054 53536
rect 21085 53533 21097 53536
rect 21131 53533 21143 53567
rect 21085 53527 21143 53533
rect 21726 53524 21732 53576
rect 21784 53564 21790 53576
rect 22005 53567 22063 53573
rect 22005 53564 22017 53567
rect 21784 53536 22017 53564
rect 21784 53524 21790 53536
rect 22005 53533 22017 53536
rect 22051 53533 22063 53567
rect 22005 53527 22063 53533
rect 22094 53524 22100 53576
rect 22152 53564 22158 53576
rect 22649 53567 22707 53573
rect 22649 53564 22661 53567
rect 22152 53536 22661 53564
rect 22152 53524 22158 53536
rect 22649 53533 22661 53536
rect 22695 53533 22707 53567
rect 22649 53527 22707 53533
rect 22830 53524 22836 53576
rect 22888 53564 22894 53576
rect 23308 53573 23336 53604
rect 24397 53601 24409 53604
rect 24443 53601 24455 53635
rect 24397 53595 24455 53601
rect 23293 53567 23351 53573
rect 23293 53564 23305 53567
rect 22888 53536 23305 53564
rect 22888 53524 22894 53536
rect 23293 53533 23305 53536
rect 23339 53533 23351 53567
rect 23293 53527 23351 53533
rect 23845 53567 23903 53573
rect 23845 53533 23857 53567
rect 23891 53564 23903 53567
rect 24486 53564 24492 53576
rect 23891 53536 24492 53564
rect 23891 53533 23903 53536
rect 23845 53527 23903 53533
rect 24486 53524 24492 53536
rect 24544 53524 24550 53576
rect 24762 53524 24768 53576
rect 24820 53564 24826 53576
rect 24949 53567 25007 53573
rect 24949 53564 24961 53567
rect 24820 53536 24961 53564
rect 24820 53524 24826 53536
rect 24949 53533 24961 53536
rect 24995 53533 25007 53567
rect 24949 53527 25007 53533
rect 7558 53496 7564 53508
rect 4448 53468 7564 53496
rect 7558 53456 7564 53468
rect 7616 53456 7622 53508
rect 18417 53499 18475 53505
rect 18417 53465 18429 53499
rect 18463 53496 18475 53499
rect 18506 53496 18512 53508
rect 18463 53468 18512 53496
rect 18463 53465 18475 53468
rect 18417 53459 18475 53465
rect 18506 53456 18512 53468
rect 18564 53456 18570 53508
rect 20441 53499 20499 53505
rect 20441 53465 20453 53499
rect 20487 53496 20499 53499
rect 20622 53496 20628 53508
rect 20487 53468 20628 53496
rect 20487 53465 20499 53468
rect 20441 53459 20499 53465
rect 20622 53456 20628 53468
rect 20680 53456 20686 53508
rect 14458 53388 14464 53440
rect 14516 53388 14522 53440
rect 15746 53388 15752 53440
rect 15804 53388 15810 53440
rect 16850 53388 16856 53440
rect 16908 53388 16914 53440
rect 17402 53388 17408 53440
rect 17460 53388 17466 53440
rect 19610 53388 19616 53440
rect 19668 53388 19674 53440
rect 20898 53388 20904 53440
rect 20956 53428 20962 53440
rect 21821 53431 21879 53437
rect 21821 53428 21833 53431
rect 20956 53400 21833 53428
rect 20956 53388 20962 53400
rect 21821 53397 21833 53400
rect 21867 53397 21879 53431
rect 21821 53391 21879 53397
rect 22462 53388 22468 53440
rect 22520 53388 22526 53440
rect 23934 53388 23940 53440
rect 23992 53388 23998 53440
rect 25038 53388 25044 53440
rect 25096 53388 25102 53440
rect 1104 53338 25852 53360
rect 1104 53286 7950 53338
rect 8002 53286 8014 53338
rect 8066 53286 8078 53338
rect 8130 53286 8142 53338
rect 8194 53286 8206 53338
rect 8258 53286 17950 53338
rect 18002 53286 18014 53338
rect 18066 53286 18078 53338
rect 18130 53286 18142 53338
rect 18194 53286 18206 53338
rect 18258 53286 25852 53338
rect 1104 53264 25852 53286
rect 2133 53227 2191 53233
rect 2133 53193 2145 53227
rect 2179 53224 2191 53227
rect 2774 53224 2780 53236
rect 2179 53196 2780 53224
rect 2179 53193 2191 53196
rect 2133 53187 2191 53193
rect 1765 53091 1823 53097
rect 1765 53057 1777 53091
rect 1811 53088 1823 53091
rect 2148 53088 2176 53187
rect 2774 53184 2780 53196
rect 2832 53184 2838 53236
rect 5166 53184 5172 53236
rect 5224 53224 5230 53236
rect 5718 53224 5724 53236
rect 5224 53196 5724 53224
rect 5224 53184 5230 53196
rect 5718 53184 5724 53196
rect 5776 53184 5782 53236
rect 17310 53184 17316 53236
rect 17368 53184 17374 53236
rect 19150 53184 19156 53236
rect 19208 53224 19214 53236
rect 19521 53227 19579 53233
rect 19521 53224 19533 53227
rect 19208 53196 19533 53224
rect 19208 53184 19214 53196
rect 19521 53193 19533 53196
rect 19567 53193 19579 53227
rect 19521 53187 19579 53193
rect 19702 53184 19708 53236
rect 19760 53184 19766 53236
rect 20990 53184 20996 53236
rect 21048 53184 21054 53236
rect 21726 53184 21732 53236
rect 21784 53224 21790 53236
rect 21821 53227 21879 53233
rect 21821 53224 21833 53227
rect 21784 53196 21833 53224
rect 21784 53184 21790 53196
rect 21821 53193 21833 53196
rect 21867 53193 21879 53227
rect 21821 53187 21879 53193
rect 22094 53184 22100 53236
rect 22152 53224 22158 53236
rect 22281 53227 22339 53233
rect 22281 53224 22293 53227
rect 22152 53196 22293 53224
rect 22152 53184 22158 53196
rect 22281 53193 22293 53196
rect 22327 53193 22339 53227
rect 22281 53187 22339 53193
rect 22554 53184 22560 53236
rect 22612 53184 22618 53236
rect 23017 53227 23075 53233
rect 23017 53193 23029 53227
rect 23063 53224 23075 53227
rect 23290 53224 23296 53236
rect 23063 53196 23296 53224
rect 23063 53193 23075 53196
rect 23017 53187 23075 53193
rect 23290 53184 23296 53196
rect 23348 53184 23354 53236
rect 3973 53159 4031 53165
rect 3973 53125 3985 53159
rect 4019 53156 4031 53159
rect 4430 53156 4436 53168
rect 4019 53128 4436 53156
rect 4019 53125 4031 53128
rect 3973 53119 4031 53125
rect 4430 53116 4436 53128
rect 4488 53116 4494 53168
rect 5813 53159 5871 53165
rect 5813 53125 5825 53159
rect 5859 53156 5871 53159
rect 6270 53156 6276 53168
rect 5859 53128 6276 53156
rect 5859 53125 5871 53128
rect 5813 53119 5871 53125
rect 6270 53116 6276 53128
rect 6328 53116 6334 53168
rect 9125 53159 9183 53165
rect 9125 53125 9137 53159
rect 9171 53156 9183 53159
rect 9214 53156 9220 53168
rect 9171 53128 9220 53156
rect 9171 53125 9183 53128
rect 9125 53119 9183 53125
rect 9214 53116 9220 53128
rect 9272 53116 9278 53168
rect 10962 53156 10968 53168
rect 9416 53128 10968 53156
rect 1811 53060 2176 53088
rect 2961 53091 3019 53097
rect 1811 53057 1823 53060
rect 1765 53051 1823 53057
rect 2961 53057 2973 53091
rect 3007 53057 3019 53091
rect 2961 53051 3019 53057
rect 4801 53091 4859 53097
rect 4801 53057 4813 53091
rect 4847 53088 4859 53091
rect 6454 53088 6460 53100
rect 4847 53060 6460 53088
rect 4847 53057 4859 53060
rect 4801 53051 4859 53057
rect 2976 53020 3004 53051
rect 6454 53048 6460 53060
rect 6512 53048 6518 53100
rect 8113 53091 8171 53097
rect 8113 53057 8125 53091
rect 8159 53088 8171 53091
rect 9416 53088 9444 53128
rect 10962 53116 10968 53128
rect 11020 53116 11026 53168
rect 13630 53116 13636 53168
rect 13688 53156 13694 53168
rect 13817 53159 13875 53165
rect 13817 53156 13829 53159
rect 13688 53128 13829 53156
rect 13688 53116 13694 53128
rect 13817 53125 13829 53128
rect 13863 53125 13875 53159
rect 13817 53119 13875 53125
rect 20714 53116 20720 53168
rect 20772 53156 20778 53168
rect 21177 53159 21235 53165
rect 21177 53156 21189 53159
rect 20772 53128 21189 53156
rect 20772 53116 20778 53128
rect 21177 53125 21189 53128
rect 21223 53125 21235 53159
rect 21177 53119 21235 53125
rect 8159 53060 9444 53088
rect 8159 53057 8171 53060
rect 8113 53051 8171 53057
rect 9766 53048 9772 53100
rect 9824 53048 9830 53100
rect 11882 53048 11888 53100
rect 11940 53048 11946 53100
rect 14366 53048 14372 53100
rect 14424 53088 14430 53100
rect 14645 53091 14703 53097
rect 14645 53088 14657 53091
rect 14424 53060 14657 53088
rect 14424 53048 14430 53060
rect 14645 53057 14657 53060
rect 14691 53088 14703 53091
rect 14921 53091 14979 53097
rect 14921 53088 14933 53091
rect 14691 53060 14933 53088
rect 14691 53057 14703 53060
rect 14645 53051 14703 53057
rect 14921 53057 14933 53060
rect 14967 53057 14979 53091
rect 14921 53051 14979 53057
rect 15838 53048 15844 53100
rect 15896 53088 15902 53100
rect 16117 53091 16175 53097
rect 16117 53088 16129 53091
rect 15896 53060 16129 53088
rect 15896 53048 15902 53060
rect 16117 53057 16129 53060
rect 16163 53088 16175 53091
rect 16393 53091 16451 53097
rect 16393 53088 16405 53091
rect 16163 53060 16405 53088
rect 16163 53057 16175 53060
rect 16117 53051 16175 53057
rect 16393 53057 16405 53060
rect 16439 53057 16451 53091
rect 16393 53051 16451 53057
rect 18782 53048 18788 53100
rect 18840 53088 18846 53100
rect 19061 53091 19119 53097
rect 19061 53088 19073 53091
rect 18840 53060 19073 53088
rect 18840 53048 18846 53060
rect 19061 53057 19073 53060
rect 19107 53088 19119 53091
rect 19337 53091 19395 53097
rect 19337 53088 19349 53091
rect 19107 53060 19349 53088
rect 19107 53057 19119 53060
rect 19061 53051 19119 53057
rect 19337 53057 19349 53060
rect 19383 53057 19395 53091
rect 19337 53051 19395 53057
rect 20254 53048 20260 53100
rect 20312 53088 20318 53100
rect 20533 53091 20591 53097
rect 20533 53088 20545 53091
rect 20312 53060 20545 53088
rect 20312 53048 20318 53060
rect 20533 53057 20545 53060
rect 20579 53088 20591 53091
rect 20809 53091 20867 53097
rect 20809 53088 20821 53091
rect 20579 53060 20821 53088
rect 20579 53057 20591 53060
rect 20533 53051 20591 53057
rect 20809 53057 20821 53060
rect 20855 53057 20867 53091
rect 23308 53088 23336 53184
rect 23477 53091 23535 53097
rect 23477 53088 23489 53091
rect 23308 53060 23489 53088
rect 20809 53051 20867 53057
rect 23477 53057 23489 53060
rect 23523 53057 23535 53091
rect 23477 53051 23535 53057
rect 23658 53048 23664 53100
rect 23716 53088 23722 53100
rect 24121 53091 24179 53097
rect 24121 53088 24133 53091
rect 23716 53060 24133 53088
rect 23716 53048 23722 53060
rect 24121 53057 24133 53060
rect 24167 53088 24179 53091
rect 24397 53091 24455 53097
rect 24397 53088 24409 53091
rect 24167 53060 24409 53088
rect 24167 53057 24179 53060
rect 24121 53051 24179 53057
rect 24397 53057 24409 53060
rect 24443 53057 24455 53091
rect 24397 53051 24455 53057
rect 24765 53091 24823 53097
rect 24765 53057 24777 53091
rect 24811 53088 24823 53091
rect 25038 53088 25044 53100
rect 24811 53060 25044 53088
rect 24811 53057 24823 53060
rect 24765 53051 24823 53057
rect 25038 53048 25044 53060
rect 25096 53048 25102 53100
rect 5534 53020 5540 53032
rect 2976 52992 5540 53020
rect 5534 52980 5540 52992
rect 5592 52980 5598 53032
rect 10410 52980 10416 53032
rect 10468 52980 10474 53032
rect 11790 52980 11796 53032
rect 11848 53020 11854 53032
rect 12345 53023 12403 53029
rect 12345 53020 12357 53023
rect 11848 52992 12357 53020
rect 11848 52980 11854 52992
rect 12345 52989 12357 52992
rect 12391 52989 12403 53023
rect 12345 52983 12403 52989
rect 3418 52912 3424 52964
rect 3476 52952 3482 52964
rect 9582 52952 9588 52964
rect 3476 52924 9588 52952
rect 3476 52912 3482 52924
rect 9582 52912 9588 52924
rect 9640 52912 9646 52964
rect 13998 52912 14004 52964
rect 14056 52912 14062 52964
rect 1581 52887 1639 52893
rect 1581 52853 1593 52887
rect 1627 52884 1639 52887
rect 4062 52884 4068 52896
rect 1627 52856 4068 52884
rect 1627 52853 1639 52856
rect 1581 52847 1639 52853
rect 4062 52844 4068 52856
rect 4120 52844 4126 52896
rect 14461 52887 14519 52893
rect 14461 52853 14473 52887
rect 14507 52884 14519 52887
rect 14642 52884 14648 52896
rect 14507 52856 14648 52884
rect 14507 52853 14519 52856
rect 14461 52847 14519 52853
rect 14642 52844 14648 52856
rect 14700 52844 14706 52896
rect 15930 52844 15936 52896
rect 15988 52844 15994 52896
rect 18598 52844 18604 52896
rect 18656 52884 18662 52896
rect 18877 52887 18935 52893
rect 18877 52884 18889 52887
rect 18656 52856 18889 52884
rect 18656 52844 18662 52856
rect 18877 52853 18889 52856
rect 18923 52853 18935 52887
rect 18877 52847 18935 52853
rect 20346 52844 20352 52896
rect 20404 52844 20410 52896
rect 22554 52844 22560 52896
rect 22612 52884 22618 52896
rect 23293 52887 23351 52893
rect 23293 52884 23305 52887
rect 22612 52856 23305 52884
rect 22612 52844 22618 52856
rect 23293 52853 23305 52856
rect 23339 52853 23351 52887
rect 23293 52847 23351 52853
rect 23934 52844 23940 52896
rect 23992 52844 23998 52896
rect 24854 52844 24860 52896
rect 24912 52884 24918 52896
rect 25225 52887 25283 52893
rect 25225 52884 25237 52887
rect 24912 52856 25237 52884
rect 24912 52844 24918 52856
rect 25225 52853 25237 52856
rect 25271 52853 25283 52887
rect 25225 52847 25283 52853
rect 1104 52794 25852 52816
rect 1104 52742 2950 52794
rect 3002 52742 3014 52794
rect 3066 52742 3078 52794
rect 3130 52742 3142 52794
rect 3194 52742 3206 52794
rect 3258 52742 12950 52794
rect 13002 52742 13014 52794
rect 13066 52742 13078 52794
rect 13130 52742 13142 52794
rect 13194 52742 13206 52794
rect 13258 52742 22950 52794
rect 23002 52742 23014 52794
rect 23066 52742 23078 52794
rect 23130 52742 23142 52794
rect 23194 52742 23206 52794
rect 23258 52742 25852 52794
rect 1104 52720 25852 52742
rect 2222 52640 2228 52692
rect 2280 52680 2286 52692
rect 3418 52680 3424 52692
rect 2280 52652 3424 52680
rect 2280 52640 2286 52652
rect 3418 52640 3424 52652
rect 3476 52640 3482 52692
rect 12618 52640 12624 52692
rect 12676 52640 12682 52692
rect 13630 52640 13636 52692
rect 13688 52680 13694 52692
rect 14093 52683 14151 52689
rect 14093 52680 14105 52683
rect 13688 52652 14105 52680
rect 13688 52640 13694 52652
rect 14093 52649 14105 52652
rect 14139 52649 14151 52683
rect 14093 52643 14151 52649
rect 24581 52683 24639 52689
rect 24581 52649 24593 52683
rect 24627 52680 24639 52683
rect 24762 52680 24768 52692
rect 24627 52652 24768 52680
rect 24627 52649 24639 52652
rect 24581 52643 24639 52649
rect 24762 52640 24768 52652
rect 24820 52640 24826 52692
rect 1854 52572 1860 52624
rect 1912 52612 1918 52624
rect 3510 52612 3516 52624
rect 1912 52584 3516 52612
rect 1912 52572 1918 52584
rect 3510 52572 3516 52584
rect 3568 52572 3574 52624
rect 25130 52572 25136 52624
rect 25188 52612 25194 52624
rect 25225 52615 25283 52621
rect 25225 52612 25237 52615
rect 25188 52584 25237 52612
rect 25188 52572 25194 52584
rect 25225 52581 25237 52584
rect 25271 52581 25283 52615
rect 25225 52575 25283 52581
rect 3237 52547 3295 52553
rect 3237 52513 3249 52547
rect 3283 52544 3295 52547
rect 3694 52544 3700 52556
rect 3283 52516 3700 52544
rect 3283 52513 3295 52516
rect 3237 52507 3295 52513
rect 3694 52504 3700 52516
rect 3752 52504 3758 52556
rect 6549 52547 6607 52553
rect 6549 52513 6561 52547
rect 6595 52544 6607 52547
rect 6638 52544 6644 52556
rect 6595 52516 6644 52544
rect 6595 52513 6607 52516
rect 6549 52507 6607 52513
rect 6638 52504 6644 52516
rect 6696 52504 6702 52556
rect 7742 52504 7748 52556
rect 7800 52504 7806 52556
rect 10686 52504 10692 52556
rect 10744 52544 10750 52556
rect 11241 52547 11299 52553
rect 11241 52544 11253 52547
rect 10744 52516 11253 52544
rect 10744 52504 10750 52516
rect 11241 52513 11253 52516
rect 11287 52513 11299 52547
rect 11241 52507 11299 52513
rect 13630 52504 13636 52556
rect 13688 52504 13694 52556
rect 2225 52479 2283 52485
rect 2225 52445 2237 52479
rect 2271 52476 2283 52479
rect 4798 52476 4804 52488
rect 2271 52448 4804 52476
rect 2271 52445 2283 52448
rect 2225 52439 2283 52445
rect 4798 52436 4804 52448
rect 4856 52436 4862 52488
rect 5445 52479 5503 52485
rect 5445 52445 5457 52479
rect 5491 52476 5503 52479
rect 5626 52476 5632 52488
rect 5491 52448 5632 52476
rect 5491 52445 5503 52448
rect 5445 52439 5503 52445
rect 5626 52436 5632 52448
rect 5684 52436 5690 52488
rect 7190 52436 7196 52488
rect 7248 52436 7254 52488
rect 10778 52436 10784 52488
rect 10836 52436 10842 52488
rect 12802 52436 12808 52488
rect 12860 52436 12866 52488
rect 24762 52436 24768 52488
rect 24820 52476 24826 52488
rect 25041 52479 25099 52485
rect 25041 52476 25053 52479
rect 24820 52448 25053 52476
rect 24820 52436 24826 52448
rect 25041 52445 25053 52448
rect 25087 52445 25099 52479
rect 25041 52439 25099 52445
rect 13354 52368 13360 52420
rect 13412 52408 13418 52420
rect 13449 52411 13507 52417
rect 13449 52408 13461 52411
rect 13412 52380 13461 52408
rect 13412 52368 13418 52380
rect 13449 52377 13461 52380
rect 13495 52377 13507 52411
rect 13449 52371 13507 52377
rect 1104 52250 25852 52272
rect 1104 52198 7950 52250
rect 8002 52198 8014 52250
rect 8066 52198 8078 52250
rect 8130 52198 8142 52250
rect 8194 52198 8206 52250
rect 8258 52198 17950 52250
rect 18002 52198 18014 52250
rect 18066 52198 18078 52250
rect 18130 52198 18142 52250
rect 18194 52198 18206 52250
rect 18258 52198 25852 52250
rect 1104 52176 25852 52198
rect 5534 52096 5540 52148
rect 5592 52136 5598 52148
rect 7009 52139 7067 52145
rect 7009 52136 7021 52139
rect 5592 52108 7021 52136
rect 5592 52096 5598 52108
rect 7009 52105 7021 52108
rect 7055 52105 7067 52139
rect 7009 52099 7067 52105
rect 11701 52139 11759 52145
rect 11701 52105 11713 52139
rect 11747 52136 11759 52139
rect 11882 52136 11888 52148
rect 11747 52108 11888 52136
rect 11747 52105 11759 52108
rect 11701 52099 11759 52105
rect 11882 52096 11888 52108
rect 11940 52096 11946 52148
rect 12342 52096 12348 52148
rect 12400 52096 12406 52148
rect 13265 52139 13323 52145
rect 13265 52105 13277 52139
rect 13311 52136 13323 52139
rect 13354 52136 13360 52148
rect 13311 52108 13360 52136
rect 13311 52105 13323 52108
rect 13265 52099 13323 52105
rect 13354 52096 13360 52108
rect 13412 52096 13418 52148
rect 25314 52096 25320 52148
rect 25372 52096 25378 52148
rect 6917 52071 6975 52077
rect 6917 52037 6929 52071
rect 6963 52068 6975 52071
rect 9214 52068 9220 52080
rect 6963 52040 9220 52068
rect 6963 52037 6975 52040
rect 6917 52031 6975 52037
rect 9214 52028 9220 52040
rect 9272 52028 9278 52080
rect 2961 52003 3019 52009
rect 2961 51969 2973 52003
rect 3007 52000 3019 52003
rect 4522 52000 4528 52012
rect 3007 51972 4528 52000
rect 3007 51969 3019 51972
rect 2961 51963 3019 51969
rect 4522 51960 4528 51972
rect 4580 51960 4586 52012
rect 4801 52003 4859 52009
rect 4801 51969 4813 52003
rect 4847 52000 4859 52003
rect 4982 52000 4988 52012
rect 4847 51972 4988 52000
rect 4847 51969 4859 51972
rect 4801 51963 4859 51969
rect 4982 51960 4988 51972
rect 5040 51960 5046 52012
rect 7374 51960 7380 52012
rect 7432 52000 7438 52012
rect 7837 52003 7895 52009
rect 7837 52000 7849 52003
rect 7432 51972 7849 52000
rect 7432 51960 7438 51972
rect 7837 51969 7849 51972
rect 7883 51969 7895 52003
rect 7837 51963 7895 51969
rect 9858 51960 9864 52012
rect 9916 51960 9922 52012
rect 11882 51960 11888 52012
rect 11940 51960 11946 52012
rect 11974 51960 11980 52012
rect 12032 52000 12038 52012
rect 12529 52003 12587 52009
rect 12529 52000 12541 52003
rect 12032 51972 12541 52000
rect 12032 51960 12038 51972
rect 12529 51969 12541 51972
rect 12575 51969 12587 52003
rect 12529 51963 12587 51969
rect 3326 51892 3332 51944
rect 3384 51892 3390 51944
rect 4890 51892 4896 51944
rect 4948 51932 4954 51944
rect 5077 51935 5135 51941
rect 5077 51932 5089 51935
rect 4948 51904 5089 51932
rect 4948 51892 4954 51904
rect 5077 51901 5089 51904
rect 5123 51901 5135 51935
rect 5077 51895 5135 51901
rect 8478 51892 8484 51944
rect 8536 51892 8542 51944
rect 9674 51892 9680 51944
rect 9732 51932 9738 51944
rect 10137 51935 10195 51941
rect 10137 51932 10149 51935
rect 9732 51904 10149 51932
rect 9732 51892 9738 51904
rect 10137 51901 10149 51904
rect 10183 51901 10195 51935
rect 10137 51895 10195 51901
rect 25498 51756 25504 51808
rect 25556 51756 25562 51808
rect 1104 51706 25852 51728
rect 1104 51654 2950 51706
rect 3002 51654 3014 51706
rect 3066 51654 3078 51706
rect 3130 51654 3142 51706
rect 3194 51654 3206 51706
rect 3258 51654 12950 51706
rect 13002 51654 13014 51706
rect 13066 51654 13078 51706
rect 13130 51654 13142 51706
rect 13194 51654 13206 51706
rect 13258 51654 22950 51706
rect 23002 51654 23014 51706
rect 23066 51654 23078 51706
rect 23130 51654 23142 51706
rect 23194 51654 23206 51706
rect 23258 51654 25852 51706
rect 1104 51632 25852 51654
rect 9950 51552 9956 51604
rect 10008 51592 10014 51604
rect 10229 51595 10287 51601
rect 10229 51592 10241 51595
rect 10008 51564 10241 51592
rect 10008 51552 10014 51564
rect 10229 51561 10241 51564
rect 10275 51561 10287 51595
rect 10229 51555 10287 51561
rect 2866 51416 2872 51468
rect 2924 51416 2930 51468
rect 5718 51416 5724 51468
rect 5776 51416 5782 51468
rect 7006 51416 7012 51468
rect 7064 51456 7070 51468
rect 7561 51459 7619 51465
rect 7561 51456 7573 51459
rect 7064 51428 7573 51456
rect 7064 51416 7070 51428
rect 7561 51425 7573 51428
rect 7607 51425 7619 51459
rect 7561 51419 7619 51425
rect 2225 51391 2283 51397
rect 2225 51357 2237 51391
rect 2271 51357 2283 51391
rect 2225 51351 2283 51357
rect 5445 51391 5503 51397
rect 5445 51357 5457 51391
rect 5491 51388 5503 51391
rect 6730 51388 6736 51400
rect 5491 51360 6736 51388
rect 5491 51357 5503 51360
rect 5445 51351 5503 51357
rect 2240 51320 2268 51351
rect 6730 51348 6736 51360
rect 6788 51348 6794 51400
rect 7098 51348 7104 51400
rect 7156 51348 7162 51400
rect 9306 51348 9312 51400
rect 9364 51388 9370 51400
rect 10413 51391 10471 51397
rect 10413 51388 10425 51391
rect 9364 51360 10425 51388
rect 9364 51348 9370 51360
rect 10413 51357 10425 51360
rect 10459 51357 10471 51391
rect 10413 51351 10471 51357
rect 25041 51391 25099 51397
rect 25041 51357 25053 51391
rect 25087 51388 25099 51391
rect 25498 51388 25504 51400
rect 25087 51360 25504 51388
rect 25087 51357 25099 51360
rect 25041 51351 25099 51357
rect 25498 51348 25504 51360
rect 25556 51348 25562 51400
rect 5534 51320 5540 51332
rect 2240 51292 5540 51320
rect 5534 51280 5540 51292
rect 5592 51280 5598 51332
rect 24946 51212 24952 51264
rect 25004 51252 25010 51264
rect 25225 51255 25283 51261
rect 25225 51252 25237 51255
rect 25004 51224 25237 51252
rect 25004 51212 25010 51224
rect 25225 51221 25237 51224
rect 25271 51221 25283 51255
rect 25225 51215 25283 51221
rect 1104 51162 25852 51184
rect 1104 51110 7950 51162
rect 8002 51110 8014 51162
rect 8066 51110 8078 51162
rect 8130 51110 8142 51162
rect 8194 51110 8206 51162
rect 8258 51110 17950 51162
rect 18002 51110 18014 51162
rect 18066 51110 18078 51162
rect 18130 51110 18142 51162
rect 18194 51110 18206 51162
rect 18258 51110 25852 51162
rect 1104 51088 25852 51110
rect 4338 51008 4344 51060
rect 4396 51008 4402 51060
rect 5534 51008 5540 51060
rect 5592 51048 5598 51060
rect 6917 51051 6975 51057
rect 6917 51048 6929 51051
rect 5592 51020 6929 51048
rect 5592 51008 5598 51020
rect 6917 51017 6929 51020
rect 6963 51017 6975 51051
rect 6917 51011 6975 51017
rect 4356 50980 4384 51008
rect 9585 50983 9643 50989
rect 4356 50952 7788 50980
rect 2501 50915 2559 50921
rect 2501 50881 2513 50915
rect 2547 50912 2559 50915
rect 4154 50912 4160 50924
rect 2547 50884 4160 50912
rect 2547 50881 2559 50884
rect 2501 50875 2559 50881
rect 4154 50872 4160 50884
rect 4212 50872 4218 50924
rect 4338 50872 4344 50924
rect 4396 50872 4402 50924
rect 6825 50915 6883 50921
rect 6825 50881 6837 50915
rect 6871 50912 6883 50915
rect 7650 50912 7656 50924
rect 6871 50884 7656 50912
rect 6871 50881 6883 50884
rect 6825 50875 6883 50881
rect 7650 50872 7656 50884
rect 7708 50872 7714 50924
rect 7760 50921 7788 50952
rect 9585 50949 9597 50983
rect 9631 50980 9643 50983
rect 10778 50980 10784 50992
rect 9631 50952 10784 50980
rect 9631 50949 9643 50952
rect 9585 50943 9643 50949
rect 10778 50940 10784 50952
rect 10836 50940 10842 50992
rect 7745 50915 7803 50921
rect 7745 50881 7757 50915
rect 7791 50881 7803 50915
rect 7745 50875 7803 50881
rect 9398 50872 9404 50924
rect 9456 50872 9462 50924
rect 24765 50915 24823 50921
rect 24765 50881 24777 50915
rect 24811 50912 24823 50915
rect 25038 50912 25044 50924
rect 24811 50884 25044 50912
rect 24811 50881 24823 50884
rect 24765 50875 24823 50881
rect 25038 50872 25044 50884
rect 25096 50872 25102 50924
rect 2774 50804 2780 50856
rect 2832 50804 2838 50856
rect 4246 50804 4252 50856
rect 4304 50844 4310 50856
rect 4617 50847 4675 50853
rect 4617 50844 4629 50847
rect 4304 50816 4629 50844
rect 4304 50804 4310 50816
rect 4617 50813 4629 50816
rect 4663 50813 4675 50847
rect 4617 50807 4675 50813
rect 7466 50804 7472 50856
rect 7524 50804 7530 50856
rect 24302 50668 24308 50720
rect 24360 50708 24366 50720
rect 25225 50711 25283 50717
rect 25225 50708 25237 50711
rect 24360 50680 25237 50708
rect 24360 50668 24366 50680
rect 25225 50677 25237 50680
rect 25271 50677 25283 50711
rect 25225 50671 25283 50677
rect 1104 50618 25852 50640
rect 1104 50566 2950 50618
rect 3002 50566 3014 50618
rect 3066 50566 3078 50618
rect 3130 50566 3142 50618
rect 3194 50566 3206 50618
rect 3258 50566 12950 50618
rect 13002 50566 13014 50618
rect 13066 50566 13078 50618
rect 13130 50566 13142 50618
rect 13194 50566 13206 50618
rect 13258 50566 22950 50618
rect 23002 50566 23014 50618
rect 23066 50566 23078 50618
rect 23130 50566 23142 50618
rect 23194 50566 23206 50618
rect 23258 50566 25852 50618
rect 1104 50544 25852 50566
rect 6822 50464 6828 50516
rect 6880 50464 6886 50516
rect 9122 50464 9128 50516
rect 9180 50504 9186 50516
rect 9217 50507 9275 50513
rect 9217 50504 9229 50507
rect 9180 50476 9229 50504
rect 9180 50464 9186 50476
rect 9217 50473 9229 50476
rect 9263 50473 9275 50507
rect 9217 50467 9275 50473
rect 21450 50396 21456 50448
rect 21508 50436 21514 50448
rect 25133 50439 25191 50445
rect 25133 50436 25145 50439
rect 21508 50408 25145 50436
rect 21508 50396 21514 50408
rect 25133 50405 25145 50408
rect 25179 50405 25191 50439
rect 25133 50399 25191 50405
rect 3237 50371 3295 50377
rect 3237 50337 3249 50371
rect 3283 50368 3295 50371
rect 3418 50368 3424 50380
rect 3283 50340 3424 50368
rect 3283 50337 3295 50340
rect 3237 50331 3295 50337
rect 3418 50328 3424 50340
rect 3476 50328 3482 50380
rect 2225 50303 2283 50309
rect 2225 50269 2237 50303
rect 2271 50300 2283 50303
rect 4706 50300 4712 50312
rect 2271 50272 4712 50300
rect 2271 50269 2283 50272
rect 2225 50263 2283 50269
rect 4706 50260 4712 50272
rect 4764 50260 4770 50312
rect 5810 50260 5816 50312
rect 5868 50300 5874 50312
rect 7009 50303 7067 50309
rect 7009 50300 7021 50303
rect 5868 50272 7021 50300
rect 5868 50260 5874 50272
rect 7009 50269 7021 50272
rect 7055 50269 7067 50303
rect 7009 50263 7067 50269
rect 8386 50260 8392 50312
rect 8444 50300 8450 50312
rect 9401 50303 9459 50309
rect 9401 50300 9413 50303
rect 8444 50272 9413 50300
rect 8444 50260 8450 50272
rect 9401 50269 9413 50272
rect 9447 50269 9459 50303
rect 9401 50263 9459 50269
rect 24673 50303 24731 50309
rect 24673 50269 24685 50303
rect 24719 50300 24731 50303
rect 25314 50300 25320 50312
rect 24719 50272 25320 50300
rect 24719 50269 24731 50272
rect 24673 50263 24731 50269
rect 25314 50260 25320 50272
rect 25372 50260 25378 50312
rect 24486 50124 24492 50176
rect 24544 50164 24550 50176
rect 24765 50167 24823 50173
rect 24765 50164 24777 50167
rect 24544 50136 24777 50164
rect 24544 50124 24550 50136
rect 24765 50133 24777 50136
rect 24811 50133 24823 50167
rect 24765 50127 24823 50133
rect 1104 50074 25852 50096
rect 1104 50022 7950 50074
rect 8002 50022 8014 50074
rect 8066 50022 8078 50074
rect 8130 50022 8142 50074
rect 8194 50022 8206 50074
rect 8258 50022 17950 50074
rect 18002 50022 18014 50074
rect 18066 50022 18078 50074
rect 18130 50022 18142 50074
rect 18194 50022 18206 50074
rect 18258 50022 25852 50074
rect 1104 50000 25852 50022
rect 6365 49963 6423 49969
rect 6365 49960 6377 49963
rect 3988 49932 6377 49960
rect 3145 49895 3203 49901
rect 3145 49861 3157 49895
rect 3191 49892 3203 49895
rect 3510 49892 3516 49904
rect 3191 49864 3516 49892
rect 3191 49861 3203 49864
rect 3145 49855 3203 49861
rect 3510 49852 3516 49864
rect 3568 49852 3574 49904
rect 2133 49827 2191 49833
rect 2133 49793 2145 49827
rect 2179 49824 2191 49827
rect 3602 49824 3608 49836
rect 2179 49796 3608 49824
rect 2179 49793 2191 49796
rect 2133 49787 2191 49793
rect 3602 49784 3608 49796
rect 3660 49784 3666 49836
rect 3988 49833 4016 49932
rect 6365 49929 6377 49932
rect 6411 49960 6423 49963
rect 6822 49960 6828 49972
rect 6411 49932 6828 49960
rect 6411 49929 6423 49932
rect 6365 49923 6423 49929
rect 6822 49920 6828 49932
rect 6880 49920 6886 49972
rect 6549 49895 6607 49901
rect 6549 49892 6561 49895
rect 5474 49864 6561 49892
rect 6549 49861 6561 49864
rect 6595 49892 6607 49895
rect 8478 49892 8484 49904
rect 6595 49864 8484 49892
rect 6595 49861 6607 49864
rect 6549 49855 6607 49861
rect 8478 49852 8484 49864
rect 8536 49852 8542 49904
rect 9401 49895 9459 49901
rect 9401 49861 9413 49895
rect 9447 49892 9459 49895
rect 9766 49892 9772 49904
rect 9447 49864 9772 49892
rect 9447 49861 9459 49864
rect 9401 49855 9459 49861
rect 9766 49852 9772 49864
rect 9824 49852 9830 49904
rect 3973 49827 4031 49833
rect 3973 49793 3985 49827
rect 4019 49793 4031 49827
rect 3973 49787 4031 49793
rect 7834 49784 7840 49836
rect 7892 49824 7898 49836
rect 9217 49827 9275 49833
rect 9217 49824 9229 49827
rect 7892 49796 9229 49824
rect 7892 49784 7898 49796
rect 9217 49793 9229 49796
rect 9263 49793 9275 49827
rect 9217 49787 9275 49793
rect 21634 49784 21640 49836
rect 21692 49824 21698 49836
rect 24765 49827 24823 49833
rect 24765 49824 24777 49827
rect 21692 49796 24777 49824
rect 21692 49784 21698 49796
rect 24765 49793 24777 49796
rect 24811 49793 24823 49827
rect 24765 49787 24823 49793
rect 5997 49759 6055 49765
rect 5997 49725 6009 49759
rect 6043 49756 6055 49759
rect 8754 49756 8760 49768
rect 6043 49728 8760 49756
rect 6043 49725 6055 49728
rect 5997 49719 6055 49725
rect 8754 49716 8760 49728
rect 8812 49716 8818 49768
rect 24486 49716 24492 49768
rect 24544 49716 24550 49768
rect 4062 49580 4068 49632
rect 4120 49620 4126 49632
rect 4230 49623 4288 49629
rect 4230 49620 4242 49623
rect 4120 49592 4242 49620
rect 4120 49580 4126 49592
rect 4230 49589 4242 49592
rect 4276 49589 4288 49623
rect 4230 49583 4288 49589
rect 1104 49530 25852 49552
rect 1104 49478 2950 49530
rect 3002 49478 3014 49530
rect 3066 49478 3078 49530
rect 3130 49478 3142 49530
rect 3194 49478 3206 49530
rect 3258 49478 12950 49530
rect 13002 49478 13014 49530
rect 13066 49478 13078 49530
rect 13130 49478 13142 49530
rect 13194 49478 13206 49530
rect 13258 49478 22950 49530
rect 23002 49478 23014 49530
rect 23066 49478 23078 49530
rect 23130 49478 23142 49530
rect 23194 49478 23206 49530
rect 23258 49478 25852 49530
rect 1104 49456 25852 49478
rect 11609 49419 11667 49425
rect 11609 49385 11621 49419
rect 11655 49416 11667 49419
rect 11974 49416 11980 49428
rect 11655 49388 11980 49416
rect 11655 49385 11667 49388
rect 11609 49379 11667 49385
rect 11974 49376 11980 49388
rect 12032 49376 12038 49428
rect 12713 49419 12771 49425
rect 12713 49385 12725 49419
rect 12759 49416 12771 49419
rect 12802 49416 12808 49428
rect 12759 49388 12808 49416
rect 12759 49385 12771 49388
rect 12713 49379 12771 49385
rect 12802 49376 12808 49388
rect 12860 49376 12866 49428
rect 1486 49240 1492 49292
rect 1544 49280 1550 49292
rect 2041 49283 2099 49289
rect 2041 49280 2053 49283
rect 1544 49252 2053 49280
rect 1544 49240 1550 49252
rect 2041 49249 2053 49252
rect 2087 49249 2099 49283
rect 2041 49243 2099 49249
rect 1765 49215 1823 49221
rect 1765 49181 1777 49215
rect 1811 49181 1823 49215
rect 1765 49175 1823 49181
rect 1780 49076 1808 49175
rect 10686 49172 10692 49224
rect 10744 49212 10750 49224
rect 11793 49215 11851 49221
rect 11793 49212 11805 49215
rect 10744 49184 11805 49212
rect 10744 49172 10750 49184
rect 11793 49181 11805 49184
rect 11839 49181 11851 49215
rect 11793 49175 11851 49181
rect 12897 49215 12955 49221
rect 12897 49181 12909 49215
rect 12943 49212 12955 49215
rect 13446 49212 13452 49224
rect 12943 49184 13452 49212
rect 12943 49181 12955 49184
rect 12897 49175 12955 49181
rect 13446 49172 13452 49184
rect 13504 49172 13510 49224
rect 24857 49215 24915 49221
rect 24857 49181 24869 49215
rect 24903 49212 24915 49215
rect 25314 49212 25320 49224
rect 24903 49184 25320 49212
rect 24903 49181 24915 49184
rect 24857 49175 24915 49181
rect 25314 49172 25320 49184
rect 25372 49172 25378 49224
rect 22066 49116 25176 49144
rect 3329 49079 3387 49085
rect 3329 49076 3341 49079
rect 1780 49048 3341 49076
rect 3329 49045 3341 49048
rect 3375 49076 3387 49079
rect 10502 49076 10508 49088
rect 3375 49048 10508 49076
rect 3375 49045 3387 49048
rect 3329 49039 3387 49045
rect 10502 49036 10508 49048
rect 10560 49036 10566 49088
rect 18782 49036 18788 49088
rect 18840 49076 18846 49088
rect 22066 49076 22094 49116
rect 25148 49085 25176 49116
rect 18840 49048 22094 49076
rect 25133 49079 25191 49085
rect 18840 49036 18846 49048
rect 25133 49045 25145 49079
rect 25179 49045 25191 49079
rect 25133 49039 25191 49045
rect 1104 48986 25852 49008
rect 1104 48934 7950 48986
rect 8002 48934 8014 48986
rect 8066 48934 8078 48986
rect 8130 48934 8142 48986
rect 8194 48934 8206 48986
rect 8258 48934 17950 48986
rect 18002 48934 18014 48986
rect 18066 48934 18078 48986
rect 18130 48934 18142 48986
rect 18194 48934 18206 48986
rect 18258 48934 25852 48986
rect 1104 48912 25852 48934
rect 24489 48671 24547 48677
rect 24489 48637 24501 48671
rect 24535 48637 24547 48671
rect 24489 48631 24547 48637
rect 24504 48532 24532 48631
rect 24670 48628 24676 48680
rect 24728 48668 24734 48680
rect 24765 48671 24823 48677
rect 24765 48668 24777 48671
rect 24728 48640 24777 48668
rect 24728 48628 24734 48640
rect 24765 48637 24777 48640
rect 24811 48637 24823 48671
rect 24765 48631 24823 48637
rect 24762 48532 24768 48544
rect 24504 48504 24768 48532
rect 24762 48492 24768 48504
rect 24820 48492 24826 48544
rect 1104 48442 25852 48464
rect 1104 48390 2950 48442
rect 3002 48390 3014 48442
rect 3066 48390 3078 48442
rect 3130 48390 3142 48442
rect 3194 48390 3206 48442
rect 3258 48390 12950 48442
rect 13002 48390 13014 48442
rect 13066 48390 13078 48442
rect 13130 48390 13142 48442
rect 13194 48390 13206 48442
rect 13258 48390 22950 48442
rect 23002 48390 23014 48442
rect 23066 48390 23078 48442
rect 23130 48390 23142 48442
rect 23194 48390 23206 48442
rect 23258 48390 25852 48442
rect 1104 48368 25852 48390
rect 11698 48220 11704 48272
rect 11756 48260 11762 48272
rect 12710 48260 12716 48272
rect 11756 48232 12716 48260
rect 11756 48220 11762 48232
rect 12710 48220 12716 48232
rect 12768 48220 12774 48272
rect 18141 48263 18199 48269
rect 18141 48229 18153 48263
rect 18187 48260 18199 48263
rect 18414 48260 18420 48272
rect 18187 48232 18420 48260
rect 18187 48229 18199 48232
rect 18141 48223 18199 48229
rect 18414 48220 18420 48232
rect 18472 48220 18478 48272
rect 17129 48127 17187 48133
rect 17129 48093 17141 48127
rect 17175 48124 17187 48127
rect 18690 48124 18696 48136
rect 17175 48096 18696 48124
rect 17175 48093 17187 48096
rect 17129 48087 17187 48093
rect 18690 48084 18696 48096
rect 18748 48084 18754 48136
rect 16022 47948 16028 48000
rect 16080 47988 16086 48000
rect 17773 47991 17831 47997
rect 17773 47988 17785 47991
rect 16080 47960 17785 47988
rect 16080 47948 16086 47960
rect 17773 47957 17785 47960
rect 17819 47957 17831 47991
rect 17773 47951 17831 47957
rect 24762 47948 24768 48000
rect 24820 47988 24826 48000
rect 25225 47991 25283 47997
rect 25225 47988 25237 47991
rect 24820 47960 25237 47988
rect 24820 47948 24826 47960
rect 25225 47957 25237 47960
rect 25271 47957 25283 47991
rect 25225 47951 25283 47957
rect 25498 47948 25504 48000
rect 25556 47948 25562 48000
rect 1104 47898 25852 47920
rect 1104 47846 7950 47898
rect 8002 47846 8014 47898
rect 8066 47846 8078 47898
rect 8130 47846 8142 47898
rect 8194 47846 8206 47898
rect 8258 47846 17950 47898
rect 18002 47846 18014 47898
rect 18066 47846 18078 47898
rect 18130 47846 18142 47898
rect 18194 47846 18206 47898
rect 18258 47846 25852 47898
rect 1104 47824 25852 47846
rect 9214 47744 9220 47796
rect 9272 47744 9278 47796
rect 15930 47744 15936 47796
rect 15988 47784 15994 47796
rect 17221 47787 17279 47793
rect 17221 47784 17233 47787
rect 15988 47756 17233 47784
rect 15988 47744 15994 47756
rect 17221 47753 17233 47756
rect 17267 47753 17279 47787
rect 17221 47747 17279 47753
rect 17402 47744 17408 47796
rect 17460 47784 17466 47796
rect 18417 47787 18475 47793
rect 18417 47784 18429 47787
rect 17460 47756 18429 47784
rect 17460 47744 17466 47756
rect 18417 47753 18429 47756
rect 18463 47753 18475 47787
rect 18417 47747 18475 47753
rect 18506 47744 18512 47796
rect 18564 47784 18570 47796
rect 19058 47784 19064 47796
rect 18564 47756 19064 47784
rect 18564 47744 18570 47756
rect 19058 47744 19064 47756
rect 19116 47784 19122 47796
rect 19245 47787 19303 47793
rect 19245 47784 19257 47787
rect 19116 47756 19257 47784
rect 19116 47744 19122 47756
rect 19245 47753 19257 47756
rect 19291 47753 19303 47787
rect 19245 47747 19303 47753
rect 18966 47716 18972 47728
rect 18432 47688 18972 47716
rect 18432 47660 18460 47688
rect 18966 47676 18972 47688
rect 19024 47676 19030 47728
rect 19153 47719 19211 47725
rect 19153 47685 19165 47719
rect 19199 47716 19211 47719
rect 19426 47716 19432 47728
rect 19199 47688 19432 47716
rect 19199 47685 19211 47688
rect 19153 47679 19211 47685
rect 9401 47651 9459 47657
rect 9401 47617 9413 47651
rect 9447 47648 9459 47651
rect 11698 47648 11704 47660
rect 9447 47620 11704 47648
rect 9447 47617 9459 47620
rect 9401 47611 9459 47617
rect 11698 47608 11704 47620
rect 11756 47608 11762 47660
rect 17313 47651 17371 47657
rect 17313 47617 17325 47651
rect 17359 47648 17371 47651
rect 18414 47648 18420 47660
rect 17359 47620 18420 47648
rect 17359 47617 17371 47620
rect 17313 47611 17371 47617
rect 18414 47608 18420 47620
rect 18472 47608 18478 47660
rect 18506 47608 18512 47660
rect 18564 47648 18570 47660
rect 19168 47648 19196 47679
rect 19426 47676 19432 47688
rect 19484 47676 19490 47728
rect 18564 47620 19196 47648
rect 24489 47651 24547 47657
rect 18564 47608 18570 47620
rect 24489 47617 24501 47651
rect 24535 47648 24547 47651
rect 25498 47648 25504 47660
rect 24535 47620 25504 47648
rect 24535 47617 24547 47620
rect 24489 47611 24547 47617
rect 25498 47608 25504 47620
rect 25556 47608 25562 47660
rect 17402 47540 17408 47592
rect 17460 47540 17466 47592
rect 18690 47540 18696 47592
rect 18748 47540 18754 47592
rect 23290 47540 23296 47592
rect 23348 47580 23354 47592
rect 24765 47583 24823 47589
rect 24765 47580 24777 47583
rect 23348 47552 24777 47580
rect 23348 47540 23354 47552
rect 24765 47549 24777 47552
rect 24811 47549 24823 47583
rect 24765 47543 24823 47549
rect 11422 47404 11428 47456
rect 11480 47444 11486 47456
rect 11977 47447 12035 47453
rect 11977 47444 11989 47447
rect 11480 47416 11989 47444
rect 11480 47404 11486 47416
rect 11977 47413 11989 47416
rect 12023 47413 12035 47447
rect 11977 47407 12035 47413
rect 16574 47404 16580 47456
rect 16632 47444 16638 47456
rect 16853 47447 16911 47453
rect 16853 47444 16865 47447
rect 16632 47416 16865 47444
rect 16632 47404 16638 47416
rect 16853 47413 16865 47416
rect 16899 47413 16911 47447
rect 16853 47407 16911 47413
rect 17494 47404 17500 47456
rect 17552 47444 17558 47456
rect 18049 47447 18107 47453
rect 18049 47444 18061 47447
rect 17552 47416 18061 47444
rect 17552 47404 17558 47416
rect 18049 47413 18061 47416
rect 18095 47413 18107 47447
rect 18049 47407 18107 47413
rect 1104 47354 25852 47376
rect 1104 47302 2950 47354
rect 3002 47302 3014 47354
rect 3066 47302 3078 47354
rect 3130 47302 3142 47354
rect 3194 47302 3206 47354
rect 3258 47302 12950 47354
rect 13002 47302 13014 47354
rect 13066 47302 13078 47354
rect 13130 47302 13142 47354
rect 13194 47302 13206 47354
rect 13258 47302 22950 47354
rect 23002 47302 23014 47354
rect 23066 47302 23078 47354
rect 23130 47302 23142 47354
rect 23194 47302 23206 47354
rect 23258 47302 25852 47354
rect 1104 47280 25852 47302
rect 18141 47175 18199 47181
rect 18141 47141 18153 47175
rect 18187 47172 18199 47175
rect 18322 47172 18328 47184
rect 18187 47144 18328 47172
rect 18187 47141 18199 47144
rect 18141 47135 18199 47141
rect 18322 47132 18328 47144
rect 18380 47132 18386 47184
rect 10137 47107 10195 47113
rect 10137 47073 10149 47107
rect 10183 47104 10195 47107
rect 12158 47104 12164 47116
rect 10183 47076 12164 47104
rect 10183 47073 10195 47076
rect 10137 47067 10195 47073
rect 12158 47064 12164 47076
rect 12216 47064 12222 47116
rect 15749 47107 15807 47113
rect 15749 47073 15761 47107
rect 15795 47104 15807 47107
rect 16758 47104 16764 47116
rect 15795 47076 16764 47104
rect 15795 47073 15807 47076
rect 15749 47067 15807 47073
rect 16758 47064 16764 47076
rect 16816 47064 16822 47116
rect 17497 47107 17555 47113
rect 17497 47073 17509 47107
rect 17543 47104 17555 47107
rect 17586 47104 17592 47116
rect 17543 47076 17592 47104
rect 17543 47073 17555 47076
rect 17497 47067 17555 47073
rect 17586 47064 17592 47076
rect 17644 47064 17650 47116
rect 18598 47064 18604 47116
rect 18656 47064 18662 47116
rect 18785 47107 18843 47113
rect 18785 47073 18797 47107
rect 18831 47073 18843 47107
rect 18785 47067 18843 47073
rect 12345 47039 12403 47045
rect 12345 47036 12357 47039
rect 11900 47008 12357 47036
rect 4062 46928 4068 46980
rect 4120 46968 4126 46980
rect 9674 46968 9680 46980
rect 4120 46940 9680 46968
rect 4120 46928 4126 46940
rect 9674 46928 9680 46940
rect 9732 46928 9738 46980
rect 10413 46971 10471 46977
rect 10413 46937 10425 46971
rect 10459 46968 10471 46971
rect 10459 46940 10824 46968
rect 10459 46937 10471 46940
rect 10413 46931 10471 46937
rect 10796 46900 10824 46940
rect 11422 46928 11428 46980
rect 11480 46928 11486 46980
rect 11146 46900 11152 46912
rect 10796 46872 11152 46900
rect 11146 46860 11152 46872
rect 11204 46860 11210 46912
rect 11330 46860 11336 46912
rect 11388 46900 11394 46912
rect 11900 46909 11928 47008
rect 12345 47005 12357 47008
rect 12391 47005 12403 47039
rect 12345 46999 12403 47005
rect 18506 46996 18512 47048
rect 18564 46996 18570 47048
rect 18800 47036 18828 47067
rect 19429 47039 19487 47045
rect 19429 47036 19441 47039
rect 18800 47008 19441 47036
rect 19429 47005 19441 47008
rect 19475 47036 19487 47039
rect 19978 47036 19984 47048
rect 19475 47008 19984 47036
rect 19475 47005 19487 47008
rect 19429 46999 19487 47005
rect 19978 46996 19984 47008
rect 20036 46996 20042 47048
rect 20438 46996 20444 47048
rect 20496 47036 20502 47048
rect 20533 47039 20591 47045
rect 20533 47036 20545 47039
rect 20496 47008 20545 47036
rect 20496 46996 20502 47008
rect 20533 47005 20545 47008
rect 20579 47005 20591 47039
rect 20533 46999 20591 47005
rect 23201 47039 23259 47045
rect 23201 47005 23213 47039
rect 23247 47005 23259 47039
rect 23201 46999 23259 47005
rect 23477 47039 23535 47045
rect 23477 47005 23489 47039
rect 23523 47036 23535 47039
rect 23750 47036 23756 47048
rect 23523 47008 23756 47036
rect 23523 47005 23535 47008
rect 23477 46999 23535 47005
rect 16022 46928 16028 46980
rect 16080 46928 16086 46980
rect 17250 46940 17816 46968
rect 17788 46912 17816 46940
rect 18414 46928 18420 46980
rect 18472 46968 18478 46980
rect 20073 46971 20131 46977
rect 20073 46968 20085 46971
rect 18472 46940 20085 46968
rect 18472 46928 18478 46940
rect 20073 46937 20085 46940
rect 20119 46937 20131 46971
rect 23216 46968 23244 46999
rect 23750 46996 23756 47008
rect 23808 46996 23814 47048
rect 24394 46968 24400 46980
rect 23216 46940 24400 46968
rect 20073 46931 20131 46937
rect 24394 46928 24400 46940
rect 24452 46928 24458 46980
rect 24578 46928 24584 46980
rect 24636 46968 24642 46980
rect 25225 46971 25283 46977
rect 25225 46968 25237 46971
rect 24636 46940 25237 46968
rect 24636 46928 24642 46940
rect 25225 46937 25237 46940
rect 25271 46937 25283 46971
rect 25225 46931 25283 46937
rect 11885 46903 11943 46909
rect 11885 46900 11897 46903
rect 11388 46872 11897 46900
rect 11388 46860 11394 46872
rect 11885 46869 11897 46872
rect 11931 46869 11943 46903
rect 11885 46863 11943 46869
rect 12434 46860 12440 46912
rect 12492 46900 12498 46912
rect 12989 46903 13047 46909
rect 12989 46900 13001 46903
rect 12492 46872 13001 46900
rect 12492 46860 12498 46872
rect 12989 46869 13001 46872
rect 13035 46869 13047 46903
rect 12989 46863 13047 46869
rect 14182 46860 14188 46912
rect 14240 46900 14246 46912
rect 14277 46903 14335 46909
rect 14277 46900 14289 46903
rect 14240 46872 14289 46900
rect 14240 46860 14246 46872
rect 14277 46869 14289 46872
rect 14323 46900 14335 46903
rect 16390 46900 16396 46912
rect 14323 46872 16396 46900
rect 14323 46869 14335 46872
rect 14277 46863 14335 46869
rect 16390 46860 16396 46872
rect 16448 46860 16454 46912
rect 17770 46860 17776 46912
rect 17828 46860 17834 46912
rect 21174 46860 21180 46912
rect 21232 46860 21238 46912
rect 23842 46860 23848 46912
rect 23900 46900 23906 46912
rect 25409 46903 25467 46909
rect 25409 46900 25421 46903
rect 23900 46872 25421 46900
rect 23900 46860 23906 46872
rect 25409 46869 25421 46872
rect 25455 46869 25467 46903
rect 25409 46863 25467 46869
rect 1104 46810 25852 46832
rect 1104 46758 7950 46810
rect 8002 46758 8014 46810
rect 8066 46758 8078 46810
rect 8130 46758 8142 46810
rect 8194 46758 8206 46810
rect 8258 46758 17950 46810
rect 18002 46758 18014 46810
rect 18066 46758 18078 46810
rect 18130 46758 18142 46810
rect 18194 46758 18206 46810
rect 18258 46758 25852 46810
rect 1104 46736 25852 46758
rect 7285 46699 7343 46705
rect 7285 46665 7297 46699
rect 7331 46696 7343 46699
rect 7466 46696 7472 46708
rect 7331 46668 7472 46696
rect 7331 46665 7343 46668
rect 7285 46659 7343 46665
rect 7466 46656 7472 46668
rect 7524 46656 7530 46708
rect 11146 46656 11152 46708
rect 11204 46656 11210 46708
rect 11701 46699 11759 46705
rect 11701 46665 11713 46699
rect 11747 46696 11759 46699
rect 11882 46696 11888 46708
rect 11747 46668 11888 46696
rect 11747 46665 11759 46668
rect 11701 46659 11759 46665
rect 11882 46656 11888 46668
rect 11940 46656 11946 46708
rect 16301 46699 16359 46705
rect 16301 46665 16313 46699
rect 16347 46696 16359 46699
rect 16942 46696 16948 46708
rect 16347 46668 16948 46696
rect 16347 46665 16359 46668
rect 16301 46659 16359 46665
rect 16942 46656 16948 46668
rect 17000 46696 17006 46708
rect 17402 46696 17408 46708
rect 17000 46668 17408 46696
rect 17000 46656 17006 46668
rect 17402 46656 17408 46668
rect 17460 46656 17466 46708
rect 17770 46696 17776 46708
rect 17512 46668 17776 46696
rect 14182 46628 14188 46640
rect 13846 46600 14188 46628
rect 14182 46588 14188 46600
rect 14240 46588 14246 46640
rect 16390 46628 16396 46640
rect 16054 46600 16396 46628
rect 16390 46588 16396 46600
rect 16448 46628 16454 46640
rect 17512 46628 17540 46668
rect 17770 46656 17776 46668
rect 17828 46656 17834 46708
rect 18601 46699 18659 46705
rect 18601 46665 18613 46699
rect 18647 46696 18659 46699
rect 18690 46696 18696 46708
rect 18647 46668 18696 46696
rect 18647 46665 18659 46668
rect 18601 46659 18659 46665
rect 18690 46656 18696 46668
rect 18748 46656 18754 46708
rect 19429 46699 19487 46705
rect 19429 46665 19441 46699
rect 19475 46696 19487 46699
rect 19610 46696 19616 46708
rect 19475 46668 19616 46696
rect 19475 46665 19487 46668
rect 19429 46659 19487 46665
rect 19610 46656 19616 46668
rect 19668 46696 19674 46708
rect 20073 46699 20131 46705
rect 20073 46696 20085 46699
rect 19668 46668 20085 46696
rect 19668 46656 19674 46668
rect 20073 46665 20085 46668
rect 20119 46665 20131 46699
rect 20073 46659 20131 46665
rect 20165 46699 20223 46705
rect 20165 46665 20177 46699
rect 20211 46696 20223 46699
rect 20346 46696 20352 46708
rect 20211 46668 20352 46696
rect 20211 46665 20223 46668
rect 20165 46659 20223 46665
rect 20346 46656 20352 46668
rect 20404 46656 20410 46708
rect 20714 46656 20720 46708
rect 20772 46696 20778 46708
rect 21545 46699 21603 46705
rect 21545 46696 21557 46699
rect 20772 46668 21557 46696
rect 20772 46656 20778 46668
rect 21545 46665 21557 46668
rect 21591 46696 21603 46699
rect 22373 46699 22431 46705
rect 22373 46696 22385 46699
rect 21591 46668 22385 46696
rect 21591 46665 21603 46668
rect 21545 46659 21603 46665
rect 22373 46665 22385 46668
rect 22419 46665 22431 46699
rect 22373 46659 22431 46665
rect 22462 46656 22468 46708
rect 22520 46656 22526 46708
rect 16448 46600 17618 46628
rect 16448 46588 16454 46600
rect 7469 46563 7527 46569
rect 7469 46529 7481 46563
rect 7515 46560 7527 46563
rect 9490 46560 9496 46572
rect 7515 46532 9496 46560
rect 7515 46529 7527 46532
rect 7469 46523 7527 46529
rect 9490 46520 9496 46532
rect 9548 46520 9554 46572
rect 10505 46563 10563 46569
rect 10505 46529 10517 46563
rect 10551 46529 10563 46563
rect 10505 46523 10563 46529
rect 10520 46492 10548 46523
rect 10594 46520 10600 46572
rect 10652 46560 10658 46572
rect 11885 46563 11943 46569
rect 11885 46560 11897 46563
rect 10652 46532 11897 46560
rect 10652 46520 10658 46532
rect 11885 46529 11897 46532
rect 11931 46529 11943 46563
rect 11885 46523 11943 46529
rect 16758 46520 16764 46572
rect 16816 46560 16822 46572
rect 16853 46563 16911 46569
rect 16853 46560 16865 46563
rect 16816 46532 16865 46560
rect 16816 46520 16822 46532
rect 16853 46529 16865 46532
rect 16899 46529 16911 46563
rect 16853 46523 16911 46529
rect 10870 46492 10876 46504
rect 10520 46464 10876 46492
rect 10870 46452 10876 46464
rect 10928 46452 10934 46504
rect 12158 46452 12164 46504
rect 12216 46492 12222 46504
rect 12345 46495 12403 46501
rect 12345 46492 12357 46495
rect 12216 46464 12357 46492
rect 12216 46452 12222 46464
rect 12345 46461 12357 46464
rect 12391 46461 12403 46495
rect 12345 46455 12403 46461
rect 12621 46495 12679 46501
rect 12621 46461 12633 46495
rect 12667 46492 12679 46495
rect 14274 46492 14280 46504
rect 12667 46464 14280 46492
rect 12667 46461 12679 46464
rect 12621 46455 12679 46461
rect 14274 46452 14280 46464
rect 14332 46452 14338 46504
rect 14550 46452 14556 46504
rect 14608 46452 14614 46504
rect 14829 46495 14887 46501
rect 14829 46461 14841 46495
rect 14875 46492 14887 46495
rect 16482 46492 16488 46504
rect 14875 46464 16488 46492
rect 14875 46461 14887 46464
rect 14829 46455 14887 46461
rect 16482 46452 16488 46464
rect 16540 46452 16546 46504
rect 17129 46495 17187 46501
rect 17129 46461 17141 46495
rect 17175 46492 17187 46495
rect 18874 46492 18880 46504
rect 17175 46464 18880 46492
rect 17175 46461 17187 46464
rect 17129 46455 17187 46461
rect 18874 46452 18880 46464
rect 18932 46452 18938 46504
rect 20346 46452 20352 46504
rect 20404 46452 20410 46504
rect 22462 46452 22468 46504
rect 22520 46492 22526 46504
rect 22557 46495 22615 46501
rect 22557 46492 22569 46495
rect 22520 46464 22569 46492
rect 22520 46452 22526 46464
rect 22557 46461 22569 46464
rect 22603 46461 22615 46495
rect 22557 46455 22615 46461
rect 24489 46495 24547 46501
rect 24489 46461 24501 46495
rect 24535 46492 24547 46495
rect 24578 46492 24584 46504
rect 24535 46464 24584 46492
rect 24535 46461 24547 46464
rect 24489 46455 24547 46461
rect 24578 46452 24584 46464
rect 24636 46452 24642 46504
rect 24762 46452 24768 46504
rect 24820 46452 24826 46504
rect 14090 46316 14096 46368
rect 14148 46316 14154 46368
rect 18782 46316 18788 46368
rect 18840 46356 18846 46368
rect 18969 46359 19027 46365
rect 18969 46356 18981 46359
rect 18840 46328 18981 46356
rect 18840 46316 18846 46328
rect 18969 46325 18981 46328
rect 19015 46356 19027 46359
rect 19153 46359 19211 46365
rect 19153 46356 19165 46359
rect 19015 46328 19165 46356
rect 19015 46325 19027 46328
rect 18969 46319 19027 46325
rect 19153 46325 19165 46328
rect 19199 46325 19211 46359
rect 19153 46319 19211 46325
rect 19705 46359 19763 46365
rect 19705 46325 19717 46359
rect 19751 46356 19763 46359
rect 19794 46356 19800 46368
rect 19751 46328 19800 46356
rect 19751 46325 19763 46328
rect 19705 46319 19763 46325
rect 19794 46316 19800 46328
rect 19852 46316 19858 46368
rect 22005 46359 22063 46365
rect 22005 46325 22017 46359
rect 22051 46356 22063 46359
rect 22738 46356 22744 46368
rect 22051 46328 22744 46356
rect 22051 46325 22063 46328
rect 22005 46319 22063 46325
rect 22738 46316 22744 46328
rect 22796 46316 22802 46368
rect 24213 46359 24271 46365
rect 24213 46325 24225 46359
rect 24259 46356 24271 46359
rect 24486 46356 24492 46368
rect 24259 46328 24492 46356
rect 24259 46325 24271 46328
rect 24213 46319 24271 46325
rect 24486 46316 24492 46328
rect 24544 46316 24550 46368
rect 1104 46266 25852 46288
rect 1104 46214 2950 46266
rect 3002 46214 3014 46266
rect 3066 46214 3078 46266
rect 3130 46214 3142 46266
rect 3194 46214 3206 46266
rect 3258 46214 12950 46266
rect 13002 46214 13014 46266
rect 13066 46214 13078 46266
rect 13130 46214 13142 46266
rect 13194 46214 13206 46266
rect 13258 46214 22950 46266
rect 23002 46214 23014 46266
rect 23066 46214 23078 46266
rect 23130 46214 23142 46266
rect 23194 46214 23206 46266
rect 23258 46214 25852 46266
rect 1104 46192 25852 46214
rect 5626 46112 5632 46164
rect 5684 46152 5690 46164
rect 8113 46155 8171 46161
rect 8113 46152 8125 46155
rect 5684 46124 8125 46152
rect 5684 46112 5690 46124
rect 8113 46121 8125 46124
rect 8159 46121 8171 46155
rect 8113 46115 8171 46121
rect 9125 46155 9183 46161
rect 9125 46121 9137 46155
rect 9171 46152 9183 46155
rect 9306 46152 9312 46164
rect 9171 46124 9312 46152
rect 9171 46121 9183 46124
rect 9125 46115 9183 46121
rect 9306 46112 9312 46124
rect 9364 46112 9370 46164
rect 10686 46112 10692 46164
rect 10744 46112 10750 46164
rect 14182 46112 14188 46164
rect 14240 46112 14246 46164
rect 16482 46112 16488 46164
rect 16540 46112 16546 46164
rect 22005 46155 22063 46161
rect 22005 46121 22017 46155
rect 22051 46152 22063 46155
rect 22186 46152 22192 46164
rect 22051 46124 22192 46152
rect 22051 46121 22063 46124
rect 22005 46115 22063 46121
rect 22186 46112 22192 46124
rect 22244 46112 22250 46164
rect 7650 46044 7656 46096
rect 7708 46084 7714 46096
rect 10045 46087 10103 46093
rect 10045 46084 10057 46087
rect 7708 46056 10057 46084
rect 7708 46044 7714 46056
rect 10045 46053 10057 46056
rect 10091 46053 10103 46087
rect 16853 46087 16911 46093
rect 16853 46084 16865 46087
rect 10045 46047 10103 46053
rect 16500 46056 16865 46084
rect 16500 46028 16528 46056
rect 16853 46053 16865 46056
rect 16899 46053 16911 46087
rect 16853 46047 16911 46053
rect 11330 45976 11336 46028
rect 11388 45976 11394 46028
rect 11885 46019 11943 46025
rect 11885 45985 11897 46019
rect 11931 46016 11943 46019
rect 12158 46016 12164 46028
rect 11931 45988 12164 46016
rect 11931 45985 11943 45988
rect 11885 45979 11943 45985
rect 12158 45976 12164 45988
rect 12216 45976 12222 46028
rect 16482 45976 16488 46028
rect 16540 45976 16546 46028
rect 16758 45976 16764 46028
rect 16816 46016 16822 46028
rect 17129 46019 17187 46025
rect 17129 46016 17141 46019
rect 16816 45988 17141 46016
rect 16816 45976 16822 45988
rect 17129 45985 17141 45988
rect 17175 45985 17187 46019
rect 17129 45979 17187 45985
rect 17405 46019 17463 46025
rect 17405 45985 17417 46019
rect 17451 46016 17463 46019
rect 18414 46016 18420 46028
rect 17451 45988 18420 46016
rect 17451 45985 17463 45988
rect 17405 45979 17463 45985
rect 18414 45976 18420 45988
rect 18472 45976 18478 46028
rect 19797 46019 19855 46025
rect 19797 45985 19809 46019
rect 19843 46016 19855 46019
rect 21174 46016 21180 46028
rect 19843 45988 21180 46016
rect 19843 45985 19855 45988
rect 19797 45979 19855 45985
rect 21174 45976 21180 45988
rect 21232 45976 21238 46028
rect 21818 45976 21824 46028
rect 21876 46016 21882 46028
rect 22833 46019 22891 46025
rect 22833 46016 22845 46019
rect 21876 45988 22845 46016
rect 21876 45976 21882 45988
rect 22833 45985 22845 45988
rect 22879 45985 22891 46019
rect 22833 45979 22891 45985
rect 7006 45908 7012 45960
rect 7064 45948 7070 45960
rect 9309 45951 9367 45957
rect 9309 45948 9321 45951
rect 7064 45920 9321 45948
rect 7064 45908 7070 45920
rect 9309 45917 9321 45920
rect 9355 45917 9367 45951
rect 9309 45911 9367 45917
rect 10229 45951 10287 45957
rect 10229 45917 10241 45951
rect 10275 45917 10287 45951
rect 10229 45911 10287 45917
rect 11057 45951 11115 45957
rect 11057 45917 11069 45951
rect 11103 45948 11115 45951
rect 11514 45948 11520 45960
rect 11103 45920 11520 45948
rect 11103 45917 11115 45920
rect 11057 45911 11115 45917
rect 8021 45883 8079 45889
rect 8021 45849 8033 45883
rect 8067 45880 8079 45883
rect 10244 45880 10272 45911
rect 11514 45908 11520 45920
rect 11572 45908 11578 45960
rect 15841 45951 15899 45957
rect 15841 45917 15853 45951
rect 15887 45948 15899 45951
rect 15887 45920 16574 45948
rect 15887 45917 15899 45920
rect 15841 45911 15899 45917
rect 12161 45883 12219 45889
rect 8067 45852 8616 45880
rect 10244 45852 11376 45880
rect 8067 45849 8079 45852
rect 8021 45843 8079 45849
rect 8588 45821 8616 45852
rect 8573 45815 8631 45821
rect 8573 45781 8585 45815
rect 8619 45812 8631 45815
rect 8846 45812 8852 45824
rect 8619 45784 8852 45812
rect 8619 45781 8631 45784
rect 8573 45775 8631 45781
rect 8846 45772 8852 45784
rect 8904 45772 8910 45824
rect 11146 45772 11152 45824
rect 11204 45772 11210 45824
rect 11348 45812 11376 45852
rect 12161 45849 12173 45883
rect 12207 45880 12219 45883
rect 12434 45880 12440 45892
rect 12207 45852 12440 45880
rect 12207 45849 12219 45852
rect 12161 45843 12219 45849
rect 12434 45840 12440 45852
rect 12492 45840 12498 45892
rect 14182 45880 14188 45892
rect 13386 45852 14188 45880
rect 14182 45840 14188 45852
rect 14240 45840 14246 45892
rect 13170 45812 13176 45824
rect 11348 45784 13176 45812
rect 13170 45772 13176 45784
rect 13228 45772 13234 45824
rect 13633 45815 13691 45821
rect 13633 45781 13645 45815
rect 13679 45812 13691 45815
rect 13722 45812 13728 45824
rect 13679 45784 13728 45812
rect 13679 45781 13691 45784
rect 13633 45775 13691 45781
rect 13722 45772 13728 45784
rect 13780 45772 13786 45824
rect 16546 45812 16574 45920
rect 19518 45908 19524 45960
rect 19576 45908 19582 45960
rect 22186 45908 22192 45960
rect 22244 45948 22250 45960
rect 22649 45951 22707 45957
rect 22649 45948 22661 45951
rect 22244 45920 22661 45948
rect 22244 45908 22250 45920
rect 22649 45917 22661 45920
rect 22695 45917 22707 45951
rect 22649 45911 22707 45917
rect 22741 45951 22799 45957
rect 22741 45917 22753 45951
rect 22787 45948 22799 45951
rect 23934 45948 23940 45960
rect 22787 45920 23940 45948
rect 22787 45917 22799 45920
rect 22741 45911 22799 45917
rect 23934 45908 23940 45920
rect 23992 45908 23998 45960
rect 24026 45908 24032 45960
rect 24084 45948 24090 45960
rect 24581 45951 24639 45957
rect 24581 45948 24593 45951
rect 24084 45920 24593 45948
rect 24084 45908 24090 45920
rect 24581 45917 24593 45920
rect 24627 45917 24639 45951
rect 24581 45911 24639 45917
rect 18782 45880 18788 45892
rect 18630 45852 18788 45880
rect 18782 45840 18788 45852
rect 18840 45840 18846 45892
rect 21022 45852 21680 45880
rect 16758 45812 16764 45824
rect 16546 45784 16764 45812
rect 16758 45772 16764 45784
rect 16816 45772 16822 45824
rect 18690 45772 18696 45824
rect 18748 45812 18754 45824
rect 18877 45815 18935 45821
rect 18877 45812 18889 45815
rect 18748 45784 18889 45812
rect 18748 45772 18754 45784
rect 18877 45781 18889 45784
rect 18923 45781 18935 45815
rect 18877 45775 18935 45781
rect 19886 45772 19892 45824
rect 19944 45812 19950 45824
rect 21652 45821 21680 45852
rect 21269 45815 21327 45821
rect 21269 45812 21281 45815
rect 19944 45784 21281 45812
rect 19944 45772 19950 45784
rect 21269 45781 21281 45784
rect 21315 45781 21327 45815
rect 21269 45775 21327 45781
rect 21637 45815 21695 45821
rect 21637 45781 21649 45815
rect 21683 45812 21695 45815
rect 21726 45812 21732 45824
rect 21683 45784 21732 45812
rect 21683 45781 21695 45784
rect 21637 45775 21695 45781
rect 21726 45772 21732 45784
rect 21784 45772 21790 45824
rect 22281 45815 22339 45821
rect 22281 45781 22293 45815
rect 22327 45812 22339 45815
rect 22830 45812 22836 45824
rect 22327 45784 22836 45812
rect 22327 45781 22339 45784
rect 22281 45775 22339 45781
rect 22830 45772 22836 45784
rect 22888 45772 22894 45824
rect 23842 45772 23848 45824
rect 23900 45812 23906 45824
rect 23937 45815 23995 45821
rect 23937 45812 23949 45815
rect 23900 45784 23949 45812
rect 23900 45772 23906 45784
rect 23937 45781 23949 45784
rect 23983 45781 23995 45815
rect 23937 45775 23995 45781
rect 24210 45772 24216 45824
rect 24268 45772 24274 45824
rect 25222 45772 25228 45824
rect 25280 45772 25286 45824
rect 1104 45722 25852 45744
rect 1104 45670 7950 45722
rect 8002 45670 8014 45722
rect 8066 45670 8078 45722
rect 8130 45670 8142 45722
rect 8194 45670 8206 45722
rect 8258 45670 17950 45722
rect 18002 45670 18014 45722
rect 18066 45670 18078 45722
rect 18130 45670 18142 45722
rect 18194 45670 18206 45722
rect 18258 45670 25852 45722
rect 1104 45648 25852 45670
rect 4062 45568 4068 45620
rect 4120 45608 4126 45620
rect 8938 45608 8944 45620
rect 4120 45580 8944 45608
rect 4120 45568 4126 45580
rect 8938 45568 8944 45580
rect 8996 45568 9002 45620
rect 10226 45568 10232 45620
rect 10284 45608 10290 45620
rect 11885 45611 11943 45617
rect 11885 45608 11897 45611
rect 10284 45580 11897 45608
rect 10284 45568 10290 45580
rect 11885 45577 11897 45580
rect 11931 45577 11943 45611
rect 11885 45571 11943 45577
rect 19978 45568 19984 45620
rect 20036 45568 20042 45620
rect 21726 45608 21732 45620
rect 20272 45580 21732 45608
rect 8754 45500 8760 45552
rect 8812 45540 8818 45552
rect 9306 45540 9312 45552
rect 8812 45512 9312 45540
rect 8812 45500 8818 45512
rect 9306 45500 9312 45512
rect 9364 45540 9370 45552
rect 9401 45543 9459 45549
rect 9401 45540 9413 45543
rect 9364 45512 9413 45540
rect 9364 45500 9370 45512
rect 9401 45509 9413 45512
rect 9447 45509 9459 45543
rect 11422 45540 11428 45552
rect 10626 45512 11428 45540
rect 9401 45503 9459 45509
rect 11422 45500 11428 45512
rect 11480 45500 11486 45552
rect 13170 45500 13176 45552
rect 13228 45540 13234 45552
rect 13630 45540 13636 45552
rect 13228 45512 13636 45540
rect 13228 45500 13234 45512
rect 13630 45500 13636 45512
rect 13688 45500 13694 45552
rect 14550 45540 14556 45552
rect 14384 45512 14556 45540
rect 6822 45432 6828 45484
rect 6880 45472 6886 45484
rect 9125 45475 9183 45481
rect 9125 45472 9137 45475
rect 6880 45444 9137 45472
rect 6880 45432 6886 45444
rect 9125 45441 9137 45444
rect 9171 45441 9183 45475
rect 9125 45435 9183 45441
rect 9140 45268 9168 45435
rect 11790 45432 11796 45484
rect 11848 45472 11854 45484
rect 12253 45475 12311 45481
rect 12253 45472 12265 45475
rect 11848 45444 12265 45472
rect 11848 45432 11854 45444
rect 12253 45441 12265 45444
rect 12299 45441 12311 45475
rect 12253 45435 12311 45441
rect 13538 45432 13544 45484
rect 13596 45432 13602 45484
rect 14384 45416 14412 45512
rect 14550 45500 14556 45512
rect 14608 45500 14614 45552
rect 16482 45540 16488 45552
rect 15870 45512 16488 45540
rect 16482 45500 16488 45512
rect 16540 45500 16546 45552
rect 20272 45540 20300 45580
rect 21726 45568 21732 45580
rect 21784 45568 21790 45620
rect 19734 45512 20300 45540
rect 20898 45500 20904 45552
rect 20956 45500 20962 45552
rect 22278 45540 22284 45552
rect 22112 45512 22284 45540
rect 16853 45475 16911 45481
rect 16853 45441 16865 45475
rect 16899 45472 16911 45475
rect 16942 45472 16948 45484
rect 16899 45444 16948 45472
rect 16899 45441 16911 45444
rect 16853 45435 16911 45441
rect 16942 45432 16948 45444
rect 17000 45432 17006 45484
rect 22112 45481 22140 45512
rect 22278 45500 22284 45512
rect 22336 45500 22342 45552
rect 23842 45540 23848 45552
rect 23598 45512 23848 45540
rect 23842 45500 23848 45512
rect 23900 45500 23906 45552
rect 20809 45475 20867 45481
rect 20809 45441 20821 45475
rect 20855 45441 20867 45475
rect 20809 45435 20867 45441
rect 22097 45475 22155 45481
rect 22097 45441 22109 45475
rect 22143 45441 22155 45475
rect 25222 45472 25228 45484
rect 22097 45435 22155 45441
rect 23768 45444 25228 45472
rect 13633 45407 13691 45413
rect 13633 45373 13645 45407
rect 13679 45373 13691 45407
rect 13633 45367 13691 45373
rect 13725 45407 13783 45413
rect 13725 45373 13737 45407
rect 13771 45404 13783 45407
rect 13814 45404 13820 45416
rect 13771 45376 13820 45404
rect 13771 45373 13783 45376
rect 13725 45367 13783 45373
rect 11054 45336 11060 45348
rect 10428 45308 11060 45336
rect 10428 45268 10456 45308
rect 11054 45296 11060 45308
rect 11112 45336 11118 45348
rect 11149 45339 11207 45345
rect 11149 45336 11161 45339
rect 11112 45308 11161 45336
rect 11112 45296 11118 45308
rect 11149 45305 11161 45308
rect 11195 45305 11207 45339
rect 11149 45299 11207 45305
rect 13173 45339 13231 45345
rect 13173 45305 13185 45339
rect 13219 45336 13231 45339
rect 13446 45336 13452 45348
rect 13219 45308 13452 45336
rect 13219 45305 13231 45308
rect 13173 45299 13231 45305
rect 13446 45296 13452 45308
rect 13504 45296 13510 45348
rect 9140 45240 10456 45268
rect 10870 45228 10876 45280
rect 10928 45268 10934 45280
rect 12066 45268 12072 45280
rect 10928 45240 12072 45268
rect 10928 45228 10934 45240
rect 12066 45228 12072 45240
rect 12124 45228 12130 45280
rect 13648 45268 13676 45367
rect 13814 45364 13820 45376
rect 13872 45404 13878 45416
rect 14090 45404 14096 45416
rect 13872 45376 14096 45404
rect 13872 45364 13878 45376
rect 14090 45364 14096 45376
rect 14148 45364 14154 45416
rect 14366 45364 14372 45416
rect 14424 45364 14430 45416
rect 14645 45407 14703 45413
rect 14645 45373 14657 45407
rect 14691 45404 14703 45407
rect 17497 45407 17555 45413
rect 17497 45404 17509 45407
rect 14691 45376 17509 45404
rect 14691 45373 14703 45376
rect 14645 45367 14703 45373
rect 17497 45373 17509 45376
rect 17543 45373 17555 45407
rect 17497 45367 17555 45373
rect 18233 45407 18291 45413
rect 18233 45373 18245 45407
rect 18279 45373 18291 45407
rect 18233 45367 18291 45373
rect 15286 45268 15292 45280
rect 13648 45240 15292 45268
rect 15286 45228 15292 45240
rect 15344 45228 15350 45280
rect 16117 45271 16175 45277
rect 16117 45237 16129 45271
rect 16163 45268 16175 45271
rect 16298 45268 16304 45280
rect 16163 45240 16304 45268
rect 16163 45237 16175 45240
rect 16117 45231 16175 45237
rect 16298 45228 16304 45240
rect 16356 45228 16362 45280
rect 16482 45228 16488 45280
rect 16540 45228 16546 45280
rect 18248 45268 18276 45367
rect 18506 45364 18512 45416
rect 18564 45364 18570 45416
rect 19242 45364 19248 45416
rect 19300 45404 19306 45416
rect 20824 45404 20852 45435
rect 19300 45376 20852 45404
rect 21085 45407 21143 45413
rect 19300 45364 19306 45376
rect 21085 45373 21097 45407
rect 21131 45404 21143 45407
rect 21266 45404 21272 45416
rect 21131 45376 21272 45404
rect 21131 45373 21143 45376
rect 21085 45367 21143 45373
rect 21266 45364 21272 45376
rect 21324 45364 21330 45416
rect 22373 45407 22431 45413
rect 22373 45373 22385 45407
rect 22419 45404 22431 45407
rect 23768 45404 23796 45444
rect 25222 45432 25228 45444
rect 25280 45432 25286 45484
rect 22419 45376 23796 45404
rect 22419 45373 22431 45376
rect 22373 45367 22431 45373
rect 23842 45364 23848 45416
rect 23900 45404 23906 45416
rect 24121 45407 24179 45413
rect 24121 45404 24133 45407
rect 23900 45376 24133 45404
rect 23900 45364 23906 45376
rect 24121 45373 24133 45376
rect 24167 45373 24179 45407
rect 24121 45367 24179 45373
rect 24486 45364 24492 45416
rect 24544 45364 24550 45416
rect 24762 45364 24768 45416
rect 24820 45364 24826 45416
rect 21284 45336 21312 45364
rect 21284 45308 22094 45336
rect 19610 45268 19616 45280
rect 18248 45240 19616 45268
rect 19610 45228 19616 45240
rect 19668 45228 19674 45280
rect 20254 45228 20260 45280
rect 20312 45268 20318 45280
rect 20441 45271 20499 45277
rect 20441 45268 20453 45271
rect 20312 45240 20453 45268
rect 20312 45228 20318 45240
rect 20441 45237 20453 45240
rect 20487 45237 20499 45271
rect 20441 45231 20499 45237
rect 21545 45271 21603 45277
rect 21545 45237 21557 45271
rect 21591 45268 21603 45271
rect 21726 45268 21732 45280
rect 21591 45240 21732 45268
rect 21591 45237 21603 45240
rect 21545 45231 21603 45237
rect 21726 45228 21732 45240
rect 21784 45228 21790 45280
rect 22066 45268 22094 45308
rect 23845 45271 23903 45277
rect 23845 45268 23857 45271
rect 22066 45240 23857 45268
rect 23845 45237 23857 45240
rect 23891 45237 23903 45271
rect 23845 45231 23903 45237
rect 1104 45178 25852 45200
rect 1104 45126 2950 45178
rect 3002 45126 3014 45178
rect 3066 45126 3078 45178
rect 3130 45126 3142 45178
rect 3194 45126 3206 45178
rect 3258 45126 12950 45178
rect 13002 45126 13014 45178
rect 13066 45126 13078 45178
rect 13130 45126 13142 45178
rect 13194 45126 13206 45178
rect 13258 45126 22950 45178
rect 23002 45126 23014 45178
rect 23066 45126 23078 45178
rect 23130 45126 23142 45178
rect 23194 45126 23206 45178
rect 23258 45126 25852 45178
rect 1104 45104 25852 45126
rect 6454 45024 6460 45076
rect 6512 45064 6518 45076
rect 7837 45067 7895 45073
rect 7837 45064 7849 45067
rect 6512 45036 7849 45064
rect 6512 45024 6518 45036
rect 7837 45033 7849 45036
rect 7883 45033 7895 45067
rect 7837 45027 7895 45033
rect 8389 45067 8447 45073
rect 8389 45033 8401 45067
rect 8435 45064 8447 45067
rect 9398 45064 9404 45076
rect 8435 45036 9404 45064
rect 8435 45033 8447 45036
rect 8389 45027 8447 45033
rect 9398 45024 9404 45036
rect 9456 45024 9462 45076
rect 9858 45024 9864 45076
rect 9916 45064 9922 45076
rect 11241 45067 11299 45073
rect 11241 45064 11253 45067
rect 9916 45036 11253 45064
rect 9916 45024 9922 45036
rect 11241 45033 11253 45036
rect 11287 45033 11299 45067
rect 11241 45027 11299 45033
rect 18874 45024 18880 45076
rect 18932 45024 18938 45076
rect 20346 45024 20352 45076
rect 20404 45064 20410 45076
rect 21453 45067 21511 45073
rect 21453 45064 21465 45067
rect 20404 45036 21465 45064
rect 20404 45024 20410 45036
rect 21453 45033 21465 45036
rect 21499 45033 21511 45067
rect 21453 45027 21511 45033
rect 21726 45024 21732 45076
rect 21784 45064 21790 45076
rect 21821 45067 21879 45073
rect 21821 45064 21833 45067
rect 21784 45036 21833 45064
rect 21784 45024 21790 45036
rect 21821 45033 21833 45036
rect 21867 45064 21879 45067
rect 23842 45064 23848 45076
rect 21867 45036 23848 45064
rect 21867 45033 21879 45036
rect 21821 45027 21879 45033
rect 23842 45024 23848 45036
rect 23900 45024 23906 45076
rect 10318 44956 10324 45008
rect 10376 44996 10382 45008
rect 12437 44999 12495 45005
rect 12437 44996 12449 44999
rect 10376 44968 12449 44996
rect 10376 44956 10382 44968
rect 12437 44965 12449 44968
rect 12483 44965 12495 44999
rect 12437 44959 12495 44965
rect 7282 44888 7288 44940
rect 7340 44928 7346 44940
rect 9401 44931 9459 44937
rect 9401 44928 9413 44931
rect 7340 44900 9413 44928
rect 7340 44888 7346 44900
rect 9401 44897 9413 44900
rect 9447 44897 9459 44931
rect 9401 44891 9459 44897
rect 11422 44888 11428 44940
rect 11480 44928 11486 44940
rect 11885 44931 11943 44937
rect 11885 44928 11897 44931
rect 11480 44900 11897 44928
rect 11480 44888 11486 44900
rect 11885 44897 11897 44900
rect 11931 44928 11943 44931
rect 14090 44928 14096 44940
rect 11931 44900 14096 44928
rect 11931 44897 11943 44900
rect 11885 44891 11943 44897
rect 14090 44888 14096 44900
rect 14148 44888 14154 44940
rect 14366 44888 14372 44940
rect 14424 44928 14430 44940
rect 15105 44931 15163 44937
rect 15105 44928 15117 44931
rect 14424 44900 15117 44928
rect 14424 44888 14430 44900
rect 15105 44897 15117 44900
rect 15151 44928 15163 44931
rect 16850 44928 16856 44940
rect 15151 44900 16856 44928
rect 15151 44897 15163 44900
rect 15105 44891 15163 44897
rect 16850 44888 16856 44900
rect 16908 44888 16914 44940
rect 19981 44931 20039 44937
rect 19981 44897 19993 44931
rect 20027 44928 20039 44931
rect 21542 44928 21548 44940
rect 20027 44900 21548 44928
rect 20027 44897 20039 44900
rect 19981 44891 20039 44897
rect 21542 44888 21548 44900
rect 21600 44888 21606 44940
rect 22557 44931 22615 44937
rect 22557 44897 22569 44931
rect 22603 44928 22615 44931
rect 25225 44931 25283 44937
rect 25225 44928 25237 44931
rect 22603 44900 25237 44928
rect 22603 44897 22615 44900
rect 22557 44891 22615 44897
rect 25225 44897 25237 44900
rect 25271 44897 25283 44931
rect 25225 44891 25283 44897
rect 7650 44820 7656 44872
rect 7708 44860 7714 44872
rect 8573 44863 8631 44869
rect 8573 44860 8585 44863
rect 7708 44832 8585 44860
rect 7708 44820 7714 44832
rect 8573 44829 8585 44832
rect 8619 44829 8631 44863
rect 8573 44823 8631 44829
rect 13081 44863 13139 44869
rect 13081 44829 13093 44863
rect 13127 44860 13139 44863
rect 13814 44860 13820 44872
rect 13127 44832 13820 44860
rect 13127 44829 13139 44832
rect 13081 44823 13139 44829
rect 13814 44820 13820 44832
rect 13872 44820 13878 44872
rect 16482 44820 16488 44872
rect 16540 44860 16546 44872
rect 18233 44863 18291 44869
rect 16540 44832 17448 44860
rect 16540 44820 16546 44832
rect 7745 44795 7803 44801
rect 7745 44761 7757 44795
rect 7791 44761 7803 44795
rect 7745 44755 7803 44761
rect 9217 44795 9275 44801
rect 9217 44761 9229 44795
rect 9263 44792 9275 44795
rect 11149 44795 11207 44801
rect 9263 44764 9812 44792
rect 9263 44761 9275 44764
rect 9217 44755 9275 44761
rect 6457 44727 6515 44733
rect 6457 44693 6469 44727
rect 6503 44724 6515 44727
rect 6638 44724 6644 44736
rect 6503 44696 6644 44724
rect 6503 44693 6515 44696
rect 6457 44687 6515 44693
rect 6638 44684 6644 44696
rect 6696 44684 6702 44736
rect 7098 44684 7104 44736
rect 7156 44724 7162 44736
rect 7285 44727 7343 44733
rect 7285 44724 7297 44727
rect 7156 44696 7297 44724
rect 7156 44684 7162 44696
rect 7285 44693 7297 44696
rect 7331 44724 7343 44727
rect 7760 44724 7788 44755
rect 9784 44736 9812 44764
rect 11149 44761 11161 44795
rect 11195 44792 11207 44795
rect 12253 44795 12311 44801
rect 11195 44764 11652 44792
rect 11195 44761 11207 44764
rect 11149 44755 11207 44761
rect 11624 44736 11652 44764
rect 12253 44761 12265 44795
rect 12299 44792 12311 44795
rect 12713 44795 12771 44801
rect 12713 44792 12725 44795
rect 12299 44764 12725 44792
rect 12299 44761 12311 44764
rect 12253 44755 12311 44761
rect 12713 44761 12725 44764
rect 12759 44792 12771 44795
rect 14182 44792 14188 44804
rect 12759 44764 14188 44792
rect 12759 44761 12771 44764
rect 12713 44755 12771 44761
rect 14182 44752 14188 44764
rect 14240 44752 14246 44804
rect 15378 44752 15384 44804
rect 15436 44752 15442 44804
rect 16758 44752 16764 44804
rect 16816 44792 16822 44804
rect 17310 44792 17316 44804
rect 16816 44764 17316 44792
rect 16816 44752 16822 44764
rect 7331 44696 7788 44724
rect 7331 44693 7343 44696
rect 7285 44687 7343 44693
rect 9766 44684 9772 44736
rect 9824 44684 9830 44736
rect 11606 44684 11612 44736
rect 11664 44684 11670 44736
rect 12802 44684 12808 44736
rect 12860 44724 12866 44736
rect 16868 44733 16896 44764
rect 17310 44752 17316 44764
rect 17368 44752 17374 44804
rect 13725 44727 13783 44733
rect 13725 44724 13737 44727
rect 12860 44696 13737 44724
rect 12860 44684 12866 44696
rect 13725 44693 13737 44696
rect 13771 44693 13783 44727
rect 13725 44687 13783 44693
rect 16853 44727 16911 44733
rect 16853 44693 16865 44727
rect 16899 44693 16911 44727
rect 16853 44687 16911 44693
rect 17221 44727 17279 44733
rect 17221 44693 17233 44727
rect 17267 44724 17279 44727
rect 17420 44724 17448 44832
rect 18233 44829 18245 44863
rect 18279 44860 18291 44863
rect 18874 44860 18880 44872
rect 18279 44832 18880 44860
rect 18279 44829 18291 44832
rect 18233 44823 18291 44829
rect 18874 44820 18880 44832
rect 18932 44820 18938 44872
rect 19705 44863 19763 44869
rect 19705 44829 19717 44863
rect 19751 44829 19763 44863
rect 19705 44823 19763 44829
rect 18782 44724 18788 44736
rect 17267 44696 18788 44724
rect 17267 44693 17279 44696
rect 17221 44687 17279 44693
rect 18782 44684 18788 44696
rect 18840 44684 18846 44736
rect 19334 44684 19340 44736
rect 19392 44684 19398 44736
rect 19610 44684 19616 44736
rect 19668 44724 19674 44736
rect 19720 44724 19748 44823
rect 22278 44820 22284 44872
rect 22336 44820 22342 44872
rect 24118 44820 24124 44872
rect 24176 44860 24182 44872
rect 24581 44863 24639 44869
rect 24581 44860 24593 44863
rect 24176 44832 24593 44860
rect 24176 44820 24182 44832
rect 24581 44829 24593 44832
rect 24627 44829 24639 44863
rect 24581 44823 24639 44829
rect 21726 44792 21732 44804
rect 21206 44764 21732 44792
rect 21726 44752 21732 44764
rect 21784 44752 21790 44804
rect 23842 44792 23848 44804
rect 23782 44764 23848 44792
rect 23842 44752 23848 44764
rect 23900 44752 23906 44804
rect 22278 44724 22284 44736
rect 19668 44696 22284 44724
rect 19668 44684 19674 44696
rect 22278 44684 22284 44696
rect 22336 44684 22342 44736
rect 23382 44684 23388 44736
rect 23440 44724 23446 44736
rect 24026 44724 24032 44736
rect 23440 44696 24032 44724
rect 23440 44684 23446 44696
rect 24026 44684 24032 44696
rect 24084 44684 24090 44736
rect 1104 44634 25852 44656
rect 1104 44582 7950 44634
rect 8002 44582 8014 44634
rect 8066 44582 8078 44634
rect 8130 44582 8142 44634
rect 8194 44582 8206 44634
rect 8258 44582 17950 44634
rect 18002 44582 18014 44634
rect 18066 44582 18078 44634
rect 18130 44582 18142 44634
rect 18194 44582 18206 44634
rect 18258 44582 25852 44634
rect 1104 44560 25852 44582
rect 5810 44480 5816 44532
rect 5868 44480 5874 44532
rect 6730 44480 6736 44532
rect 6788 44480 6794 44532
rect 7190 44480 7196 44532
rect 7248 44520 7254 44532
rect 9033 44523 9091 44529
rect 9033 44520 9045 44523
rect 7248 44492 9045 44520
rect 7248 44480 7254 44492
rect 9033 44489 9045 44492
rect 9079 44489 9091 44523
rect 9033 44483 9091 44489
rect 10962 44480 10968 44532
rect 11020 44520 11026 44532
rect 11057 44523 11115 44529
rect 11057 44520 11069 44523
rect 11020 44492 11069 44520
rect 11020 44480 11026 44492
rect 11057 44489 11069 44492
rect 11103 44489 11115 44523
rect 11057 44483 11115 44489
rect 11146 44480 11152 44532
rect 11204 44520 11210 44532
rect 11885 44523 11943 44529
rect 11885 44520 11897 44523
rect 11204 44492 11897 44520
rect 11204 44480 11210 44492
rect 11885 44489 11897 44492
rect 11931 44489 11943 44523
rect 11885 44483 11943 44489
rect 12434 44480 12440 44532
rect 12492 44520 12498 44532
rect 13722 44520 13728 44532
rect 12492 44492 13728 44520
rect 12492 44480 12498 44492
rect 7558 44412 7564 44464
rect 7616 44412 7622 44464
rect 12158 44412 12164 44464
rect 12216 44452 12222 44464
rect 13372 44461 13400 44492
rect 13722 44480 13728 44492
rect 13780 44480 13786 44532
rect 15197 44523 15255 44529
rect 15197 44489 15209 44523
rect 15243 44520 15255 44523
rect 16482 44520 16488 44532
rect 15243 44492 16488 44520
rect 15243 44489 15255 44492
rect 15197 44483 15255 44489
rect 13357 44455 13415 44461
rect 12216 44424 13124 44452
rect 12216 44412 12222 44424
rect 5997 44387 6055 44393
rect 5997 44353 6009 44387
rect 6043 44384 6055 44387
rect 6546 44384 6552 44396
rect 6043 44356 6552 44384
rect 6043 44353 6055 44356
rect 5997 44347 6055 44353
rect 6546 44344 6552 44356
rect 6604 44344 6610 44396
rect 6638 44344 6644 44396
rect 6696 44344 6702 44396
rect 7377 44387 7435 44393
rect 7377 44353 7389 44387
rect 7423 44384 7435 44387
rect 7742 44384 7748 44396
rect 7423 44356 7748 44384
rect 7423 44353 7435 44356
rect 7377 44347 7435 44353
rect 7742 44344 7748 44356
rect 7800 44344 7806 44396
rect 8941 44387 8999 44393
rect 8941 44353 8953 44387
rect 8987 44384 8999 44387
rect 9214 44384 9220 44396
rect 8987 44356 9220 44384
rect 8987 44353 8999 44356
rect 8941 44347 8999 44353
rect 9214 44344 9220 44356
rect 9272 44344 9278 44396
rect 9861 44387 9919 44393
rect 9861 44353 9873 44387
rect 9907 44384 9919 44387
rect 10226 44384 10232 44396
rect 9907 44356 10232 44384
rect 9907 44353 9919 44356
rect 9861 44347 9919 44353
rect 10226 44344 10232 44356
rect 10284 44344 10290 44396
rect 13096 44393 13124 44424
rect 13357 44421 13369 44455
rect 13403 44421 13415 44455
rect 15212 44452 15240 44483
rect 16482 44480 16488 44492
rect 16540 44480 16546 44532
rect 18506 44480 18512 44532
rect 18564 44520 18570 44532
rect 20809 44523 20867 44529
rect 20809 44520 20821 44523
rect 18564 44492 20821 44520
rect 18564 44480 18570 44492
rect 20809 44489 20821 44492
rect 20855 44489 20867 44523
rect 20809 44483 20867 44489
rect 18782 44452 18788 44464
rect 14582 44438 15240 44452
rect 13357 44415 13415 44421
rect 14568 44424 15240 44438
rect 18354 44424 18788 44452
rect 10965 44387 11023 44393
rect 10965 44353 10977 44387
rect 11011 44384 11023 44387
rect 12253 44387 12311 44393
rect 11011 44356 11652 44384
rect 11011 44353 11023 44356
rect 10965 44347 11023 44353
rect 11624 44260 11652 44356
rect 12253 44353 12265 44387
rect 12299 44384 12311 44387
rect 13081 44387 13139 44393
rect 12299 44356 13032 44384
rect 12299 44353 12311 44356
rect 12253 44347 12311 44353
rect 12345 44319 12403 44325
rect 12345 44316 12357 44319
rect 11716 44288 12357 44316
rect 7374 44208 7380 44260
rect 7432 44248 7438 44260
rect 7432 44220 10364 44248
rect 7432 44208 7438 44220
rect 7742 44140 7748 44192
rect 7800 44180 7806 44192
rect 7837 44183 7895 44189
rect 7837 44180 7849 44183
rect 7800 44152 7849 44180
rect 7800 44140 7806 44152
rect 7837 44149 7849 44152
rect 7883 44149 7895 44183
rect 7837 44143 7895 44149
rect 9214 44140 9220 44192
rect 9272 44180 9278 44192
rect 10336 44189 10364 44220
rect 11606 44208 11612 44260
rect 11664 44208 11670 44260
rect 9401 44183 9459 44189
rect 9401 44180 9413 44183
rect 9272 44152 9413 44180
rect 9272 44140 9278 44152
rect 9401 44149 9413 44152
rect 9447 44149 9459 44183
rect 9401 44143 9459 44149
rect 10321 44183 10379 44189
rect 10321 44149 10333 44183
rect 10367 44149 10379 44183
rect 10321 44143 10379 44149
rect 10410 44140 10416 44192
rect 10468 44180 10474 44192
rect 11716 44180 11744 44288
rect 12345 44285 12357 44288
rect 12391 44285 12403 44319
rect 12345 44279 12403 44285
rect 12437 44319 12495 44325
rect 12437 44285 12449 44319
rect 12483 44285 12495 44319
rect 12437 44279 12495 44285
rect 12066 44208 12072 44260
rect 12124 44248 12130 44260
rect 12452 44248 12480 44279
rect 12124 44220 12480 44248
rect 12124 44208 12130 44220
rect 10468 44152 11744 44180
rect 13004 44180 13032 44356
rect 13081 44353 13093 44387
rect 13127 44353 13139 44387
rect 13081 44347 13139 44353
rect 14090 44276 14096 44328
rect 14148 44316 14154 44328
rect 14568 44316 14596 44424
rect 18782 44412 18788 44424
rect 18840 44412 18846 44464
rect 23842 44452 23848 44464
rect 23782 44424 23848 44452
rect 23842 44412 23848 44424
rect 23900 44412 23906 44464
rect 16850 44344 16856 44396
rect 16908 44344 16914 44396
rect 19061 44387 19119 44393
rect 19061 44353 19073 44387
rect 19107 44384 19119 44387
rect 19886 44384 19892 44396
rect 19107 44356 19892 44384
rect 19107 44353 19119 44356
rect 19061 44347 19119 44353
rect 19886 44344 19892 44356
rect 19944 44344 19950 44396
rect 20070 44344 20076 44396
rect 20128 44384 20134 44396
rect 20165 44387 20223 44393
rect 20165 44384 20177 44387
rect 20128 44356 20177 44384
rect 20128 44344 20134 44356
rect 20165 44353 20177 44356
rect 20211 44353 20223 44387
rect 20165 44347 20223 44353
rect 24302 44344 24308 44396
rect 24360 44384 24366 44396
rect 24765 44387 24823 44393
rect 24765 44384 24777 44387
rect 24360 44356 24777 44384
rect 24360 44344 24366 44356
rect 24765 44353 24777 44356
rect 24811 44353 24823 44387
rect 24765 44347 24823 44353
rect 14148 44288 14596 44316
rect 17129 44319 17187 44325
rect 14148 44276 14154 44288
rect 17129 44285 17141 44319
rect 17175 44316 17187 44319
rect 18506 44316 18512 44328
rect 17175 44288 18512 44316
rect 17175 44285 17187 44288
rect 17129 44279 17187 44285
rect 18506 44276 18512 44288
rect 18564 44316 18570 44328
rect 18690 44316 18696 44328
rect 18564 44288 18696 44316
rect 18564 44276 18570 44288
rect 18690 44276 18696 44288
rect 18748 44276 18754 44328
rect 22278 44276 22284 44328
rect 22336 44276 22342 44328
rect 22557 44319 22615 44325
rect 22557 44285 22569 44319
rect 22603 44316 22615 44319
rect 22646 44316 22652 44328
rect 22603 44288 22652 44316
rect 22603 44285 22615 44288
rect 22557 44279 22615 44285
rect 22646 44276 22652 44288
rect 22704 44276 22710 44328
rect 24489 44319 24547 44325
rect 24489 44285 24501 44319
rect 24535 44316 24547 44319
rect 24578 44316 24584 44328
rect 24535 44288 24584 44316
rect 24535 44285 24547 44288
rect 24489 44279 24547 44285
rect 24578 44276 24584 44288
rect 24636 44276 24642 44328
rect 14366 44180 14372 44192
rect 13004 44152 14372 44180
rect 10468 44140 10474 44152
rect 14366 44140 14372 44152
rect 14424 44140 14430 44192
rect 14458 44140 14464 44192
rect 14516 44180 14522 44192
rect 14826 44180 14832 44192
rect 14516 44152 14832 44180
rect 14516 44140 14522 44152
rect 14826 44140 14832 44152
rect 14884 44140 14890 44192
rect 16206 44140 16212 44192
rect 16264 44180 16270 44192
rect 16758 44180 16764 44192
rect 16264 44152 16764 44180
rect 16264 44140 16270 44152
rect 16758 44140 16764 44152
rect 16816 44140 16822 44192
rect 18601 44183 18659 44189
rect 18601 44149 18613 44183
rect 18647 44180 18659 44183
rect 18874 44180 18880 44192
rect 18647 44152 18880 44180
rect 18647 44149 18659 44152
rect 18601 44143 18659 44149
rect 18874 44140 18880 44152
rect 18932 44140 18938 44192
rect 19518 44140 19524 44192
rect 19576 44180 19582 44192
rect 19705 44183 19763 44189
rect 19705 44180 19717 44183
rect 19576 44152 19717 44180
rect 19576 44140 19582 44152
rect 19705 44149 19717 44152
rect 19751 44149 19763 44183
rect 19705 44143 19763 44149
rect 20806 44140 20812 44192
rect 20864 44180 20870 44192
rect 21910 44180 21916 44192
rect 20864 44152 21916 44180
rect 20864 44140 20870 44152
rect 21910 44140 21916 44152
rect 21968 44140 21974 44192
rect 24026 44140 24032 44192
rect 24084 44140 24090 44192
rect 1104 44090 25852 44112
rect 1104 44038 2950 44090
rect 3002 44038 3014 44090
rect 3066 44038 3078 44090
rect 3130 44038 3142 44090
rect 3194 44038 3206 44090
rect 3258 44038 12950 44090
rect 13002 44038 13014 44090
rect 13066 44038 13078 44090
rect 13130 44038 13142 44090
rect 13194 44038 13206 44090
rect 13258 44038 22950 44090
rect 23002 44038 23014 44090
rect 23066 44038 23078 44090
rect 23130 44038 23142 44090
rect 23194 44038 23206 44090
rect 23258 44038 25852 44090
rect 1104 44016 25852 44038
rect 4982 43936 4988 43988
rect 5040 43976 5046 43988
rect 6733 43979 6791 43985
rect 6733 43976 6745 43979
rect 5040 43948 6745 43976
rect 5040 43936 5046 43948
rect 6733 43945 6745 43948
rect 6779 43945 6791 43979
rect 6733 43939 6791 43945
rect 8386 43936 8392 43988
rect 8444 43936 8450 43988
rect 9950 43976 9956 43988
rect 8496 43948 9956 43976
rect 7193 43911 7251 43917
rect 7193 43877 7205 43911
rect 7239 43908 7251 43911
rect 8496 43908 8524 43948
rect 9950 43936 9956 43948
rect 10008 43936 10014 43988
rect 10502 43936 10508 43988
rect 10560 43976 10566 43988
rect 10873 43979 10931 43985
rect 10873 43976 10885 43979
rect 10560 43948 10885 43976
rect 10560 43936 10566 43948
rect 10873 43945 10885 43948
rect 10919 43945 10931 43979
rect 10873 43939 10931 43945
rect 11333 43979 11391 43985
rect 11333 43945 11345 43979
rect 11379 43976 11391 43979
rect 11422 43976 11428 43988
rect 11379 43948 11428 43976
rect 11379 43945 11391 43948
rect 11333 43939 11391 43945
rect 7239 43880 8524 43908
rect 7239 43877 7251 43880
rect 7193 43871 7251 43877
rect 6641 43775 6699 43781
rect 6641 43741 6653 43775
rect 6687 43772 6699 43775
rect 7208 43772 7236 43871
rect 9125 43843 9183 43849
rect 9125 43809 9137 43843
rect 9171 43840 9183 43843
rect 10870 43840 10876 43852
rect 9171 43812 10876 43840
rect 9171 43809 9183 43812
rect 9125 43803 9183 43809
rect 10870 43800 10876 43812
rect 10928 43800 10934 43852
rect 6687 43744 7236 43772
rect 8573 43775 8631 43781
rect 6687 43741 6699 43744
rect 6641 43735 6699 43741
rect 8573 43741 8585 43775
rect 8619 43772 8631 43775
rect 9030 43772 9036 43784
rect 8619 43744 9036 43772
rect 8619 43741 8631 43744
rect 8573 43735 8631 43741
rect 9030 43732 9036 43744
rect 9088 43732 9094 43784
rect 11348 43772 11376 43939
rect 11422 43936 11428 43948
rect 11480 43936 11486 43988
rect 21542 43936 21548 43988
rect 21600 43936 21606 43988
rect 15378 43868 15384 43920
rect 15436 43908 15442 43920
rect 15436 43880 17632 43908
rect 15436 43868 15442 43880
rect 17604 43852 17632 43880
rect 17678 43868 17684 43920
rect 17736 43908 17742 43920
rect 18141 43911 18199 43917
rect 18141 43908 18153 43911
rect 17736 43880 18153 43908
rect 17736 43868 17742 43880
rect 18141 43877 18153 43880
rect 18187 43908 18199 43911
rect 21634 43908 21640 43920
rect 18187 43880 21640 43908
rect 18187 43877 18199 43880
rect 18141 43871 18199 43877
rect 21634 43868 21640 43880
rect 21692 43868 21698 43920
rect 25130 43908 25136 43920
rect 21744 43880 25136 43908
rect 17494 43800 17500 43852
rect 17552 43800 17558 43852
rect 17586 43800 17592 43852
rect 17644 43800 17650 43852
rect 18325 43843 18383 43849
rect 18325 43809 18337 43843
rect 18371 43840 18383 43843
rect 21744 43840 21772 43880
rect 25130 43868 25136 43880
rect 25188 43868 25194 43920
rect 18371 43812 21772 43840
rect 18371 43809 18383 43812
rect 18325 43803 18383 43809
rect 10534 43744 11376 43772
rect 13814 43732 13820 43784
rect 13872 43772 13878 43784
rect 14277 43775 14335 43781
rect 14277 43772 14289 43775
rect 13872 43744 14289 43772
rect 13872 43732 13878 43744
rect 14277 43741 14289 43744
rect 14323 43741 14335 43775
rect 14277 43735 14335 43741
rect 15381 43775 15439 43781
rect 15381 43741 15393 43775
rect 15427 43772 15439 43775
rect 16298 43772 16304 43784
rect 15427 43744 16304 43772
rect 15427 43741 15439 43744
rect 15381 43735 15439 43741
rect 16298 43732 16304 43744
rect 16356 43732 16362 43784
rect 17402 43732 17408 43784
rect 17460 43772 17466 43784
rect 18340 43772 18368 43803
rect 22554 43800 22560 43852
rect 22612 43800 22618 43852
rect 22741 43843 22799 43849
rect 22741 43809 22753 43843
rect 22787 43840 22799 43843
rect 24486 43840 24492 43852
rect 22787 43812 24492 43840
rect 22787 43809 22799 43812
rect 22741 43803 22799 43809
rect 24486 43800 24492 43812
rect 24544 43800 24550 43852
rect 17460 43744 18368 43772
rect 19429 43775 19487 43781
rect 17460 43732 17466 43744
rect 19429 43741 19441 43775
rect 19475 43772 19487 43775
rect 20622 43772 20628 43784
rect 19475 43744 20628 43772
rect 19475 43741 19487 43744
rect 19429 43735 19487 43741
rect 20622 43732 20628 43744
rect 20680 43732 20686 43784
rect 20901 43775 20959 43781
rect 20901 43741 20913 43775
rect 20947 43772 20959 43775
rect 21174 43772 21180 43784
rect 20947 43744 21180 43772
rect 20947 43741 20959 43744
rect 20901 43735 20959 43741
rect 21174 43732 21180 43744
rect 21232 43732 21238 43784
rect 21266 43732 21272 43784
rect 21324 43772 21330 43784
rect 23293 43775 23351 43781
rect 23293 43772 23305 43775
rect 21324 43744 23305 43772
rect 21324 43732 21330 43744
rect 23293 43741 23305 43744
rect 23339 43741 23351 43775
rect 23293 43735 23351 43741
rect 24210 43732 24216 43784
rect 24268 43772 24274 43784
rect 24762 43772 24768 43784
rect 24268 43744 24768 43772
rect 24268 43732 24274 43744
rect 24762 43732 24768 43744
rect 24820 43772 24826 43784
rect 25317 43775 25375 43781
rect 25317 43772 25329 43775
rect 24820 43744 25329 43772
rect 24820 43732 24826 43744
rect 25317 43741 25329 43744
rect 25363 43741 25375 43775
rect 25317 43735 25375 43741
rect 9401 43707 9459 43713
rect 9401 43673 9413 43707
rect 9447 43673 9459 43707
rect 15838 43704 15844 43716
rect 9401 43667 9459 43673
rect 10796 43676 15844 43704
rect 9416 43636 9444 43667
rect 10796 43636 10824 43676
rect 15838 43664 15844 43676
rect 15896 43664 15902 43716
rect 20441 43707 20499 43713
rect 20441 43673 20453 43707
rect 20487 43704 20499 43707
rect 20487 43676 20944 43704
rect 20487 43673 20499 43676
rect 20441 43667 20499 43673
rect 20916 43648 20944 43676
rect 21910 43664 21916 43716
rect 21968 43704 21974 43716
rect 22465 43707 22523 43713
rect 22465 43704 22477 43707
rect 21968 43676 22477 43704
rect 21968 43664 21974 43676
rect 22465 43673 22477 43676
rect 22511 43673 22523 43707
rect 22465 43667 22523 43673
rect 23842 43664 23848 43716
rect 23900 43704 23906 43716
rect 23900 43676 24256 43704
rect 23900 43664 23906 43676
rect 24228 43648 24256 43676
rect 9416 43608 10824 43636
rect 14921 43639 14979 43645
rect 14921 43605 14933 43639
rect 14967 43636 14979 43639
rect 15010 43636 15016 43648
rect 14967 43608 15016 43636
rect 14967 43605 14979 43608
rect 14921 43599 14979 43605
rect 15010 43596 15016 43608
rect 15068 43596 15074 43648
rect 16022 43596 16028 43648
rect 16080 43596 16086 43648
rect 17037 43639 17095 43645
rect 17037 43605 17049 43639
rect 17083 43636 17095 43639
rect 17218 43636 17224 43648
rect 17083 43608 17224 43636
rect 17083 43605 17095 43608
rect 17037 43599 17095 43605
rect 17218 43596 17224 43608
rect 17276 43596 17282 43648
rect 18782 43596 18788 43648
rect 18840 43636 18846 43648
rect 19242 43636 19248 43648
rect 18840 43608 19248 43636
rect 18840 43596 18846 43608
rect 19242 43596 19248 43608
rect 19300 43596 19306 43648
rect 19334 43596 19340 43648
rect 19392 43636 19398 43648
rect 20073 43639 20131 43645
rect 20073 43636 20085 43639
rect 19392 43608 20085 43636
rect 19392 43596 19398 43608
rect 20073 43605 20085 43608
rect 20119 43605 20131 43639
rect 20073 43599 20131 43605
rect 20530 43596 20536 43648
rect 20588 43596 20594 43648
rect 20898 43596 20904 43648
rect 20956 43596 20962 43648
rect 22097 43639 22155 43645
rect 22097 43605 22109 43639
rect 22143 43636 22155 43639
rect 22186 43636 22192 43648
rect 22143 43608 22192 43636
rect 22143 43605 22155 43608
rect 22097 43599 22155 43605
rect 22186 43596 22192 43608
rect 22244 43596 22250 43648
rect 23934 43596 23940 43648
rect 23992 43596 23998 43648
rect 24210 43596 24216 43648
rect 24268 43636 24274 43648
rect 24489 43639 24547 43645
rect 24489 43636 24501 43639
rect 24268 43608 24501 43636
rect 24268 43596 24274 43608
rect 24489 43605 24501 43608
rect 24535 43636 24547 43639
rect 24673 43639 24731 43645
rect 24673 43636 24685 43639
rect 24535 43608 24685 43636
rect 24535 43605 24547 43608
rect 24489 43599 24547 43605
rect 24673 43605 24685 43608
rect 24719 43605 24731 43639
rect 24673 43599 24731 43605
rect 25133 43639 25191 43645
rect 25133 43605 25145 43639
rect 25179 43636 25191 43639
rect 25222 43636 25228 43648
rect 25179 43608 25228 43636
rect 25179 43605 25191 43608
rect 25133 43599 25191 43605
rect 25222 43596 25228 43608
rect 25280 43596 25286 43648
rect 1104 43546 25852 43568
rect 1104 43494 7950 43546
rect 8002 43494 8014 43546
rect 8066 43494 8078 43546
rect 8130 43494 8142 43546
rect 8194 43494 8206 43546
rect 8258 43494 17950 43546
rect 18002 43494 18014 43546
rect 18066 43494 18078 43546
rect 18130 43494 18142 43546
rect 18194 43494 18206 43546
rect 18258 43494 25852 43546
rect 1104 43472 25852 43494
rect 7745 43435 7803 43441
rect 7745 43401 7757 43435
rect 7791 43432 7803 43435
rect 7834 43432 7840 43444
rect 7791 43404 7840 43432
rect 7791 43401 7803 43404
rect 7745 43395 7803 43401
rect 7834 43392 7840 43404
rect 7892 43392 7898 43444
rect 9125 43435 9183 43441
rect 9125 43401 9137 43435
rect 9171 43432 9183 43435
rect 10410 43432 10416 43444
rect 9171 43404 10416 43432
rect 9171 43401 9183 43404
rect 9125 43395 9183 43401
rect 10410 43392 10416 43404
rect 10468 43392 10474 43444
rect 13722 43392 13728 43444
rect 13780 43432 13786 43444
rect 13780 43404 14596 43432
rect 13780 43392 13786 43404
rect 4614 43324 4620 43376
rect 4672 43364 4678 43376
rect 8665 43367 8723 43373
rect 8665 43364 8677 43367
rect 4672 43336 8677 43364
rect 4672 43324 4678 43336
rect 8665 43333 8677 43336
rect 8711 43333 8723 43367
rect 8665 43327 8723 43333
rect 9493 43367 9551 43373
rect 9493 43333 9505 43367
rect 9539 43364 9551 43367
rect 9582 43364 9588 43376
rect 9539 43336 9588 43364
rect 9539 43333 9551 43336
rect 9493 43327 9551 43333
rect 9582 43324 9588 43336
rect 9640 43324 9646 43376
rect 12802 43324 12808 43376
rect 12860 43324 12866 43376
rect 14090 43364 14096 43376
rect 14030 43336 14096 43364
rect 14090 43324 14096 43336
rect 14148 43324 14154 43376
rect 14568 43364 14596 43404
rect 14642 43392 14648 43444
rect 14700 43432 14706 43444
rect 15197 43435 15255 43441
rect 15197 43432 15209 43435
rect 14700 43404 15209 43432
rect 14700 43392 14706 43404
rect 15197 43401 15209 43404
rect 15243 43401 15255 43435
rect 15197 43395 15255 43401
rect 17313 43435 17371 43441
rect 17313 43401 17325 43435
rect 17359 43432 17371 43435
rect 17678 43432 17684 43444
rect 17359 43404 17684 43432
rect 17359 43401 17371 43404
rect 17313 43395 17371 43401
rect 17678 43392 17684 43404
rect 17736 43392 17742 43444
rect 22370 43392 22376 43444
rect 22428 43432 22434 43444
rect 22465 43435 22523 43441
rect 22465 43432 22477 43435
rect 22428 43404 22477 43432
rect 22428 43392 22434 43404
rect 22465 43401 22477 43404
rect 22511 43401 22523 43435
rect 22465 43395 22523 43401
rect 23293 43435 23351 43441
rect 23293 43401 23305 43435
rect 23339 43432 23351 43435
rect 24578 43432 24584 43444
rect 23339 43404 24584 43432
rect 23339 43401 23351 43404
rect 23293 43395 23351 43401
rect 24578 43392 24584 43404
rect 24636 43392 24642 43444
rect 14568 43336 16574 43364
rect 1302 43256 1308 43308
rect 1360 43296 1366 43308
rect 1673 43299 1731 43305
rect 1673 43296 1685 43299
rect 1360 43268 1685 43296
rect 1360 43256 1366 43268
rect 1673 43265 1685 43268
rect 1719 43296 1731 43299
rect 2133 43299 2191 43305
rect 2133 43296 2145 43299
rect 1719 43268 2145 43296
rect 1719 43265 1731 43268
rect 1673 43259 1731 43265
rect 2133 43265 2145 43268
rect 2179 43265 2191 43299
rect 2133 43259 2191 43265
rect 7650 43256 7656 43308
rect 7708 43296 7714 43308
rect 7929 43299 7987 43305
rect 7929 43296 7941 43299
rect 7708 43268 7941 43296
rect 7708 43256 7714 43268
rect 7929 43265 7941 43268
rect 7975 43265 7987 43299
rect 7929 43259 7987 43265
rect 8481 43299 8539 43305
rect 8481 43265 8493 43299
rect 8527 43265 8539 43299
rect 8481 43259 8539 43265
rect 8496 43228 8524 43259
rect 9306 43256 9312 43308
rect 9364 43296 9370 43308
rect 10137 43299 10195 43305
rect 10137 43296 10149 43299
rect 9364 43268 10149 43296
rect 9364 43256 9370 43268
rect 7484 43200 8524 43228
rect 1857 43163 1915 43169
rect 1857 43129 1869 43163
rect 1903 43160 1915 43163
rect 3510 43160 3516 43172
rect 1903 43132 3516 43160
rect 1903 43129 1915 43132
rect 1857 43123 1915 43129
rect 3510 43120 3516 43132
rect 3568 43120 3574 43172
rect 7484 43104 7512 43200
rect 8938 43188 8944 43240
rect 8996 43228 9002 43240
rect 9692 43237 9720 43268
rect 10137 43265 10149 43268
rect 10183 43296 10195 43299
rect 10226 43296 10232 43308
rect 10183 43268 10232 43296
rect 10183 43265 10195 43268
rect 10137 43259 10195 43265
rect 10226 43256 10232 43268
rect 10284 43256 10290 43308
rect 15289 43299 15347 43305
rect 15289 43265 15301 43299
rect 15335 43296 15347 43299
rect 15930 43296 15936 43308
rect 15335 43268 15936 43296
rect 15335 43265 15347 43268
rect 15289 43259 15347 43265
rect 15930 43256 15936 43268
rect 15988 43256 15994 43308
rect 16546 43296 16574 43336
rect 16850 43324 16856 43376
rect 16908 43364 16914 43376
rect 16908 43336 18276 43364
rect 16908 43324 16914 43336
rect 18248 43308 18276 43336
rect 19242 43324 19248 43376
rect 19300 43324 19306 43376
rect 21361 43367 21419 43373
rect 21361 43333 21373 43367
rect 21407 43364 21419 43367
rect 22278 43364 22284 43376
rect 21407 43336 22284 43364
rect 21407 43333 21419 43336
rect 21361 43327 21419 43333
rect 22278 43324 22284 43336
rect 22336 43364 22342 43376
rect 22336 43336 23520 43364
rect 22336 43324 22342 43336
rect 16546 43268 17632 43296
rect 9585 43231 9643 43237
rect 9585 43228 9597 43231
rect 8996 43200 9597 43228
rect 8996 43188 9002 43200
rect 9585 43197 9597 43200
rect 9631 43197 9643 43231
rect 9585 43191 9643 43197
rect 9677 43231 9735 43237
rect 9677 43197 9689 43231
rect 9723 43197 9735 43231
rect 9677 43191 9735 43197
rect 12529 43231 12587 43237
rect 12529 43197 12541 43231
rect 12575 43228 12587 43231
rect 14642 43228 14648 43240
rect 12575 43200 14648 43228
rect 12575 43197 12587 43200
rect 12529 43191 12587 43197
rect 14642 43188 14648 43200
rect 14700 43188 14706 43240
rect 17604 43237 17632 43268
rect 18230 43256 18236 43308
rect 18288 43256 18294 43308
rect 20162 43256 20168 43308
rect 20220 43296 20226 43308
rect 20530 43296 20536 43308
rect 20220 43268 20536 43296
rect 20220 43256 20226 43268
rect 20530 43256 20536 43268
rect 20588 43256 20594 43308
rect 21910 43256 21916 43308
rect 21968 43296 21974 43308
rect 22373 43299 22431 43305
rect 22373 43296 22385 43299
rect 21968 43268 22385 43296
rect 21968 43256 21974 43268
rect 22373 43265 22385 43268
rect 22419 43296 22431 43299
rect 23017 43299 23075 43305
rect 23017 43296 23029 43299
rect 22419 43268 23029 43296
rect 22419 43265 22431 43268
rect 22373 43259 22431 43265
rect 23017 43265 23029 43268
rect 23063 43265 23075 43299
rect 23017 43259 23075 43265
rect 23492 43240 23520 43336
rect 24118 43324 24124 43376
rect 24176 43364 24182 43376
rect 24176 43336 24334 43364
rect 24176 43324 24182 43336
rect 25130 43256 25136 43308
rect 25188 43296 25194 43308
rect 25590 43296 25596 43308
rect 25188 43268 25596 43296
rect 25188 43256 25194 43268
rect 25590 43256 25596 43268
rect 25648 43256 25654 43308
rect 15381 43231 15439 43237
rect 15381 43197 15393 43231
rect 15427 43197 15439 43231
rect 17405 43231 17463 43237
rect 17405 43228 17417 43231
rect 15381 43191 15439 43197
rect 16546 43200 17417 43228
rect 14090 43120 14096 43172
rect 14148 43160 14154 43172
rect 14277 43163 14335 43169
rect 14277 43160 14289 43163
rect 14148 43132 14289 43160
rect 14148 43120 14154 43132
rect 14277 43129 14289 43132
rect 14323 43129 14335 43163
rect 14277 43123 14335 43129
rect 14734 43120 14740 43172
rect 14792 43160 14798 43172
rect 15396 43160 15424 43191
rect 14792 43132 15424 43160
rect 15841 43163 15899 43169
rect 14792 43120 14798 43132
rect 15841 43129 15853 43163
rect 15887 43160 15899 43163
rect 16114 43160 16120 43172
rect 15887 43132 16120 43160
rect 15887 43129 15899 43132
rect 15841 43123 15899 43129
rect 16114 43120 16120 43132
rect 16172 43120 16178 43172
rect 7466 43052 7472 43104
rect 7524 43052 7530 43104
rect 14829 43095 14887 43101
rect 14829 43061 14841 43095
rect 14875 43092 14887 43095
rect 14918 43092 14924 43104
rect 14875 43064 14924 43092
rect 14875 43061 14887 43064
rect 14829 43055 14887 43061
rect 14918 43052 14924 43064
rect 14976 43052 14982 43104
rect 15930 43052 15936 43104
rect 15988 43092 15994 43104
rect 16025 43095 16083 43101
rect 16025 43092 16037 43095
rect 15988 43064 16037 43092
rect 15988 43052 15994 43064
rect 16025 43061 16037 43064
rect 16071 43061 16083 43095
rect 16025 43055 16083 43061
rect 16390 43052 16396 43104
rect 16448 43092 16454 43104
rect 16546 43092 16574 43200
rect 17405 43197 17417 43200
rect 17451 43197 17463 43231
rect 17405 43191 17463 43197
rect 17589 43231 17647 43237
rect 17589 43197 17601 43231
rect 17635 43228 17647 43231
rect 18509 43231 18567 43237
rect 17635 43200 18000 43228
rect 17635 43197 17647 43200
rect 17589 43191 17647 43197
rect 16448 43064 16574 43092
rect 16448 43052 16454 43064
rect 16942 43052 16948 43104
rect 17000 43052 17006 43104
rect 17972 43092 18000 43200
rect 18509 43197 18521 43231
rect 18555 43228 18567 43231
rect 19518 43228 19524 43240
rect 18555 43200 19524 43228
rect 18555 43197 18567 43200
rect 18509 43191 18567 43197
rect 19518 43188 19524 43200
rect 19576 43188 19582 43240
rect 22554 43188 22560 43240
rect 22612 43188 22618 43240
rect 23474 43188 23480 43240
rect 23532 43228 23538 43240
rect 23569 43231 23627 43237
rect 23569 43228 23581 43231
rect 23532 43200 23581 43228
rect 23532 43188 23538 43200
rect 23569 43197 23581 43200
rect 23615 43197 23627 43231
rect 23569 43191 23627 43197
rect 23842 43188 23848 43240
rect 23900 43188 23906 43240
rect 25406 43160 25412 43172
rect 24872 43132 25412 43160
rect 19518 43092 19524 43104
rect 17972 43064 19524 43092
rect 19518 43052 19524 43064
rect 19576 43052 19582 43104
rect 19981 43095 20039 43101
rect 19981 43061 19993 43095
rect 20027 43092 20039 43095
rect 20070 43092 20076 43104
rect 20027 43064 20076 43092
rect 20027 43061 20039 43064
rect 19981 43055 20039 43061
rect 20070 43052 20076 43064
rect 20128 43052 20134 43104
rect 22005 43095 22063 43101
rect 22005 43061 22017 43095
rect 22051 43092 22063 43095
rect 24872 43092 24900 43132
rect 25406 43120 25412 43132
rect 25464 43120 25470 43172
rect 22051 43064 24900 43092
rect 22051 43061 22063 43064
rect 22005 43055 22063 43061
rect 25314 43052 25320 43104
rect 25372 43052 25378 43104
rect 1104 43002 25852 43024
rect 1104 42950 2950 43002
rect 3002 42950 3014 43002
rect 3066 42950 3078 43002
rect 3130 42950 3142 43002
rect 3194 42950 3206 43002
rect 3258 42950 12950 43002
rect 13002 42950 13014 43002
rect 13066 42950 13078 43002
rect 13130 42950 13142 43002
rect 13194 42950 13206 43002
rect 13258 42950 22950 43002
rect 23002 42950 23014 43002
rect 23066 42950 23078 43002
rect 23130 42950 23142 43002
rect 23194 42950 23206 43002
rect 23258 42950 25852 43002
rect 1104 42928 25852 42950
rect 8938 42848 8944 42900
rect 8996 42848 9002 42900
rect 9217 42891 9275 42897
rect 9217 42857 9229 42891
rect 9263 42888 9275 42891
rect 9582 42888 9588 42900
rect 9263 42860 9588 42888
rect 9263 42857 9275 42860
rect 9217 42851 9275 42857
rect 9582 42848 9588 42860
rect 9640 42848 9646 42900
rect 9674 42848 9680 42900
rect 9732 42888 9738 42900
rect 11238 42888 11244 42900
rect 9732 42860 11244 42888
rect 9732 42848 9738 42860
rect 11238 42848 11244 42860
rect 11296 42888 11302 42900
rect 16390 42888 16396 42900
rect 11296 42860 16396 42888
rect 11296 42848 11302 42860
rect 16390 42848 16396 42860
rect 16448 42848 16454 42900
rect 16853 42891 16911 42897
rect 16853 42857 16865 42891
rect 16899 42888 16911 42891
rect 19242 42888 19248 42900
rect 16899 42860 19248 42888
rect 16899 42857 16911 42860
rect 16853 42851 16911 42857
rect 12989 42823 13047 42829
rect 12989 42820 13001 42823
rect 12268 42792 13001 42820
rect 4522 42712 4528 42764
rect 4580 42752 4586 42764
rect 4985 42755 5043 42761
rect 4985 42752 4997 42755
rect 4580 42724 4997 42752
rect 4580 42712 4586 42724
rect 4985 42721 4997 42724
rect 5031 42721 5043 42755
rect 4985 42715 5043 42721
rect 8478 42712 8484 42764
rect 8536 42752 8542 42764
rect 9401 42755 9459 42761
rect 9401 42752 9413 42755
rect 8536 42724 9413 42752
rect 8536 42712 8542 42724
rect 9401 42721 9413 42724
rect 9447 42721 9459 42755
rect 9401 42715 9459 42721
rect 10870 42712 10876 42764
rect 10928 42752 10934 42764
rect 12158 42752 12164 42764
rect 10928 42724 12164 42752
rect 10928 42712 10934 42724
rect 12158 42712 12164 42724
rect 12216 42712 12222 42764
rect 7837 42687 7895 42693
rect 7837 42653 7849 42687
rect 7883 42684 7895 42687
rect 8294 42684 8300 42696
rect 7883 42656 8300 42684
rect 7883 42653 7895 42656
rect 7837 42647 7895 42653
rect 8294 42644 8300 42656
rect 8352 42644 8358 42696
rect 9766 42644 9772 42696
rect 9824 42644 9830 42696
rect 12268 42670 12296 42792
rect 12989 42789 13001 42792
rect 13035 42820 13047 42823
rect 13998 42820 14004 42832
rect 13035 42792 14004 42820
rect 13035 42789 13047 42792
rect 12989 42783 13047 42789
rect 13998 42780 14004 42792
rect 14056 42780 14062 42832
rect 16485 42823 16543 42829
rect 16485 42789 16497 42823
rect 16531 42820 16543 42823
rect 16574 42820 16580 42832
rect 16531 42792 16580 42820
rect 16531 42789 16543 42792
rect 16485 42783 16543 42789
rect 16574 42780 16580 42792
rect 16632 42780 16638 42832
rect 12342 42712 12348 42764
rect 12400 42752 12406 42764
rect 12621 42755 12679 42761
rect 12621 42752 12633 42755
rect 12400 42724 12633 42752
rect 12400 42712 12406 42724
rect 12621 42721 12633 42724
rect 12667 42752 12679 42755
rect 13814 42752 13820 42764
rect 12667 42724 13820 42752
rect 12667 42721 12679 42724
rect 12621 42715 12679 42721
rect 13814 42712 13820 42724
rect 13872 42712 13878 42764
rect 14642 42712 14648 42764
rect 14700 42752 14706 42764
rect 14737 42755 14795 42761
rect 14737 42752 14749 42755
rect 14700 42724 14749 42752
rect 14700 42712 14706 42724
rect 14737 42721 14749 42724
rect 14783 42752 14795 42755
rect 16850 42752 16856 42764
rect 14783 42724 16856 42752
rect 14783 42721 14795 42724
rect 14737 42715 14795 42721
rect 16850 42712 16856 42724
rect 16908 42712 16914 42764
rect 16114 42644 16120 42696
rect 16172 42684 16178 42696
rect 16482 42684 16488 42696
rect 16172 42656 16488 42684
rect 16172 42644 16178 42656
rect 16482 42644 16488 42656
rect 16540 42684 16546 42696
rect 16960 42684 16988 42860
rect 19242 42848 19248 42860
rect 19300 42848 19306 42900
rect 19876 42891 19934 42897
rect 19876 42857 19888 42891
rect 19922 42888 19934 42891
rect 23934 42888 23940 42900
rect 19922 42860 23940 42888
rect 19922 42857 19934 42860
rect 19876 42851 19934 42857
rect 23934 42848 23940 42860
rect 23992 42848 23998 42900
rect 24118 42848 24124 42900
rect 24176 42888 24182 42900
rect 24946 42888 24952 42900
rect 24176 42860 24952 42888
rect 24176 42848 24182 42860
rect 24946 42848 24952 42860
rect 25004 42848 25010 42900
rect 22370 42780 22376 42832
rect 22428 42820 22434 42832
rect 24026 42820 24032 42832
rect 22428 42792 24032 42820
rect 22428 42780 22434 42792
rect 17586 42712 17592 42764
rect 17644 42752 17650 42764
rect 22002 42752 22008 42764
rect 17644 42724 22008 42752
rect 17644 42712 17650 42724
rect 22002 42712 22008 42724
rect 22060 42712 22066 42764
rect 22480 42761 22508 42792
rect 24026 42780 24032 42792
rect 24084 42780 24090 42832
rect 22465 42755 22523 42761
rect 22465 42721 22477 42755
rect 22511 42721 22523 42755
rect 22465 42715 22523 42721
rect 23014 42712 23020 42764
rect 23072 42752 23078 42764
rect 23477 42755 23535 42761
rect 23477 42752 23489 42755
rect 23072 42724 23489 42752
rect 23072 42712 23078 42724
rect 23477 42721 23489 42724
rect 23523 42721 23535 42755
rect 23477 42715 23535 42721
rect 16540 42656 16988 42684
rect 16540 42644 16546 42656
rect 18230 42644 18236 42696
rect 18288 42684 18294 42696
rect 18693 42687 18751 42693
rect 18693 42684 18705 42687
rect 18288 42656 18705 42684
rect 18288 42644 18294 42656
rect 18693 42653 18705 42656
rect 18739 42684 18751 42687
rect 18782 42684 18788 42696
rect 18739 42656 18788 42684
rect 18739 42653 18751 42656
rect 18693 42647 18751 42653
rect 18782 42644 18788 42656
rect 18840 42644 18846 42696
rect 19610 42644 19616 42696
rect 19668 42644 19674 42696
rect 22925 42687 22983 42693
rect 22925 42653 22937 42687
rect 22971 42684 22983 42687
rect 23198 42684 23204 42696
rect 22971 42656 23204 42684
rect 22971 42653 22983 42656
rect 22925 42647 22983 42653
rect 23198 42644 23204 42656
rect 23256 42644 23262 42696
rect 24673 42687 24731 42693
rect 24673 42653 24685 42687
rect 24719 42684 24731 42687
rect 25130 42684 25136 42696
rect 24719 42656 25136 42684
rect 24719 42653 24731 42656
rect 24673 42647 24731 42653
rect 25130 42644 25136 42656
rect 25188 42684 25194 42696
rect 25314 42684 25320 42696
rect 25188 42656 25320 42684
rect 25188 42644 25194 42656
rect 25314 42644 25320 42656
rect 25372 42644 25378 42696
rect 4801 42619 4859 42625
rect 4801 42585 4813 42619
rect 4847 42616 4859 42619
rect 10413 42619 10471 42625
rect 4847 42588 5396 42616
rect 4847 42585 4859 42588
rect 4801 42579 4859 42585
rect 5368 42557 5396 42588
rect 10413 42585 10425 42619
rect 10459 42616 10471 42619
rect 11149 42619 11207 42625
rect 11149 42616 11161 42619
rect 10459 42588 11161 42616
rect 10459 42585 10471 42588
rect 10413 42579 10471 42585
rect 11149 42585 11161 42588
rect 11195 42585 11207 42619
rect 11149 42579 11207 42585
rect 15010 42576 15016 42628
rect 15068 42576 15074 42628
rect 17126 42576 17132 42628
rect 17184 42616 17190 42628
rect 17681 42619 17739 42625
rect 17681 42616 17693 42619
rect 17184 42588 17693 42616
rect 17184 42576 17190 42588
rect 17681 42585 17693 42588
rect 17727 42616 17739 42619
rect 17957 42619 18015 42625
rect 17957 42616 17969 42619
rect 17727 42588 17969 42616
rect 17727 42585 17739 42588
rect 17681 42579 17739 42585
rect 17957 42585 17969 42588
rect 18003 42616 18015 42619
rect 20162 42616 20168 42628
rect 18003 42588 20168 42616
rect 18003 42585 18015 42588
rect 17957 42579 18015 42585
rect 20162 42576 20168 42588
rect 20220 42576 20226 42628
rect 20898 42576 20904 42628
rect 20956 42576 20962 42628
rect 22281 42619 22339 42625
rect 22281 42585 22293 42619
rect 22327 42616 22339 42619
rect 22738 42616 22744 42628
rect 22327 42588 22744 42616
rect 22327 42585 22339 42588
rect 22281 42579 22339 42585
rect 22738 42576 22744 42588
rect 22796 42576 22802 42628
rect 5353 42551 5411 42557
rect 5353 42517 5365 42551
rect 5399 42548 5411 42551
rect 6730 42548 6736 42560
rect 5399 42520 6736 42548
rect 5399 42517 5411 42520
rect 5353 42511 5411 42517
rect 6730 42508 6736 42520
rect 6788 42508 6794 42560
rect 7834 42508 7840 42560
rect 7892 42548 7898 42560
rect 8481 42551 8539 42557
rect 8481 42548 8493 42551
rect 7892 42520 8493 42548
rect 7892 42508 7898 42520
rect 8481 42517 8493 42520
rect 8527 42517 8539 42551
rect 8481 42511 8539 42517
rect 20622 42508 20628 42560
rect 20680 42548 20686 42560
rect 21361 42551 21419 42557
rect 21361 42548 21373 42551
rect 20680 42520 21373 42548
rect 20680 42508 20686 42520
rect 21361 42517 21373 42520
rect 21407 42517 21419 42551
rect 21361 42511 21419 42517
rect 21542 42508 21548 42560
rect 21600 42548 21606 42560
rect 21821 42551 21879 42557
rect 21821 42548 21833 42551
rect 21600 42520 21833 42548
rect 21600 42508 21606 42520
rect 21821 42517 21833 42520
rect 21867 42517 21879 42551
rect 21821 42511 21879 42517
rect 22002 42508 22008 42560
rect 22060 42548 22066 42560
rect 22189 42551 22247 42557
rect 22189 42548 22201 42551
rect 22060 42520 22201 42548
rect 22060 42508 22066 42520
rect 22189 42517 22201 42520
rect 22235 42517 22247 42551
rect 22189 42511 22247 42517
rect 23750 42508 23756 42560
rect 23808 42548 23814 42560
rect 25317 42551 25375 42557
rect 25317 42548 25329 42551
rect 23808 42520 25329 42548
rect 23808 42508 23814 42520
rect 25317 42517 25329 42520
rect 25363 42517 25375 42551
rect 25317 42511 25375 42517
rect 1104 42458 25852 42480
rect 1104 42406 7950 42458
rect 8002 42406 8014 42458
rect 8066 42406 8078 42458
rect 8130 42406 8142 42458
rect 8194 42406 8206 42458
rect 8258 42406 17950 42458
rect 18002 42406 18014 42458
rect 18066 42406 18078 42458
rect 18130 42406 18142 42458
rect 18194 42406 18206 42458
rect 18258 42406 25852 42458
rect 1104 42384 25852 42406
rect 4338 42304 4344 42356
rect 4396 42344 4402 42356
rect 5813 42347 5871 42353
rect 5813 42344 5825 42347
rect 4396 42316 5825 42344
rect 4396 42304 4402 42316
rect 5813 42313 5825 42316
rect 5859 42313 5871 42347
rect 5813 42307 5871 42313
rect 9490 42304 9496 42356
rect 9548 42344 9554 42356
rect 9769 42347 9827 42353
rect 9769 42344 9781 42347
rect 9548 42316 9781 42344
rect 9548 42304 9554 42316
rect 9769 42313 9781 42316
rect 9815 42313 9827 42347
rect 9769 42307 9827 42313
rect 11054 42304 11060 42356
rect 11112 42304 11118 42356
rect 11698 42304 11704 42356
rect 11756 42304 11762 42356
rect 12897 42347 12955 42353
rect 12897 42313 12909 42347
rect 12943 42344 12955 42347
rect 13538 42344 13544 42356
rect 12943 42316 13544 42344
rect 12943 42313 12955 42316
rect 12897 42307 12955 42313
rect 13538 42304 13544 42316
rect 13596 42304 13602 42356
rect 15286 42304 15292 42356
rect 15344 42304 15350 42356
rect 15749 42347 15807 42353
rect 15749 42313 15761 42347
rect 15795 42344 15807 42347
rect 16942 42344 16948 42356
rect 15795 42316 16948 42344
rect 15795 42313 15807 42316
rect 15749 42307 15807 42313
rect 16942 42304 16948 42316
rect 17000 42304 17006 42356
rect 17129 42347 17187 42353
rect 17129 42313 17141 42347
rect 17175 42313 17187 42347
rect 17129 42307 17187 42313
rect 17589 42347 17647 42353
rect 17589 42313 17601 42347
rect 17635 42344 17647 42347
rect 18233 42347 18291 42353
rect 18233 42344 18245 42347
rect 17635 42316 18245 42344
rect 17635 42313 17647 42316
rect 17589 42307 17647 42313
rect 18233 42313 18245 42316
rect 18279 42344 18291 42347
rect 18598 42344 18604 42356
rect 18279 42316 18604 42344
rect 18279 42313 18291 42316
rect 18233 42307 18291 42313
rect 7834 42236 7840 42288
rect 7892 42236 7898 42288
rect 8478 42236 8484 42288
rect 8536 42236 8542 42288
rect 10229 42279 10287 42285
rect 10229 42245 10241 42279
rect 10275 42276 10287 42279
rect 12158 42276 12164 42288
rect 10275 42248 12164 42276
rect 10275 42245 10287 42248
rect 10229 42239 10287 42245
rect 12158 42236 12164 42248
rect 12216 42236 12222 42288
rect 13357 42279 13415 42285
rect 13357 42245 13369 42279
rect 13403 42276 13415 42279
rect 13446 42276 13452 42288
rect 13403 42248 13452 42276
rect 13403 42245 13415 42248
rect 13357 42239 13415 42245
rect 13446 42236 13452 42248
rect 13504 42236 13510 42288
rect 14366 42236 14372 42288
rect 14424 42276 14430 42288
rect 17144 42276 17172 42307
rect 18598 42304 18604 42316
rect 18656 42304 18662 42356
rect 22002 42304 22008 42356
rect 22060 42344 22066 42356
rect 22186 42344 22192 42356
rect 22060 42316 22192 42344
rect 22060 42304 22066 42316
rect 22186 42304 22192 42316
rect 22244 42304 22250 42356
rect 22646 42304 22652 42356
rect 22704 42344 22710 42356
rect 23017 42347 23075 42353
rect 23017 42344 23029 42347
rect 22704 42316 23029 42344
rect 22704 42304 22710 42316
rect 23017 42313 23029 42316
rect 23063 42313 23075 42347
rect 23017 42307 23075 42313
rect 24486 42304 24492 42356
rect 24544 42344 24550 42356
rect 25225 42347 25283 42353
rect 25225 42344 25237 42347
rect 24544 42316 25237 42344
rect 24544 42304 24550 42316
rect 25225 42313 25237 42316
rect 25271 42313 25283 42347
rect 25225 42307 25283 42313
rect 19061 42279 19119 42285
rect 14424 42248 17172 42276
rect 17420 42248 18736 42276
rect 14424 42236 14430 42248
rect 5353 42211 5411 42217
rect 5353 42177 5365 42211
rect 5399 42208 5411 42211
rect 5721 42211 5779 42217
rect 5721 42208 5733 42211
rect 5399 42180 5733 42208
rect 5399 42177 5411 42180
rect 5353 42171 5411 42177
rect 5721 42177 5733 42180
rect 5767 42208 5779 42211
rect 5902 42208 5908 42220
rect 5767 42180 5908 42208
rect 5767 42177 5779 42180
rect 5721 42171 5779 42177
rect 5902 42168 5908 42180
rect 5960 42168 5966 42220
rect 6822 42168 6828 42220
rect 6880 42208 6886 42220
rect 7561 42211 7619 42217
rect 7561 42208 7573 42211
rect 6880 42180 7573 42208
rect 6880 42168 6886 42180
rect 7561 42177 7573 42180
rect 7607 42177 7619 42211
rect 7561 42171 7619 42177
rect 10134 42168 10140 42220
rect 10192 42168 10198 42220
rect 10502 42168 10508 42220
rect 10560 42208 10566 42220
rect 12069 42211 12127 42217
rect 12069 42208 12081 42211
rect 10560 42180 12081 42208
rect 10560 42168 10566 42180
rect 12069 42177 12081 42180
rect 12115 42177 12127 42211
rect 12069 42171 12127 42177
rect 13265 42211 13323 42217
rect 13265 42177 13277 42211
rect 13311 42208 13323 42211
rect 14093 42211 14151 42217
rect 14093 42208 14105 42211
rect 13311 42180 14105 42208
rect 13311 42177 13323 42180
rect 13265 42171 13323 42177
rect 14093 42177 14105 42180
rect 14139 42177 14151 42211
rect 14093 42171 14151 42177
rect 15657 42211 15715 42217
rect 15657 42177 15669 42211
rect 15703 42208 15715 42211
rect 17420 42208 17448 42248
rect 15703 42180 17448 42208
rect 15703 42177 15715 42180
rect 15657 42171 15715 42177
rect 17494 42168 17500 42220
rect 17552 42168 17558 42220
rect 9309 42143 9367 42149
rect 9309 42109 9321 42143
rect 9355 42140 9367 42143
rect 9766 42140 9772 42152
rect 9355 42112 9772 42140
rect 9355 42109 9367 42112
rect 9309 42103 9367 42109
rect 9766 42100 9772 42112
rect 9824 42100 9830 42152
rect 10318 42100 10324 42152
rect 10376 42100 10382 42152
rect 12161 42143 12219 42149
rect 12161 42109 12173 42143
rect 12207 42109 12219 42143
rect 12161 42103 12219 42109
rect 10226 42032 10232 42084
rect 10284 42072 10290 42084
rect 12176 42072 12204 42103
rect 12342 42100 12348 42152
rect 12400 42100 12406 42152
rect 13541 42143 13599 42149
rect 13541 42109 13553 42143
rect 13587 42140 13599 42143
rect 14826 42140 14832 42152
rect 13587 42112 14832 42140
rect 13587 42109 13599 42112
rect 13541 42103 13599 42109
rect 14826 42100 14832 42112
rect 14884 42140 14890 42152
rect 15841 42143 15899 42149
rect 15841 42140 15853 42143
rect 14884 42112 15853 42140
rect 14884 42100 14890 42112
rect 15841 42109 15853 42112
rect 15887 42109 15899 42143
rect 15841 42103 15899 42109
rect 17681 42143 17739 42149
rect 17681 42109 17693 42143
rect 17727 42109 17739 42143
rect 18708 42140 18736 42248
rect 19061 42245 19073 42279
rect 19107 42276 19119 42279
rect 19334 42276 19340 42288
rect 19107 42248 19340 42276
rect 19107 42245 19119 42248
rect 19061 42239 19119 42245
rect 19334 42236 19340 42248
rect 19392 42236 19398 42288
rect 20898 42276 20904 42288
rect 20286 42248 20904 42276
rect 20898 42236 20904 42248
rect 20956 42236 20962 42288
rect 23750 42236 23756 42288
rect 23808 42236 23814 42288
rect 24210 42236 24216 42288
rect 24268 42236 24274 42288
rect 18782 42168 18788 42220
rect 18840 42168 18846 42220
rect 21453 42211 21511 42217
rect 21453 42177 21465 42211
rect 21499 42177 21511 42211
rect 21453 42171 21511 42177
rect 22373 42211 22431 42217
rect 22373 42177 22385 42211
rect 22419 42208 22431 42211
rect 22462 42208 22468 42220
rect 22419 42180 22468 42208
rect 22419 42177 22431 42180
rect 22373 42171 22431 42177
rect 19426 42140 19432 42152
rect 18708 42112 19432 42140
rect 17681 42103 17739 42109
rect 15102 42072 15108 42084
rect 10284 42044 10916 42072
rect 12176 42044 15108 42072
rect 10284 42032 10290 42044
rect 10778 41964 10784 42016
rect 10836 41964 10842 42016
rect 10888 42004 10916 42044
rect 15102 42032 15108 42044
rect 15160 42032 15166 42084
rect 16853 42075 16911 42081
rect 16853 42072 16865 42075
rect 16546 42044 16865 42072
rect 16546 42004 16574 42044
rect 16853 42041 16865 42044
rect 16899 42072 16911 42075
rect 17696 42072 17724 42103
rect 19426 42100 19432 42112
rect 19484 42100 19490 42152
rect 20088 42112 21312 42140
rect 16899 42044 17724 42072
rect 16899 42041 16911 42044
rect 16853 42035 16911 42041
rect 10888 41976 16574 42004
rect 17770 41964 17776 42016
rect 17828 42004 17834 42016
rect 20088 42004 20116 42112
rect 20533 42075 20591 42081
rect 20533 42041 20545 42075
rect 20579 42072 20591 42075
rect 21174 42072 21180 42084
rect 20579 42044 21180 42072
rect 20579 42041 20591 42044
rect 20533 42035 20591 42041
rect 21174 42032 21180 42044
rect 21232 42032 21238 42084
rect 21284 42081 21312 42112
rect 21269 42075 21327 42081
rect 21269 42041 21281 42075
rect 21315 42041 21327 42075
rect 21468 42072 21496 42171
rect 22462 42168 22468 42180
rect 22520 42208 22526 42220
rect 22646 42208 22652 42220
rect 22520 42180 22652 42208
rect 22520 42168 22526 42180
rect 22646 42168 22652 42180
rect 22704 42168 22710 42220
rect 22005 42143 22063 42149
rect 22005 42109 22017 42143
rect 22051 42140 22063 42143
rect 22051 42112 23428 42140
rect 22051 42109 22063 42112
rect 22005 42103 22063 42109
rect 21913 42075 21971 42081
rect 21913 42072 21925 42075
rect 21468 42044 21925 42072
rect 21269 42035 21327 42041
rect 21913 42041 21925 42044
rect 21959 42072 21971 42075
rect 22094 42072 22100 42084
rect 21959 42044 22100 42072
rect 21959 42041 21971 42044
rect 21913 42035 21971 42041
rect 22094 42032 22100 42044
rect 22152 42032 22158 42084
rect 17828 41976 20116 42004
rect 17828 41964 17834 41976
rect 20898 41964 20904 42016
rect 20956 42004 20962 42016
rect 22204 42004 22232 42112
rect 20956 41976 22232 42004
rect 20956 41964 20962 41976
rect 22462 41964 22468 42016
rect 22520 42004 22526 42016
rect 23290 42004 23296 42016
rect 22520 41976 23296 42004
rect 22520 41964 22526 41976
rect 23290 41964 23296 41976
rect 23348 41964 23354 42016
rect 23400 42004 23428 42112
rect 23474 42100 23480 42152
rect 23532 42100 23538 42152
rect 24210 42004 24216 42016
rect 23400 41976 24216 42004
rect 24210 41964 24216 41976
rect 24268 41964 24274 42016
rect 1104 41914 25852 41936
rect 1104 41862 2950 41914
rect 3002 41862 3014 41914
rect 3066 41862 3078 41914
rect 3130 41862 3142 41914
rect 3194 41862 3206 41914
rect 3258 41862 12950 41914
rect 13002 41862 13014 41914
rect 13066 41862 13078 41914
rect 13130 41862 13142 41914
rect 13194 41862 13206 41914
rect 13258 41862 22950 41914
rect 23002 41862 23014 41914
rect 23066 41862 23078 41914
rect 23130 41862 23142 41914
rect 23194 41862 23206 41914
rect 23258 41862 25852 41914
rect 1104 41840 25852 41862
rect 4154 41760 4160 41812
rect 4212 41760 4218 41812
rect 4798 41760 4804 41812
rect 4856 41800 4862 41812
rect 4893 41803 4951 41809
rect 4893 41800 4905 41803
rect 4856 41772 4905 41800
rect 4856 41760 4862 41772
rect 4893 41769 4905 41772
rect 4939 41769 4951 41803
rect 6454 41800 6460 41812
rect 4893 41763 4951 41769
rect 6012 41772 6460 41800
rect 6012 41673 6040 41772
rect 6454 41760 6460 41772
rect 6512 41800 6518 41812
rect 6822 41800 6828 41812
rect 6512 41772 6828 41800
rect 6512 41760 6518 41772
rect 6822 41760 6828 41772
rect 6880 41800 6886 41812
rect 8021 41803 8079 41809
rect 8021 41800 8033 41803
rect 6880 41772 8033 41800
rect 6880 41760 6886 41772
rect 8021 41769 8033 41772
rect 8067 41800 8079 41803
rect 8478 41800 8484 41812
rect 8067 41772 8484 41800
rect 8067 41769 8079 41772
rect 8021 41763 8079 41769
rect 8478 41760 8484 41772
rect 8536 41760 8542 41812
rect 8757 41803 8815 41809
rect 8757 41769 8769 41803
rect 8803 41800 8815 41803
rect 8938 41800 8944 41812
rect 8803 41772 8944 41800
rect 8803 41769 8815 41772
rect 8757 41763 8815 41769
rect 8938 41760 8944 41772
rect 8996 41760 9002 41812
rect 11514 41760 11520 41812
rect 11572 41760 11578 41812
rect 22462 41800 22468 41812
rect 17420 41772 22468 41800
rect 7745 41735 7803 41741
rect 7745 41701 7757 41735
rect 7791 41732 7803 41735
rect 8294 41732 8300 41744
rect 7791 41704 8300 41732
rect 7791 41701 7803 41704
rect 7745 41695 7803 41701
rect 8294 41692 8300 41704
rect 8352 41732 8358 41744
rect 10318 41732 10324 41744
rect 8352 41704 10324 41732
rect 8352 41692 8358 41704
rect 10318 41692 10324 41704
rect 10376 41692 10382 41744
rect 12802 41732 12808 41744
rect 10980 41704 12808 41732
rect 5997 41667 6055 41673
rect 5997 41633 6009 41667
rect 6043 41633 6055 41667
rect 5997 41627 6055 41633
rect 6273 41667 6331 41673
rect 6273 41633 6285 41667
rect 6319 41664 6331 41667
rect 7282 41664 7288 41676
rect 6319 41636 7288 41664
rect 6319 41633 6331 41636
rect 6273 41627 6331 41633
rect 7282 41624 7288 41636
rect 7340 41624 7346 41676
rect 8938 41624 8944 41676
rect 8996 41664 9002 41676
rect 9585 41667 9643 41673
rect 9585 41664 9597 41667
rect 8996 41636 9597 41664
rect 8996 41624 9002 41636
rect 9585 41633 9597 41636
rect 9631 41633 9643 41667
rect 9585 41627 9643 41633
rect 9769 41667 9827 41673
rect 9769 41633 9781 41667
rect 9815 41664 9827 41667
rect 10778 41664 10784 41676
rect 9815 41636 10784 41664
rect 9815 41633 9827 41636
rect 9769 41627 9827 41633
rect 8297 41599 8355 41605
rect 8297 41596 8309 41599
rect 7406 41568 8309 41596
rect 8297 41565 8309 41568
rect 8343 41596 8355 41599
rect 8386 41596 8392 41608
rect 8343 41568 8392 41596
rect 8343 41565 8355 41568
rect 8297 41559 8355 41565
rect 8386 41556 8392 41568
rect 8444 41596 8450 41608
rect 8662 41596 8668 41608
rect 8444 41568 8668 41596
rect 8444 41556 8450 41568
rect 8662 41556 8668 41568
rect 8720 41596 8726 41608
rect 9490 41596 9496 41608
rect 8720 41568 9496 41596
rect 8720 41556 8726 41568
rect 9490 41556 9496 41568
rect 9548 41556 9554 41608
rect 9600 41596 9628 41627
rect 10778 41624 10784 41636
rect 10836 41624 10842 41676
rect 10870 41624 10876 41676
rect 10928 41624 10934 41676
rect 10980 41596 11008 41704
rect 12802 41692 12808 41704
rect 12860 41692 12866 41744
rect 12066 41624 12072 41676
rect 12124 41624 12130 41676
rect 14829 41667 14887 41673
rect 14829 41664 14841 41667
rect 12406 41636 14841 41664
rect 11422 41596 11428 41608
rect 9600 41568 11008 41596
rect 11072 41568 11428 41596
rect 3605 41531 3663 41537
rect 3605 41497 3617 41531
rect 3651 41528 3663 41531
rect 4062 41528 4068 41540
rect 3651 41500 4068 41528
rect 3651 41497 3663 41500
rect 3605 41491 3663 41497
rect 4062 41488 4068 41500
rect 4120 41488 4126 41540
rect 4801 41531 4859 41537
rect 4801 41497 4813 41531
rect 4847 41528 4859 41531
rect 5258 41528 5264 41540
rect 4847 41500 5264 41528
rect 4847 41497 4859 41500
rect 4801 41491 4859 41497
rect 5258 41488 5264 41500
rect 5316 41488 5322 41540
rect 11072 41528 11100 41568
rect 11422 41556 11428 41568
rect 11480 41596 11486 41608
rect 12406 41596 12434 41636
rect 14829 41633 14841 41636
rect 14875 41664 14887 41667
rect 15657 41667 15715 41673
rect 15657 41664 15669 41667
rect 14875 41636 15669 41664
rect 14875 41633 14887 41636
rect 14829 41627 14887 41633
rect 15657 41633 15669 41636
rect 15703 41633 15715 41667
rect 15657 41627 15715 41633
rect 15749 41667 15807 41673
rect 15749 41633 15761 41667
rect 15795 41633 15807 41667
rect 15749 41627 15807 41633
rect 11480 41568 12434 41596
rect 11480 41556 11486 41568
rect 12526 41556 12532 41608
rect 12584 41596 12590 41608
rect 12713 41599 12771 41605
rect 12713 41596 12725 41599
rect 12584 41568 12725 41596
rect 12584 41556 12590 41568
rect 12713 41565 12725 41568
rect 12759 41565 12771 41599
rect 15764 41596 15792 41627
rect 16298 41624 16304 41676
rect 16356 41664 16362 41676
rect 16945 41667 17003 41673
rect 16945 41664 16957 41667
rect 16356 41636 16957 41664
rect 16356 41624 16362 41636
rect 16945 41633 16957 41636
rect 16991 41633 17003 41667
rect 16945 41627 17003 41633
rect 12713 41559 12771 41565
rect 14660 41568 15792 41596
rect 8496 41500 11100 41528
rect 3970 41420 3976 41472
rect 4028 41460 4034 41472
rect 8496 41469 8524 41500
rect 8481 41463 8539 41469
rect 8481 41460 8493 41463
rect 4028 41432 8493 41460
rect 4028 41420 4034 41432
rect 8481 41429 8493 41432
rect 8527 41429 8539 41463
rect 8481 41423 8539 41429
rect 9122 41420 9128 41472
rect 9180 41420 9186 41472
rect 9508 41469 9536 41500
rect 11146 41488 11152 41540
rect 11204 41528 11210 41540
rect 11885 41531 11943 41537
rect 11885 41528 11897 41531
rect 11204 41500 11897 41528
rect 11204 41488 11210 41500
rect 11885 41497 11897 41500
rect 11931 41497 11943 41531
rect 11885 41491 11943 41497
rect 11977 41531 12035 41537
rect 11977 41497 11989 41531
rect 12023 41528 12035 41531
rect 14458 41528 14464 41540
rect 12023 41500 14464 41528
rect 12023 41497 12035 41500
rect 11977 41491 12035 41497
rect 14458 41488 14464 41500
rect 14516 41488 14522 41540
rect 9493 41463 9551 41469
rect 9493 41429 9505 41463
rect 9539 41429 9551 41463
rect 9493 41423 9551 41429
rect 10321 41463 10379 41469
rect 10321 41429 10333 41463
rect 10367 41460 10379 41463
rect 10594 41460 10600 41472
rect 10367 41432 10600 41460
rect 10367 41429 10379 41432
rect 10321 41423 10379 41429
rect 10594 41420 10600 41432
rect 10652 41420 10658 41472
rect 10686 41420 10692 41472
rect 10744 41420 10750 41472
rect 10781 41463 10839 41469
rect 10781 41429 10793 41463
rect 10827 41460 10839 41463
rect 11790 41460 11796 41472
rect 10827 41432 11796 41460
rect 10827 41429 10839 41432
rect 10781 41423 10839 41429
rect 11790 41420 11796 41432
rect 11848 41420 11854 41472
rect 13354 41420 13360 41472
rect 13412 41420 13418 41472
rect 14182 41420 14188 41472
rect 14240 41460 14246 41472
rect 14660 41469 14688 41568
rect 16666 41556 16672 41608
rect 16724 41596 16730 41608
rect 16853 41599 16911 41605
rect 16853 41596 16865 41599
rect 16724 41568 16865 41596
rect 16724 41556 16730 41568
rect 16853 41565 16865 41568
rect 16899 41565 16911 41599
rect 16853 41559 16911 41565
rect 15565 41531 15623 41537
rect 15565 41497 15577 41531
rect 15611 41528 15623 41531
rect 16114 41528 16120 41540
rect 15611 41500 16120 41528
rect 15611 41497 15623 41500
rect 15565 41491 15623 41497
rect 16114 41488 16120 41500
rect 16172 41528 16178 41540
rect 17420 41528 17448 41772
rect 22462 41760 22468 41772
rect 22520 41760 22526 41812
rect 22649 41803 22707 41809
rect 22649 41769 22661 41803
rect 22695 41800 22707 41803
rect 22695 41772 23796 41800
rect 22695 41769 22707 41772
rect 22649 41763 22707 41769
rect 17494 41692 17500 41744
rect 17552 41732 17558 41744
rect 20346 41732 20352 41744
rect 17552 41704 20352 41732
rect 17552 41692 17558 41704
rect 20346 41692 20352 41704
rect 20404 41732 20410 41744
rect 21361 41735 21419 41741
rect 20404 41704 20760 41732
rect 20404 41692 20410 41704
rect 18322 41624 18328 41676
rect 18380 41664 18386 41676
rect 18601 41667 18659 41673
rect 18601 41664 18613 41667
rect 18380 41636 18613 41664
rect 18380 41624 18386 41636
rect 18601 41633 18613 41636
rect 18647 41633 18659 41667
rect 18601 41627 18659 41633
rect 18693 41667 18751 41673
rect 18693 41633 18705 41667
rect 18739 41633 18751 41667
rect 18693 41627 18751 41633
rect 17497 41599 17555 41605
rect 17497 41565 17509 41599
rect 17543 41596 17555 41599
rect 17586 41596 17592 41608
rect 17543 41568 17592 41596
rect 17543 41565 17555 41568
rect 17497 41559 17555 41565
rect 16172 41500 17448 41528
rect 16172 41488 16178 41500
rect 14645 41463 14703 41469
rect 14645 41460 14657 41463
rect 14240 41432 14657 41460
rect 14240 41420 14246 41432
rect 14645 41429 14657 41432
rect 14691 41429 14703 41463
rect 14645 41423 14703 41429
rect 15197 41463 15255 41469
rect 15197 41429 15209 41463
rect 15243 41460 15255 41463
rect 15286 41460 15292 41472
rect 15243 41432 15292 41460
rect 15243 41429 15255 41432
rect 15197 41423 15255 41429
rect 15286 41420 15292 41432
rect 15344 41420 15350 41472
rect 16390 41420 16396 41472
rect 16448 41420 16454 41472
rect 16761 41463 16819 41469
rect 16761 41429 16773 41463
rect 16807 41460 16819 41463
rect 17512 41460 17540 41559
rect 17586 41556 17592 41568
rect 17644 41556 17650 41608
rect 18506 41556 18512 41608
rect 18564 41596 18570 41608
rect 18708 41596 18736 41627
rect 20162 41624 20168 41676
rect 20220 41664 20226 41676
rect 20622 41664 20628 41676
rect 20220 41636 20628 41664
rect 20220 41624 20226 41636
rect 20622 41624 20628 41636
rect 20680 41624 20686 41676
rect 18564 41568 18736 41596
rect 20073 41599 20131 41605
rect 18564 41556 18570 41568
rect 20073 41565 20085 41599
rect 20119 41596 20131 41599
rect 20254 41596 20260 41608
rect 20119 41568 20260 41596
rect 20119 41565 20131 41568
rect 20073 41559 20131 41565
rect 20254 41556 20260 41568
rect 20312 41556 20318 41608
rect 20732 41596 20760 41704
rect 21361 41701 21373 41735
rect 21407 41732 21419 41735
rect 22922 41732 22928 41744
rect 21407 41704 22928 41732
rect 21407 41701 21419 41704
rect 21361 41695 21419 41701
rect 22922 41692 22928 41704
rect 22980 41692 22986 41744
rect 23198 41692 23204 41744
rect 23256 41732 23262 41744
rect 23474 41732 23480 41744
rect 23256 41704 23480 41732
rect 23256 41692 23262 41704
rect 23474 41692 23480 41704
rect 23532 41692 23538 41744
rect 23768 41732 23796 41772
rect 23842 41760 23848 41812
rect 23900 41800 23906 41812
rect 25225 41803 25283 41809
rect 25225 41800 25237 41803
rect 23900 41772 25237 41800
rect 23900 41760 23906 41772
rect 25225 41769 25237 41772
rect 25271 41769 25283 41803
rect 25225 41763 25283 41769
rect 25038 41732 25044 41744
rect 23768 41704 25044 41732
rect 25038 41692 25044 41704
rect 25096 41692 25102 41744
rect 22005 41667 22063 41673
rect 22005 41633 22017 41667
rect 22051 41664 22063 41667
rect 22370 41664 22376 41676
rect 22051 41636 22376 41664
rect 22051 41633 22063 41636
rect 22005 41627 22063 41633
rect 22370 41624 22376 41636
rect 22428 41624 22434 41676
rect 22738 41624 22744 41676
rect 22796 41664 22802 41676
rect 23109 41667 23167 41673
rect 23109 41664 23121 41667
rect 22796 41636 23121 41664
rect 22796 41624 22802 41636
rect 23109 41633 23121 41636
rect 23155 41633 23167 41667
rect 23109 41627 23167 41633
rect 23293 41667 23351 41673
rect 23293 41633 23305 41667
rect 23339 41664 23351 41667
rect 23658 41664 23664 41676
rect 23339 41636 23664 41664
rect 23339 41633 23351 41636
rect 23293 41627 23351 41633
rect 23658 41624 23664 41636
rect 23716 41664 23722 41676
rect 23716 41636 24624 41664
rect 23716 41624 23722 41636
rect 24596 41608 24624 41636
rect 24029 41599 24087 41605
rect 20732 41568 23888 41596
rect 18322 41488 18328 41540
rect 18380 41528 18386 41540
rect 19337 41531 19395 41537
rect 19337 41528 19349 41531
rect 18380 41500 19349 41528
rect 18380 41488 18386 41500
rect 16807 41432 17540 41460
rect 18141 41463 18199 41469
rect 16807 41429 16819 41432
rect 16761 41423 16819 41429
rect 18141 41429 18153 41463
rect 18187 41460 18199 41463
rect 18414 41460 18420 41472
rect 18187 41432 18420 41460
rect 18187 41429 18199 41432
rect 18141 41423 18199 41429
rect 18414 41420 18420 41432
rect 18472 41420 18478 41472
rect 18524 41469 18552 41500
rect 19337 41497 19349 41500
rect 19383 41528 19395 41531
rect 20622 41528 20628 41540
rect 19383 41500 20628 41528
rect 19383 41497 19395 41500
rect 19337 41491 19395 41497
rect 20622 41488 20628 41500
rect 20680 41488 20686 41540
rect 20714 41488 20720 41540
rect 20772 41528 20778 41540
rect 21821 41531 21879 41537
rect 21821 41528 21833 41531
rect 20772 41500 21833 41528
rect 20772 41488 20778 41500
rect 21821 41497 21833 41500
rect 21867 41497 21879 41531
rect 21821 41491 21879 41497
rect 18509 41463 18567 41469
rect 18509 41429 18521 41463
rect 18555 41429 18567 41463
rect 18509 41423 18567 41429
rect 18966 41420 18972 41472
rect 19024 41460 19030 41472
rect 19150 41460 19156 41472
rect 19024 41432 19156 41460
rect 19024 41420 19030 41432
rect 19150 41420 19156 41432
rect 19208 41420 19214 41472
rect 19610 41420 19616 41472
rect 19668 41420 19674 41472
rect 19978 41420 19984 41472
rect 20036 41420 20042 41472
rect 21726 41420 21732 41472
rect 21784 41420 21790 41472
rect 22738 41420 22744 41472
rect 22796 41460 22802 41472
rect 23860 41469 23888 41568
rect 24029 41565 24041 41599
rect 24075 41596 24087 41599
rect 24118 41596 24124 41608
rect 24075 41568 24124 41596
rect 24075 41565 24087 41568
rect 24029 41559 24087 41565
rect 24118 41556 24124 41568
rect 24176 41556 24182 41608
rect 24578 41556 24584 41608
rect 24636 41556 24642 41608
rect 23017 41463 23075 41469
rect 23017 41460 23029 41463
rect 22796 41432 23029 41460
rect 22796 41420 22802 41432
rect 23017 41429 23029 41432
rect 23063 41429 23075 41463
rect 23017 41423 23075 41429
rect 23845 41463 23903 41469
rect 23845 41429 23857 41463
rect 23891 41429 23903 41463
rect 23845 41423 23903 41429
rect 1104 41370 25852 41392
rect 1104 41318 7950 41370
rect 8002 41318 8014 41370
rect 8066 41318 8078 41370
rect 8130 41318 8142 41370
rect 8194 41318 8206 41370
rect 8258 41318 17950 41370
rect 18002 41318 18014 41370
rect 18066 41318 18078 41370
rect 18130 41318 18142 41370
rect 18194 41318 18206 41370
rect 18258 41318 25852 41370
rect 1104 41296 25852 41318
rect 3602 41216 3608 41268
rect 3660 41216 3666 41268
rect 4706 41216 4712 41268
rect 4764 41216 4770 41268
rect 10781 41259 10839 41265
rect 10781 41256 10793 41259
rect 7944 41228 10793 41256
rect 1302 41080 1308 41132
rect 1360 41120 1366 41132
rect 1765 41123 1823 41129
rect 1765 41120 1777 41123
rect 1360 41092 1777 41120
rect 1360 41080 1366 41092
rect 1765 41089 1777 41092
rect 1811 41120 1823 41123
rect 2041 41123 2099 41129
rect 2041 41120 2053 41123
rect 1811 41092 2053 41120
rect 1811 41089 1823 41092
rect 1765 41083 1823 41089
rect 2041 41089 2053 41092
rect 2087 41089 2099 41123
rect 2041 41083 2099 41089
rect 3513 41123 3571 41129
rect 3513 41089 3525 41123
rect 3559 41120 3571 41123
rect 3973 41123 4031 41129
rect 3973 41120 3985 41123
rect 3559 41092 3985 41120
rect 3559 41089 3571 41092
rect 3513 41083 3571 41089
rect 3973 41089 3985 41092
rect 4019 41120 4031 41123
rect 4522 41120 4528 41132
rect 4019 41092 4528 41120
rect 4019 41089 4031 41092
rect 3973 41083 4031 41089
rect 4522 41080 4528 41092
rect 4580 41080 4586 41132
rect 4617 41123 4675 41129
rect 4617 41089 4629 41123
rect 4663 41120 4675 41123
rect 5074 41120 5080 41132
rect 4663 41092 5080 41120
rect 4663 41089 4675 41092
rect 4617 41083 4675 41089
rect 5074 41080 5080 41092
rect 5132 41080 5138 41132
rect 7944 41129 7972 41228
rect 10781 41225 10793 41228
rect 10827 41256 10839 41259
rect 10870 41256 10876 41268
rect 10827 41228 10876 41256
rect 10827 41225 10839 41228
rect 10781 41219 10839 41225
rect 10870 41216 10876 41228
rect 10928 41216 10934 41268
rect 11054 41216 11060 41268
rect 11112 41216 11118 41268
rect 13173 41259 13231 41265
rect 13173 41256 13185 41259
rect 11716 41228 13185 41256
rect 11716 41197 11744 41228
rect 13173 41225 13185 41228
rect 13219 41256 13231 41259
rect 17126 41256 17132 41268
rect 13219 41228 17132 41256
rect 13219 41225 13231 41228
rect 13173 41219 13231 41225
rect 17126 41216 17132 41228
rect 17184 41216 17190 41268
rect 19794 41216 19800 41268
rect 19852 41216 19858 41268
rect 20898 41216 20904 41268
rect 20956 41256 20962 41268
rect 20956 41228 21496 41256
rect 20956 41216 20962 41228
rect 11701 41191 11759 41197
rect 11701 41188 11713 41191
rect 11072 41160 11713 41188
rect 11072 41132 11100 41160
rect 11701 41157 11713 41160
rect 11747 41157 11759 41191
rect 11701 41151 11759 41157
rect 16114 41148 16120 41200
rect 16172 41148 16178 41200
rect 18966 41188 18972 41200
rect 18446 41160 18972 41188
rect 18966 41148 18972 41160
rect 19024 41188 19030 41200
rect 19242 41188 19248 41200
rect 19024 41160 19248 41188
rect 19024 41148 19030 41160
rect 19242 41148 19248 41160
rect 19300 41148 19306 41200
rect 19705 41191 19763 41197
rect 19705 41157 19717 41191
rect 19751 41188 19763 41191
rect 20441 41191 20499 41197
rect 20441 41188 20453 41191
rect 19751 41160 20453 41188
rect 19751 41157 19763 41160
rect 19705 41151 19763 41157
rect 20441 41157 20453 41160
rect 20487 41188 20499 41191
rect 21468 41188 21496 41228
rect 21818 41216 21824 41268
rect 21876 41256 21882 41268
rect 22005 41259 22063 41265
rect 22005 41256 22017 41259
rect 21876 41228 22017 41256
rect 21876 41216 21882 41228
rect 22005 41225 22017 41228
rect 22051 41225 22063 41259
rect 22005 41219 22063 41225
rect 22756 41228 24440 41256
rect 22756 41188 22784 41228
rect 23198 41188 23204 41200
rect 20487 41160 21220 41188
rect 21468 41160 22784 41188
rect 22848 41160 23204 41188
rect 20487 41157 20499 41160
rect 20441 41151 20499 41157
rect 7929 41123 7987 41129
rect 7929 41089 7941 41123
rect 7975 41089 7987 41123
rect 10870 41120 10876 41132
rect 10442 41092 10876 41120
rect 7929 41083 7987 41089
rect 10870 41080 10876 41092
rect 10928 41080 10934 41132
rect 11054 41080 11060 41132
rect 11112 41080 11118 41132
rect 11974 41080 11980 41132
rect 12032 41120 12038 41132
rect 12250 41120 12256 41132
rect 12032 41092 12256 41120
rect 12032 41080 12038 41092
rect 12250 41080 12256 41092
rect 12308 41120 12314 41132
rect 12529 41123 12587 41129
rect 12529 41120 12541 41123
rect 12308 41092 12541 41120
rect 12308 41080 12314 41092
rect 12529 41089 12541 41092
rect 12575 41120 12587 41123
rect 13817 41123 13875 41129
rect 13817 41120 13829 41123
rect 12575 41092 13829 41120
rect 12575 41089 12587 41092
rect 12529 41083 12587 41089
rect 13817 41089 13829 41092
rect 13863 41089 13875 41123
rect 13817 41083 13875 41089
rect 15194 41080 15200 41132
rect 15252 41120 15258 41132
rect 15933 41123 15991 41129
rect 15933 41120 15945 41123
rect 15252 41092 15945 41120
rect 15252 41080 15258 41092
rect 15933 41089 15945 41092
rect 15979 41120 15991 41123
rect 16482 41120 16488 41132
rect 15979 41092 16488 41120
rect 15979 41089 15991 41092
rect 15933 41083 15991 41089
rect 16482 41080 16488 41092
rect 16540 41080 16546 41132
rect 16850 41080 16856 41132
rect 16908 41120 16914 41132
rect 16945 41123 17003 41129
rect 16945 41120 16957 41123
rect 16908 41092 16957 41120
rect 16908 41080 16914 41092
rect 16945 41089 16957 41092
rect 16991 41089 17003 41123
rect 16945 41083 17003 41089
rect 20898 41080 20904 41132
rect 20956 41120 20962 41132
rect 21085 41123 21143 41129
rect 21085 41120 21097 41123
rect 20956 41092 21097 41120
rect 20956 41080 20962 41092
rect 21085 41089 21097 41092
rect 21131 41089 21143 41123
rect 21192 41120 21220 41160
rect 22094 41120 22100 41132
rect 21192 41092 22100 41120
rect 21085 41083 21143 41089
rect 22094 41080 22100 41092
rect 22152 41080 22158 41132
rect 22848 41129 22876 41160
rect 23198 41148 23204 41160
rect 23256 41148 23262 41200
rect 24412 41188 24440 41228
rect 24578 41216 24584 41268
rect 24636 41216 24642 41268
rect 25222 41188 25228 41200
rect 24412 41160 25228 41188
rect 25222 41148 25228 41160
rect 25280 41148 25286 41200
rect 22833 41123 22891 41129
rect 22833 41089 22845 41123
rect 22879 41089 22891 41123
rect 22833 41083 22891 41089
rect 24210 41080 24216 41132
rect 24268 41120 24274 41132
rect 24394 41120 24400 41132
rect 24268 41092 24400 41120
rect 24268 41080 24274 41092
rect 24394 41080 24400 41092
rect 24452 41080 24458 41132
rect 25314 41080 25320 41132
rect 25372 41080 25378 41132
rect 8478 41012 8484 41064
rect 8536 41052 8542 41064
rect 9033 41055 9091 41061
rect 9033 41052 9045 41055
rect 8536 41024 9045 41052
rect 8536 41012 8542 41024
rect 9033 41021 9045 41024
rect 9079 41021 9091 41055
rect 9033 41015 9091 41021
rect 9309 41055 9367 41061
rect 9309 41021 9321 41055
rect 9355 41052 9367 41055
rect 13354 41052 13360 41064
rect 9355 41024 13360 41052
rect 9355 41021 9367 41024
rect 9309 41015 9367 41021
rect 13354 41012 13360 41024
rect 13412 41012 13418 41064
rect 14093 41055 14151 41061
rect 14093 41021 14105 41055
rect 14139 41052 14151 41055
rect 16022 41052 16028 41064
rect 14139 41024 16028 41052
rect 14139 41021 14151 41024
rect 14093 41015 14151 41021
rect 16022 41012 16028 41024
rect 16080 41012 16086 41064
rect 17221 41055 17279 41061
rect 17221 41021 17233 41055
rect 17267 41052 17279 41055
rect 18598 41052 18604 41064
rect 17267 41024 18604 41052
rect 17267 41021 17279 41024
rect 17221 41015 17279 41021
rect 18598 41012 18604 41024
rect 18656 41012 18662 41064
rect 19886 41012 19892 41064
rect 19944 41012 19950 41064
rect 20990 41012 20996 41064
rect 21048 41052 21054 41064
rect 21177 41055 21235 41061
rect 21177 41052 21189 41055
rect 21048 41024 21189 41052
rect 21048 41012 21054 41024
rect 21177 41021 21189 41024
rect 21223 41021 21235 41055
rect 21177 41015 21235 41021
rect 21361 41055 21419 41061
rect 21361 41021 21373 41055
rect 21407 41052 21419 41055
rect 23109 41055 23167 41061
rect 21407 41024 21588 41052
rect 21407 41021 21419 41024
rect 21361 41015 21419 41021
rect 15565 40987 15623 40993
rect 15565 40953 15577 40987
rect 15611 40984 15623 40987
rect 16482 40984 16488 40996
rect 15611 40956 16488 40984
rect 15611 40953 15623 40956
rect 15565 40947 15623 40953
rect 16482 40944 16488 40956
rect 16540 40944 16546 40996
rect 21192 40984 21220 41015
rect 21450 40984 21456 40996
rect 18248 40956 20852 40984
rect 21192 40956 21456 40984
rect 1581 40919 1639 40925
rect 1581 40885 1593 40919
rect 1627 40916 1639 40919
rect 3602 40916 3608 40928
rect 1627 40888 3608 40916
rect 1627 40885 1639 40888
rect 1581 40879 1639 40885
rect 3602 40876 3608 40888
rect 3660 40876 3666 40928
rect 5074 40876 5080 40928
rect 5132 40876 5138 40928
rect 8570 40876 8576 40928
rect 8628 40876 8634 40928
rect 10870 40876 10876 40928
rect 10928 40916 10934 40928
rect 11333 40919 11391 40925
rect 11333 40916 11345 40919
rect 10928 40888 11345 40916
rect 10928 40876 10934 40888
rect 11333 40885 11345 40888
rect 11379 40916 11391 40919
rect 12342 40916 12348 40928
rect 11379 40888 12348 40916
rect 11379 40885 11391 40888
rect 11333 40879 11391 40885
rect 12342 40876 12348 40888
rect 12400 40876 12406 40928
rect 12989 40919 13047 40925
rect 12989 40885 13001 40919
rect 13035 40916 13047 40919
rect 13814 40916 13820 40928
rect 13035 40888 13820 40916
rect 13035 40885 13047 40888
rect 12989 40879 13047 40885
rect 13814 40876 13820 40888
rect 13872 40876 13878 40928
rect 16574 40876 16580 40928
rect 16632 40916 16638 40928
rect 17862 40916 17868 40928
rect 16632 40888 17868 40916
rect 16632 40876 16638 40888
rect 17862 40876 17868 40888
rect 17920 40916 17926 40928
rect 18248 40916 18276 40956
rect 17920 40888 18276 40916
rect 18693 40919 18751 40925
rect 17920 40876 17926 40888
rect 18693 40885 18705 40919
rect 18739 40916 18751 40919
rect 18782 40916 18788 40928
rect 18739 40888 18788 40916
rect 18739 40885 18751 40888
rect 18693 40879 18751 40885
rect 18782 40876 18788 40888
rect 18840 40876 18846 40928
rect 18966 40876 18972 40928
rect 19024 40876 19030 40928
rect 19334 40876 19340 40928
rect 19392 40876 19398 40928
rect 20438 40876 20444 40928
rect 20496 40916 20502 40928
rect 20717 40919 20775 40925
rect 20717 40916 20729 40919
rect 20496 40888 20729 40916
rect 20496 40876 20502 40888
rect 20717 40885 20729 40888
rect 20763 40885 20775 40919
rect 20824 40916 20852 40956
rect 21450 40944 21456 40956
rect 21508 40944 21514 40996
rect 21560 40916 21588 41024
rect 23109 41021 23121 41055
rect 23155 41052 23167 41055
rect 24946 41052 24952 41064
rect 23155 41024 24952 41052
rect 23155 41021 23167 41024
rect 23109 41015 23167 41021
rect 24946 41012 24952 41024
rect 25004 41012 25010 41064
rect 20824 40888 21588 40916
rect 20717 40879 20775 40885
rect 21726 40876 21732 40928
rect 21784 40916 21790 40928
rect 21910 40916 21916 40928
rect 21784 40888 21916 40916
rect 21784 40876 21790 40888
rect 21910 40876 21916 40888
rect 21968 40876 21974 40928
rect 22557 40919 22615 40925
rect 22557 40885 22569 40919
rect 22603 40916 22615 40919
rect 24118 40916 24124 40928
rect 22603 40888 24124 40916
rect 22603 40885 22615 40888
rect 22557 40879 22615 40885
rect 24118 40876 24124 40888
rect 24176 40876 24182 40928
rect 25133 40919 25191 40925
rect 25133 40885 25145 40919
rect 25179 40916 25191 40919
rect 25498 40916 25504 40928
rect 25179 40888 25504 40916
rect 25179 40885 25191 40888
rect 25133 40879 25191 40885
rect 25498 40876 25504 40888
rect 25556 40876 25562 40928
rect 1104 40826 25852 40848
rect 1104 40774 2950 40826
rect 3002 40774 3014 40826
rect 3066 40774 3078 40826
rect 3130 40774 3142 40826
rect 3194 40774 3206 40826
rect 3258 40774 12950 40826
rect 13002 40774 13014 40826
rect 13066 40774 13078 40826
rect 13130 40774 13142 40826
rect 13194 40774 13206 40826
rect 13258 40774 22950 40826
rect 23002 40774 23014 40826
rect 23066 40774 23078 40826
rect 23130 40774 23142 40826
rect 23194 40774 23206 40826
rect 23258 40774 25852 40826
rect 1104 40752 25852 40774
rect 7282 40672 7288 40724
rect 7340 40712 7346 40724
rect 7340 40684 7880 40712
rect 7340 40672 7346 40684
rect 7852 40656 7880 40684
rect 8662 40672 8668 40724
rect 8720 40672 8726 40724
rect 10226 40672 10232 40724
rect 10284 40712 10290 40724
rect 10413 40715 10471 40721
rect 10413 40712 10425 40715
rect 10284 40684 10425 40712
rect 10284 40672 10290 40684
rect 10413 40681 10425 40684
rect 10459 40712 10471 40715
rect 11054 40712 11060 40724
rect 10459 40684 11060 40712
rect 10459 40681 10471 40684
rect 10413 40675 10471 40681
rect 11054 40672 11060 40684
rect 11112 40672 11118 40724
rect 11790 40672 11796 40724
rect 11848 40712 11854 40724
rect 14277 40715 14335 40721
rect 14277 40712 14289 40715
rect 11848 40684 14289 40712
rect 11848 40672 11854 40684
rect 14277 40681 14289 40684
rect 14323 40681 14335 40715
rect 14277 40675 14335 40681
rect 15838 40672 15844 40724
rect 15896 40712 15902 40724
rect 16117 40715 16175 40721
rect 16117 40712 16129 40715
rect 15896 40684 16129 40712
rect 15896 40672 15902 40684
rect 16117 40681 16129 40684
rect 16163 40681 16175 40715
rect 16117 40675 16175 40681
rect 18598 40672 18604 40724
rect 18656 40672 18662 40724
rect 20901 40715 20959 40721
rect 20901 40681 20913 40715
rect 20947 40712 20959 40715
rect 22186 40712 22192 40724
rect 20947 40684 22192 40712
rect 20947 40681 20959 40684
rect 20901 40675 20959 40681
rect 22186 40672 22192 40684
rect 22244 40672 22250 40724
rect 23845 40715 23903 40721
rect 23845 40712 23857 40715
rect 22296 40684 23857 40712
rect 7834 40604 7840 40656
rect 7892 40644 7898 40656
rect 8205 40647 8263 40653
rect 8205 40644 8217 40647
rect 7892 40616 8217 40644
rect 7892 40604 7898 40616
rect 8205 40613 8217 40616
rect 8251 40613 8263 40647
rect 8205 40607 8263 40613
rect 10870 40604 10876 40656
rect 10928 40604 10934 40656
rect 11425 40647 11483 40653
rect 11425 40613 11437 40647
rect 11471 40644 11483 40647
rect 12618 40644 12624 40656
rect 11471 40616 12624 40644
rect 11471 40613 11483 40616
rect 11425 40607 11483 40613
rect 12618 40604 12624 40616
rect 12676 40604 12682 40656
rect 13725 40647 13783 40653
rect 13725 40644 13737 40647
rect 13096 40616 13737 40644
rect 6733 40579 6791 40585
rect 6733 40545 6745 40579
rect 6779 40576 6791 40579
rect 7374 40576 7380 40588
rect 6779 40548 7380 40576
rect 6779 40545 6791 40548
rect 6733 40539 6791 40545
rect 7374 40536 7380 40548
rect 7432 40536 7438 40588
rect 8754 40536 8760 40588
rect 8812 40576 8818 40588
rect 11977 40579 12035 40585
rect 11977 40576 11989 40579
rect 8812 40548 11989 40576
rect 8812 40536 8818 40548
rect 11977 40545 11989 40548
rect 12023 40545 12035 40579
rect 12894 40576 12900 40588
rect 11977 40539 12035 40545
rect 12406 40548 12900 40576
rect 6454 40468 6460 40520
rect 6512 40468 6518 40520
rect 8478 40468 8484 40520
rect 8536 40508 8542 40520
rect 9861 40511 9919 40517
rect 9861 40508 9873 40511
rect 8536 40480 9873 40508
rect 8536 40468 8542 40480
rect 9861 40477 9873 40480
rect 9907 40477 9919 40511
rect 9861 40471 9919 40477
rect 11793 40511 11851 40517
rect 11793 40477 11805 40511
rect 11839 40508 11851 40511
rect 12406 40508 12434 40548
rect 12894 40536 12900 40548
rect 12952 40536 12958 40588
rect 13096 40585 13124 40616
rect 13725 40613 13737 40616
rect 13771 40644 13783 40647
rect 16574 40644 16580 40656
rect 13771 40616 16580 40644
rect 13771 40613 13783 40616
rect 13725 40607 13783 40613
rect 16574 40604 16580 40616
rect 16632 40604 16638 40656
rect 16761 40647 16819 40653
rect 16761 40613 16773 40647
rect 16807 40644 16819 40647
rect 17586 40644 17592 40656
rect 16807 40616 17592 40644
rect 16807 40613 16819 40616
rect 16761 40607 16819 40613
rect 17586 40604 17592 40616
rect 17644 40604 17650 40656
rect 22002 40644 22008 40656
rect 21468 40616 22008 40644
rect 21468 40588 21496 40616
rect 22002 40604 22008 40616
rect 22060 40604 22066 40656
rect 22094 40604 22100 40656
rect 22152 40644 22158 40656
rect 22296 40644 22324 40684
rect 23845 40681 23857 40684
rect 23891 40681 23903 40715
rect 23845 40675 23903 40681
rect 22152 40616 22324 40644
rect 22152 40604 22158 40616
rect 23566 40604 23572 40656
rect 23624 40644 23630 40656
rect 23934 40644 23940 40656
rect 23624 40616 23940 40644
rect 23624 40604 23630 40616
rect 23934 40604 23940 40616
rect 23992 40604 23998 40656
rect 24026 40604 24032 40656
rect 24084 40604 24090 40656
rect 13081 40579 13139 40585
rect 13081 40545 13093 40579
rect 13127 40545 13139 40579
rect 13081 40539 13139 40545
rect 13265 40579 13323 40585
rect 13265 40545 13277 40579
rect 13311 40545 13323 40579
rect 13265 40539 13323 40545
rect 11839 40480 12434 40508
rect 11839 40477 11851 40480
rect 11793 40471 11851 40477
rect 12710 40468 12716 40520
rect 12768 40508 12774 40520
rect 12989 40511 13047 40517
rect 12989 40508 13001 40511
rect 12768 40480 13001 40508
rect 12768 40468 12774 40480
rect 12989 40477 13001 40480
rect 13035 40477 13047 40511
rect 13280 40508 13308 40539
rect 13354 40536 13360 40588
rect 13412 40576 13418 40588
rect 14829 40579 14887 40585
rect 14829 40576 14841 40579
rect 13412 40548 14841 40576
rect 13412 40536 13418 40548
rect 14829 40545 14841 40548
rect 14875 40545 14887 40579
rect 14829 40539 14887 40545
rect 17218 40536 17224 40588
rect 17276 40536 17282 40588
rect 17310 40536 17316 40588
rect 17368 40536 17374 40588
rect 21450 40536 21456 40588
rect 21508 40536 21514 40588
rect 21542 40536 21548 40588
rect 21600 40576 21606 40588
rect 22925 40579 22983 40585
rect 22925 40576 22937 40579
rect 21600 40548 22937 40576
rect 21600 40536 21606 40548
rect 22925 40545 22937 40548
rect 22971 40545 22983 40579
rect 22925 40539 22983 40545
rect 23109 40579 23167 40585
rect 23109 40545 23121 40579
rect 23155 40576 23167 40579
rect 23382 40576 23388 40588
rect 23155 40548 23388 40576
rect 23155 40545 23167 40548
rect 23109 40539 23167 40545
rect 23382 40536 23388 40548
rect 23440 40536 23446 40588
rect 24044 40576 24072 40604
rect 23481 40548 24072 40576
rect 13722 40508 13728 40520
rect 13280 40480 13728 40508
rect 12989 40471 13047 40477
rect 13722 40468 13728 40480
rect 13780 40468 13786 40520
rect 14737 40511 14795 40517
rect 14737 40477 14749 40511
rect 14783 40508 14795 40511
rect 15286 40508 15292 40520
rect 14783 40480 15292 40508
rect 14783 40477 14795 40480
rect 14737 40471 14795 40477
rect 15286 40468 15292 40480
rect 15344 40468 15350 40520
rect 15473 40511 15531 40517
rect 15473 40477 15485 40511
rect 15519 40508 15531 40511
rect 15746 40508 15752 40520
rect 15519 40480 15752 40508
rect 15519 40477 15531 40480
rect 15473 40471 15531 40477
rect 15746 40468 15752 40480
rect 15804 40468 15810 40520
rect 17862 40468 17868 40520
rect 17920 40508 17926 40520
rect 17957 40511 18015 40517
rect 17957 40508 17969 40511
rect 17920 40480 17969 40508
rect 17920 40468 17926 40480
rect 17957 40477 17969 40480
rect 18003 40477 18015 40511
rect 17957 40471 18015 40477
rect 20622 40468 20628 40520
rect 20680 40508 20686 40520
rect 21361 40511 21419 40517
rect 21361 40508 21373 40511
rect 20680 40480 21373 40508
rect 20680 40468 20686 40480
rect 21361 40477 21373 40480
rect 21407 40477 21419 40511
rect 21361 40471 21419 40477
rect 8662 40440 8668 40452
rect 7958 40412 8668 40440
rect 8662 40400 8668 40412
rect 8720 40400 8726 40452
rect 9125 40443 9183 40449
rect 9125 40409 9137 40443
rect 9171 40440 9183 40443
rect 10226 40440 10232 40452
rect 9171 40412 10232 40440
rect 9171 40409 9183 40412
rect 9125 40403 9183 40409
rect 10226 40400 10232 40412
rect 10284 40400 10290 40452
rect 13538 40440 13544 40452
rect 12636 40412 13544 40440
rect 8478 40332 8484 40384
rect 8536 40332 8542 40384
rect 8680 40372 8708 40400
rect 9398 40372 9404 40384
rect 8680 40344 9404 40372
rect 9398 40332 9404 40344
rect 9456 40332 9462 40384
rect 9674 40332 9680 40384
rect 9732 40372 9738 40384
rect 10597 40375 10655 40381
rect 10597 40372 10609 40375
rect 9732 40344 10609 40372
rect 9732 40332 9738 40344
rect 10597 40341 10609 40344
rect 10643 40372 10655 40375
rect 11057 40375 11115 40381
rect 11057 40372 11069 40375
rect 10643 40344 11069 40372
rect 10643 40341 10655 40344
rect 10597 40335 10655 40341
rect 11057 40341 11069 40344
rect 11103 40372 11115 40375
rect 11885 40375 11943 40381
rect 11885 40372 11897 40375
rect 11103 40344 11897 40372
rect 11103 40341 11115 40344
rect 11057 40335 11115 40341
rect 11885 40341 11897 40344
rect 11931 40372 11943 40375
rect 12066 40372 12072 40384
rect 11931 40344 12072 40372
rect 11931 40341 11943 40344
rect 11885 40335 11943 40341
rect 12066 40332 12072 40344
rect 12124 40332 12130 40384
rect 12636 40381 12664 40412
rect 13538 40400 13544 40412
rect 13596 40400 13602 40452
rect 13814 40400 13820 40452
rect 13872 40440 13878 40452
rect 19702 40440 19708 40452
rect 13872 40412 19708 40440
rect 13872 40400 13878 40412
rect 19702 40400 19708 40412
rect 19760 40440 19766 40452
rect 20530 40440 20536 40452
rect 19760 40412 20536 40440
rect 19760 40400 19766 40412
rect 20530 40400 20536 40412
rect 20588 40400 20594 40452
rect 21376 40440 21404 40471
rect 22002 40468 22008 40520
rect 22060 40508 22066 40520
rect 22646 40508 22652 40520
rect 22060 40480 22652 40508
rect 22060 40468 22066 40480
rect 22646 40468 22652 40480
rect 22704 40468 22710 40520
rect 22830 40468 22836 40520
rect 22888 40468 22894 40520
rect 23481 40508 23509 40548
rect 22940 40480 23509 40508
rect 23569 40511 23627 40517
rect 22940 40452 22968 40480
rect 23569 40477 23581 40511
rect 23615 40508 23627 40511
rect 24026 40508 24032 40520
rect 23615 40480 24032 40508
rect 23615 40477 23627 40480
rect 23569 40471 23627 40477
rect 24026 40468 24032 40480
rect 24084 40468 24090 40520
rect 24210 40468 24216 40520
rect 24268 40508 24274 40520
rect 24486 40508 24492 40520
rect 24268 40480 24492 40508
rect 24268 40468 24274 40480
rect 24486 40468 24492 40480
rect 24544 40508 24550 40520
rect 24581 40511 24639 40517
rect 24581 40508 24593 40511
rect 24544 40480 24593 40508
rect 24544 40468 24550 40480
rect 24581 40477 24593 40480
rect 24627 40477 24639 40511
rect 24581 40471 24639 40477
rect 24854 40468 24860 40520
rect 24912 40468 24918 40520
rect 21913 40443 21971 40449
rect 21913 40440 21925 40443
rect 21376 40412 21925 40440
rect 21913 40409 21925 40412
rect 21959 40440 21971 40443
rect 22922 40440 22928 40452
rect 21959 40412 22928 40440
rect 21959 40409 21971 40412
rect 21913 40403 21971 40409
rect 22922 40400 22928 40412
rect 22980 40400 22986 40452
rect 23382 40400 23388 40452
rect 23440 40440 23446 40452
rect 24872 40440 24900 40468
rect 23440 40412 24900 40440
rect 23440 40400 23446 40412
rect 12621 40375 12679 40381
rect 12621 40341 12633 40375
rect 12667 40341 12679 40375
rect 12621 40335 12679 40341
rect 12894 40332 12900 40384
rect 12952 40372 12958 40384
rect 13832 40372 13860 40400
rect 12952 40344 13860 40372
rect 14645 40375 14703 40381
rect 12952 40332 12958 40344
rect 14645 40341 14657 40375
rect 14691 40372 14703 40375
rect 15010 40372 15016 40384
rect 14691 40344 15016 40372
rect 14691 40341 14703 40344
rect 14645 40335 14703 40341
rect 15010 40332 15016 40344
rect 15068 40332 15074 40384
rect 16850 40332 16856 40384
rect 16908 40372 16914 40384
rect 17129 40375 17187 40381
rect 17129 40372 17141 40375
rect 16908 40344 17141 40372
rect 16908 40332 16914 40344
rect 17129 40341 17141 40344
rect 17175 40341 17187 40375
rect 17129 40335 17187 40341
rect 21269 40375 21327 40381
rect 21269 40341 21281 40375
rect 21315 40372 21327 40375
rect 21358 40372 21364 40384
rect 21315 40344 21364 40372
rect 21315 40341 21327 40344
rect 21269 40335 21327 40341
rect 21358 40332 21364 40344
rect 21416 40372 21422 40384
rect 21818 40372 21824 40384
rect 21416 40344 21824 40372
rect 21416 40332 21422 40344
rect 21818 40332 21824 40344
rect 21876 40372 21882 40384
rect 22189 40375 22247 40381
rect 22189 40372 22201 40375
rect 21876 40344 22201 40372
rect 21876 40332 21882 40344
rect 22189 40341 22201 40344
rect 22235 40372 22247 40375
rect 22370 40372 22376 40384
rect 22235 40344 22376 40372
rect 22235 40341 22247 40344
rect 22189 40335 22247 40341
rect 22370 40332 22376 40344
rect 22428 40332 22434 40384
rect 22465 40375 22523 40381
rect 22465 40341 22477 40375
rect 22511 40372 22523 40375
rect 23566 40372 23572 40384
rect 22511 40344 23572 40372
rect 22511 40341 22523 40344
rect 22465 40335 22523 40341
rect 23566 40332 23572 40344
rect 23624 40332 23630 40384
rect 24854 40332 24860 40384
rect 24912 40372 24918 40384
rect 25225 40375 25283 40381
rect 25225 40372 25237 40375
rect 24912 40344 25237 40372
rect 24912 40332 24918 40344
rect 25225 40341 25237 40344
rect 25271 40341 25283 40375
rect 25225 40335 25283 40341
rect 1104 40282 25852 40304
rect 1104 40230 7950 40282
rect 8002 40230 8014 40282
rect 8066 40230 8078 40282
rect 8130 40230 8142 40282
rect 8194 40230 8206 40282
rect 8258 40230 17950 40282
rect 18002 40230 18014 40282
rect 18066 40230 18078 40282
rect 18130 40230 18142 40282
rect 18194 40230 18206 40282
rect 18258 40230 25852 40282
rect 1104 40208 25852 40230
rect 7006 40128 7012 40180
rect 7064 40168 7070 40180
rect 7469 40171 7527 40177
rect 7469 40168 7481 40171
rect 7064 40140 7481 40168
rect 7064 40128 7070 40140
rect 7469 40137 7481 40140
rect 7515 40137 7527 40171
rect 7469 40131 7527 40137
rect 7837 40171 7895 40177
rect 7837 40137 7849 40171
rect 7883 40168 7895 40171
rect 8846 40168 8852 40180
rect 7883 40140 8852 40168
rect 7883 40137 7895 40140
rect 7837 40131 7895 40137
rect 8846 40128 8852 40140
rect 8904 40128 8910 40180
rect 9674 40128 9680 40180
rect 9732 40168 9738 40180
rect 11701 40171 11759 40177
rect 11701 40168 11713 40171
rect 9732 40140 11713 40168
rect 9732 40128 9738 40140
rect 11701 40137 11713 40140
rect 11747 40137 11759 40171
rect 11701 40131 11759 40137
rect 12066 40128 12072 40180
rect 12124 40128 12130 40180
rect 14384 40140 14596 40168
rect 6825 40103 6883 40109
rect 6825 40069 6837 40103
rect 6871 40100 6883 40103
rect 8386 40100 8392 40112
rect 6871 40072 8392 40100
rect 6871 40069 6883 40072
rect 6825 40063 6883 40069
rect 8386 40060 8392 40072
rect 8444 40060 8450 40112
rect 8570 40060 8576 40112
rect 8628 40100 8634 40112
rect 8941 40103 8999 40109
rect 8941 40100 8953 40103
rect 8628 40072 8953 40100
rect 8628 40060 8634 40072
rect 8941 40069 8953 40072
rect 8987 40069 8999 40103
rect 8941 40063 8999 40069
rect 9490 40060 9496 40112
rect 9548 40060 9554 40112
rect 10594 40060 10600 40112
rect 10652 40100 10658 40112
rect 10689 40103 10747 40109
rect 10689 40100 10701 40103
rect 10652 40072 10701 40100
rect 10652 40060 10658 40072
rect 10689 40069 10701 40072
rect 10735 40100 10747 40103
rect 10778 40100 10784 40112
rect 10735 40072 10784 40100
rect 10735 40069 10747 40072
rect 10689 40063 10747 40069
rect 10778 40060 10784 40072
rect 10836 40060 10842 40112
rect 14384 40044 14412 40140
rect 14568 40100 14596 40140
rect 14734 40128 14740 40180
rect 14792 40128 14798 40180
rect 15102 40128 15108 40180
rect 15160 40168 15166 40180
rect 15565 40171 15623 40177
rect 15565 40168 15577 40171
rect 15160 40140 15577 40168
rect 15160 40128 15166 40140
rect 15565 40137 15577 40140
rect 15611 40137 15623 40171
rect 15565 40131 15623 40137
rect 18230 40128 18236 40180
rect 18288 40128 18294 40180
rect 19334 40128 19340 40180
rect 19392 40168 19398 40180
rect 19889 40171 19947 40177
rect 19889 40168 19901 40171
rect 19392 40140 19901 40168
rect 19392 40128 19398 40140
rect 19889 40137 19901 40140
rect 19935 40137 19947 40171
rect 19889 40131 19947 40137
rect 19978 40128 19984 40180
rect 20036 40168 20042 40180
rect 20625 40171 20683 40177
rect 20625 40168 20637 40171
rect 20036 40140 20637 40168
rect 20036 40128 20042 40140
rect 20625 40137 20637 40140
rect 20671 40137 20683 40171
rect 20625 40131 20683 40137
rect 20993 40171 21051 40177
rect 20993 40137 21005 40171
rect 21039 40168 21051 40171
rect 22094 40168 22100 40180
rect 21039 40140 22100 40168
rect 21039 40137 21051 40140
rect 20993 40131 21051 40137
rect 22094 40128 22100 40140
rect 22152 40168 22158 40180
rect 22152 40140 22197 40168
rect 22152 40128 22158 40140
rect 22370 40128 22376 40180
rect 22428 40128 22434 40180
rect 22646 40128 22652 40180
rect 22704 40168 22710 40180
rect 25133 40171 25191 40177
rect 25133 40168 25145 40171
rect 22704 40140 25145 40168
rect 22704 40128 22710 40140
rect 25133 40137 25145 40140
rect 25179 40137 25191 40171
rect 25133 40131 25191 40137
rect 14568 40072 15148 40100
rect 7929 40035 7987 40041
rect 7929 40001 7941 40035
rect 7975 40032 7987 40035
rect 11149 40035 11207 40041
rect 7975 40004 8616 40032
rect 7975 40001 7987 40004
rect 7929 39995 7987 40001
rect 8588 39976 8616 40004
rect 11149 40001 11161 40035
rect 11195 40032 11207 40035
rect 11330 40032 11336 40044
rect 11195 40004 11336 40032
rect 11195 40001 11207 40004
rect 11149 39995 11207 40001
rect 11330 39992 11336 40004
rect 11388 40032 11394 40044
rect 12710 40032 12716 40044
rect 11388 40004 12716 40032
rect 11388 39992 11394 40004
rect 7742 39924 7748 39976
rect 7800 39964 7806 39976
rect 8021 39967 8079 39973
rect 8021 39964 8033 39967
rect 7800 39936 8033 39964
rect 7800 39924 7806 39936
rect 8021 39933 8033 39936
rect 8067 39933 8079 39967
rect 8021 39927 8079 39933
rect 8570 39924 8576 39976
rect 8628 39924 8634 39976
rect 8662 39924 8668 39976
rect 8720 39924 8726 39976
rect 12176 39973 12204 40004
rect 12710 39992 12716 40004
rect 12768 39992 12774 40044
rect 14366 39992 14372 40044
rect 14424 39992 14430 40044
rect 15120 40041 15148 40072
rect 15286 40060 15292 40112
rect 15344 40100 15350 40112
rect 15933 40103 15991 40109
rect 15933 40100 15945 40103
rect 15344 40072 15945 40100
rect 15344 40060 15350 40072
rect 15933 40069 15945 40072
rect 15979 40069 15991 40103
rect 15933 40063 15991 40069
rect 16574 40060 16580 40112
rect 16632 40100 16638 40112
rect 18601 40103 18659 40109
rect 18601 40100 18613 40103
rect 16632 40072 18613 40100
rect 16632 40060 16638 40072
rect 18601 40069 18613 40072
rect 18647 40069 18659 40103
rect 22462 40100 22468 40112
rect 18601 40063 18659 40069
rect 19444 40072 22468 40100
rect 15105 40035 15163 40041
rect 15105 40001 15117 40035
rect 15151 40032 15163 40035
rect 15194 40032 15200 40044
rect 15151 40004 15200 40032
rect 15151 40001 15163 40004
rect 15105 39995 15163 40001
rect 15194 39992 15200 40004
rect 15252 39992 15258 40044
rect 16025 40035 16083 40041
rect 16025 40001 16037 40035
rect 16071 40032 16083 40035
rect 16071 40004 16436 40032
rect 16071 40001 16083 40004
rect 16025 39995 16083 40001
rect 12161 39967 12219 39973
rect 12161 39933 12173 39967
rect 12207 39933 12219 39967
rect 12161 39927 12219 39933
rect 12253 39967 12311 39973
rect 12253 39933 12265 39967
rect 12299 39933 12311 39967
rect 12253 39927 12311 39933
rect 12989 39967 13047 39973
rect 12989 39933 13001 39967
rect 13035 39933 13047 39967
rect 12989 39927 13047 39933
rect 13265 39967 13323 39973
rect 13265 39933 13277 39967
rect 13311 39964 13323 39967
rect 13311 39936 15424 39964
rect 13311 39933 13323 39936
rect 13265 39927 13323 39933
rect 12268 39896 12296 39927
rect 11532 39868 12296 39896
rect 11532 39840 11560 39868
rect 11333 39831 11391 39837
rect 11333 39797 11345 39831
rect 11379 39828 11391 39831
rect 11514 39828 11520 39840
rect 11379 39800 11520 39828
rect 11379 39797 11391 39800
rect 11333 39791 11391 39797
rect 11514 39788 11520 39800
rect 11572 39788 11578 39840
rect 13004 39828 13032 39927
rect 15396 39896 15424 39936
rect 16114 39924 16120 39976
rect 16172 39924 16178 39976
rect 16408 39964 16436 40004
rect 16482 39992 16488 40044
rect 16540 40032 16546 40044
rect 16853 40035 16911 40041
rect 16853 40032 16865 40035
rect 16540 40004 16865 40032
rect 16540 39992 16546 40004
rect 16853 40001 16865 40004
rect 16899 40001 16911 40035
rect 16853 39995 16911 40001
rect 16666 39964 16672 39976
rect 16408 39936 16672 39964
rect 16666 39924 16672 39936
rect 16724 39964 16730 39976
rect 17770 39964 17776 39976
rect 16724 39936 17776 39964
rect 16724 39924 16730 39936
rect 17770 39924 17776 39936
rect 17828 39924 17834 39976
rect 18414 39924 18420 39976
rect 18472 39964 18478 39976
rect 18693 39967 18751 39973
rect 18693 39964 18705 39967
rect 18472 39936 18705 39964
rect 18472 39924 18478 39936
rect 18693 39933 18705 39936
rect 18739 39933 18751 39967
rect 18693 39927 18751 39933
rect 18874 39924 18880 39976
rect 18932 39924 18938 39976
rect 19444 39905 19472 40072
rect 22462 40060 22468 40072
rect 22520 40060 22526 40112
rect 24394 40060 24400 40112
rect 24452 40060 24458 40112
rect 19797 40035 19855 40041
rect 19797 40001 19809 40035
rect 19843 40001 19855 40035
rect 22281 40035 22339 40041
rect 22281 40032 22293 40035
rect 19797 39995 19855 40001
rect 21836 40004 22293 40032
rect 17497 39899 17555 39905
rect 17497 39896 17509 39899
rect 15396 39868 17509 39896
rect 17497 39865 17509 39868
rect 17543 39865 17555 39899
rect 17497 39859 17555 39865
rect 19429 39899 19487 39905
rect 19429 39865 19441 39899
rect 19475 39865 19487 39899
rect 19429 39859 19487 39865
rect 14642 39828 14648 39840
rect 13004 39800 14648 39828
rect 14642 39788 14648 39800
rect 14700 39788 14706 39840
rect 19242 39788 19248 39840
rect 19300 39828 19306 39840
rect 19812 39828 19840 39995
rect 21836 39976 21864 40004
rect 22281 40001 22293 40004
rect 22327 40032 22339 40035
rect 22922 40032 22928 40044
rect 22327 40004 22928 40032
rect 22327 40001 22339 40004
rect 22281 39995 22339 40001
rect 22922 39992 22928 40004
rect 22980 39992 22986 40044
rect 20070 39924 20076 39976
rect 20128 39924 20134 39976
rect 21085 39967 21143 39973
rect 21085 39933 21097 39967
rect 21131 39933 21143 39967
rect 21085 39927 21143 39933
rect 19300 39800 19840 39828
rect 21100 39828 21128 39927
rect 21266 39924 21272 39976
rect 21324 39924 21330 39976
rect 21818 39924 21824 39976
rect 21876 39924 21882 39976
rect 22370 39924 22376 39976
rect 22428 39964 22434 39976
rect 23385 39967 23443 39973
rect 23385 39964 23397 39967
rect 22428 39936 23397 39964
rect 22428 39924 22434 39936
rect 23385 39933 23397 39936
rect 23431 39933 23443 39967
rect 23385 39927 23443 39933
rect 23661 39967 23719 39973
rect 23661 39933 23673 39967
rect 23707 39964 23719 39967
rect 25222 39964 25228 39976
rect 23707 39936 25228 39964
rect 23707 39933 23719 39936
rect 23661 39927 23719 39933
rect 25222 39924 25228 39936
rect 25280 39924 25286 39976
rect 25314 39896 25320 39908
rect 24872 39868 25320 39896
rect 21910 39828 21916 39840
rect 21100 39800 21916 39828
rect 19300 39788 19306 39800
rect 21910 39788 21916 39800
rect 21968 39788 21974 39840
rect 22830 39788 22836 39840
rect 22888 39788 22894 39840
rect 23109 39831 23167 39837
rect 23109 39797 23121 39831
rect 23155 39828 23167 39831
rect 24872 39828 24900 39868
rect 25314 39856 25320 39868
rect 25372 39856 25378 39908
rect 23155 39800 24900 39828
rect 23155 39797 23167 39800
rect 23109 39791 23167 39797
rect 1104 39738 25852 39760
rect 1104 39686 2950 39738
rect 3002 39686 3014 39738
rect 3066 39686 3078 39738
rect 3130 39686 3142 39738
rect 3194 39686 3206 39738
rect 3258 39686 12950 39738
rect 13002 39686 13014 39738
rect 13066 39686 13078 39738
rect 13130 39686 13142 39738
rect 13194 39686 13206 39738
rect 13258 39686 22950 39738
rect 23002 39686 23014 39738
rect 23066 39686 23078 39738
rect 23130 39686 23142 39738
rect 23194 39686 23206 39738
rect 23258 39686 25852 39738
rect 1104 39664 25852 39686
rect 5902 39584 5908 39636
rect 5960 39624 5966 39636
rect 5960 39596 7328 39624
rect 5960 39584 5966 39596
rect 6454 39488 6460 39500
rect 5184 39460 6460 39488
rect 5184 39432 5212 39460
rect 6454 39448 6460 39460
rect 6512 39448 6518 39500
rect 6917 39491 6975 39497
rect 6917 39457 6929 39491
rect 6963 39457 6975 39491
rect 7300 39488 7328 39596
rect 7374 39584 7380 39636
rect 7432 39624 7438 39636
rect 8113 39627 8171 39633
rect 8113 39624 8125 39627
rect 7432 39596 8125 39624
rect 7432 39584 7438 39596
rect 8113 39593 8125 39596
rect 8159 39593 8171 39627
rect 8113 39587 8171 39593
rect 8478 39584 8484 39636
rect 8536 39584 8542 39636
rect 8570 39584 8576 39636
rect 8628 39624 8634 39636
rect 9769 39627 9827 39633
rect 9769 39624 9781 39627
rect 8628 39596 9781 39624
rect 8628 39584 8634 39596
rect 9769 39593 9781 39596
rect 9815 39593 9827 39627
rect 9769 39587 9827 39593
rect 11228 39627 11286 39633
rect 11228 39593 11240 39627
rect 11274 39624 11286 39627
rect 11882 39624 11888 39636
rect 11274 39596 11888 39624
rect 11274 39593 11286 39596
rect 11228 39587 11286 39593
rect 11882 39584 11888 39596
rect 11940 39624 11946 39636
rect 11940 39596 12434 39624
rect 11940 39584 11946 39596
rect 8662 39516 8668 39568
rect 8720 39556 8726 39568
rect 12406 39556 12434 39596
rect 12526 39584 12532 39636
rect 12584 39624 12590 39636
rect 12713 39627 12771 39633
rect 12713 39624 12725 39627
rect 12584 39596 12725 39624
rect 12584 39584 12590 39596
rect 12713 39593 12725 39596
rect 12759 39624 12771 39627
rect 13354 39624 13360 39636
rect 12759 39596 13360 39624
rect 12759 39593 12771 39596
rect 12713 39587 12771 39593
rect 13354 39584 13360 39596
rect 13412 39584 13418 39636
rect 13814 39624 13820 39636
rect 13464 39596 13820 39624
rect 13464 39556 13492 39596
rect 13814 39584 13820 39596
rect 13872 39624 13878 39636
rect 14182 39624 14188 39636
rect 13872 39596 14188 39624
rect 13872 39584 13878 39596
rect 14182 39584 14188 39596
rect 14240 39584 14246 39636
rect 14461 39627 14519 39633
rect 14461 39593 14473 39627
rect 14507 39624 14519 39627
rect 16850 39624 16856 39636
rect 14507 39596 16856 39624
rect 14507 39593 14519 39596
rect 14461 39587 14519 39593
rect 16850 39584 16856 39596
rect 16908 39584 16914 39636
rect 21361 39627 21419 39633
rect 21361 39593 21373 39627
rect 21407 39624 21419 39627
rect 22738 39624 22744 39636
rect 21407 39596 22744 39624
rect 21407 39593 21419 39596
rect 21361 39587 21419 39593
rect 22738 39584 22744 39596
rect 22796 39584 22802 39636
rect 8720 39528 11008 39556
rect 12406 39528 13492 39556
rect 8720 39516 8726 39528
rect 8570 39488 8576 39500
rect 7300 39460 8576 39488
rect 6917 39451 6975 39457
rect 5166 39380 5172 39432
rect 5224 39380 5230 39432
rect 6932 39420 6960 39451
rect 8570 39448 8576 39460
rect 8628 39448 8634 39500
rect 9122 39448 9128 39500
rect 9180 39488 9186 39500
rect 10980 39497 11008 39528
rect 13630 39516 13636 39568
rect 13688 39556 13694 39568
rect 15657 39559 15715 39565
rect 15657 39556 15669 39559
rect 13688 39528 15669 39556
rect 13688 39516 13694 39528
rect 15657 39525 15669 39528
rect 15703 39525 15715 39559
rect 15657 39519 15715 39525
rect 19150 39516 19156 39568
rect 19208 39556 19214 39568
rect 20441 39559 20499 39565
rect 20441 39556 20453 39559
rect 19208 39528 20453 39556
rect 19208 39516 19214 39528
rect 20441 39525 20453 39528
rect 20487 39556 20499 39559
rect 21082 39556 21088 39568
rect 20487 39528 21088 39556
rect 20487 39525 20499 39528
rect 20441 39519 20499 39525
rect 21082 39516 21088 39528
rect 21140 39516 21146 39568
rect 21726 39516 21732 39568
rect 21784 39556 21790 39568
rect 21784 39528 21956 39556
rect 21784 39516 21790 39528
rect 10229 39491 10287 39497
rect 10229 39488 10241 39491
rect 9180 39460 10241 39488
rect 9180 39448 9186 39460
rect 10229 39457 10241 39460
rect 10275 39457 10287 39491
rect 10229 39451 10287 39457
rect 10321 39491 10379 39497
rect 10321 39457 10333 39491
rect 10367 39457 10379 39491
rect 10321 39451 10379 39457
rect 10965 39491 11023 39497
rect 10965 39457 10977 39491
rect 11011 39488 11023 39491
rect 11974 39488 11980 39500
rect 11011 39460 11980 39488
rect 11011 39457 11023 39460
rect 10965 39451 11023 39457
rect 7469 39423 7527 39429
rect 7469 39420 7481 39423
rect 6932 39392 7481 39420
rect 7469 39389 7481 39392
rect 7515 39420 7527 39423
rect 8754 39420 8760 39432
rect 7515 39392 8760 39420
rect 7515 39389 7527 39392
rect 7469 39383 7527 39389
rect 8754 39380 8760 39392
rect 8812 39380 8818 39432
rect 9306 39380 9312 39432
rect 9364 39420 9370 39432
rect 10336 39420 10364 39451
rect 11974 39448 11980 39460
rect 12032 39448 12038 39500
rect 12710 39448 12716 39500
rect 12768 39488 12774 39500
rect 13906 39488 13912 39500
rect 12768 39460 13912 39488
rect 12768 39448 12774 39460
rect 13906 39448 13912 39460
rect 13964 39448 13970 39500
rect 15105 39491 15163 39497
rect 15105 39457 15117 39491
rect 15151 39488 15163 39491
rect 15378 39488 15384 39500
rect 15151 39460 15384 39488
rect 15151 39457 15163 39460
rect 15105 39451 15163 39457
rect 15378 39448 15384 39460
rect 15436 39448 15442 39500
rect 15562 39448 15568 39500
rect 15620 39488 15626 39500
rect 16301 39491 16359 39497
rect 15620 39460 16252 39488
rect 15620 39448 15626 39460
rect 9364 39392 10364 39420
rect 9364 39380 9370 39392
rect 12342 39380 12348 39432
rect 12400 39420 12406 39432
rect 13357 39423 13415 39429
rect 13357 39420 13369 39423
rect 12400 39392 13369 39420
rect 12400 39380 12406 39392
rect 13357 39389 13369 39392
rect 13403 39420 13415 39423
rect 13630 39420 13636 39432
rect 13403 39392 13636 39420
rect 13403 39389 13415 39392
rect 13357 39383 13415 39389
rect 13630 39380 13636 39392
rect 13688 39420 13694 39432
rect 14366 39420 14372 39432
rect 13688 39392 14372 39420
rect 13688 39380 13694 39392
rect 14366 39380 14372 39392
rect 14424 39380 14430 39432
rect 16224 39420 16252 39460
rect 16301 39457 16313 39491
rect 16347 39488 16359 39491
rect 18598 39488 18604 39500
rect 16347 39460 18604 39488
rect 16347 39457 16359 39460
rect 16301 39451 16359 39457
rect 18598 39448 18604 39460
rect 18656 39448 18662 39500
rect 18782 39488 18788 39500
rect 18708 39460 18788 39488
rect 17681 39423 17739 39429
rect 17681 39420 17693 39423
rect 16224 39392 17693 39420
rect 17681 39389 17693 39392
rect 17727 39420 17739 39423
rect 18708 39420 18736 39460
rect 18782 39448 18788 39460
rect 18840 39488 18846 39500
rect 19981 39491 20039 39497
rect 19981 39488 19993 39491
rect 18840 39460 19993 39488
rect 18840 39448 18846 39460
rect 19981 39457 19993 39460
rect 20027 39457 20039 39491
rect 19981 39451 20039 39457
rect 21818 39448 21824 39500
rect 21876 39448 21882 39500
rect 21928 39497 21956 39528
rect 21913 39491 21971 39497
rect 21913 39457 21925 39491
rect 21959 39457 21971 39491
rect 21913 39451 21971 39457
rect 23201 39491 23259 39497
rect 23201 39457 23213 39491
rect 23247 39488 23259 39491
rect 23658 39488 23664 39500
rect 23247 39460 23664 39488
rect 23247 39457 23259 39460
rect 23201 39451 23259 39457
rect 23658 39448 23664 39460
rect 23716 39448 23722 39500
rect 25038 39448 25044 39500
rect 25096 39448 25102 39500
rect 25130 39448 25136 39500
rect 25188 39448 25194 39500
rect 17727 39392 18736 39420
rect 19889 39423 19947 39429
rect 17727 39389 17739 39392
rect 17681 39383 17739 39389
rect 19889 39389 19901 39423
rect 19935 39420 19947 39423
rect 20438 39420 20444 39432
rect 19935 39392 20444 39420
rect 19935 39389 19947 39392
rect 19889 39383 19947 39389
rect 20438 39380 20444 39392
rect 20496 39380 20502 39432
rect 20622 39380 20628 39432
rect 20680 39420 20686 39432
rect 23017 39423 23075 39429
rect 23017 39420 23029 39423
rect 20680 39392 23029 39420
rect 20680 39380 20686 39392
rect 23017 39389 23029 39392
rect 23063 39389 23075 39423
rect 23017 39383 23075 39389
rect 5442 39312 5448 39364
rect 5500 39312 5506 39364
rect 8662 39352 8668 39364
rect 6670 39324 8668 39352
rect 6454 39244 6460 39296
rect 6512 39284 6518 39296
rect 6748 39284 6776 39324
rect 8662 39312 8668 39324
rect 8720 39352 8726 39364
rect 9398 39352 9404 39364
rect 8720 39324 9404 39352
rect 8720 39312 8726 39324
rect 9398 39312 9404 39324
rect 9456 39312 9462 39364
rect 10137 39355 10195 39361
rect 10137 39321 10149 39355
rect 10183 39352 10195 39355
rect 14921 39355 14979 39361
rect 14921 39352 14933 39355
rect 10183 39324 11192 39352
rect 10183 39321 10195 39324
rect 10137 39315 10195 39321
rect 6512 39256 6776 39284
rect 9125 39287 9183 39293
rect 6512 39244 6518 39256
rect 9125 39253 9137 39287
rect 9171 39284 9183 39287
rect 10042 39284 10048 39296
rect 9171 39256 10048 39284
rect 9171 39253 9183 39256
rect 9125 39247 9183 39253
rect 10042 39244 10048 39256
rect 10100 39244 10106 39296
rect 11164 39284 11192 39324
rect 14108 39324 14933 39352
rect 12986 39284 12992 39296
rect 11164 39256 12992 39284
rect 12986 39244 12992 39256
rect 13044 39244 13050 39296
rect 13078 39244 13084 39296
rect 13136 39244 13142 39296
rect 13541 39287 13599 39293
rect 13541 39253 13553 39287
rect 13587 39284 13599 39287
rect 13814 39284 13820 39296
rect 13587 39256 13820 39284
rect 13587 39253 13599 39256
rect 13541 39247 13599 39253
rect 13814 39244 13820 39256
rect 13872 39244 13878 39296
rect 13998 39244 14004 39296
rect 14056 39284 14062 39296
rect 14108 39293 14136 39324
rect 14921 39321 14933 39324
rect 14967 39321 14979 39355
rect 14921 39315 14979 39321
rect 16117 39355 16175 39361
rect 16117 39321 16129 39355
rect 16163 39352 16175 39355
rect 16163 39324 19472 39352
rect 16163 39321 16175 39324
rect 16117 39315 16175 39321
rect 14093 39287 14151 39293
rect 14093 39284 14105 39287
rect 14056 39256 14105 39284
rect 14056 39244 14062 39256
rect 14093 39253 14105 39256
rect 14139 39253 14151 39287
rect 14093 39247 14151 39253
rect 14826 39244 14832 39296
rect 14884 39244 14890 39296
rect 15194 39244 15200 39296
rect 15252 39284 15258 39296
rect 16025 39287 16083 39293
rect 16025 39284 16037 39287
rect 15252 39256 16037 39284
rect 15252 39244 15258 39256
rect 16025 39253 16037 39256
rect 16071 39253 16083 39287
rect 16025 39247 16083 39253
rect 17218 39244 17224 39296
rect 17276 39284 17282 39296
rect 19444 39293 19472 39324
rect 19978 39312 19984 39364
rect 20036 39352 20042 39364
rect 21358 39352 21364 39364
rect 20036 39324 21364 39352
rect 20036 39312 20042 39324
rect 21358 39312 21364 39324
rect 21416 39352 21422 39364
rect 21729 39355 21787 39361
rect 21729 39352 21741 39355
rect 21416 39324 21741 39352
rect 21416 39312 21422 39324
rect 21729 39321 21741 39324
rect 21775 39321 21787 39355
rect 21729 39315 21787 39321
rect 22925 39355 22983 39361
rect 22925 39321 22937 39355
rect 22971 39352 22983 39355
rect 23753 39355 23811 39361
rect 23753 39352 23765 39355
rect 22971 39324 23765 39352
rect 22971 39321 22983 39324
rect 22925 39315 22983 39321
rect 23753 39321 23765 39324
rect 23799 39321 23811 39355
rect 24949 39355 25007 39361
rect 24949 39352 24961 39355
rect 23753 39315 23811 39321
rect 23860 39324 24961 39352
rect 18325 39287 18383 39293
rect 18325 39284 18337 39287
rect 17276 39256 18337 39284
rect 17276 39244 17282 39256
rect 18325 39253 18337 39256
rect 18371 39253 18383 39287
rect 18325 39247 18383 39253
rect 19429 39287 19487 39293
rect 19429 39253 19441 39287
rect 19475 39253 19487 39287
rect 19429 39247 19487 39253
rect 19797 39287 19855 39293
rect 19797 39253 19809 39287
rect 19843 39284 19855 39287
rect 20070 39284 20076 39296
rect 19843 39256 20076 39284
rect 19843 39253 19855 39256
rect 19797 39247 19855 39253
rect 20070 39244 20076 39256
rect 20128 39244 20134 39296
rect 22557 39287 22615 39293
rect 22557 39253 22569 39287
rect 22603 39284 22615 39287
rect 23860 39284 23888 39324
rect 24949 39321 24961 39324
rect 24995 39321 25007 39355
rect 24949 39315 25007 39321
rect 22603 39256 23888 39284
rect 24581 39287 24639 39293
rect 22603 39253 22615 39256
rect 22557 39247 22615 39253
rect 24581 39253 24593 39287
rect 24627 39284 24639 39287
rect 24762 39284 24768 39296
rect 24627 39256 24768 39284
rect 24627 39253 24639 39256
rect 24581 39247 24639 39253
rect 24762 39244 24768 39256
rect 24820 39244 24826 39296
rect 1104 39194 25852 39216
rect 1104 39142 7950 39194
rect 8002 39142 8014 39194
rect 8066 39142 8078 39194
rect 8130 39142 8142 39194
rect 8194 39142 8206 39194
rect 8258 39142 17950 39194
rect 18002 39142 18014 39194
rect 18066 39142 18078 39194
rect 18130 39142 18142 39194
rect 18194 39142 18206 39194
rect 18258 39142 25852 39194
rect 1104 39120 25852 39142
rect 5442 39040 5448 39092
rect 5500 39080 5506 39092
rect 5997 39083 6055 39089
rect 5997 39080 6009 39083
rect 5500 39052 6009 39080
rect 5500 39040 5506 39052
rect 5997 39049 6009 39052
rect 6043 39049 6055 39083
rect 5997 39043 6055 39049
rect 6546 39040 6552 39092
rect 6604 39040 6610 39092
rect 8386 39040 8392 39092
rect 8444 39080 8450 39092
rect 9493 39083 9551 39089
rect 9493 39080 9505 39083
rect 8444 39052 9505 39080
rect 8444 39040 8450 39052
rect 9493 39049 9505 39052
rect 9539 39049 9551 39083
rect 9493 39043 9551 39049
rect 10413 39083 10471 39089
rect 10413 39049 10425 39083
rect 10459 39080 10471 39083
rect 10686 39080 10692 39092
rect 10459 39052 10692 39080
rect 10459 39049 10471 39052
rect 10413 39043 10471 39049
rect 10686 39040 10692 39052
rect 10744 39040 10750 39092
rect 12158 39040 12164 39092
rect 12216 39080 12222 39092
rect 12253 39083 12311 39089
rect 12253 39080 12265 39083
rect 12216 39052 12265 39080
rect 12216 39040 12222 39052
rect 12253 39049 12265 39052
rect 12299 39049 12311 39083
rect 12253 39043 12311 39049
rect 12618 39040 12624 39092
rect 12676 39080 12682 39092
rect 12713 39083 12771 39089
rect 12713 39080 12725 39083
rect 12676 39052 12725 39080
rect 12676 39040 12682 39052
rect 12713 39049 12725 39052
rect 12759 39049 12771 39083
rect 16114 39080 16120 39092
rect 12713 39043 12771 39049
rect 12820 39052 16120 39080
rect 5810 39012 5816 39024
rect 5368 38984 5816 39012
rect 5368 38953 5396 38984
rect 5810 38972 5816 38984
rect 5868 39012 5874 39024
rect 5868 38984 7144 39012
rect 5868 38972 5874 38984
rect 5353 38947 5411 38953
rect 5353 38913 5365 38947
rect 5399 38913 5411 38947
rect 5353 38907 5411 38913
rect 5442 38904 5448 38956
rect 5500 38944 5506 38956
rect 6917 38947 6975 38953
rect 6917 38944 6929 38947
rect 5500 38916 6929 38944
rect 5500 38904 5506 38916
rect 6917 38913 6929 38916
rect 6963 38913 6975 38947
rect 6917 38907 6975 38913
rect 7116 38885 7144 38984
rect 8938 38972 8944 39024
rect 8996 39012 9002 39024
rect 9582 39012 9588 39024
rect 8996 38984 9588 39012
rect 8996 38972 9002 38984
rect 9582 38972 9588 38984
rect 9640 38972 9646 39024
rect 10962 38972 10968 39024
rect 11020 39012 11026 39024
rect 12820 39012 12848 39052
rect 16114 39040 16120 39052
rect 16172 39040 16178 39092
rect 18598 39040 18604 39092
rect 18656 39040 18662 39092
rect 19426 39040 19432 39092
rect 19484 39040 19490 39092
rect 20990 39040 20996 39092
rect 21048 39040 21054 39092
rect 21082 39040 21088 39092
rect 21140 39040 21146 39092
rect 21913 39083 21971 39089
rect 21913 39049 21925 39083
rect 21959 39080 21971 39083
rect 22097 39083 22155 39089
rect 22097 39080 22109 39083
rect 21959 39052 22109 39080
rect 21959 39049 21971 39052
rect 21913 39043 21971 39049
rect 22097 39049 22109 39052
rect 22143 39080 22155 39083
rect 22830 39080 22836 39092
rect 22143 39052 22836 39080
rect 22143 39049 22155 39052
rect 22097 39043 22155 39049
rect 22830 39040 22836 39052
rect 22888 39080 22894 39092
rect 22888 39052 23980 39080
rect 22888 39040 22894 39052
rect 11020 38984 12848 39012
rect 11020 38972 11026 38984
rect 14642 38972 14648 39024
rect 14700 39012 14706 39024
rect 15470 39012 15476 39024
rect 14700 38984 15476 39012
rect 14700 38972 14706 38984
rect 15470 38972 15476 38984
rect 15528 39012 15534 39024
rect 17129 39015 17187 39021
rect 15528 38984 16896 39012
rect 15528 38972 15534 38984
rect 7742 38904 7748 38956
rect 7800 38904 7806 38956
rect 7834 38904 7840 38956
rect 7892 38944 7898 38956
rect 10781 38947 10839 38953
rect 7892 38916 9812 38944
rect 7892 38904 7898 38916
rect 7009 38879 7067 38885
rect 7009 38845 7021 38879
rect 7055 38845 7067 38879
rect 7009 38839 7067 38845
rect 7101 38879 7159 38885
rect 7101 38845 7113 38879
rect 7147 38845 7159 38879
rect 7101 38839 7159 38845
rect 7024 38808 7052 38839
rect 9582 38836 9588 38888
rect 9640 38836 9646 38888
rect 9784 38885 9812 38916
rect 10781 38913 10793 38947
rect 10827 38944 10839 38947
rect 11698 38944 11704 38956
rect 10827 38916 11704 38944
rect 10827 38913 10839 38916
rect 10781 38907 10839 38913
rect 11698 38904 11704 38916
rect 11756 38904 11762 38956
rect 12621 38947 12679 38953
rect 12621 38913 12633 38947
rect 12667 38944 12679 38947
rect 12710 38944 12716 38956
rect 12667 38916 12716 38944
rect 12667 38913 12679 38916
rect 12621 38907 12679 38913
rect 12710 38904 12716 38916
rect 12768 38944 12774 38956
rect 13078 38944 13084 38956
rect 12768 38916 13084 38944
rect 12768 38904 12774 38916
rect 13078 38904 13084 38916
rect 13136 38904 13142 38956
rect 13449 38947 13507 38953
rect 13449 38913 13461 38947
rect 13495 38944 13507 38947
rect 14734 38944 14740 38956
rect 13495 38916 14740 38944
rect 13495 38913 13507 38916
rect 13449 38907 13507 38913
rect 14734 38904 14740 38916
rect 14792 38904 14798 38956
rect 15289 38947 15347 38953
rect 15289 38913 15301 38947
rect 15335 38944 15347 38947
rect 16666 38944 16672 38956
rect 15335 38916 16672 38944
rect 15335 38913 15347 38916
rect 15289 38907 15347 38913
rect 16666 38904 16672 38916
rect 16724 38904 16730 38956
rect 16868 38953 16896 38984
rect 17129 38981 17141 39015
rect 17175 39012 17187 39015
rect 17218 39012 17224 39024
rect 17175 38984 17224 39012
rect 17175 38981 17187 38984
rect 17129 38975 17187 38981
rect 17218 38972 17224 38984
rect 17276 38972 17282 39024
rect 18877 39015 18935 39021
rect 18877 39012 18889 39015
rect 18354 38984 18889 39012
rect 18877 38981 18889 38984
rect 18923 39012 18935 39015
rect 18966 39012 18972 39024
rect 18923 38984 18972 39012
rect 18923 38981 18935 38984
rect 18877 38975 18935 38981
rect 18966 38972 18972 38984
rect 19024 38972 19030 39024
rect 19797 39015 19855 39021
rect 19797 38981 19809 39015
rect 19843 39012 19855 39015
rect 19886 39012 19892 39024
rect 19843 38984 19892 39012
rect 19843 38981 19855 38984
rect 19797 38975 19855 38981
rect 19886 38972 19892 38984
rect 19944 38972 19950 39024
rect 23952 39012 23980 39052
rect 25222 39040 25228 39092
rect 25280 39040 25286 39092
rect 24394 39012 24400 39024
rect 23874 38984 24400 39012
rect 24394 38972 24400 38984
rect 24452 39012 24458 39024
rect 24452 38984 24992 39012
rect 24452 38972 24458 38984
rect 16853 38947 16911 38953
rect 16853 38913 16865 38947
rect 16899 38913 16911 38947
rect 16853 38907 16911 38913
rect 19518 38904 19524 38956
rect 19576 38944 19582 38956
rect 19576 38916 20024 38944
rect 19576 38904 19582 38916
rect 9769 38879 9827 38885
rect 9769 38845 9781 38879
rect 9815 38876 9827 38879
rect 9815 38848 10272 38876
rect 9815 38845 9827 38848
rect 9769 38839 9827 38845
rect 8938 38808 8944 38820
rect 7024 38780 8944 38808
rect 8938 38768 8944 38780
rect 8996 38768 9002 38820
rect 9125 38811 9183 38817
rect 9125 38777 9137 38811
rect 9171 38808 9183 38811
rect 10134 38808 10140 38820
rect 9171 38780 10140 38808
rect 9171 38777 9183 38780
rect 9125 38771 9183 38777
rect 10134 38768 10140 38780
rect 10192 38768 10198 38820
rect 10244 38808 10272 38848
rect 10870 38836 10876 38888
rect 10928 38836 10934 38888
rect 10965 38879 11023 38885
rect 10965 38845 10977 38879
rect 11011 38876 11023 38879
rect 12526 38876 12532 38888
rect 11011 38848 12532 38876
rect 11011 38845 11023 38848
rect 10965 38839 11023 38845
rect 12526 38836 12532 38848
rect 12584 38836 12590 38888
rect 12805 38879 12863 38885
rect 12805 38845 12817 38879
rect 12851 38845 12863 38879
rect 12805 38839 12863 38845
rect 12820 38808 12848 38839
rect 12986 38836 12992 38888
rect 13044 38876 13050 38888
rect 15102 38876 15108 38888
rect 13044 38848 15108 38876
rect 13044 38836 13050 38848
rect 15102 38836 15108 38848
rect 15160 38836 15166 38888
rect 15378 38836 15384 38888
rect 15436 38836 15442 38888
rect 15565 38879 15623 38885
rect 15565 38845 15577 38879
rect 15611 38876 15623 38879
rect 15746 38876 15752 38888
rect 15611 38848 15752 38876
rect 15611 38845 15623 38848
rect 15565 38839 15623 38845
rect 15746 38836 15752 38848
rect 15804 38836 15810 38888
rect 19996 38885 20024 38916
rect 24486 38904 24492 38956
rect 24544 38944 24550 38956
rect 24581 38947 24639 38953
rect 24581 38944 24593 38947
rect 24544 38916 24593 38944
rect 24544 38904 24550 38916
rect 24581 38913 24593 38916
rect 24627 38913 24639 38947
rect 24581 38907 24639 38913
rect 19889 38879 19947 38885
rect 19889 38845 19901 38879
rect 19935 38845 19947 38879
rect 19889 38839 19947 38845
rect 19981 38879 20039 38885
rect 19981 38845 19993 38879
rect 20027 38845 20039 38879
rect 19981 38839 20039 38845
rect 10244 38780 12848 38808
rect 13814 38768 13820 38820
rect 13872 38808 13878 38820
rect 15654 38808 15660 38820
rect 13872 38780 15660 38808
rect 13872 38768 13878 38780
rect 15654 38768 15660 38780
rect 15712 38768 15718 38820
rect 19904 38808 19932 38839
rect 21266 38836 21272 38888
rect 21324 38836 21330 38888
rect 22370 38836 22376 38888
rect 22428 38836 22434 38888
rect 22649 38879 22707 38885
rect 22649 38845 22661 38879
rect 22695 38876 22707 38879
rect 24854 38876 24860 38888
rect 22695 38848 24860 38876
rect 22695 38845 22707 38848
rect 22649 38839 22707 38845
rect 24854 38836 24860 38848
rect 24912 38836 24918 38888
rect 20530 38808 20536 38820
rect 19904 38780 20536 38808
rect 20530 38768 20536 38780
rect 20588 38808 20594 38820
rect 22002 38808 22008 38820
rect 20588 38780 22008 38808
rect 20588 38768 20594 38780
rect 22002 38768 22008 38780
rect 22060 38768 22066 38820
rect 6822 38700 6828 38752
rect 6880 38740 6886 38752
rect 8389 38743 8447 38749
rect 8389 38740 8401 38743
rect 6880 38712 8401 38740
rect 6880 38700 6886 38712
rect 8389 38709 8401 38712
rect 8435 38709 8447 38743
rect 8389 38703 8447 38709
rect 8849 38743 8907 38749
rect 8849 38709 8861 38743
rect 8895 38740 8907 38743
rect 9582 38740 9588 38752
rect 8895 38712 9588 38740
rect 8895 38709 8907 38712
rect 8849 38703 8907 38709
rect 9582 38700 9588 38712
rect 9640 38740 9646 38752
rect 12158 38740 12164 38752
rect 9640 38712 12164 38740
rect 9640 38700 9646 38712
rect 12158 38700 12164 38712
rect 12216 38740 12222 38752
rect 13998 38740 14004 38752
rect 12216 38712 14004 38740
rect 12216 38700 12222 38712
rect 13998 38700 14004 38712
rect 14056 38700 14062 38752
rect 14090 38700 14096 38752
rect 14148 38700 14154 38752
rect 14182 38700 14188 38752
rect 14240 38740 14246 38752
rect 14921 38743 14979 38749
rect 14921 38740 14933 38743
rect 14240 38712 14933 38740
rect 14240 38700 14246 38712
rect 14921 38709 14933 38712
rect 14967 38709 14979 38743
rect 14921 38703 14979 38709
rect 15378 38700 15384 38752
rect 15436 38740 15442 38752
rect 15930 38740 15936 38752
rect 15436 38712 15936 38740
rect 15436 38700 15442 38712
rect 15930 38700 15936 38712
rect 15988 38700 15994 38752
rect 20625 38743 20683 38749
rect 20625 38709 20637 38743
rect 20671 38740 20683 38743
rect 21358 38740 21364 38752
rect 20671 38712 21364 38740
rect 20671 38709 20683 38712
rect 20625 38703 20683 38709
rect 21358 38700 21364 38712
rect 21416 38700 21422 38752
rect 24026 38700 24032 38752
rect 24084 38740 24090 38752
rect 24121 38743 24179 38749
rect 24121 38740 24133 38743
rect 24084 38712 24133 38740
rect 24084 38700 24090 38712
rect 24121 38709 24133 38712
rect 24167 38709 24179 38743
rect 24121 38703 24179 38709
rect 24854 38700 24860 38752
rect 24912 38740 24918 38752
rect 24964 38740 24992 38984
rect 24912 38712 24992 38740
rect 24912 38700 24918 38712
rect 1104 38650 25852 38672
rect 1104 38598 2950 38650
rect 3002 38598 3014 38650
rect 3066 38598 3078 38650
rect 3130 38598 3142 38650
rect 3194 38598 3206 38650
rect 3258 38598 12950 38650
rect 13002 38598 13014 38650
rect 13066 38598 13078 38650
rect 13130 38598 13142 38650
rect 13194 38598 13206 38650
rect 13258 38598 22950 38650
rect 23002 38598 23014 38650
rect 23066 38598 23078 38650
rect 23130 38598 23142 38650
rect 23194 38598 23206 38650
rect 23258 38598 25852 38650
rect 1104 38576 25852 38598
rect 6086 38496 6092 38548
rect 6144 38536 6150 38548
rect 6144 38508 7236 38536
rect 6144 38496 6150 38508
rect 5166 38360 5172 38412
rect 5224 38400 5230 38412
rect 5445 38403 5503 38409
rect 5445 38400 5457 38403
rect 5224 38372 5457 38400
rect 5224 38360 5230 38372
rect 5445 38369 5457 38372
rect 5491 38400 5503 38403
rect 7208 38400 7236 38508
rect 7558 38496 7564 38548
rect 7616 38536 7622 38548
rect 7653 38539 7711 38545
rect 7653 38536 7665 38539
rect 7616 38508 7665 38536
rect 7616 38496 7622 38508
rect 7653 38505 7665 38508
rect 7699 38505 7711 38539
rect 7653 38499 7711 38505
rect 10413 38539 10471 38545
rect 10413 38505 10425 38539
rect 10459 38536 10471 38539
rect 10502 38536 10508 38548
rect 10459 38508 10508 38536
rect 10459 38505 10471 38508
rect 10413 38499 10471 38505
rect 10502 38496 10508 38508
rect 10560 38496 10566 38548
rect 12240 38539 12298 38545
rect 12240 38505 12252 38539
rect 12286 38536 12298 38539
rect 14090 38536 14096 38548
rect 12286 38508 14096 38536
rect 12286 38505 12298 38508
rect 12240 38499 12298 38505
rect 14090 38496 14096 38508
rect 14148 38496 14154 38548
rect 15102 38496 15108 38548
rect 15160 38536 15166 38548
rect 16209 38539 16267 38545
rect 15160 38508 15976 38536
rect 15160 38496 15166 38508
rect 9214 38428 9220 38480
rect 9272 38468 9278 38480
rect 9272 38440 12112 38468
rect 9272 38428 9278 38440
rect 8205 38403 8263 38409
rect 8205 38400 8217 38403
rect 5491 38372 7144 38400
rect 7208 38372 8217 38400
rect 5491 38369 5503 38372
rect 5445 38363 5503 38369
rect 1302 38292 1308 38344
rect 1360 38332 1366 38344
rect 1765 38335 1823 38341
rect 1765 38332 1777 38335
rect 1360 38304 1777 38332
rect 1360 38292 1366 38304
rect 1765 38301 1777 38304
rect 1811 38332 1823 38335
rect 2041 38335 2099 38341
rect 2041 38332 2053 38335
rect 1811 38304 2053 38332
rect 1811 38301 1823 38304
rect 1765 38295 1823 38301
rect 2041 38301 2053 38304
rect 2087 38301 2099 38335
rect 7116 38332 7144 38372
rect 8205 38369 8217 38372
rect 8251 38369 8263 38403
rect 8205 38363 8263 38369
rect 9674 38360 9680 38412
rect 9732 38360 9738 38412
rect 9769 38403 9827 38409
rect 9769 38369 9781 38403
rect 9815 38369 9827 38403
rect 9769 38363 9827 38369
rect 8665 38335 8723 38341
rect 8665 38332 8677 38335
rect 7116 38304 8677 38332
rect 2041 38295 2099 38301
rect 8665 38301 8677 38304
rect 8711 38301 8723 38335
rect 9784 38332 9812 38363
rect 9858 38360 9864 38412
rect 9916 38400 9922 38412
rect 10962 38400 10968 38412
rect 9916 38372 10968 38400
rect 9916 38360 9922 38372
rect 10962 38360 10968 38372
rect 11020 38360 11026 38412
rect 11974 38360 11980 38412
rect 12032 38360 12038 38412
rect 12084 38400 12112 38440
rect 13354 38428 13360 38480
rect 13412 38468 13418 38480
rect 13725 38471 13783 38477
rect 13725 38468 13737 38471
rect 13412 38440 13737 38468
rect 13412 38428 13418 38440
rect 13725 38437 13737 38440
rect 13771 38437 13783 38471
rect 15841 38471 15899 38477
rect 15841 38468 15853 38471
rect 13725 38431 13783 38437
rect 13832 38440 15853 38468
rect 12618 38400 12624 38412
rect 12084 38372 12624 38400
rect 12618 38360 12624 38372
rect 12676 38400 12682 38412
rect 13832 38400 13860 38440
rect 15841 38437 15853 38440
rect 15887 38437 15899 38471
rect 15948 38468 15976 38508
rect 16209 38505 16221 38539
rect 16255 38536 16267 38539
rect 16574 38536 16580 38548
rect 16255 38508 16580 38536
rect 16255 38505 16267 38508
rect 16209 38499 16267 38505
rect 16574 38496 16580 38508
rect 16632 38496 16638 38548
rect 17405 38539 17463 38545
rect 17405 38536 17417 38539
rect 16684 38508 17417 38536
rect 16684 38468 16712 38508
rect 17405 38505 17417 38508
rect 17451 38505 17463 38539
rect 17405 38499 17463 38505
rect 18690 38496 18696 38548
rect 18748 38536 18754 38548
rect 18785 38539 18843 38545
rect 18785 38536 18797 38539
rect 18748 38508 18797 38536
rect 18748 38496 18754 38508
rect 18785 38505 18797 38508
rect 18831 38505 18843 38539
rect 18785 38499 18843 38505
rect 21542 38496 21548 38548
rect 21600 38536 21606 38548
rect 24670 38536 24676 38548
rect 21600 38508 24676 38536
rect 21600 38496 21606 38508
rect 24670 38496 24676 38508
rect 24728 38496 24734 38548
rect 18506 38468 18512 38480
rect 15948 38440 16712 38468
rect 16868 38440 18512 38468
rect 15841 38431 15899 38437
rect 12676 38372 13860 38400
rect 14277 38403 14335 38409
rect 12676 38360 12682 38372
rect 14277 38369 14289 38403
rect 14323 38400 14335 38403
rect 14826 38400 14832 38412
rect 14323 38372 14832 38400
rect 14323 38369 14335 38372
rect 14277 38363 14335 38369
rect 14826 38360 14832 38372
rect 14884 38360 14890 38412
rect 15856 38400 15884 38431
rect 16868 38409 16896 38440
rect 18506 38428 18512 38440
rect 18564 38428 18570 38480
rect 22094 38428 22100 38480
rect 22152 38468 22158 38480
rect 24121 38471 24179 38477
rect 24121 38468 24133 38471
rect 22152 38440 24133 38468
rect 22152 38428 22158 38440
rect 24121 38437 24133 38440
rect 24167 38437 24179 38471
rect 24121 38431 24179 38437
rect 24578 38428 24584 38480
rect 24636 38428 24642 38480
rect 16669 38403 16727 38409
rect 16669 38400 16681 38403
rect 15856 38372 16681 38400
rect 16669 38369 16681 38372
rect 16715 38369 16727 38403
rect 16669 38363 16727 38369
rect 16853 38403 16911 38409
rect 16853 38369 16865 38403
rect 16899 38369 16911 38403
rect 16853 38363 16911 38369
rect 17494 38360 17500 38412
rect 17552 38400 17558 38412
rect 17957 38403 18015 38409
rect 17957 38400 17969 38403
rect 17552 38372 17969 38400
rect 17552 38360 17558 38372
rect 17957 38369 17969 38372
rect 18003 38369 18015 38403
rect 17957 38363 18015 38369
rect 18414 38360 18420 38412
rect 18472 38400 18478 38412
rect 21542 38400 21548 38412
rect 18472 38372 21548 38400
rect 18472 38360 18478 38372
rect 21542 38360 21548 38372
rect 21600 38360 21606 38412
rect 22278 38360 22284 38412
rect 22336 38400 22342 38412
rect 23201 38403 23259 38409
rect 23201 38400 23213 38403
rect 22336 38372 23213 38400
rect 22336 38360 22342 38372
rect 23201 38369 23213 38372
rect 23247 38369 23259 38403
rect 23201 38363 23259 38369
rect 23293 38403 23351 38409
rect 23293 38369 23305 38403
rect 23339 38400 23351 38403
rect 24026 38400 24032 38412
rect 23339 38372 24032 38400
rect 23339 38369 23351 38372
rect 23293 38363 23351 38369
rect 8665 38295 8723 38301
rect 8772 38304 9812 38332
rect 5721 38267 5779 38273
rect 5721 38233 5733 38267
rect 5767 38264 5779 38267
rect 5994 38264 6000 38276
rect 5767 38236 6000 38264
rect 5767 38233 5779 38236
rect 5721 38227 5779 38233
rect 5994 38224 6000 38236
rect 6052 38224 6058 38276
rect 6454 38224 6460 38276
rect 6512 38224 6518 38276
rect 7006 38224 7012 38276
rect 7064 38264 7070 38276
rect 8772 38264 8800 38304
rect 10042 38292 10048 38344
rect 10100 38332 10106 38344
rect 10781 38335 10839 38341
rect 10781 38332 10793 38335
rect 10100 38304 10793 38332
rect 10100 38292 10106 38304
rect 10781 38301 10793 38304
rect 10827 38301 10839 38335
rect 10781 38295 10839 38301
rect 15838 38292 15844 38344
rect 15896 38332 15902 38344
rect 17126 38332 17132 38344
rect 15896 38304 17132 38332
rect 15896 38292 15902 38304
rect 17126 38292 17132 38304
rect 17184 38332 17190 38344
rect 18601 38335 18659 38341
rect 18601 38332 18613 38335
rect 17184 38304 18613 38332
rect 17184 38292 17190 38304
rect 18601 38301 18613 38304
rect 18647 38332 18659 38335
rect 19429 38335 19487 38341
rect 19429 38332 19441 38335
rect 18647 38304 19441 38332
rect 18647 38301 18659 38304
rect 18601 38295 18659 38301
rect 19429 38301 19441 38304
rect 19475 38332 19487 38335
rect 20993 38335 21051 38341
rect 20993 38332 21005 38335
rect 19475 38304 21005 38332
rect 19475 38301 19487 38304
rect 19429 38295 19487 38301
rect 20993 38301 21005 38304
rect 21039 38332 21051 38335
rect 21361 38335 21419 38341
rect 21361 38332 21373 38335
rect 21039 38304 21373 38332
rect 21039 38301 21051 38304
rect 20993 38295 21051 38301
rect 21361 38301 21373 38304
rect 21407 38301 21419 38335
rect 23109 38335 23167 38341
rect 23109 38332 23121 38335
rect 21361 38295 21419 38301
rect 22066 38304 23121 38332
rect 22066 38276 22094 38304
rect 23109 38301 23121 38304
rect 23155 38301 23167 38335
rect 23308 38332 23336 38363
rect 24026 38360 24032 38372
rect 24084 38360 24090 38412
rect 24394 38360 24400 38412
rect 24452 38400 24458 38412
rect 25133 38403 25191 38409
rect 25133 38400 25145 38403
rect 24452 38372 25145 38400
rect 24452 38360 24458 38372
rect 25133 38369 25145 38372
rect 25179 38369 25191 38403
rect 25133 38363 25191 38369
rect 23109 38295 23167 38301
rect 23216 38304 23336 38332
rect 23216 38276 23244 38304
rect 23474 38292 23480 38344
rect 23532 38332 23538 38344
rect 24949 38335 25007 38341
rect 24949 38332 24961 38335
rect 23532 38304 24961 38332
rect 23532 38292 23538 38304
rect 24949 38301 24961 38304
rect 24995 38301 25007 38335
rect 24949 38295 25007 38301
rect 25041 38335 25099 38341
rect 25041 38301 25053 38335
rect 25087 38332 25099 38335
rect 25406 38332 25412 38344
rect 25087 38304 25412 38332
rect 25087 38301 25099 38304
rect 25041 38295 25099 38301
rect 25406 38292 25412 38304
rect 25464 38292 25470 38344
rect 7064 38236 8800 38264
rect 9585 38267 9643 38273
rect 7064 38224 7070 38236
rect 9585 38233 9597 38267
rect 9631 38264 9643 38267
rect 11238 38264 11244 38276
rect 9631 38236 11244 38264
rect 9631 38233 9643 38236
rect 9585 38227 9643 38233
rect 11238 38224 11244 38236
rect 11296 38224 11302 38276
rect 13630 38264 13636 38276
rect 13478 38236 13636 38264
rect 13630 38224 13636 38236
rect 13688 38224 13694 38276
rect 17494 38264 17500 38276
rect 15304 38236 17500 38264
rect 1581 38199 1639 38205
rect 1581 38165 1593 38199
rect 1627 38196 1639 38199
rect 3878 38196 3884 38208
rect 1627 38168 3884 38196
rect 1627 38165 1639 38168
rect 1581 38159 1639 38165
rect 3878 38156 3884 38168
rect 3936 38156 3942 38208
rect 7193 38199 7251 38205
rect 7193 38165 7205 38199
rect 7239 38196 7251 38199
rect 7742 38196 7748 38208
rect 7239 38168 7748 38196
rect 7239 38165 7251 38168
rect 7193 38159 7251 38165
rect 7742 38156 7748 38168
rect 7800 38156 7806 38208
rect 7834 38156 7840 38208
rect 7892 38196 7898 38208
rect 8021 38199 8079 38205
rect 8021 38196 8033 38199
rect 7892 38168 8033 38196
rect 7892 38156 7898 38168
rect 8021 38165 8033 38168
rect 8067 38165 8079 38199
rect 8021 38159 8079 38165
rect 8113 38199 8171 38205
rect 8113 38165 8125 38199
rect 8159 38196 8171 38199
rect 9217 38199 9275 38205
rect 9217 38196 9229 38199
rect 8159 38168 9229 38196
rect 8159 38165 8171 38168
rect 8113 38159 8171 38165
rect 9217 38165 9229 38168
rect 9263 38165 9275 38199
rect 9217 38159 9275 38165
rect 9858 38156 9864 38208
rect 9916 38196 9922 38208
rect 10686 38196 10692 38208
rect 9916 38168 10692 38196
rect 9916 38156 9922 38168
rect 10686 38156 10692 38168
rect 10744 38196 10750 38208
rect 10873 38199 10931 38205
rect 10873 38196 10885 38199
rect 10744 38168 10885 38196
rect 10744 38156 10750 38168
rect 10873 38165 10885 38168
rect 10919 38165 10931 38199
rect 10873 38159 10931 38165
rect 10962 38156 10968 38208
rect 11020 38196 11026 38208
rect 15304 38196 15332 38236
rect 17494 38224 17500 38236
rect 17552 38224 17558 38276
rect 17773 38267 17831 38273
rect 17773 38233 17785 38267
rect 17819 38264 17831 38267
rect 18782 38264 18788 38276
rect 17819 38236 18788 38264
rect 17819 38233 17831 38236
rect 17773 38227 17831 38233
rect 18782 38224 18788 38236
rect 18840 38224 18846 38276
rect 20162 38224 20168 38276
rect 20220 38224 20226 38276
rect 22002 38224 22008 38276
rect 22060 38236 22094 38276
rect 22189 38267 22247 38273
rect 22060 38224 22066 38236
rect 22189 38233 22201 38267
rect 22235 38264 22247 38267
rect 22370 38264 22376 38276
rect 22235 38236 22376 38264
rect 22235 38233 22247 38236
rect 22189 38227 22247 38233
rect 22370 38224 22376 38236
rect 22428 38264 22434 38276
rect 22830 38264 22836 38276
rect 22428 38236 22836 38264
rect 22428 38224 22434 38236
rect 22830 38224 22836 38236
rect 22888 38224 22894 38276
rect 23198 38224 23204 38276
rect 23256 38224 23262 38276
rect 24029 38267 24087 38273
rect 24029 38233 24041 38267
rect 24075 38264 24087 38267
rect 24670 38264 24676 38276
rect 24075 38236 24676 38264
rect 24075 38233 24087 38236
rect 24029 38227 24087 38233
rect 24670 38224 24676 38236
rect 24728 38224 24734 38276
rect 11020 38168 15332 38196
rect 11020 38156 11026 38168
rect 15378 38156 15384 38208
rect 15436 38156 15442 38208
rect 16574 38156 16580 38208
rect 16632 38156 16638 38208
rect 17865 38199 17923 38205
rect 17865 38165 17877 38199
rect 17911 38196 17923 38199
rect 18414 38196 18420 38208
rect 17911 38168 18420 38196
rect 17911 38165 17923 38168
rect 17865 38159 17923 38165
rect 18414 38156 18420 38168
rect 18472 38156 18478 38208
rect 18874 38156 18880 38208
rect 18932 38196 18938 38208
rect 18969 38199 19027 38205
rect 18969 38196 18981 38199
rect 18932 38168 18981 38196
rect 18932 38156 18938 38168
rect 18969 38165 18981 38168
rect 19015 38196 19027 38199
rect 19058 38196 19064 38208
rect 19015 38168 19064 38196
rect 19015 38165 19027 38168
rect 18969 38159 19027 38165
rect 19058 38156 19064 38168
rect 19116 38156 19122 38208
rect 22738 38156 22744 38208
rect 22796 38156 22802 38208
rect 22922 38156 22928 38208
rect 22980 38196 22986 38208
rect 23845 38199 23903 38205
rect 23845 38196 23857 38199
rect 22980 38168 23857 38196
rect 22980 38156 22986 38168
rect 23845 38165 23857 38168
rect 23891 38196 23903 38199
rect 25590 38196 25596 38208
rect 23891 38168 25596 38196
rect 23891 38165 23903 38168
rect 23845 38159 23903 38165
rect 25590 38156 25596 38168
rect 25648 38156 25654 38208
rect 1104 38106 25852 38128
rect 1104 38054 7950 38106
rect 8002 38054 8014 38106
rect 8066 38054 8078 38106
rect 8130 38054 8142 38106
rect 8194 38054 8206 38106
rect 8258 38054 17950 38106
rect 18002 38054 18014 38106
rect 18066 38054 18078 38106
rect 18130 38054 18142 38106
rect 18194 38054 18206 38106
rect 18258 38054 25852 38106
rect 1104 38032 25852 38054
rect 5994 37952 6000 38004
rect 6052 37952 6058 38004
rect 6638 37952 6644 38004
rect 6696 37992 6702 38004
rect 6696 37964 8984 37992
rect 6696 37952 6702 37964
rect 6822 37884 6828 37936
rect 6880 37884 6886 37936
rect 8202 37924 8208 37936
rect 8050 37896 8208 37924
rect 8202 37884 8208 37896
rect 8260 37924 8266 37936
rect 8662 37924 8668 37936
rect 8260 37896 8668 37924
rect 8260 37884 8266 37896
rect 8662 37884 8668 37896
rect 8720 37924 8726 37936
rect 8849 37927 8907 37933
rect 8849 37924 8861 37927
rect 8720 37896 8861 37924
rect 8720 37884 8726 37896
rect 8849 37893 8861 37896
rect 8895 37893 8907 37927
rect 8956 37924 8984 37964
rect 9030 37952 9036 38004
rect 9088 37992 9094 38004
rect 9401 37995 9459 38001
rect 9401 37992 9413 37995
rect 9088 37964 9413 37992
rect 9088 37952 9094 37964
rect 9401 37961 9413 37964
rect 9447 37961 9459 37995
rect 9401 37955 9459 37961
rect 9490 37952 9496 38004
rect 9548 37992 9554 38004
rect 10594 37992 10600 38004
rect 9548 37964 10600 37992
rect 9548 37952 9554 37964
rect 10594 37952 10600 37964
rect 10652 37992 10658 38004
rect 10962 37992 10968 38004
rect 10652 37964 10968 37992
rect 10652 37952 10658 37964
rect 10962 37952 10968 37964
rect 11020 37952 11026 38004
rect 11333 37995 11391 38001
rect 11333 37961 11345 37995
rect 11379 37992 11391 37995
rect 11422 37992 11428 38004
rect 11379 37964 11428 37992
rect 11379 37961 11391 37964
rect 11333 37955 11391 37961
rect 11422 37952 11428 37964
rect 11480 37952 11486 38004
rect 11698 37952 11704 38004
rect 11756 37952 11762 38004
rect 13630 37952 13636 38004
rect 13688 37992 13694 38004
rect 13909 37995 13967 38001
rect 13909 37992 13921 37995
rect 13688 37964 13921 37992
rect 13688 37952 13694 37964
rect 13909 37961 13921 37964
rect 13955 37992 13967 37995
rect 13998 37992 14004 38004
rect 13955 37964 14004 37992
rect 13955 37961 13967 37964
rect 13909 37955 13967 37961
rect 13998 37952 14004 37964
rect 14056 37952 14062 38004
rect 15378 37952 15384 38004
rect 15436 37952 15442 38004
rect 16574 37952 16580 38004
rect 16632 37992 16638 38004
rect 16853 37995 16911 38001
rect 16853 37992 16865 37995
rect 16632 37964 16865 37992
rect 16632 37952 16638 37964
rect 16853 37961 16865 37964
rect 16899 37961 16911 37995
rect 16853 37955 16911 37961
rect 17494 37952 17500 38004
rect 17552 37952 17558 38004
rect 18325 37995 18383 38001
rect 18325 37961 18337 37995
rect 18371 37992 18383 37995
rect 18690 37992 18696 38004
rect 18371 37964 18696 37992
rect 18371 37961 18383 37964
rect 18325 37955 18383 37961
rect 18690 37952 18696 37964
rect 18748 37952 18754 38004
rect 19610 37952 19616 38004
rect 19668 37992 19674 38004
rect 21085 37995 21143 38001
rect 21085 37992 21097 37995
rect 19668 37964 21097 37992
rect 19668 37952 19674 37964
rect 21085 37961 21097 37964
rect 21131 37961 21143 37995
rect 21085 37955 21143 37961
rect 22002 37952 22008 38004
rect 22060 37952 22066 38004
rect 22094 37952 22100 38004
rect 22152 37992 22158 38004
rect 22373 37995 22431 38001
rect 22373 37992 22385 37995
rect 22152 37964 22385 37992
rect 22152 37952 22158 37964
rect 22373 37961 22385 37964
rect 22419 37961 22431 37995
rect 22373 37955 22431 37961
rect 22646 37952 22652 38004
rect 22704 37992 22710 38004
rect 23017 37995 23075 38001
rect 23017 37992 23029 37995
rect 22704 37964 23029 37992
rect 22704 37952 22710 37964
rect 23017 37961 23029 37964
rect 23063 37961 23075 37995
rect 24210 37992 24216 38004
rect 23017 37955 23075 37961
rect 23584 37964 24216 37992
rect 10413 37927 10471 37933
rect 10413 37924 10425 37927
rect 8956 37896 10425 37924
rect 8849 37887 8907 37893
rect 10413 37893 10425 37896
rect 10459 37924 10471 37927
rect 10502 37924 10508 37936
rect 10459 37896 10508 37924
rect 10459 37893 10471 37896
rect 10413 37887 10471 37893
rect 5353 37859 5411 37865
rect 5353 37825 5365 37859
rect 5399 37825 5411 37859
rect 8864 37856 8892 37887
rect 10502 37884 10508 37896
rect 10560 37884 10566 37936
rect 10686 37884 10692 37936
rect 10744 37884 10750 37936
rect 11514 37884 11520 37936
rect 11572 37924 11578 37936
rect 20993 37927 21051 37933
rect 20993 37924 21005 37927
rect 11572 37896 15608 37924
rect 11572 37884 11578 37896
rect 9033 37859 9091 37865
rect 9033 37856 9045 37859
rect 8864 37828 9045 37856
rect 5353 37819 5411 37825
rect 9033 37825 9045 37828
rect 9079 37825 9091 37859
rect 9033 37819 9091 37825
rect 5368 37652 5396 37819
rect 9398 37816 9404 37868
rect 9456 37856 9462 37868
rect 9769 37859 9827 37865
rect 9769 37856 9781 37859
rect 9456 37828 9781 37856
rect 9456 37816 9462 37828
rect 9769 37825 9781 37828
rect 9815 37825 9827 37859
rect 9769 37819 9827 37825
rect 9861 37859 9919 37865
rect 9861 37825 9873 37859
rect 9907 37856 9919 37859
rect 11330 37856 11336 37868
rect 9907 37828 11336 37856
rect 9907 37825 9919 37828
rect 9861 37819 9919 37825
rect 11330 37816 11336 37828
rect 11388 37816 11394 37868
rect 12897 37859 12955 37865
rect 12897 37825 12909 37859
rect 12943 37856 12955 37859
rect 13817 37859 13875 37865
rect 13817 37856 13829 37859
rect 12943 37828 13829 37856
rect 12943 37825 12955 37828
rect 12897 37819 12955 37825
rect 13817 37825 13829 37828
rect 13863 37856 13875 37859
rect 15102 37856 15108 37868
rect 13863 37828 15108 37856
rect 13863 37825 13875 37828
rect 13817 37819 13875 37825
rect 15102 37816 15108 37828
rect 15160 37816 15166 37868
rect 6546 37748 6552 37800
rect 6604 37748 6610 37800
rect 7190 37748 7196 37800
rect 7248 37788 7254 37800
rect 8573 37791 8631 37797
rect 8573 37788 8585 37791
rect 7248 37760 8585 37788
rect 7248 37748 7254 37760
rect 8573 37757 8585 37760
rect 8619 37757 8631 37791
rect 8573 37751 8631 37757
rect 9953 37791 10011 37797
rect 9953 37757 9965 37791
rect 9999 37757 10011 37791
rect 9953 37751 10011 37757
rect 8588 37720 8616 37751
rect 8588 37692 9536 37720
rect 8570 37652 8576 37664
rect 5368 37624 8576 37652
rect 8570 37612 8576 37624
rect 8628 37612 8634 37664
rect 9508 37652 9536 37692
rect 9582 37680 9588 37732
rect 9640 37720 9646 37732
rect 9968 37720 9996 37751
rect 11422 37748 11428 37800
rect 11480 37788 11486 37800
rect 12989 37791 13047 37797
rect 12989 37788 13001 37791
rect 11480 37760 13001 37788
rect 11480 37748 11486 37760
rect 12989 37757 13001 37760
rect 13035 37757 13047 37791
rect 12989 37751 13047 37757
rect 13173 37791 13231 37797
rect 13173 37757 13185 37791
rect 13219 37788 13231 37791
rect 13630 37788 13636 37800
rect 13219 37760 13636 37788
rect 13219 37757 13231 37760
rect 13173 37751 13231 37757
rect 13630 37748 13636 37760
rect 13688 37748 13694 37800
rect 15286 37748 15292 37800
rect 15344 37788 15350 37800
rect 15473 37791 15531 37797
rect 15473 37788 15485 37791
rect 15344 37760 15485 37788
rect 15344 37748 15350 37760
rect 15473 37757 15485 37760
rect 15519 37757 15531 37791
rect 15473 37751 15531 37757
rect 11514 37720 11520 37732
rect 9640 37692 9996 37720
rect 10520 37692 11520 37720
rect 9640 37680 9646 37692
rect 10520 37652 10548 37692
rect 11514 37680 11520 37692
rect 11572 37680 11578 37732
rect 11698 37680 11704 37732
rect 11756 37720 11762 37732
rect 15013 37723 15071 37729
rect 15013 37720 15025 37723
rect 11756 37692 15025 37720
rect 11756 37680 11762 37692
rect 15013 37689 15025 37692
rect 15059 37689 15071 37723
rect 15013 37683 15071 37689
rect 9508 37624 10548 37652
rect 12250 37612 12256 37664
rect 12308 37612 12314 37664
rect 12526 37612 12532 37664
rect 12584 37612 12590 37664
rect 12710 37612 12716 37664
rect 12768 37652 12774 37664
rect 13541 37655 13599 37661
rect 13541 37652 13553 37655
rect 12768 37624 13553 37652
rect 12768 37612 12774 37624
rect 13541 37621 13553 37624
rect 13587 37621 13599 37655
rect 13541 37615 13599 37621
rect 14274 37612 14280 37664
rect 14332 37652 14338 37664
rect 14645 37655 14703 37661
rect 14645 37652 14657 37655
rect 14332 37624 14657 37652
rect 14332 37612 14338 37624
rect 14645 37621 14657 37624
rect 14691 37652 14703 37655
rect 15378 37652 15384 37664
rect 14691 37624 15384 37652
rect 14691 37621 14703 37624
rect 14645 37615 14703 37621
rect 15378 37612 15384 37624
rect 15436 37612 15442 37664
rect 15580 37652 15608 37896
rect 17420 37896 21005 37924
rect 16206 37816 16212 37868
rect 16264 37856 16270 37868
rect 17420 37856 17448 37896
rect 20993 37893 21005 37896
rect 21039 37893 21051 37927
rect 20993 37887 21051 37893
rect 21910 37884 21916 37936
rect 21968 37924 21974 37936
rect 22465 37927 22523 37933
rect 22465 37924 22477 37927
rect 21968 37896 22477 37924
rect 21968 37884 21974 37896
rect 22465 37893 22477 37896
rect 22511 37924 22523 37927
rect 22922 37924 22928 37936
rect 22511 37896 22928 37924
rect 22511 37893 22523 37896
rect 22465 37887 22523 37893
rect 22922 37884 22928 37896
rect 22980 37884 22986 37936
rect 23293 37927 23351 37933
rect 23293 37893 23305 37927
rect 23339 37924 23351 37927
rect 23382 37924 23388 37936
rect 23339 37896 23388 37924
rect 23339 37893 23351 37896
rect 23293 37887 23351 37893
rect 23382 37884 23388 37896
rect 23440 37884 23446 37936
rect 16264 37828 17448 37856
rect 18417 37859 18475 37865
rect 16264 37816 16270 37828
rect 18417 37825 18429 37859
rect 18463 37856 18475 37859
rect 18874 37856 18880 37868
rect 18463 37828 18880 37856
rect 18463 37825 18475 37828
rect 18417 37819 18475 37825
rect 18874 37816 18880 37828
rect 18932 37816 18938 37868
rect 19334 37816 19340 37868
rect 19392 37856 19398 37868
rect 19521 37859 19579 37865
rect 19521 37856 19533 37859
rect 19392 37828 19533 37856
rect 19392 37816 19398 37828
rect 19521 37825 19533 37828
rect 19567 37825 19579 37859
rect 19521 37819 19579 37825
rect 19613 37859 19671 37865
rect 19613 37825 19625 37859
rect 19659 37856 19671 37859
rect 20257 37859 20315 37865
rect 20257 37856 20269 37859
rect 19659 37828 20269 37856
rect 19659 37825 19671 37828
rect 19613 37819 19671 37825
rect 20257 37825 20269 37828
rect 20303 37856 20315 37859
rect 20438 37856 20444 37868
rect 20303 37828 20444 37856
rect 20303 37825 20315 37828
rect 20257 37819 20315 37825
rect 20438 37816 20444 37828
rect 20496 37816 20502 37868
rect 21450 37856 21456 37868
rect 21100 37828 21456 37856
rect 15657 37791 15715 37797
rect 15657 37757 15669 37791
rect 15703 37788 15715 37791
rect 15746 37788 15752 37800
rect 15703 37760 15752 37788
rect 15703 37757 15715 37760
rect 15657 37751 15715 37757
rect 15746 37748 15752 37760
rect 15804 37748 15810 37800
rect 18509 37791 18567 37797
rect 18509 37757 18521 37791
rect 18555 37757 18567 37791
rect 18509 37751 18567 37757
rect 19797 37791 19855 37797
rect 19797 37757 19809 37791
rect 19843 37788 19855 37791
rect 21100 37788 21128 37828
rect 21450 37816 21456 37828
rect 21508 37816 21514 37868
rect 23584 37856 23612 37964
rect 24210 37952 24216 37964
rect 24268 37952 24274 38004
rect 24854 37884 24860 37936
rect 24912 37884 24918 37936
rect 22664 37828 23612 37856
rect 19843 37760 21128 37788
rect 19843 37757 19855 37760
rect 19797 37751 19855 37757
rect 16022 37680 16028 37732
rect 16080 37720 16086 37732
rect 17957 37723 18015 37729
rect 17957 37720 17969 37723
rect 16080 37692 17969 37720
rect 16080 37680 16086 37692
rect 17957 37689 17969 37692
rect 18003 37689 18015 37723
rect 17957 37683 18015 37689
rect 18414 37680 18420 37732
rect 18472 37720 18478 37732
rect 18524 37720 18552 37751
rect 21174 37748 21180 37800
rect 21232 37748 21238 37800
rect 22664 37797 22692 37828
rect 22649 37791 22707 37797
rect 22649 37757 22661 37791
rect 22695 37757 22707 37791
rect 22649 37751 22707 37757
rect 22830 37748 22836 37800
rect 22888 37788 22894 37800
rect 23569 37791 23627 37797
rect 23569 37788 23581 37791
rect 22888 37760 23581 37788
rect 22888 37748 22894 37760
rect 23569 37757 23581 37760
rect 23615 37757 23627 37791
rect 23569 37751 23627 37757
rect 23842 37748 23848 37800
rect 23900 37748 23906 37800
rect 18472 37692 18552 37720
rect 19153 37723 19211 37729
rect 18472 37680 18478 37692
rect 19153 37689 19165 37723
rect 19199 37720 19211 37723
rect 20714 37720 20720 37732
rect 19199 37692 20720 37720
rect 19199 37689 19211 37692
rect 19153 37683 19211 37689
rect 20714 37680 20720 37692
rect 20772 37680 20778 37732
rect 22186 37680 22192 37732
rect 22244 37720 22250 37732
rect 23198 37720 23204 37732
rect 22244 37692 23204 37720
rect 22244 37680 22250 37692
rect 23198 37680 23204 37692
rect 23256 37680 23262 37732
rect 17405 37655 17463 37661
rect 17405 37652 17417 37655
rect 15580 37624 17417 37652
rect 17405 37621 17417 37624
rect 17451 37652 17463 37655
rect 17862 37652 17868 37664
rect 17451 37624 17868 37652
rect 17451 37621 17463 37624
rect 17405 37615 17463 37621
rect 17862 37612 17868 37624
rect 17920 37612 17926 37664
rect 18690 37612 18696 37664
rect 18748 37652 18754 37664
rect 19058 37652 19064 37664
rect 18748 37624 19064 37652
rect 18748 37612 18754 37624
rect 19058 37612 19064 37624
rect 19116 37612 19122 37664
rect 20254 37612 20260 37664
rect 20312 37652 20318 37664
rect 20625 37655 20683 37661
rect 20625 37652 20637 37655
rect 20312 37624 20637 37652
rect 20312 37612 20318 37624
rect 20625 37621 20637 37624
rect 20671 37621 20683 37655
rect 20625 37615 20683 37621
rect 21910 37612 21916 37664
rect 21968 37652 21974 37664
rect 22370 37652 22376 37664
rect 21968 37624 22376 37652
rect 21968 37612 21974 37624
rect 22370 37612 22376 37624
rect 22428 37652 22434 37664
rect 23382 37652 23388 37664
rect 22428 37624 23388 37652
rect 22428 37612 22434 37624
rect 23382 37612 23388 37624
rect 23440 37612 23446 37664
rect 23934 37612 23940 37664
rect 23992 37652 23998 37664
rect 24486 37652 24492 37664
rect 23992 37624 24492 37652
rect 23992 37612 23998 37624
rect 24486 37612 24492 37624
rect 24544 37652 24550 37664
rect 25317 37655 25375 37661
rect 25317 37652 25329 37655
rect 24544 37624 25329 37652
rect 24544 37612 24550 37624
rect 25317 37621 25329 37624
rect 25363 37621 25375 37655
rect 25317 37615 25375 37621
rect 1104 37562 25852 37584
rect 1104 37510 2950 37562
rect 3002 37510 3014 37562
rect 3066 37510 3078 37562
rect 3130 37510 3142 37562
rect 3194 37510 3206 37562
rect 3258 37510 12950 37562
rect 13002 37510 13014 37562
rect 13066 37510 13078 37562
rect 13130 37510 13142 37562
rect 13194 37510 13206 37562
rect 13258 37510 22950 37562
rect 23002 37510 23014 37562
rect 23066 37510 23078 37562
rect 23130 37510 23142 37562
rect 23194 37510 23206 37562
rect 23258 37510 25852 37562
rect 1104 37488 25852 37510
rect 6181 37451 6239 37457
rect 6181 37417 6193 37451
rect 6227 37448 6239 37451
rect 6454 37448 6460 37460
rect 6227 37420 6460 37448
rect 6227 37417 6239 37420
rect 6181 37411 6239 37417
rect 6454 37408 6460 37420
rect 6512 37408 6518 37460
rect 6914 37408 6920 37460
rect 6972 37448 6978 37460
rect 6972 37420 8524 37448
rect 6972 37408 6978 37420
rect 6638 37380 6644 37392
rect 5460 37352 6644 37380
rect 4341 37315 4399 37321
rect 4341 37281 4353 37315
rect 4387 37312 4399 37315
rect 5460 37312 5488 37352
rect 6638 37340 6644 37352
rect 6696 37340 6702 37392
rect 8496 37380 8524 37420
rect 8570 37408 8576 37460
rect 8628 37448 8634 37460
rect 9306 37448 9312 37460
rect 8628 37420 9312 37448
rect 8628 37408 8634 37420
rect 9306 37408 9312 37420
rect 9364 37408 9370 37460
rect 9677 37451 9735 37457
rect 9677 37417 9689 37451
rect 9723 37448 9735 37451
rect 9723 37420 10088 37448
rect 9723 37417 9735 37420
rect 9677 37411 9735 37417
rect 9858 37380 9864 37392
rect 8496 37352 9864 37380
rect 9858 37340 9864 37352
rect 9916 37340 9922 37392
rect 9953 37383 10011 37389
rect 9953 37349 9965 37383
rect 9999 37349 10011 37383
rect 9953 37343 10011 37349
rect 4387 37284 5488 37312
rect 4387 37281 4399 37284
rect 4341 37275 4399 37281
rect 5626 37272 5632 37324
rect 5684 37312 5690 37324
rect 6546 37312 6552 37324
rect 5684 37284 6552 37312
rect 5684 37272 5690 37284
rect 6546 37272 6552 37284
rect 6604 37312 6610 37324
rect 6825 37315 6883 37321
rect 6825 37312 6837 37315
rect 6604 37284 6837 37312
rect 6604 37272 6610 37284
rect 6825 37281 6837 37284
rect 6871 37281 6883 37315
rect 6825 37275 6883 37281
rect 7101 37315 7159 37321
rect 7101 37281 7113 37315
rect 7147 37312 7159 37315
rect 8570 37312 8576 37324
rect 7147 37284 8576 37312
rect 7147 37281 7159 37284
rect 7101 37275 7159 37281
rect 8570 37272 8576 37284
rect 8628 37272 8634 37324
rect 4065 37247 4123 37253
rect 4065 37213 4077 37247
rect 4111 37213 4123 37247
rect 4065 37207 4123 37213
rect 4080 37176 4108 37207
rect 8202 37204 8208 37256
rect 8260 37204 8266 37256
rect 9968 37244 9996 37343
rect 10060 37312 10088 37420
rect 10410 37408 10416 37460
rect 10468 37448 10474 37460
rect 10962 37448 10968 37460
rect 10468 37420 10968 37448
rect 10468 37408 10474 37420
rect 10962 37408 10968 37420
rect 11020 37448 11026 37460
rect 11057 37451 11115 37457
rect 11057 37448 11069 37451
rect 11020 37420 11069 37448
rect 11020 37408 11026 37420
rect 11057 37417 11069 37420
rect 11103 37417 11115 37451
rect 11057 37411 11115 37417
rect 12250 37408 12256 37460
rect 12308 37448 12314 37460
rect 13078 37448 13084 37460
rect 12308 37420 13084 37448
rect 12308 37408 12314 37420
rect 13078 37408 13084 37420
rect 13136 37408 13142 37460
rect 13814 37408 13820 37460
rect 13872 37448 13878 37460
rect 16298 37448 16304 37460
rect 13872 37420 16304 37448
rect 13872 37408 13878 37420
rect 16298 37408 16304 37420
rect 16356 37408 16362 37460
rect 18690 37408 18696 37460
rect 18748 37408 18754 37460
rect 19242 37408 19248 37460
rect 19300 37408 19306 37460
rect 19334 37408 19340 37460
rect 19392 37408 19398 37460
rect 20898 37408 20904 37460
rect 20956 37448 20962 37460
rect 21269 37451 21327 37457
rect 21269 37448 21281 37451
rect 20956 37420 21281 37448
rect 20956 37408 20962 37420
rect 21269 37417 21281 37420
rect 21315 37448 21327 37451
rect 21634 37448 21640 37460
rect 21315 37420 21640 37448
rect 21315 37417 21327 37420
rect 21269 37411 21327 37417
rect 21634 37408 21640 37420
rect 21692 37408 21698 37460
rect 22094 37408 22100 37460
rect 22152 37448 22158 37460
rect 22741 37451 22799 37457
rect 22741 37448 22753 37451
rect 22152 37420 22753 37448
rect 22152 37408 22158 37420
rect 22741 37417 22753 37420
rect 22787 37417 22799 37451
rect 22741 37411 22799 37417
rect 23842 37408 23848 37460
rect 23900 37448 23906 37460
rect 24029 37451 24087 37457
rect 24029 37448 24041 37451
rect 23900 37420 24041 37448
rect 23900 37408 23906 37420
rect 24029 37417 24041 37420
rect 24075 37417 24087 37451
rect 24029 37411 24087 37417
rect 16482 37340 16488 37392
rect 16540 37380 16546 37392
rect 18708 37380 18736 37408
rect 19260 37380 19288 37408
rect 23658 37380 23664 37392
rect 16540 37352 16712 37380
rect 16540 37340 16546 37352
rect 10318 37312 10324 37324
rect 10060 37284 10324 37312
rect 10318 37272 10324 37284
rect 10376 37312 10382 37324
rect 10594 37312 10600 37324
rect 10376 37284 10600 37312
rect 10376 37272 10382 37284
rect 10594 37272 10600 37284
rect 10652 37272 10658 37324
rect 10962 37272 10968 37324
rect 11020 37312 11026 37324
rect 11885 37315 11943 37321
rect 11885 37312 11897 37315
rect 11020 37284 11897 37312
rect 11020 37272 11026 37284
rect 11885 37281 11897 37284
rect 11931 37281 11943 37315
rect 11885 37275 11943 37281
rect 13078 37272 13084 37324
rect 13136 37321 13142 37324
rect 13136 37315 13185 37321
rect 13136 37281 13139 37315
rect 13173 37281 13185 37315
rect 13136 37275 13185 37281
rect 13136 37272 13142 37275
rect 13354 37272 13360 37324
rect 13412 37312 13418 37324
rect 13909 37315 13967 37321
rect 13909 37312 13921 37315
rect 13412 37284 13921 37312
rect 13412 37272 13418 37284
rect 13909 37281 13921 37284
rect 13955 37312 13967 37315
rect 15473 37315 15531 37321
rect 15473 37312 15485 37315
rect 13955 37284 15485 37312
rect 13955 37281 13967 37284
rect 13909 37275 13967 37281
rect 15473 37281 15485 37284
rect 15519 37281 15531 37315
rect 15473 37275 15531 37281
rect 16390 37272 16396 37324
rect 16448 37312 16454 37324
rect 16684 37321 16712 37352
rect 17788 37352 18920 37380
rect 19260 37352 23664 37380
rect 17788 37321 17816 37352
rect 16577 37315 16635 37321
rect 16577 37312 16589 37315
rect 16448 37284 16589 37312
rect 16448 37272 16454 37284
rect 16577 37281 16589 37284
rect 16623 37281 16635 37315
rect 16577 37275 16635 37281
rect 16669 37315 16727 37321
rect 16669 37281 16681 37315
rect 16715 37281 16727 37315
rect 16669 37275 16727 37281
rect 17773 37315 17831 37321
rect 17773 37281 17785 37315
rect 17819 37281 17831 37315
rect 17773 37275 17831 37281
rect 17862 37272 17868 37324
rect 17920 37272 17926 37324
rect 11146 37244 11152 37256
rect 9968 37216 11152 37244
rect 11146 37204 11152 37216
rect 11204 37204 11210 37256
rect 11698 37204 11704 37256
rect 11756 37204 11762 37256
rect 11793 37247 11851 37253
rect 11793 37213 11805 37247
rect 11839 37244 11851 37247
rect 14182 37244 14188 37256
rect 11839 37216 14188 37244
rect 11839 37213 11851 37216
rect 11793 37207 11851 37213
rect 14182 37204 14188 37216
rect 14240 37204 14246 37256
rect 15289 37247 15347 37253
rect 15289 37213 15301 37247
rect 15335 37244 15347 37247
rect 15378 37244 15384 37256
rect 15335 37216 15384 37244
rect 15335 37213 15347 37216
rect 15289 37207 15347 37213
rect 15378 37204 15384 37216
rect 15436 37204 15442 37256
rect 17681 37247 17739 37253
rect 17681 37213 17693 37247
rect 17727 37244 17739 37247
rect 18782 37244 18788 37256
rect 17727 37216 18788 37244
rect 17727 37213 17739 37216
rect 17681 37207 17739 37213
rect 18782 37204 18788 37216
rect 18840 37204 18846 37256
rect 6454 37176 6460 37188
rect 4080 37148 4200 37176
rect 5566 37148 6460 37176
rect 4172 37108 4200 37148
rect 6454 37136 6460 37148
rect 6512 37136 6518 37188
rect 9125 37179 9183 37185
rect 9125 37145 9137 37179
rect 9171 37176 9183 37179
rect 10321 37179 10379 37185
rect 10321 37176 10333 37179
rect 9171 37148 10333 37176
rect 9171 37145 9183 37148
rect 9125 37139 9183 37145
rect 10321 37145 10333 37148
rect 10367 37145 10379 37179
rect 10321 37139 10379 37145
rect 10413 37179 10471 37185
rect 10413 37145 10425 37179
rect 10459 37176 10471 37179
rect 10502 37176 10508 37188
rect 10459 37148 10508 37176
rect 10459 37145 10471 37148
rect 10413 37139 10471 37145
rect 10502 37136 10508 37148
rect 10560 37136 10566 37188
rect 10686 37136 10692 37188
rect 10744 37176 10750 37188
rect 10744 37148 12434 37176
rect 10744 37136 10750 37148
rect 5626 37108 5632 37120
rect 4172 37080 5632 37108
rect 5626 37068 5632 37080
rect 5684 37068 5690 37120
rect 5810 37068 5816 37120
rect 5868 37068 5874 37120
rect 11146 37068 11152 37120
rect 11204 37108 11210 37120
rect 11333 37111 11391 37117
rect 11333 37108 11345 37111
rect 11204 37080 11345 37108
rect 11204 37068 11210 37080
rect 11333 37077 11345 37080
rect 11379 37077 11391 37111
rect 12406 37108 12434 37148
rect 12802 37136 12808 37188
rect 12860 37176 12866 37188
rect 12989 37179 13047 37185
rect 12989 37176 13001 37179
rect 12860 37148 13001 37176
rect 12860 37136 12866 37148
rect 12989 37145 13001 37148
rect 13035 37145 13047 37179
rect 12989 37139 13047 37145
rect 12529 37111 12587 37117
rect 12529 37108 12541 37111
rect 12406 37080 12541 37108
rect 11333 37071 11391 37077
rect 12529 37077 12541 37080
rect 12575 37077 12587 37111
rect 12529 37071 12587 37077
rect 12710 37068 12716 37120
rect 12768 37108 12774 37120
rect 12897 37111 12955 37117
rect 12897 37108 12909 37111
rect 12768 37080 12909 37108
rect 12768 37068 12774 37080
rect 12897 37077 12909 37080
rect 12943 37077 12955 37111
rect 13004 37108 13032 37139
rect 13078 37136 13084 37188
rect 13136 37176 13142 37188
rect 16485 37179 16543 37185
rect 16485 37176 16497 37179
rect 13136 37148 16497 37176
rect 13136 37136 13142 37148
rect 16485 37145 16497 37148
rect 16531 37145 16543 37179
rect 16485 37139 16543 37145
rect 17770 37136 17776 37188
rect 17828 37176 17834 37188
rect 18892 37176 18920 37352
rect 23658 37340 23664 37352
rect 23716 37340 23722 37392
rect 19150 37272 19156 37324
rect 19208 37312 19214 37324
rect 20717 37315 20775 37321
rect 20717 37312 20729 37315
rect 19208 37284 20729 37312
rect 19208 37272 19214 37284
rect 20717 37281 20729 37284
rect 20763 37281 20775 37315
rect 22189 37315 22247 37321
rect 20717 37275 20775 37281
rect 21836 37284 22048 37312
rect 19288 37204 19294 37256
rect 19346 37244 19352 37256
rect 19346 37216 20300 37244
rect 19346 37204 19352 37216
rect 18966 37176 18972 37188
rect 17828 37148 18644 37176
rect 18892 37148 18972 37176
rect 17828 37136 17834 37148
rect 13541 37111 13599 37117
rect 13541 37108 13553 37111
rect 13004 37080 13553 37108
rect 12897 37071 12955 37077
rect 13541 37077 13553 37080
rect 13587 37077 13599 37111
rect 13541 37071 13599 37077
rect 14274 37068 14280 37120
rect 14332 37068 14338 37120
rect 14458 37068 14464 37120
rect 14516 37108 14522 37120
rect 14921 37111 14979 37117
rect 14921 37108 14933 37111
rect 14516 37080 14933 37108
rect 14516 37068 14522 37080
rect 14921 37077 14933 37080
rect 14967 37077 14979 37111
rect 14921 37071 14979 37077
rect 15381 37111 15439 37117
rect 15381 37077 15393 37111
rect 15427 37108 15439 37111
rect 15930 37108 15936 37120
rect 15427 37080 15936 37108
rect 15427 37077 15439 37080
rect 15381 37071 15439 37077
rect 15930 37068 15936 37080
rect 15988 37068 15994 37120
rect 16114 37068 16120 37120
rect 16172 37068 16178 37120
rect 17310 37068 17316 37120
rect 17368 37068 17374 37120
rect 18506 37068 18512 37120
rect 18564 37068 18570 37120
rect 18616 37108 18644 37148
rect 18966 37136 18972 37148
rect 19024 37136 19030 37188
rect 20272 37176 20300 37216
rect 20530 37204 20536 37256
rect 20588 37204 20594 37256
rect 20625 37247 20683 37253
rect 20625 37213 20637 37247
rect 20671 37244 20683 37247
rect 20898 37244 20904 37256
rect 20671 37216 20904 37244
rect 20671 37213 20683 37216
rect 20625 37207 20683 37213
rect 20898 37204 20904 37216
rect 20956 37204 20962 37256
rect 21836 37244 21864 37284
rect 21376 37216 21864 37244
rect 21376 37176 21404 37216
rect 21910 37204 21916 37256
rect 21968 37204 21974 37256
rect 22020 37244 22048 37284
rect 22189 37281 22201 37315
rect 22235 37312 22247 37315
rect 22554 37312 22560 37324
rect 22235 37284 22560 37312
rect 22235 37281 22247 37284
rect 22189 37275 22247 37281
rect 22554 37272 22560 37284
rect 22612 37312 22618 37324
rect 23106 37312 23112 37324
rect 22612 37284 23112 37312
rect 22612 37272 22618 37284
rect 23106 37272 23112 37284
rect 23164 37272 23170 37324
rect 22094 37244 22100 37256
rect 22020 37216 22100 37244
rect 22094 37204 22100 37216
rect 22152 37204 22158 37256
rect 22925 37247 22983 37253
rect 22664 37216 22876 37244
rect 22664 37176 22692 37216
rect 19306 37148 20208 37176
rect 20272 37148 21404 37176
rect 21560 37148 22692 37176
rect 19306 37108 19334 37148
rect 20180 37117 20208 37148
rect 21560 37117 21588 37148
rect 18616 37080 19334 37108
rect 20165 37111 20223 37117
rect 20165 37077 20177 37111
rect 20211 37077 20223 37111
rect 20165 37071 20223 37077
rect 21545 37111 21603 37117
rect 21545 37077 21557 37111
rect 21591 37077 21603 37111
rect 21545 37071 21603 37077
rect 21818 37068 21824 37120
rect 21876 37108 21882 37120
rect 22005 37111 22063 37117
rect 22005 37108 22017 37111
rect 21876 37080 22017 37108
rect 21876 37068 21882 37080
rect 22005 37077 22017 37080
rect 22051 37108 22063 37111
rect 22646 37108 22652 37120
rect 22051 37080 22652 37108
rect 22051 37077 22063 37080
rect 22005 37071 22063 37077
rect 22646 37068 22652 37080
rect 22704 37068 22710 37120
rect 22848 37108 22876 37216
rect 22925 37213 22937 37247
rect 22971 37213 22983 37247
rect 22925 37207 22983 37213
rect 22940 37176 22968 37207
rect 23290 37204 23296 37256
rect 23348 37244 23354 37256
rect 23385 37247 23443 37253
rect 23385 37244 23397 37247
rect 23348 37216 23397 37244
rect 23348 37204 23354 37216
rect 23385 37213 23397 37216
rect 23431 37244 23443 37247
rect 24394 37244 24400 37256
rect 23431 37216 24400 37244
rect 23431 37213 23443 37216
rect 23385 37207 23443 37213
rect 24394 37204 24400 37216
rect 24452 37204 24458 37256
rect 24581 37247 24639 37253
rect 24581 37213 24593 37247
rect 24627 37244 24639 37247
rect 24946 37244 24952 37256
rect 24627 37216 24952 37244
rect 24627 37213 24639 37216
rect 24581 37207 24639 37213
rect 24946 37204 24952 37216
rect 25004 37204 25010 37256
rect 25038 37204 25044 37256
rect 25096 37244 25102 37256
rect 25225 37247 25283 37253
rect 25225 37244 25237 37247
rect 25096 37216 25237 37244
rect 25096 37204 25102 37216
rect 25225 37213 25237 37216
rect 25271 37213 25283 37247
rect 25225 37207 25283 37213
rect 24670 37176 24676 37188
rect 22940 37148 24676 37176
rect 24670 37136 24676 37148
rect 24728 37136 24734 37188
rect 23474 37108 23480 37120
rect 22848 37080 23480 37108
rect 23474 37068 23480 37080
rect 23532 37068 23538 37120
rect 23842 37068 23848 37120
rect 23900 37108 23906 37120
rect 24578 37108 24584 37120
rect 23900 37080 24584 37108
rect 23900 37068 23906 37080
rect 24578 37068 24584 37080
rect 24636 37068 24642 37120
rect 1104 37018 25852 37040
rect 1104 36966 7950 37018
rect 8002 36966 8014 37018
rect 8066 36966 8078 37018
rect 8130 36966 8142 37018
rect 8194 36966 8206 37018
rect 8258 36966 17950 37018
rect 18002 36966 18014 37018
rect 18066 36966 18078 37018
rect 18130 36966 18142 37018
rect 18194 36966 18206 37018
rect 18258 36966 25852 37018
rect 1104 36944 25852 36966
rect 6454 36864 6460 36916
rect 6512 36904 6518 36916
rect 7282 36904 7288 36916
rect 6512 36876 7288 36904
rect 6512 36864 6518 36876
rect 7282 36864 7288 36876
rect 7340 36864 7346 36916
rect 10413 36907 10471 36913
rect 10413 36904 10425 36907
rect 9140 36876 10425 36904
rect 9140 36845 9168 36876
rect 10413 36873 10425 36876
rect 10459 36904 10471 36907
rect 11054 36904 11060 36916
rect 10459 36876 11060 36904
rect 10459 36873 10471 36876
rect 10413 36867 10471 36873
rect 11054 36864 11060 36876
rect 11112 36864 11118 36916
rect 12989 36907 13047 36913
rect 12989 36873 13001 36907
rect 13035 36904 13047 36907
rect 13078 36904 13084 36916
rect 13035 36876 13084 36904
rect 13035 36873 13047 36876
rect 12989 36867 13047 36873
rect 13078 36864 13084 36876
rect 13136 36864 13142 36916
rect 13357 36907 13415 36913
rect 13357 36873 13369 36907
rect 13403 36904 13415 36907
rect 14274 36904 14280 36916
rect 13403 36876 14280 36904
rect 13403 36873 13415 36876
rect 13357 36867 13415 36873
rect 14274 36864 14280 36876
rect 14332 36864 14338 36916
rect 14918 36864 14924 36916
rect 14976 36864 14982 36916
rect 17037 36907 17095 36913
rect 17037 36873 17049 36907
rect 17083 36904 17095 36907
rect 17126 36904 17132 36916
rect 17083 36876 17132 36904
rect 17083 36873 17095 36876
rect 17037 36867 17095 36873
rect 17126 36864 17132 36876
rect 17184 36864 17190 36916
rect 17405 36907 17463 36913
rect 17405 36873 17417 36907
rect 17451 36904 17463 36907
rect 18506 36904 18512 36916
rect 17451 36876 18512 36904
rect 17451 36873 17463 36876
rect 17405 36867 17463 36873
rect 18506 36864 18512 36876
rect 18564 36864 18570 36916
rect 18690 36864 18696 36916
rect 18748 36904 18754 36916
rect 19981 36907 20039 36913
rect 18748 36876 19932 36904
rect 18748 36864 18754 36876
rect 9125 36839 9183 36845
rect 9125 36805 9137 36839
rect 9171 36805 9183 36839
rect 9125 36799 9183 36805
rect 10778 36796 10784 36848
rect 10836 36836 10842 36848
rect 11517 36839 11575 36845
rect 11517 36836 11529 36839
rect 10836 36808 11529 36836
rect 10836 36796 10842 36808
rect 11517 36805 11529 36808
rect 11563 36836 11575 36839
rect 13449 36839 13507 36845
rect 13449 36836 13461 36839
rect 11563 36808 13461 36836
rect 11563 36805 11575 36808
rect 11517 36799 11575 36805
rect 13449 36805 13461 36808
rect 13495 36805 13507 36839
rect 13449 36799 13507 36805
rect 13556 36808 15148 36836
rect 11885 36771 11943 36777
rect 11885 36737 11897 36771
rect 11931 36737 11943 36771
rect 11885 36731 11943 36737
rect 9674 36660 9680 36712
rect 9732 36700 9738 36712
rect 9861 36703 9919 36709
rect 9861 36700 9873 36703
rect 9732 36672 9873 36700
rect 9732 36660 9738 36672
rect 9861 36669 9873 36672
rect 9907 36669 9919 36703
rect 11900 36700 11928 36731
rect 12434 36728 12440 36780
rect 12492 36768 12498 36780
rect 13354 36768 13360 36780
rect 12492 36740 13360 36768
rect 12492 36728 12498 36740
rect 13354 36728 13360 36740
rect 13412 36728 13418 36780
rect 12802 36700 12808 36712
rect 11900 36672 12808 36700
rect 9861 36663 9919 36669
rect 12802 36660 12808 36672
rect 12860 36700 12866 36712
rect 13262 36700 13268 36712
rect 12860 36672 13268 36700
rect 12860 36660 12866 36672
rect 13262 36660 13268 36672
rect 13320 36700 13326 36712
rect 13556 36700 13584 36808
rect 14090 36728 14096 36780
rect 14148 36768 14154 36780
rect 14826 36768 14832 36780
rect 14148 36740 14832 36768
rect 14148 36728 14154 36740
rect 14826 36728 14832 36740
rect 14884 36728 14890 36780
rect 13320 36672 13584 36700
rect 13633 36703 13691 36709
rect 13320 36660 13326 36672
rect 13633 36669 13645 36703
rect 13679 36700 13691 36703
rect 13814 36700 13820 36712
rect 13679 36672 13820 36700
rect 13679 36669 13691 36672
rect 13633 36663 13691 36669
rect 13814 36660 13820 36672
rect 13872 36660 13878 36712
rect 15120 36709 15148 36808
rect 17218 36796 17224 36848
rect 17276 36836 17282 36848
rect 19150 36836 19156 36848
rect 17276 36808 19156 36836
rect 17276 36796 17282 36808
rect 19150 36796 19156 36808
rect 19208 36796 19214 36848
rect 19904 36836 19932 36876
rect 19981 36873 19993 36907
rect 20027 36904 20039 36907
rect 20622 36904 20628 36916
rect 20027 36876 20628 36904
rect 20027 36873 20039 36876
rect 19981 36867 20039 36873
rect 20622 36864 20628 36876
rect 20680 36864 20686 36916
rect 21634 36904 21640 36916
rect 20732 36876 21640 36904
rect 20732 36836 20760 36876
rect 21634 36864 21640 36876
rect 21692 36904 21698 36916
rect 22189 36907 22247 36913
rect 22189 36904 22201 36907
rect 21692 36876 22201 36904
rect 21692 36864 21698 36876
rect 22189 36873 22201 36876
rect 22235 36873 22247 36907
rect 22189 36867 22247 36873
rect 22554 36864 22560 36916
rect 22612 36904 22618 36916
rect 23198 36904 23204 36916
rect 22612 36876 23204 36904
rect 22612 36864 22618 36876
rect 23198 36864 23204 36876
rect 23256 36864 23262 36916
rect 24394 36864 24400 36916
rect 24452 36904 24458 36916
rect 24581 36907 24639 36913
rect 24581 36904 24593 36907
rect 24452 36876 24593 36904
rect 24452 36864 24458 36876
rect 24581 36873 24593 36876
rect 24627 36873 24639 36907
rect 24854 36904 24860 36916
rect 24581 36867 24639 36873
rect 24688 36876 24860 36904
rect 19904 36808 20760 36836
rect 21913 36839 21971 36845
rect 21913 36805 21925 36839
rect 21959 36836 21971 36839
rect 23382 36836 23388 36848
rect 21959 36808 23388 36836
rect 21959 36805 21971 36808
rect 21913 36799 21971 36805
rect 16666 36728 16672 36780
rect 16724 36768 16730 36780
rect 17497 36771 17555 36777
rect 17497 36768 17509 36771
rect 16724 36740 17509 36768
rect 16724 36728 16730 36740
rect 17497 36737 17509 36740
rect 17543 36737 17555 36771
rect 17497 36731 17555 36737
rect 18233 36771 18291 36777
rect 18233 36737 18245 36771
rect 18279 36768 18291 36771
rect 18598 36768 18604 36780
rect 18279 36740 18604 36768
rect 18279 36737 18291 36740
rect 18233 36731 18291 36737
rect 18598 36728 18604 36740
rect 18656 36728 18662 36780
rect 18782 36728 18788 36780
rect 18840 36768 18846 36780
rect 19242 36768 19248 36780
rect 18840 36740 19248 36768
rect 18840 36728 18846 36740
rect 19242 36728 19248 36740
rect 19300 36728 19306 36780
rect 19610 36728 19616 36780
rect 19668 36768 19674 36780
rect 20349 36771 20407 36777
rect 20349 36768 20361 36771
rect 19668 36740 20361 36768
rect 19668 36728 19674 36740
rect 20349 36737 20361 36740
rect 20395 36737 20407 36771
rect 20349 36731 20407 36737
rect 20438 36728 20444 36780
rect 20496 36768 20502 36780
rect 21082 36768 21088 36780
rect 20496 36740 21088 36768
rect 20496 36728 20502 36740
rect 21082 36728 21088 36740
rect 21140 36728 21146 36780
rect 22388 36777 22416 36808
rect 23382 36796 23388 36808
rect 23440 36796 23446 36848
rect 24688 36836 24716 36876
rect 24854 36864 24860 36876
rect 24912 36864 24918 36916
rect 24412 36808 24716 36836
rect 24412 36780 24440 36808
rect 22373 36771 22431 36777
rect 22373 36737 22385 36771
rect 22419 36737 22431 36771
rect 24394 36768 24400 36780
rect 24242 36740 24400 36768
rect 22373 36731 22431 36737
rect 24394 36728 24400 36740
rect 24452 36728 24458 36780
rect 24854 36728 24860 36780
rect 24912 36768 24918 36780
rect 25317 36771 25375 36777
rect 25317 36768 25329 36771
rect 24912 36740 25329 36768
rect 24912 36728 24918 36740
rect 25317 36737 25329 36740
rect 25363 36737 25375 36771
rect 25317 36731 25375 36737
rect 15105 36703 15163 36709
rect 15105 36669 15117 36703
rect 15151 36669 15163 36703
rect 15105 36663 15163 36669
rect 17681 36703 17739 36709
rect 17681 36669 17693 36703
rect 17727 36700 17739 36703
rect 19794 36700 19800 36712
rect 17727 36672 19800 36700
rect 17727 36669 17739 36672
rect 17681 36663 17739 36669
rect 19794 36660 19800 36672
rect 19852 36660 19858 36712
rect 20625 36703 20683 36709
rect 20625 36669 20637 36703
rect 20671 36700 20683 36703
rect 21726 36700 21732 36712
rect 20671 36672 21732 36700
rect 20671 36669 20683 36672
rect 20625 36663 20683 36669
rect 21726 36660 21732 36672
rect 21784 36700 21790 36712
rect 22646 36700 22652 36712
rect 21784 36672 22652 36700
rect 21784 36660 21790 36672
rect 22646 36660 22652 36672
rect 22704 36660 22710 36712
rect 22830 36660 22836 36712
rect 22888 36660 22894 36712
rect 23106 36660 23112 36712
rect 23164 36700 23170 36712
rect 23474 36700 23480 36712
rect 23164 36672 23480 36700
rect 23164 36660 23170 36672
rect 23474 36660 23480 36672
rect 23532 36660 23538 36712
rect 11238 36592 11244 36644
rect 11296 36632 11302 36644
rect 17310 36632 17316 36644
rect 11296 36604 17316 36632
rect 11296 36592 11302 36604
rect 17310 36592 17316 36604
rect 17368 36592 17374 36644
rect 19978 36632 19984 36644
rect 18248 36604 19984 36632
rect 7190 36524 7196 36576
rect 7248 36524 7254 36576
rect 8570 36524 8576 36576
rect 8628 36564 8634 36576
rect 8665 36567 8723 36573
rect 8665 36564 8677 36567
rect 8628 36536 8677 36564
rect 8628 36524 8634 36536
rect 8665 36533 8677 36536
rect 8711 36564 8723 36567
rect 9490 36564 9496 36576
rect 8711 36536 9496 36564
rect 8711 36533 8723 36536
rect 8665 36527 8723 36533
rect 9490 36524 9496 36536
rect 9548 36524 9554 36576
rect 12434 36524 12440 36576
rect 12492 36564 12498 36576
rect 12529 36567 12587 36573
rect 12529 36564 12541 36567
rect 12492 36536 12541 36564
rect 12492 36524 12498 36536
rect 12529 36533 12541 36536
rect 12575 36533 12587 36567
rect 12529 36527 12587 36533
rect 14185 36567 14243 36573
rect 14185 36533 14197 36567
rect 14231 36564 14243 36567
rect 14366 36564 14372 36576
rect 14231 36536 14372 36564
rect 14231 36533 14243 36536
rect 14185 36527 14243 36533
rect 14366 36524 14372 36536
rect 14424 36524 14430 36576
rect 14458 36524 14464 36576
rect 14516 36524 14522 36576
rect 14826 36524 14832 36576
rect 14884 36564 14890 36576
rect 15473 36567 15531 36573
rect 15473 36564 15485 36567
rect 14884 36536 15485 36564
rect 14884 36524 14890 36536
rect 15473 36533 15485 36536
rect 15519 36564 15531 36567
rect 18248 36564 18276 36604
rect 19978 36592 19984 36604
rect 20036 36592 20042 36644
rect 25133 36635 25191 36641
rect 25133 36632 25145 36635
rect 20456 36604 22968 36632
rect 20456 36576 20484 36604
rect 15519 36536 18276 36564
rect 15519 36533 15531 36536
rect 15473 36527 15531 36533
rect 18322 36524 18328 36576
rect 18380 36564 18386 36576
rect 18877 36567 18935 36573
rect 18877 36564 18889 36567
rect 18380 36536 18889 36564
rect 18380 36524 18386 36536
rect 18877 36533 18889 36536
rect 18923 36533 18935 36567
rect 18877 36527 18935 36533
rect 19610 36524 19616 36576
rect 19668 36524 19674 36576
rect 20438 36524 20444 36576
rect 20496 36524 20502 36576
rect 21082 36524 21088 36576
rect 21140 36524 21146 36576
rect 22940 36564 22968 36604
rect 24136 36604 25145 36632
rect 24136 36564 24164 36604
rect 25133 36601 25145 36604
rect 25179 36601 25191 36635
rect 25133 36595 25191 36601
rect 22940 36536 24164 36564
rect 1104 36474 25852 36496
rect 1104 36422 2950 36474
rect 3002 36422 3014 36474
rect 3066 36422 3078 36474
rect 3130 36422 3142 36474
rect 3194 36422 3206 36474
rect 3258 36422 12950 36474
rect 13002 36422 13014 36474
rect 13066 36422 13078 36474
rect 13130 36422 13142 36474
rect 13194 36422 13206 36474
rect 13258 36422 22950 36474
rect 23002 36422 23014 36474
rect 23066 36422 23078 36474
rect 23130 36422 23142 36474
rect 23194 36422 23206 36474
rect 23258 36422 25852 36474
rect 1104 36400 25852 36422
rect 7006 36320 7012 36372
rect 7064 36320 7070 36372
rect 7282 36320 7288 36372
rect 7340 36320 7346 36372
rect 7650 36320 7656 36372
rect 7708 36360 7714 36372
rect 7745 36363 7803 36369
rect 7745 36360 7757 36363
rect 7708 36332 7757 36360
rect 7708 36320 7714 36332
rect 7745 36329 7757 36332
rect 7791 36329 7803 36363
rect 7745 36323 7803 36329
rect 8938 36320 8944 36372
rect 8996 36360 9002 36372
rect 9125 36363 9183 36369
rect 9125 36360 9137 36363
rect 8996 36332 9137 36360
rect 8996 36320 9002 36332
rect 9125 36329 9137 36332
rect 9171 36329 9183 36363
rect 9125 36323 9183 36329
rect 9950 36320 9956 36372
rect 10008 36360 10014 36372
rect 10318 36360 10324 36372
rect 10008 36332 10324 36360
rect 10008 36320 10014 36332
rect 10318 36320 10324 36332
rect 10376 36360 10382 36372
rect 10781 36363 10839 36369
rect 10781 36360 10793 36363
rect 10376 36332 10793 36360
rect 10376 36320 10382 36332
rect 10781 36329 10793 36332
rect 10827 36329 10839 36363
rect 10781 36323 10839 36329
rect 10796 36292 10824 36323
rect 11054 36320 11060 36372
rect 11112 36320 11118 36372
rect 11238 36320 11244 36372
rect 11296 36360 11302 36372
rect 12897 36363 12955 36369
rect 11296 36332 12848 36360
rect 11296 36320 11302 36332
rect 10796 36264 12756 36292
rect 5261 36227 5319 36233
rect 5261 36193 5273 36227
rect 5307 36224 5319 36227
rect 5626 36224 5632 36236
rect 5307 36196 5632 36224
rect 5307 36193 5319 36196
rect 5261 36187 5319 36193
rect 5626 36184 5632 36196
rect 5684 36184 5690 36236
rect 7650 36184 7656 36236
rect 7708 36224 7714 36236
rect 8297 36227 8355 36233
rect 8297 36224 8309 36227
rect 7708 36196 8309 36224
rect 7708 36184 7714 36196
rect 8297 36193 8309 36196
rect 8343 36193 8355 36227
rect 8297 36187 8355 36193
rect 8754 36184 8760 36236
rect 8812 36224 8818 36236
rect 9677 36227 9735 36233
rect 9677 36224 9689 36227
rect 8812 36196 9689 36224
rect 8812 36184 8818 36196
rect 9677 36193 9689 36196
rect 9723 36193 9735 36227
rect 12526 36224 12532 36236
rect 9677 36187 9735 36193
rect 10980 36196 12532 36224
rect 1762 36116 1768 36168
rect 1820 36156 1826 36168
rect 2041 36159 2099 36165
rect 2041 36156 2053 36159
rect 1820 36128 2053 36156
rect 1820 36116 1826 36128
rect 2041 36125 2053 36128
rect 2087 36125 2099 36159
rect 2041 36119 2099 36125
rect 9585 36159 9643 36165
rect 9585 36125 9597 36159
rect 9631 36156 9643 36159
rect 10980 36156 11008 36196
rect 12526 36184 12532 36196
rect 12584 36184 12590 36236
rect 9631 36128 11008 36156
rect 9631 36125 9643 36128
rect 9585 36119 9643 36125
rect 11054 36116 11060 36168
rect 11112 36156 11118 36168
rect 11517 36159 11575 36165
rect 11517 36156 11529 36159
rect 11112 36128 11529 36156
rect 11112 36116 11118 36128
rect 11517 36125 11529 36128
rect 11563 36125 11575 36159
rect 11517 36119 11575 36125
rect 5537 36091 5595 36097
rect 5537 36057 5549 36091
rect 5583 36057 5595 36091
rect 6822 36088 6828 36100
rect 6762 36060 6828 36088
rect 5537 36051 5595 36057
rect 1578 35980 1584 36032
rect 1636 35980 1642 36032
rect 5552 36020 5580 36051
rect 6822 36048 6828 36060
rect 6880 36088 6886 36100
rect 7282 36088 7288 36100
rect 6880 36060 7288 36088
rect 6880 36048 6886 36060
rect 7282 36048 7288 36060
rect 7340 36048 7346 36100
rect 8205 36091 8263 36097
rect 8205 36057 8217 36091
rect 8251 36088 8263 36091
rect 9493 36091 9551 36097
rect 8251 36060 9444 36088
rect 8251 36057 8263 36060
rect 8205 36051 8263 36057
rect 7190 36020 7196 36032
rect 5552 35992 7196 36020
rect 7190 35980 7196 35992
rect 7248 35980 7254 36032
rect 7558 35980 7564 36032
rect 7616 36020 7622 36032
rect 8113 36023 8171 36029
rect 8113 36020 8125 36023
rect 7616 35992 8125 36020
rect 7616 35980 7622 35992
rect 8113 35989 8125 35992
rect 8159 35989 8171 36023
rect 9416 36020 9444 36060
rect 9493 36057 9505 36091
rect 9539 36088 9551 36091
rect 9539 36060 11284 36088
rect 9539 36057 9551 36060
rect 9493 36051 9551 36057
rect 10226 36020 10232 36032
rect 9416 35992 10232 36020
rect 8113 35983 8171 35989
rect 10226 35980 10232 35992
rect 10284 35980 10290 36032
rect 11256 36020 11284 36060
rect 11698 36048 11704 36100
rect 11756 36088 11762 36100
rect 12253 36091 12311 36097
rect 12253 36088 12265 36091
rect 11756 36060 12265 36088
rect 11756 36048 11762 36060
rect 12253 36057 12265 36060
rect 12299 36057 12311 36091
rect 12253 36051 12311 36057
rect 12618 36020 12624 36032
rect 11256 35992 12624 36020
rect 12618 35980 12624 35992
rect 12676 35980 12682 36032
rect 12728 36020 12756 36264
rect 12820 36088 12848 36332
rect 12897 36329 12909 36363
rect 12943 36360 12955 36363
rect 13446 36360 13452 36372
rect 12943 36332 13452 36360
rect 12943 36329 12955 36332
rect 12897 36323 12955 36329
rect 13446 36320 13452 36332
rect 13504 36320 13510 36372
rect 14277 36363 14335 36369
rect 14277 36329 14289 36363
rect 14323 36360 14335 36363
rect 15194 36360 15200 36372
rect 14323 36332 15200 36360
rect 14323 36329 14335 36332
rect 14277 36323 14335 36329
rect 15194 36320 15200 36332
rect 15252 36320 15258 36372
rect 16206 36320 16212 36372
rect 16264 36320 16270 36372
rect 17034 36320 17040 36372
rect 17092 36360 17098 36372
rect 17586 36360 17592 36372
rect 17092 36332 17592 36360
rect 17092 36320 17098 36332
rect 17586 36320 17592 36332
rect 17644 36320 17650 36372
rect 22646 36320 22652 36372
rect 22704 36360 22710 36372
rect 25038 36360 25044 36372
rect 22704 36332 25044 36360
rect 22704 36320 22710 36332
rect 25038 36320 25044 36332
rect 25096 36320 25102 36372
rect 15010 36252 15016 36304
rect 15068 36292 15074 36304
rect 19429 36295 19487 36301
rect 19429 36292 19441 36295
rect 15068 36264 19441 36292
rect 15068 36252 15074 36264
rect 19429 36261 19441 36264
rect 19475 36261 19487 36295
rect 23293 36295 23351 36301
rect 19429 36255 19487 36261
rect 19904 36264 22094 36292
rect 13354 36184 13360 36236
rect 13412 36224 13418 36236
rect 13449 36227 13507 36233
rect 13449 36224 13461 36227
rect 13412 36196 13461 36224
rect 13412 36184 13418 36196
rect 13449 36193 13461 36196
rect 13495 36193 13507 36227
rect 13449 36187 13507 36193
rect 14921 36227 14979 36233
rect 14921 36193 14933 36227
rect 14967 36224 14979 36227
rect 15562 36224 15568 36236
rect 14967 36196 15568 36224
rect 14967 36193 14979 36196
rect 14921 36187 14979 36193
rect 15562 36184 15568 36196
rect 15620 36184 15626 36236
rect 16853 36227 16911 36233
rect 16853 36193 16865 36227
rect 16899 36224 16911 36227
rect 16942 36224 16948 36236
rect 16899 36196 16948 36224
rect 16899 36193 16911 36196
rect 16853 36187 16911 36193
rect 16942 36184 16948 36196
rect 17000 36184 17006 36236
rect 19904 36233 19932 36264
rect 19889 36227 19947 36233
rect 19889 36193 19901 36227
rect 19935 36193 19947 36227
rect 19889 36187 19947 36193
rect 19981 36227 20039 36233
rect 19981 36193 19993 36227
rect 20027 36193 20039 36227
rect 19981 36187 20039 36193
rect 15654 36116 15660 36168
rect 15712 36156 15718 36168
rect 19061 36159 19119 36165
rect 19061 36156 19073 36159
rect 15712 36128 19073 36156
rect 15712 36116 15718 36128
rect 19061 36125 19073 36128
rect 19107 36156 19119 36159
rect 19996 36156 20024 36187
rect 21358 36184 21364 36236
rect 21416 36184 21422 36236
rect 21453 36227 21511 36233
rect 21453 36193 21465 36227
rect 21499 36193 21511 36227
rect 21453 36187 21511 36193
rect 19107 36128 20024 36156
rect 19107 36125 19119 36128
rect 19061 36119 19119 36125
rect 21266 36116 21272 36168
rect 21324 36156 21330 36168
rect 21468 36156 21496 36187
rect 21324 36128 21496 36156
rect 21324 36116 21330 36128
rect 22066 36100 22094 36264
rect 23293 36261 23305 36295
rect 23339 36292 23351 36295
rect 24486 36292 24492 36304
rect 23339 36264 24492 36292
rect 23339 36261 23351 36264
rect 23293 36255 23351 36261
rect 24486 36252 24492 36264
rect 24544 36252 24550 36304
rect 23934 36184 23940 36236
rect 23992 36184 23998 36236
rect 25498 36224 25504 36236
rect 24044 36196 25504 36224
rect 23753 36159 23811 36165
rect 23753 36125 23765 36159
rect 23799 36156 23811 36159
rect 23842 36156 23848 36168
rect 23799 36128 23848 36156
rect 23799 36125 23811 36128
rect 23753 36119 23811 36125
rect 23842 36116 23848 36128
rect 23900 36116 23906 36168
rect 14645 36091 14703 36097
rect 12820 36060 13400 36088
rect 13372 36029 13400 36060
rect 14645 36057 14657 36091
rect 14691 36088 14703 36091
rect 15473 36091 15531 36097
rect 15473 36088 15485 36091
rect 14691 36060 15485 36088
rect 14691 36057 14703 36060
rect 14645 36051 14703 36057
rect 15473 36057 15485 36060
rect 15519 36057 15531 36091
rect 15473 36051 15531 36057
rect 16577 36091 16635 36097
rect 16577 36057 16589 36091
rect 16623 36088 16635 36091
rect 17405 36091 17463 36097
rect 17405 36088 17417 36091
rect 16623 36060 17417 36088
rect 16623 36057 16635 36060
rect 16577 36051 16635 36057
rect 17405 36057 17417 36060
rect 17451 36057 17463 36091
rect 17405 36051 17463 36057
rect 19797 36091 19855 36097
rect 19797 36057 19809 36091
rect 19843 36088 19855 36091
rect 21174 36088 21180 36100
rect 19843 36060 21180 36088
rect 19843 36057 19855 36060
rect 19797 36051 19855 36057
rect 21174 36048 21180 36060
rect 21232 36048 21238 36100
rect 22066 36060 22100 36100
rect 22094 36048 22100 36060
rect 22152 36088 22158 36100
rect 24044 36088 24072 36196
rect 25498 36184 25504 36196
rect 25556 36184 25562 36236
rect 24670 36116 24676 36168
rect 24728 36156 24734 36168
rect 25317 36159 25375 36165
rect 25317 36156 25329 36159
rect 24728 36128 25329 36156
rect 24728 36116 24734 36128
rect 25317 36125 25329 36128
rect 25363 36125 25375 36159
rect 25317 36119 25375 36125
rect 22152 36060 24072 36088
rect 22152 36048 22158 36060
rect 13265 36023 13323 36029
rect 13265 36020 13277 36023
rect 12728 35992 13277 36020
rect 13265 35989 13277 35992
rect 13311 35989 13323 36023
rect 13265 35983 13323 35989
rect 13357 36023 13415 36029
rect 13357 35989 13369 36023
rect 13403 36020 13415 36023
rect 13814 36020 13820 36032
rect 13403 35992 13820 36020
rect 13403 35989 13415 35992
rect 13357 35983 13415 35989
rect 13814 35980 13820 35992
rect 13872 35980 13878 36032
rect 14366 35980 14372 36032
rect 14424 36020 14430 36032
rect 14737 36023 14795 36029
rect 14737 36020 14749 36023
rect 14424 35992 14749 36020
rect 14424 35980 14430 35992
rect 14737 35989 14749 35992
rect 14783 35989 14795 36023
rect 14737 35983 14795 35989
rect 16666 35980 16672 36032
rect 16724 35980 16730 36032
rect 19978 35980 19984 36032
rect 20036 36020 20042 36032
rect 20901 36023 20959 36029
rect 20901 36020 20913 36023
rect 20036 35992 20913 36020
rect 20036 35980 20042 35992
rect 20901 35989 20913 35992
rect 20947 35989 20959 36023
rect 20901 35983 20959 35989
rect 20990 35980 20996 36032
rect 21048 36020 21054 36032
rect 21269 36023 21327 36029
rect 21269 36020 21281 36023
rect 21048 35992 21281 36020
rect 21048 35980 21054 35992
rect 21269 35989 21281 35992
rect 21315 35989 21327 36023
rect 21269 35983 21327 35989
rect 22646 35980 22652 36032
rect 22704 35980 22710 36032
rect 23658 35980 23664 36032
rect 23716 35980 23722 36032
rect 24394 35980 24400 36032
rect 24452 35980 24458 36032
rect 24670 35980 24676 36032
rect 24728 35980 24734 36032
rect 24854 35980 24860 36032
rect 24912 35980 24918 36032
rect 25130 35980 25136 36032
rect 25188 35980 25194 36032
rect 1104 35930 25852 35952
rect 1104 35878 7950 35930
rect 8002 35878 8014 35930
rect 8066 35878 8078 35930
rect 8130 35878 8142 35930
rect 8194 35878 8206 35930
rect 8258 35878 17950 35930
rect 18002 35878 18014 35930
rect 18066 35878 18078 35930
rect 18130 35878 18142 35930
rect 18194 35878 18206 35930
rect 18258 35878 25852 35930
rect 1104 35856 25852 35878
rect 5997 35819 6055 35825
rect 5997 35785 6009 35819
rect 6043 35816 6055 35819
rect 6086 35816 6092 35828
rect 6043 35788 6092 35816
rect 6043 35785 6055 35788
rect 5997 35779 6055 35785
rect 6086 35776 6092 35788
rect 6144 35776 6150 35828
rect 6457 35819 6515 35825
rect 6457 35785 6469 35819
rect 6503 35816 6515 35819
rect 6822 35816 6828 35828
rect 6503 35788 6828 35816
rect 6503 35785 6515 35788
rect 6457 35779 6515 35785
rect 6472 35748 6500 35779
rect 6822 35776 6828 35788
rect 6880 35776 6886 35828
rect 9861 35819 9919 35825
rect 9861 35816 9873 35819
rect 7024 35788 9873 35816
rect 5750 35720 6500 35748
rect 7024 35689 7052 35788
rect 9861 35785 9873 35788
rect 9907 35816 9919 35819
rect 13354 35816 13360 35828
rect 9907 35788 13360 35816
rect 9907 35785 9919 35788
rect 9861 35779 9919 35785
rect 13354 35776 13360 35788
rect 13412 35816 13418 35828
rect 13630 35816 13636 35828
rect 13412 35788 13636 35816
rect 13412 35776 13418 35788
rect 13630 35776 13636 35788
rect 13688 35776 13694 35828
rect 13906 35776 13912 35828
rect 13964 35816 13970 35828
rect 14093 35819 14151 35825
rect 14093 35816 14105 35819
rect 13964 35788 14105 35816
rect 13964 35776 13970 35788
rect 14093 35785 14105 35788
rect 14139 35816 14151 35819
rect 14921 35819 14979 35825
rect 14921 35816 14933 35819
rect 14139 35788 14933 35816
rect 14139 35785 14151 35788
rect 14093 35779 14151 35785
rect 14921 35785 14933 35788
rect 14967 35785 14979 35819
rect 14921 35779 14979 35785
rect 15930 35776 15936 35828
rect 15988 35816 15994 35828
rect 15988 35788 19334 35816
rect 15988 35776 15994 35788
rect 7282 35708 7288 35760
rect 7340 35748 7346 35760
rect 8110 35748 8116 35760
rect 7340 35720 8116 35748
rect 7340 35708 7346 35720
rect 8110 35708 8116 35720
rect 8168 35748 8174 35760
rect 13446 35748 13452 35760
rect 8168 35720 8878 35748
rect 13202 35720 13452 35748
rect 8168 35708 8174 35720
rect 13446 35708 13452 35720
rect 13504 35748 13510 35760
rect 13817 35751 13875 35757
rect 13817 35748 13829 35751
rect 13504 35720 13829 35748
rect 13504 35708 13510 35720
rect 13817 35717 13829 35720
rect 13863 35748 13875 35751
rect 13998 35748 14004 35760
rect 13863 35720 14004 35748
rect 13863 35717 13875 35720
rect 13817 35711 13875 35717
rect 13998 35708 14004 35720
rect 14056 35708 14062 35760
rect 18046 35748 18052 35760
rect 17696 35720 18052 35748
rect 4249 35683 4307 35689
rect 4249 35649 4261 35683
rect 4295 35649 4307 35683
rect 4249 35643 4307 35649
rect 7009 35683 7067 35689
rect 7009 35649 7021 35683
rect 7055 35649 7067 35683
rect 7009 35643 7067 35649
rect 4264 35612 4292 35643
rect 11698 35640 11704 35692
rect 11756 35640 11762 35692
rect 14829 35683 14887 35689
rect 14829 35649 14841 35683
rect 14875 35649 14887 35683
rect 14829 35643 14887 35649
rect 4525 35615 4583 35621
rect 4264 35584 4384 35612
rect 4356 35476 4384 35584
rect 4525 35581 4537 35615
rect 4571 35612 4583 35615
rect 8113 35615 8171 35621
rect 4571 35584 7052 35612
rect 4571 35581 4583 35584
rect 4525 35575 4583 35581
rect 7024 35556 7052 35584
rect 8113 35581 8125 35615
rect 8159 35581 8171 35615
rect 8113 35575 8171 35581
rect 8389 35615 8447 35621
rect 8389 35581 8401 35615
rect 8435 35612 8447 35615
rect 9766 35612 9772 35624
rect 8435 35584 9772 35612
rect 8435 35581 8447 35584
rect 8389 35575 8447 35581
rect 7006 35504 7012 35556
rect 7064 35504 7070 35556
rect 5626 35476 5632 35488
rect 4356 35448 5632 35476
rect 5626 35436 5632 35448
rect 5684 35436 5690 35488
rect 6546 35436 6552 35488
rect 6604 35476 6610 35488
rect 7653 35479 7711 35485
rect 7653 35476 7665 35479
rect 6604 35448 7665 35476
rect 6604 35436 6610 35448
rect 7653 35445 7665 35448
rect 7699 35445 7711 35479
rect 8128 35476 8156 35575
rect 9766 35572 9772 35584
rect 9824 35572 9830 35624
rect 11977 35615 12035 35621
rect 11977 35581 11989 35615
rect 12023 35612 12035 35615
rect 14734 35612 14740 35624
rect 12023 35584 14740 35612
rect 12023 35581 12035 35584
rect 11977 35575 12035 35581
rect 14734 35572 14740 35584
rect 14792 35572 14798 35624
rect 13449 35547 13507 35553
rect 13449 35513 13461 35547
rect 13495 35544 13507 35547
rect 13630 35544 13636 35556
rect 13495 35516 13636 35544
rect 13495 35513 13507 35516
rect 13449 35507 13507 35513
rect 8386 35476 8392 35488
rect 8128 35448 8392 35476
rect 7653 35439 7711 35445
rect 8386 35436 8392 35448
rect 8444 35436 8450 35488
rect 9858 35436 9864 35488
rect 9916 35476 9922 35488
rect 10137 35479 10195 35485
rect 10137 35476 10149 35479
rect 9916 35448 10149 35476
rect 9916 35436 9922 35448
rect 10137 35445 10149 35448
rect 10183 35476 10195 35479
rect 12342 35476 12348 35488
rect 10183 35448 12348 35476
rect 10183 35445 10195 35448
rect 10137 35439 10195 35445
rect 12342 35436 12348 35448
rect 12400 35436 12406 35488
rect 12526 35436 12532 35488
rect 12584 35476 12590 35488
rect 13464 35476 13492 35507
rect 13630 35504 13636 35516
rect 13688 35504 13694 35556
rect 14844 35544 14872 35643
rect 15470 35640 15476 35692
rect 15528 35680 15534 35692
rect 16482 35680 16488 35692
rect 15528 35652 16488 35680
rect 15528 35640 15534 35652
rect 16482 35640 16488 35652
rect 16540 35680 16546 35692
rect 17696 35689 17724 35720
rect 18046 35708 18052 35720
rect 18104 35708 18110 35760
rect 18690 35708 18696 35760
rect 18748 35708 18754 35760
rect 19306 35748 19334 35788
rect 20346 35776 20352 35828
rect 20404 35776 20410 35828
rect 22373 35819 22431 35825
rect 22373 35785 22385 35819
rect 22419 35816 22431 35819
rect 22646 35816 22652 35828
rect 22419 35788 22652 35816
rect 22419 35785 22431 35788
rect 22373 35779 22431 35785
rect 22646 35776 22652 35788
rect 22704 35776 22710 35828
rect 22922 35776 22928 35828
rect 22980 35816 22986 35828
rect 23474 35816 23480 35828
rect 22980 35788 23480 35816
rect 22980 35776 22986 35788
rect 23474 35776 23480 35788
rect 23532 35816 23538 35828
rect 24949 35819 25007 35825
rect 24949 35816 24961 35819
rect 23532 35788 24961 35816
rect 23532 35776 23538 35788
rect 24949 35785 24961 35788
rect 24995 35785 25007 35819
rect 24949 35779 25007 35785
rect 20257 35751 20315 35757
rect 20257 35748 20269 35751
rect 19306 35720 20269 35748
rect 20257 35717 20269 35720
rect 20303 35748 20315 35751
rect 21910 35748 21916 35760
rect 20303 35720 21916 35748
rect 20303 35717 20315 35720
rect 20257 35711 20315 35717
rect 21910 35708 21916 35720
rect 21968 35708 21974 35760
rect 22830 35708 22836 35760
rect 22888 35748 22894 35760
rect 23382 35748 23388 35760
rect 22888 35720 23388 35748
rect 22888 35708 22894 35720
rect 23216 35689 23244 35720
rect 23382 35708 23388 35720
rect 23440 35708 23446 35760
rect 25406 35748 25412 35760
rect 24702 35720 25412 35748
rect 25406 35708 25412 35720
rect 25464 35708 25470 35760
rect 17681 35683 17739 35689
rect 17681 35680 17693 35683
rect 16540 35652 17693 35680
rect 16540 35640 16546 35652
rect 17681 35649 17693 35652
rect 17727 35649 17739 35683
rect 23201 35683 23259 35689
rect 17681 35643 17739 35649
rect 19352 35652 20484 35680
rect 15010 35572 15016 35624
rect 15068 35572 15074 35624
rect 17957 35615 18015 35621
rect 17957 35581 17969 35615
rect 18003 35612 18015 35615
rect 18322 35612 18328 35624
rect 18003 35584 18328 35612
rect 18003 35581 18015 35584
rect 17957 35575 18015 35581
rect 18322 35572 18328 35584
rect 18380 35572 18386 35624
rect 18598 35572 18604 35624
rect 18656 35612 18662 35624
rect 19352 35612 19380 35652
rect 20456 35621 20484 35652
rect 23201 35649 23213 35683
rect 23247 35649 23259 35683
rect 23201 35643 23259 35649
rect 18656 35584 19380 35612
rect 19429 35615 19487 35621
rect 18656 35572 18662 35584
rect 19429 35581 19441 35615
rect 19475 35612 19487 35615
rect 20441 35615 20499 35621
rect 19475 35584 20392 35612
rect 19475 35581 19487 35584
rect 19429 35575 19487 35581
rect 15565 35547 15623 35553
rect 15565 35544 15577 35547
rect 14844 35516 15577 35544
rect 15565 35513 15577 35516
rect 15611 35544 15623 35547
rect 17310 35544 17316 35556
rect 15611 35516 17316 35544
rect 15611 35513 15623 35516
rect 15565 35507 15623 35513
rect 17310 35504 17316 35516
rect 17368 35504 17374 35556
rect 12584 35448 13492 35476
rect 12584 35436 12590 35448
rect 14182 35436 14188 35488
rect 14240 35476 14246 35488
rect 14461 35479 14519 35485
rect 14461 35476 14473 35479
rect 14240 35448 14473 35476
rect 14240 35436 14246 35448
rect 14461 35445 14473 35448
rect 14507 35445 14519 35479
rect 14461 35439 14519 35445
rect 15654 35436 15660 35488
rect 15712 35476 15718 35488
rect 16025 35479 16083 35485
rect 16025 35476 16037 35479
rect 15712 35448 16037 35476
rect 15712 35436 15718 35448
rect 16025 35445 16037 35448
rect 16071 35476 16083 35479
rect 16666 35476 16672 35488
rect 16071 35448 16672 35476
rect 16071 35445 16083 35448
rect 16025 35439 16083 35445
rect 16666 35436 16672 35448
rect 16724 35436 16730 35488
rect 19518 35436 19524 35488
rect 19576 35476 19582 35488
rect 19889 35479 19947 35485
rect 19889 35476 19901 35479
rect 19576 35448 19901 35476
rect 19576 35436 19582 35448
rect 19889 35445 19901 35448
rect 19935 35445 19947 35479
rect 20364 35476 20392 35584
rect 20441 35581 20453 35615
rect 20487 35581 20499 35615
rect 20441 35575 20499 35581
rect 22462 35572 22468 35624
rect 22520 35572 22526 35624
rect 22649 35615 22707 35621
rect 22649 35581 22661 35615
rect 22695 35612 22707 35615
rect 23106 35612 23112 35624
rect 22695 35584 23112 35612
rect 22695 35581 22707 35584
rect 22649 35575 22707 35581
rect 23106 35572 23112 35584
rect 23164 35572 23170 35624
rect 23477 35615 23535 35621
rect 23477 35581 23489 35615
rect 23523 35612 23535 35615
rect 25222 35612 25228 35624
rect 23523 35584 25228 35612
rect 23523 35581 23535 35584
rect 23477 35575 23535 35581
rect 25222 35572 25228 35584
rect 25280 35572 25286 35624
rect 20714 35476 20720 35488
rect 20364 35448 20720 35476
rect 19889 35439 19947 35445
rect 20714 35436 20720 35448
rect 20772 35436 20778 35488
rect 20990 35436 20996 35488
rect 21048 35476 21054 35488
rect 21269 35479 21327 35485
rect 21269 35476 21281 35479
rect 21048 35448 21281 35476
rect 21048 35436 21054 35448
rect 21269 35445 21281 35448
rect 21315 35445 21327 35479
rect 21269 35439 21327 35445
rect 22005 35479 22063 35485
rect 22005 35445 22017 35479
rect 22051 35476 22063 35479
rect 23658 35476 23664 35488
rect 22051 35448 23664 35476
rect 22051 35445 22063 35448
rect 22005 35439 22063 35445
rect 23658 35436 23664 35448
rect 23716 35436 23722 35488
rect 25406 35436 25412 35488
rect 25464 35436 25470 35488
rect 1104 35386 25852 35408
rect 1104 35334 2950 35386
rect 3002 35334 3014 35386
rect 3066 35334 3078 35386
rect 3130 35334 3142 35386
rect 3194 35334 3206 35386
rect 3258 35334 12950 35386
rect 13002 35334 13014 35386
rect 13066 35334 13078 35386
rect 13130 35334 13142 35386
rect 13194 35334 13206 35386
rect 13258 35334 22950 35386
rect 23002 35334 23014 35386
rect 23066 35334 23078 35386
rect 23130 35334 23142 35386
rect 23194 35334 23206 35386
rect 23258 35334 25852 35386
rect 1104 35312 25852 35334
rect 6638 35232 6644 35284
rect 6696 35272 6702 35284
rect 8021 35275 8079 35281
rect 8021 35272 8033 35275
rect 6696 35244 8033 35272
rect 6696 35232 6702 35244
rect 8021 35241 8033 35244
rect 8067 35272 8079 35275
rect 8754 35272 8760 35284
rect 8067 35244 8760 35272
rect 8067 35241 8079 35244
rect 8021 35235 8079 35241
rect 8754 35232 8760 35244
rect 8812 35232 8818 35284
rect 8846 35232 8852 35284
rect 8904 35272 8910 35284
rect 9125 35275 9183 35281
rect 9125 35272 9137 35275
rect 8904 35244 9137 35272
rect 8904 35232 8910 35244
rect 9125 35241 9137 35244
rect 9171 35241 9183 35275
rect 9125 35235 9183 35241
rect 10584 35275 10642 35281
rect 10584 35241 10596 35275
rect 10630 35272 10642 35275
rect 11054 35272 11060 35284
rect 10630 35244 11060 35272
rect 10630 35241 10642 35244
rect 10584 35235 10642 35241
rect 11054 35232 11060 35244
rect 11112 35232 11118 35284
rect 11330 35232 11336 35284
rect 11388 35272 11394 35284
rect 12805 35275 12863 35281
rect 12805 35272 12817 35275
rect 11388 35244 12817 35272
rect 11388 35232 11394 35244
rect 12805 35241 12817 35244
rect 12851 35241 12863 35275
rect 12805 35235 12863 35241
rect 13188 35244 14688 35272
rect 8110 35164 8116 35216
rect 8168 35204 8174 35216
rect 8297 35207 8355 35213
rect 8297 35204 8309 35207
rect 8168 35176 8309 35204
rect 8168 35164 8174 35176
rect 8297 35173 8309 35176
rect 8343 35173 8355 35207
rect 8297 35167 8355 35173
rect 8386 35164 8392 35216
rect 8444 35204 8450 35216
rect 9490 35204 9496 35216
rect 8444 35176 9496 35204
rect 8444 35164 8450 35176
rect 9490 35164 9496 35176
rect 9548 35204 9554 35216
rect 9548 35176 10364 35204
rect 9548 35164 9554 35176
rect 6086 35136 6092 35148
rect 5184 35108 6092 35136
rect 5184 35077 5212 35108
rect 6086 35096 6092 35108
rect 6144 35096 6150 35148
rect 6546 35096 6552 35148
rect 6604 35096 6610 35148
rect 7742 35096 7748 35148
rect 7800 35096 7806 35148
rect 5169 35071 5227 35077
rect 5169 35037 5181 35071
rect 5215 35037 5227 35071
rect 5169 35031 5227 35037
rect 5626 35028 5632 35080
rect 5684 35068 5690 35080
rect 6273 35071 6331 35077
rect 6273 35068 6285 35071
rect 5684 35040 6285 35068
rect 5684 35028 5690 35040
rect 6273 35037 6285 35040
rect 6319 35037 6331 35071
rect 7760 35068 7788 35096
rect 8128 35068 8156 35164
rect 9306 35096 9312 35148
rect 9364 35136 9370 35148
rect 10336 35145 10364 35176
rect 11698 35164 11704 35216
rect 11756 35164 11762 35216
rect 12710 35164 12716 35216
rect 12768 35204 12774 35216
rect 13188 35204 13216 35244
rect 14182 35204 14188 35216
rect 12768 35176 13216 35204
rect 13280 35176 14188 35204
rect 12768 35164 12774 35176
rect 9677 35139 9735 35145
rect 9677 35136 9689 35139
rect 9364 35108 9689 35136
rect 9364 35096 9370 35108
rect 9677 35105 9689 35108
rect 9723 35105 9735 35139
rect 9677 35099 9735 35105
rect 10321 35139 10379 35145
rect 10321 35105 10333 35139
rect 10367 35136 10379 35139
rect 11716 35136 11744 35164
rect 13280 35145 13308 35176
rect 14182 35164 14188 35176
rect 14240 35164 14246 35216
rect 14660 35204 14688 35244
rect 14734 35232 14740 35284
rect 14792 35272 14798 35284
rect 14921 35275 14979 35281
rect 14921 35272 14933 35275
rect 14792 35244 14933 35272
rect 14792 35232 14798 35244
rect 14921 35241 14933 35244
rect 14967 35241 14979 35275
rect 14921 35235 14979 35241
rect 15746 35232 15752 35284
rect 15804 35272 15810 35284
rect 17221 35275 17279 35281
rect 17221 35272 17233 35275
rect 15804 35244 17233 35272
rect 15804 35232 15810 35244
rect 17221 35241 17233 35244
rect 17267 35241 17279 35275
rect 17221 35235 17279 35241
rect 17310 35232 17316 35284
rect 17368 35272 17374 35284
rect 17368 35244 20760 35272
rect 17368 35232 17374 35244
rect 19242 35204 19248 35216
rect 14660 35176 15608 35204
rect 10367 35108 11744 35136
rect 13265 35139 13323 35145
rect 10367 35105 10379 35108
rect 10321 35099 10379 35105
rect 13265 35105 13277 35139
rect 13311 35105 13323 35139
rect 13265 35099 13323 35105
rect 13357 35139 13415 35145
rect 13357 35105 13369 35139
rect 13403 35105 13415 35139
rect 13357 35099 13415 35105
rect 8478 35068 8484 35080
rect 7682 35040 8484 35068
rect 6273 35031 6331 35037
rect 8478 35028 8484 35040
rect 8536 35068 8542 35080
rect 9858 35068 9864 35080
rect 8536 35040 9864 35068
rect 8536 35028 8542 35040
rect 9858 35028 9864 35040
rect 9916 35028 9922 35080
rect 11974 35028 11980 35080
rect 12032 35068 12038 35080
rect 13372 35068 13400 35099
rect 15470 35096 15476 35148
rect 15528 35096 15534 35148
rect 15580 35136 15608 35176
rect 17972 35176 19248 35204
rect 17972 35136 18000 35176
rect 19242 35164 19248 35176
rect 19300 35164 19306 35216
rect 20732 35204 20760 35244
rect 20990 35232 20996 35284
rect 21048 35272 21054 35284
rect 21048 35244 23704 35272
rect 21048 35232 21054 35244
rect 22002 35204 22008 35216
rect 20732 35176 22008 35204
rect 22002 35164 22008 35176
rect 22060 35164 22066 35216
rect 15580 35108 18000 35136
rect 18046 35096 18052 35148
rect 18104 35136 18110 35148
rect 18322 35136 18328 35148
rect 18104 35108 18328 35136
rect 18104 35096 18110 35108
rect 18322 35096 18328 35108
rect 18380 35136 18386 35148
rect 19429 35139 19487 35145
rect 19429 35136 19441 35139
rect 18380 35108 19441 35136
rect 18380 35096 18386 35108
rect 19429 35105 19441 35108
rect 19475 35136 19487 35139
rect 20162 35136 20168 35148
rect 19475 35108 20168 35136
rect 19475 35105 19487 35108
rect 19429 35099 19487 35105
rect 20162 35096 20168 35108
rect 20220 35096 20226 35148
rect 22281 35139 22339 35145
rect 22281 35105 22293 35139
rect 22327 35136 22339 35139
rect 23290 35136 23296 35148
rect 22327 35108 23296 35136
rect 22327 35105 22339 35108
rect 22281 35099 22339 35105
rect 23290 35096 23296 35108
rect 23348 35096 23354 35148
rect 23676 35136 23704 35244
rect 25222 35232 25228 35284
rect 25280 35232 25286 35284
rect 24394 35136 24400 35148
rect 23676 35108 24400 35136
rect 12032 35040 13400 35068
rect 12032 35028 12038 35040
rect 14274 35028 14280 35080
rect 14332 35028 14338 35080
rect 18233 35071 18291 35077
rect 9493 35003 9551 35009
rect 9493 35000 9505 35003
rect 7852 34972 9505 35000
rect 5810 34892 5816 34944
rect 5868 34892 5874 34944
rect 7282 34892 7288 34944
rect 7340 34932 7346 34944
rect 7852 34932 7880 34972
rect 9493 34969 9505 34972
rect 9539 34969 9551 35003
rect 9876 35000 9904 35028
rect 9876 34972 11086 35000
rect 9493 34963 9551 34969
rect 12342 34960 12348 35012
rect 12400 35000 12406 35012
rect 12437 35003 12495 35009
rect 12437 35000 12449 35003
rect 12400 34972 12449 35000
rect 12400 34960 12406 34972
rect 12437 34969 12449 34972
rect 12483 35000 12495 35003
rect 13446 35000 13452 35012
rect 12483 34972 13452 35000
rect 12483 34969 12495 34972
rect 12437 34963 12495 34969
rect 13446 34960 13452 34972
rect 13504 34960 13510 35012
rect 15746 34960 15752 35012
rect 15804 34960 15810 35012
rect 7340 34904 7880 34932
rect 9585 34935 9643 34941
rect 7340 34892 7346 34904
rect 9585 34901 9597 34935
rect 9631 34932 9643 34935
rect 11238 34932 11244 34944
rect 9631 34904 11244 34932
rect 9631 34901 9643 34904
rect 9585 34895 9643 34901
rect 11238 34892 11244 34904
rect 11296 34892 11302 34944
rect 12066 34892 12072 34944
rect 12124 34892 12130 34944
rect 13173 34935 13231 34941
rect 13173 34901 13185 34935
rect 13219 34932 13231 34935
rect 14918 34932 14924 34944
rect 13219 34904 14924 34932
rect 13219 34901 13231 34904
rect 13173 34895 13231 34901
rect 14918 34892 14924 34904
rect 14976 34892 14982 34944
rect 16574 34892 16580 34944
rect 16632 34932 16638 34944
rect 16868 34932 16896 35054
rect 18233 35037 18245 35071
rect 18279 35037 18291 35071
rect 23676 35054 23704 35108
rect 24394 35096 24400 35108
rect 24452 35096 24458 35148
rect 24581 35071 24639 35077
rect 24581 35068 24593 35071
rect 18233 35031 18291 35037
rect 24044 35040 24593 35068
rect 17497 34935 17555 34941
rect 17497 34932 17509 34935
rect 16632 34904 17509 34932
rect 16632 34892 16638 34904
rect 17497 34901 17509 34904
rect 17543 34901 17555 34935
rect 18248 34932 18276 35031
rect 18877 35003 18935 35009
rect 18877 34969 18889 35003
rect 18923 35000 18935 35003
rect 19705 35003 19763 35009
rect 19705 35000 19717 35003
rect 18923 34972 19717 35000
rect 18923 34969 18935 34972
rect 18877 34963 18935 34969
rect 19705 34969 19717 34972
rect 19751 34969 19763 35003
rect 20990 35000 20996 35012
rect 20930 34972 20996 35000
rect 19705 34963 19763 34969
rect 20990 34960 20996 34972
rect 21048 34960 21054 35012
rect 22186 34960 22192 35012
rect 22244 35000 22250 35012
rect 22557 35003 22615 35009
rect 22557 35000 22569 35003
rect 22244 34972 22569 35000
rect 22244 34960 22250 34972
rect 22557 34969 22569 34972
rect 22603 34969 22615 35003
rect 22557 34963 22615 34969
rect 24044 34944 24072 35040
rect 24581 35037 24593 35040
rect 24627 35037 24639 35071
rect 24581 35031 24639 35037
rect 18506 34932 18512 34944
rect 18248 34904 18512 34932
rect 17497 34895 17555 34901
rect 18506 34892 18512 34904
rect 18564 34932 18570 34944
rect 21082 34932 21088 34944
rect 18564 34904 21088 34932
rect 18564 34892 18570 34904
rect 21082 34892 21088 34904
rect 21140 34892 21146 34944
rect 21177 34935 21235 34941
rect 21177 34901 21189 34935
rect 21223 34932 21235 34935
rect 21266 34932 21272 34944
rect 21223 34904 21272 34932
rect 21223 34901 21235 34904
rect 21177 34895 21235 34901
rect 21266 34892 21272 34904
rect 21324 34892 21330 34944
rect 21637 34935 21695 34941
rect 21637 34901 21649 34935
rect 21683 34932 21695 34935
rect 22370 34932 22376 34944
rect 21683 34904 22376 34932
rect 21683 34901 21695 34904
rect 21637 34895 21695 34901
rect 22370 34892 22376 34904
rect 22428 34892 22434 34944
rect 24026 34892 24032 34944
rect 24084 34892 24090 34944
rect 1104 34842 25852 34864
rect 1104 34790 7950 34842
rect 8002 34790 8014 34842
rect 8066 34790 8078 34842
rect 8130 34790 8142 34842
rect 8194 34790 8206 34842
rect 8258 34790 17950 34842
rect 18002 34790 18014 34842
rect 18066 34790 18078 34842
rect 18130 34790 18142 34842
rect 18194 34790 18206 34842
rect 18258 34790 25852 34842
rect 1104 34768 25852 34790
rect 7469 34731 7527 34737
rect 7469 34697 7481 34731
rect 7515 34728 7527 34731
rect 7742 34728 7748 34740
rect 7515 34700 7748 34728
rect 7515 34697 7527 34700
rect 7469 34691 7527 34697
rect 7742 34688 7748 34700
rect 7800 34688 7806 34740
rect 8386 34688 8392 34740
rect 8444 34688 8450 34740
rect 9493 34731 9551 34737
rect 9493 34697 9505 34731
rect 9539 34728 9551 34731
rect 9582 34728 9588 34740
rect 9539 34700 9588 34728
rect 9539 34697 9551 34700
rect 9493 34691 9551 34697
rect 9582 34688 9588 34700
rect 9640 34688 9646 34740
rect 9858 34688 9864 34740
rect 9916 34688 9922 34740
rect 11054 34688 11060 34740
rect 11112 34728 11118 34740
rect 12437 34731 12495 34737
rect 12437 34728 12449 34731
rect 11112 34700 12449 34728
rect 11112 34688 11118 34700
rect 12437 34697 12449 34700
rect 12483 34697 12495 34731
rect 12437 34691 12495 34697
rect 12710 34688 12716 34740
rect 12768 34728 12774 34740
rect 13081 34731 13139 34737
rect 13081 34728 13093 34731
rect 12768 34700 13093 34728
rect 12768 34688 12774 34700
rect 13081 34697 13093 34700
rect 13127 34697 13139 34731
rect 13081 34691 13139 34697
rect 13538 34688 13544 34740
rect 13596 34688 13602 34740
rect 15194 34688 15200 34740
rect 15252 34728 15258 34740
rect 15565 34731 15623 34737
rect 15565 34728 15577 34731
rect 15252 34700 15577 34728
rect 15252 34688 15258 34700
rect 15565 34697 15577 34700
rect 15611 34697 15623 34731
rect 15565 34691 15623 34697
rect 15746 34688 15752 34740
rect 15804 34728 15810 34740
rect 17957 34731 18015 34737
rect 17957 34728 17969 34731
rect 15804 34700 17969 34728
rect 15804 34688 15810 34700
rect 17957 34697 17969 34700
rect 18003 34697 18015 34731
rect 17957 34691 18015 34697
rect 18782 34688 18788 34740
rect 18840 34688 18846 34740
rect 18877 34731 18935 34737
rect 18877 34697 18889 34731
rect 18923 34728 18935 34731
rect 18966 34728 18972 34740
rect 18923 34700 18972 34728
rect 18923 34697 18935 34700
rect 18877 34691 18935 34697
rect 18966 34688 18972 34700
rect 19024 34728 19030 34740
rect 19429 34731 19487 34737
rect 19429 34728 19441 34731
rect 19024 34700 19441 34728
rect 19024 34688 19030 34700
rect 19429 34697 19441 34700
rect 19475 34697 19487 34731
rect 19429 34691 19487 34697
rect 22465 34731 22523 34737
rect 22465 34697 22477 34731
rect 22511 34728 22523 34731
rect 22554 34728 22560 34740
rect 22511 34700 22560 34728
rect 22511 34697 22523 34700
rect 22465 34691 22523 34697
rect 22554 34688 22560 34700
rect 22612 34728 22618 34740
rect 23017 34731 23075 34737
rect 23017 34728 23029 34731
rect 22612 34700 23029 34728
rect 22612 34688 22618 34700
rect 23017 34697 23029 34700
rect 23063 34697 23075 34731
rect 23017 34691 23075 34697
rect 8404 34660 8432 34688
rect 7760 34632 8432 34660
rect 7760 34601 7788 34632
rect 8478 34620 8484 34672
rect 8536 34620 8542 34672
rect 15654 34660 15660 34672
rect 9324 34632 15660 34660
rect 7745 34595 7803 34601
rect 7745 34561 7757 34595
rect 7791 34561 7803 34595
rect 7745 34555 7803 34561
rect 7374 34484 7380 34536
rect 7432 34524 7438 34536
rect 9324 34524 9352 34632
rect 15654 34620 15660 34632
rect 15712 34620 15718 34672
rect 15933 34663 15991 34669
rect 15933 34629 15945 34663
rect 15979 34660 15991 34663
rect 19518 34660 19524 34672
rect 15979 34632 19524 34660
rect 15979 34629 15991 34632
rect 15933 34623 15991 34629
rect 19518 34620 19524 34632
rect 19576 34620 19582 34672
rect 21085 34663 21143 34669
rect 21085 34629 21097 34663
rect 21131 34660 21143 34663
rect 21542 34660 21548 34672
rect 21131 34632 21548 34660
rect 21131 34629 21143 34632
rect 21085 34623 21143 34629
rect 21542 34620 21548 34632
rect 21600 34620 21606 34672
rect 24305 34663 24363 34669
rect 24305 34629 24317 34663
rect 24351 34660 24363 34663
rect 24394 34660 24400 34672
rect 24351 34632 24400 34660
rect 24351 34629 24363 34632
rect 24305 34623 24363 34629
rect 24394 34620 24400 34632
rect 24452 34660 24458 34672
rect 25406 34660 25412 34672
rect 24452 34632 25412 34660
rect 24452 34620 24458 34632
rect 25406 34620 25412 34632
rect 25464 34620 25470 34672
rect 11793 34595 11851 34601
rect 11793 34561 11805 34595
rect 11839 34592 11851 34595
rect 12526 34592 12532 34604
rect 11839 34564 12532 34592
rect 11839 34561 11851 34564
rect 11793 34555 11851 34561
rect 12526 34552 12532 34564
rect 12584 34552 12590 34604
rect 13449 34595 13507 34601
rect 13449 34561 13461 34595
rect 13495 34592 13507 34595
rect 13538 34592 13544 34604
rect 13495 34564 13544 34592
rect 13495 34561 13507 34564
rect 13449 34555 13507 34561
rect 13538 34552 13544 34564
rect 13596 34592 13602 34604
rect 14185 34595 14243 34601
rect 14185 34592 14197 34595
rect 13596 34564 14197 34592
rect 13596 34552 13602 34564
rect 14185 34561 14197 34564
rect 14231 34592 14243 34595
rect 16850 34592 16856 34604
rect 14231 34564 16856 34592
rect 14231 34561 14243 34564
rect 14185 34555 14243 34561
rect 16850 34552 16856 34564
rect 16908 34552 16914 34604
rect 17313 34595 17371 34601
rect 17313 34561 17325 34595
rect 17359 34592 17371 34595
rect 20070 34592 20076 34604
rect 17359 34564 20076 34592
rect 17359 34561 17371 34564
rect 17313 34555 17371 34561
rect 20070 34552 20076 34564
rect 20128 34552 20134 34604
rect 20993 34595 21051 34601
rect 20993 34561 21005 34595
rect 21039 34592 21051 34595
rect 22373 34595 22431 34601
rect 21039 34564 21312 34592
rect 21039 34561 21051 34564
rect 20993 34555 21051 34561
rect 7432 34496 9352 34524
rect 13633 34527 13691 34533
rect 7432 34484 7438 34496
rect 13633 34493 13645 34527
rect 13679 34493 13691 34527
rect 13633 34487 13691 34493
rect 5994 34416 6000 34468
rect 6052 34456 6058 34468
rect 6822 34456 6828 34468
rect 6052 34428 6828 34456
rect 6052 34416 6058 34428
rect 6822 34416 6828 34428
rect 6880 34416 6886 34468
rect 11054 34416 11060 34468
rect 11112 34456 11118 34468
rect 12066 34456 12072 34468
rect 11112 34428 12072 34456
rect 11112 34416 11118 34428
rect 12066 34416 12072 34428
rect 12124 34456 12130 34468
rect 13648 34456 13676 34487
rect 16022 34484 16028 34536
rect 16080 34484 16086 34536
rect 16117 34527 16175 34533
rect 16117 34493 16129 34527
rect 16163 34493 16175 34527
rect 16117 34487 16175 34493
rect 18969 34527 19027 34533
rect 18969 34493 18981 34527
rect 19015 34493 19027 34527
rect 18969 34487 19027 34493
rect 19981 34527 20039 34533
rect 19981 34493 19993 34527
rect 20027 34524 20039 34527
rect 20898 34524 20904 34536
rect 20027 34496 20904 34524
rect 20027 34493 20039 34496
rect 19981 34487 20039 34493
rect 12124 34428 13676 34456
rect 12124 34416 12130 34428
rect 15746 34416 15752 34468
rect 15804 34456 15810 34468
rect 16132 34456 16160 34487
rect 15804 34428 16160 34456
rect 15804 34416 15810 34428
rect 17862 34416 17868 34468
rect 17920 34456 17926 34468
rect 18984 34456 19012 34487
rect 20898 34484 20904 34496
rect 20956 34484 20962 34536
rect 21177 34527 21235 34533
rect 21177 34493 21189 34527
rect 21223 34493 21235 34527
rect 21284 34524 21312 34564
rect 22373 34561 22385 34595
rect 22419 34561 22431 34595
rect 22373 34555 22431 34561
rect 21634 34524 21640 34536
rect 21284 34496 21640 34524
rect 21177 34487 21235 34493
rect 17920 34428 19012 34456
rect 17920 34416 17926 34428
rect 8008 34391 8066 34397
rect 8008 34357 8020 34391
rect 8054 34388 8066 34391
rect 8386 34388 8392 34400
rect 8054 34360 8392 34388
rect 8054 34357 8066 34360
rect 8008 34351 8066 34357
rect 8386 34348 8392 34360
rect 8444 34348 8450 34400
rect 15286 34348 15292 34400
rect 15344 34388 15350 34400
rect 16390 34388 16396 34400
rect 15344 34360 16396 34388
rect 15344 34348 15350 34360
rect 16390 34348 16396 34360
rect 16448 34348 16454 34400
rect 18414 34348 18420 34400
rect 18472 34348 18478 34400
rect 20622 34348 20628 34400
rect 20680 34348 20686 34400
rect 21082 34348 21088 34400
rect 21140 34388 21146 34400
rect 21192 34388 21220 34487
rect 21634 34484 21640 34496
rect 21692 34484 21698 34536
rect 22094 34484 22100 34536
rect 22152 34524 22158 34536
rect 22388 34524 22416 34555
rect 23566 34552 23572 34604
rect 23624 34592 23630 34604
rect 23937 34595 23995 34601
rect 23937 34592 23949 34595
rect 23624 34564 23949 34592
rect 23624 34552 23630 34564
rect 23937 34561 23949 34564
rect 23983 34561 23995 34595
rect 23937 34555 23995 34561
rect 25314 34552 25320 34604
rect 25372 34552 25378 34604
rect 22152 34496 22416 34524
rect 22557 34527 22615 34533
rect 22152 34484 22158 34496
rect 22557 34493 22569 34527
rect 22603 34493 22615 34527
rect 24670 34524 24676 34536
rect 22557 34487 22615 34493
rect 23768 34496 24676 34524
rect 22572 34400 22600 34487
rect 23768 34465 23796 34496
rect 24670 34484 24676 34496
rect 24728 34484 24734 34536
rect 23753 34459 23811 34465
rect 23753 34425 23765 34459
rect 23799 34425 23811 34459
rect 23753 34419 23811 34425
rect 21140 34360 21220 34388
rect 21140 34348 21146 34360
rect 22002 34348 22008 34400
rect 22060 34348 22066 34400
rect 22554 34348 22560 34400
rect 22612 34348 22618 34400
rect 23566 34348 23572 34400
rect 23624 34388 23630 34400
rect 25133 34391 25191 34397
rect 25133 34388 25145 34391
rect 23624 34360 25145 34388
rect 23624 34348 23630 34360
rect 25133 34357 25145 34360
rect 25179 34357 25191 34391
rect 25133 34351 25191 34357
rect 1104 34298 25852 34320
rect 1104 34246 2950 34298
rect 3002 34246 3014 34298
rect 3066 34246 3078 34298
rect 3130 34246 3142 34298
rect 3194 34246 3206 34298
rect 3258 34246 12950 34298
rect 13002 34246 13014 34298
rect 13066 34246 13078 34298
rect 13130 34246 13142 34298
rect 13194 34246 13206 34298
rect 13258 34246 22950 34298
rect 23002 34246 23014 34298
rect 23066 34246 23078 34298
rect 23130 34246 23142 34298
rect 23194 34246 23206 34298
rect 23258 34246 25852 34298
rect 1104 34224 25852 34246
rect 7834 34144 7840 34196
rect 7892 34144 7898 34196
rect 9766 34144 9772 34196
rect 9824 34144 9830 34196
rect 10226 34144 10232 34196
rect 10284 34144 10290 34196
rect 16298 34184 16304 34196
rect 11348 34156 16304 34184
rect 8294 34076 8300 34128
rect 8352 34116 8358 34128
rect 8352 34088 10824 34116
rect 8352 34076 8358 34088
rect 5810 34008 5816 34060
rect 5868 34008 5874 34060
rect 7098 34008 7104 34060
rect 7156 34048 7162 34060
rect 8389 34051 8447 34057
rect 8389 34048 8401 34051
rect 7156 34020 8401 34048
rect 7156 34008 7162 34020
rect 8389 34017 8401 34020
rect 8435 34017 8447 34051
rect 8389 34011 8447 34017
rect 10686 34008 10692 34060
rect 10744 34008 10750 34060
rect 10796 34057 10824 34088
rect 10781 34051 10839 34057
rect 10781 34017 10793 34051
rect 10827 34017 10839 34051
rect 10781 34011 10839 34017
rect 5534 33940 5540 33992
rect 5592 33940 5598 33992
rect 6914 33940 6920 33992
rect 6972 33980 6978 33992
rect 7742 33980 7748 33992
rect 6972 33952 7748 33980
rect 6972 33940 6978 33952
rect 7742 33940 7748 33952
rect 7800 33940 7806 33992
rect 9125 33983 9183 33989
rect 9125 33949 9137 33983
rect 9171 33980 9183 33983
rect 9582 33980 9588 33992
rect 9171 33952 9588 33980
rect 9171 33949 9183 33952
rect 9125 33943 9183 33949
rect 9582 33940 9588 33952
rect 9640 33940 9646 33992
rect 10597 33983 10655 33989
rect 10597 33949 10609 33983
rect 10643 33980 10655 33983
rect 11348 33980 11376 34156
rect 16298 34144 16304 34156
rect 16356 34144 16362 34196
rect 16390 34144 16396 34196
rect 16448 34184 16454 34196
rect 17405 34187 17463 34193
rect 16448 34156 16988 34184
rect 16448 34144 16454 34156
rect 13173 34119 13231 34125
rect 13173 34085 13185 34119
rect 13219 34116 13231 34119
rect 14274 34116 14280 34128
rect 13219 34088 14280 34116
rect 13219 34085 13231 34088
rect 13173 34079 13231 34085
rect 14274 34076 14280 34088
rect 14332 34116 14338 34128
rect 14826 34116 14832 34128
rect 14332 34088 14832 34116
rect 14332 34076 14338 34088
rect 14826 34076 14832 34088
rect 14884 34076 14890 34128
rect 16960 34116 16988 34156
rect 17405 34153 17417 34187
rect 17451 34184 17463 34187
rect 18506 34184 18512 34196
rect 17451 34156 18512 34184
rect 17451 34153 17463 34156
rect 17405 34147 17463 34153
rect 18506 34144 18512 34156
rect 18564 34144 18570 34196
rect 18616 34156 21128 34184
rect 18616 34116 18644 34156
rect 20990 34116 20996 34128
rect 16960 34088 18644 34116
rect 18708 34088 20996 34116
rect 18708 34060 18736 34088
rect 20990 34076 20996 34088
rect 21048 34076 21054 34128
rect 21100 34116 21128 34156
rect 21542 34144 21548 34196
rect 21600 34184 21606 34196
rect 21821 34187 21879 34193
rect 21821 34184 21833 34187
rect 21600 34156 21833 34184
rect 21600 34144 21606 34156
rect 21821 34153 21833 34156
rect 21867 34153 21879 34187
rect 21821 34147 21879 34153
rect 21910 34144 21916 34196
rect 21968 34184 21974 34196
rect 23842 34184 23848 34196
rect 21968 34156 23848 34184
rect 21968 34144 21974 34156
rect 23842 34144 23848 34156
rect 23900 34144 23906 34196
rect 25314 34144 25320 34196
rect 25372 34144 25378 34196
rect 25406 34144 25412 34196
rect 25464 34144 25470 34196
rect 22646 34116 22652 34128
rect 21100 34088 22652 34116
rect 22646 34076 22652 34088
rect 22704 34076 22710 34128
rect 11425 34051 11483 34057
rect 11425 34017 11437 34051
rect 11471 34048 11483 34051
rect 11698 34048 11704 34060
rect 11471 34020 11704 34048
rect 11471 34017 11483 34020
rect 11425 34011 11483 34017
rect 11698 34008 11704 34020
rect 11756 34048 11762 34060
rect 11756 34020 13768 34048
rect 11756 34008 11762 34020
rect 13740 33992 13768 34020
rect 16574 34008 16580 34060
rect 16632 34048 16638 34060
rect 17681 34051 17739 34057
rect 17681 34048 17693 34051
rect 16632 34020 17693 34048
rect 16632 34008 16638 34020
rect 17681 34017 17693 34020
rect 17727 34048 17739 34051
rect 18690 34048 18696 34060
rect 17727 34020 18696 34048
rect 17727 34017 17739 34020
rect 17681 34011 17739 34017
rect 18690 34008 18696 34020
rect 18748 34008 18754 34060
rect 21266 34048 21272 34060
rect 19812 34020 21272 34048
rect 13446 33980 13452 33992
rect 10643 33952 11376 33980
rect 12834 33952 13452 33980
rect 10643 33949 10655 33952
rect 10597 33943 10655 33949
rect 13446 33940 13452 33952
rect 13504 33940 13510 33992
rect 13722 33940 13728 33992
rect 13780 33980 13786 33992
rect 19812 33989 19840 34020
rect 21266 34008 21272 34020
rect 21324 34008 21330 34060
rect 22833 34051 22891 34057
rect 22833 34017 22845 34051
rect 22879 34048 22891 34051
rect 22922 34048 22928 34060
rect 22879 34020 22928 34048
rect 22879 34017 22891 34020
rect 22833 34011 22891 34017
rect 22922 34008 22928 34020
rect 22980 34008 22986 34060
rect 23017 34051 23075 34057
rect 23017 34017 23029 34051
rect 23063 34048 23075 34051
rect 24026 34048 24032 34060
rect 23063 34020 24032 34048
rect 23063 34017 23075 34020
rect 23017 34011 23075 34017
rect 24026 34008 24032 34020
rect 24084 34008 24090 34060
rect 15657 33983 15715 33989
rect 15657 33980 15669 33983
rect 13780 33952 15669 33980
rect 13780 33940 13786 33952
rect 15657 33949 15669 33952
rect 15703 33949 15715 33983
rect 15657 33943 15715 33949
rect 19797 33983 19855 33989
rect 19797 33949 19809 33983
rect 19843 33949 19855 33983
rect 19797 33943 19855 33949
rect 20714 33940 20720 33992
rect 20772 33980 20778 33992
rect 20901 33983 20959 33989
rect 20901 33980 20913 33983
rect 20772 33952 20913 33980
rect 20772 33940 20778 33952
rect 20901 33949 20913 33952
rect 20947 33949 20959 33983
rect 22741 33983 22799 33989
rect 22741 33980 22753 33983
rect 20901 33943 20959 33949
rect 21008 33952 22753 33980
rect 8570 33912 8576 33924
rect 7300 33884 8576 33912
rect 7300 33853 7328 33884
rect 8570 33872 8576 33884
rect 8628 33872 8634 33924
rect 11701 33915 11759 33921
rect 11701 33881 11713 33915
rect 11747 33881 11759 33915
rect 11701 33875 11759 33881
rect 7285 33847 7343 33853
rect 7285 33813 7297 33847
rect 7331 33813 7343 33847
rect 7285 33807 7343 33813
rect 7466 33804 7472 33856
rect 7524 33844 7530 33856
rect 8205 33847 8263 33853
rect 8205 33844 8217 33847
rect 7524 33816 8217 33844
rect 7524 33804 7530 33816
rect 8205 33813 8217 33816
rect 8251 33813 8263 33847
rect 8205 33807 8263 33813
rect 8297 33847 8355 33853
rect 8297 33813 8309 33847
rect 8343 33844 8355 33847
rect 10502 33844 10508 33856
rect 8343 33816 10508 33844
rect 8343 33813 8355 33816
rect 8297 33807 8355 33813
rect 10502 33804 10508 33816
rect 10560 33804 10566 33856
rect 11716 33844 11744 33875
rect 15930 33872 15936 33924
rect 15988 33872 15994 33924
rect 16574 33872 16580 33924
rect 16632 33872 16638 33924
rect 20530 33872 20536 33924
rect 20588 33912 20594 33924
rect 21008 33912 21036 33952
rect 22741 33949 22753 33952
rect 22787 33949 22799 33983
rect 22741 33943 22799 33949
rect 24762 33940 24768 33992
rect 24820 33940 24826 33992
rect 20588 33884 21036 33912
rect 21545 33915 21603 33921
rect 20588 33872 20594 33884
rect 21545 33881 21557 33915
rect 21591 33912 21603 33915
rect 21591 33884 21956 33912
rect 21591 33881 21603 33884
rect 21545 33875 21603 33881
rect 12434 33844 12440 33856
rect 11716 33816 12440 33844
rect 12434 33804 12440 33816
rect 12492 33804 12498 33856
rect 14274 33804 14280 33856
rect 14332 33844 14338 33856
rect 19521 33847 19579 33853
rect 19521 33844 19533 33847
rect 14332 33816 19533 33844
rect 14332 33804 14338 33816
rect 19521 33813 19533 33816
rect 19567 33844 19579 33847
rect 20162 33844 20168 33856
rect 19567 33816 20168 33844
rect 19567 33813 19579 33816
rect 19521 33807 19579 33813
rect 20162 33804 20168 33816
rect 20220 33804 20226 33856
rect 20438 33804 20444 33856
rect 20496 33804 20502 33856
rect 21928 33844 21956 33884
rect 22094 33844 22100 33856
rect 21928 33816 22100 33844
rect 22094 33804 22100 33816
rect 22152 33804 22158 33856
rect 22373 33847 22431 33853
rect 22373 33813 22385 33847
rect 22419 33844 22431 33847
rect 23934 33844 23940 33856
rect 22419 33816 23940 33844
rect 22419 33813 22431 33816
rect 22373 33807 22431 33813
rect 23934 33804 23940 33816
rect 23992 33804 23998 33856
rect 24578 33804 24584 33856
rect 24636 33804 24642 33856
rect 1104 33754 25852 33776
rect 1104 33702 7950 33754
rect 8002 33702 8014 33754
rect 8066 33702 8078 33754
rect 8130 33702 8142 33754
rect 8194 33702 8206 33754
rect 8258 33702 17950 33754
rect 18002 33702 18014 33754
rect 18066 33702 18078 33754
rect 18130 33702 18142 33754
rect 18194 33702 18206 33754
rect 18258 33702 25852 33754
rect 1104 33680 25852 33702
rect 7285 33643 7343 33649
rect 7285 33609 7297 33643
rect 7331 33640 7343 33643
rect 7742 33640 7748 33652
rect 7331 33612 7748 33640
rect 7331 33609 7343 33612
rect 7285 33603 7343 33609
rect 7742 33600 7748 33612
rect 7800 33600 7806 33652
rect 8846 33600 8852 33652
rect 8904 33640 8910 33652
rect 10505 33643 10563 33649
rect 10505 33640 10517 33643
rect 8904 33612 10517 33640
rect 8904 33600 8910 33612
rect 10505 33609 10517 33612
rect 10551 33640 10563 33643
rect 10962 33640 10968 33652
rect 10551 33612 10968 33640
rect 10551 33609 10563 33612
rect 10505 33603 10563 33609
rect 10962 33600 10968 33612
rect 11020 33600 11026 33652
rect 12618 33600 12624 33652
rect 12676 33640 12682 33652
rect 12805 33643 12863 33649
rect 12805 33640 12817 33643
rect 12676 33612 12817 33640
rect 12676 33600 12682 33612
rect 12805 33609 12817 33612
rect 12851 33609 12863 33643
rect 12805 33603 12863 33609
rect 13265 33643 13323 33649
rect 13265 33609 13277 33643
rect 13311 33640 13323 33643
rect 20438 33640 20444 33652
rect 13311 33612 17080 33640
rect 13311 33609 13323 33612
rect 13265 33603 13323 33609
rect 12713 33575 12771 33581
rect 12713 33541 12725 33575
rect 12759 33572 12771 33575
rect 13280 33572 13308 33603
rect 12759 33544 13308 33572
rect 12759 33541 12771 33544
rect 12713 33535 12771 33541
rect 13446 33532 13452 33584
rect 13504 33572 13510 33584
rect 13504 33544 14766 33572
rect 13504 33532 13510 33544
rect 1302 33464 1308 33516
rect 1360 33504 1366 33516
rect 1765 33507 1823 33513
rect 1765 33504 1777 33507
rect 1360 33476 1777 33504
rect 1360 33464 1366 33476
rect 1765 33473 1777 33476
rect 1811 33504 1823 33507
rect 2041 33507 2099 33513
rect 2041 33504 2053 33507
rect 1811 33476 2053 33504
rect 1811 33473 1823 33476
rect 1765 33467 1823 33473
rect 2041 33473 2053 33476
rect 2087 33473 2099 33507
rect 2041 33467 2099 33473
rect 7561 33507 7619 33513
rect 7561 33473 7573 33507
rect 7607 33504 7619 33507
rect 7650 33504 7656 33516
rect 7607 33476 7656 33504
rect 7607 33473 7619 33476
rect 7561 33467 7619 33473
rect 7650 33464 7656 33476
rect 7708 33464 7714 33516
rect 12526 33464 12532 33516
rect 12584 33504 12590 33516
rect 13173 33507 13231 33513
rect 13173 33504 13185 33507
rect 12584 33476 13185 33504
rect 12584 33464 12590 33476
rect 13173 33473 13185 33476
rect 13219 33473 13231 33507
rect 13173 33467 13231 33473
rect 13722 33464 13728 33516
rect 13780 33504 13786 33516
rect 14001 33507 14059 33513
rect 14001 33504 14013 33507
rect 13780 33476 14013 33504
rect 13780 33464 13786 33476
rect 14001 33473 14013 33476
rect 14047 33473 14059 33507
rect 14001 33467 14059 33473
rect 5534 33396 5540 33448
rect 5592 33436 5598 33448
rect 5629 33439 5687 33445
rect 5629 33436 5641 33439
rect 5592 33408 5641 33436
rect 5592 33396 5598 33408
rect 5629 33405 5641 33408
rect 5675 33405 5687 33439
rect 5629 33399 5687 33405
rect 9766 33396 9772 33448
rect 9824 33396 9830 33448
rect 13354 33396 13360 33448
rect 13412 33396 13418 33448
rect 13446 33396 13452 33448
rect 13504 33436 13510 33448
rect 13630 33436 13636 33448
rect 13504 33408 13636 33436
rect 13504 33396 13510 33408
rect 13630 33396 13636 33408
rect 13688 33396 13694 33448
rect 14277 33439 14335 33445
rect 14277 33405 14289 33439
rect 14323 33436 14335 33439
rect 16114 33436 16120 33448
rect 14323 33408 16120 33436
rect 14323 33405 14335 33408
rect 14277 33399 14335 33405
rect 16114 33396 16120 33408
rect 16172 33396 16178 33448
rect 17052 33436 17080 33612
rect 18616 33612 20444 33640
rect 18616 33581 18644 33612
rect 20438 33600 20444 33612
rect 20496 33600 20502 33652
rect 20530 33600 20536 33652
rect 20588 33600 20594 33652
rect 20898 33600 20904 33652
rect 20956 33600 20962 33652
rect 22370 33600 22376 33652
rect 22428 33600 22434 33652
rect 25038 33600 25044 33652
rect 25096 33640 25102 33652
rect 25225 33643 25283 33649
rect 25225 33640 25237 33643
rect 25096 33612 25237 33640
rect 25096 33600 25102 33612
rect 25225 33609 25237 33612
rect 25271 33609 25283 33643
rect 25225 33603 25283 33609
rect 18601 33575 18659 33581
rect 18601 33541 18613 33575
rect 18647 33541 18659 33575
rect 18601 33535 18659 33541
rect 18690 33532 18696 33584
rect 18748 33572 18754 33584
rect 18748 33544 19090 33572
rect 18748 33532 18754 33544
rect 20162 33532 20168 33584
rect 20220 33572 20226 33584
rect 20993 33575 21051 33581
rect 20993 33572 21005 33575
rect 20220 33544 21005 33572
rect 20220 33532 20226 33544
rect 20993 33541 21005 33544
rect 21039 33541 21051 33575
rect 20993 33535 21051 33541
rect 21450 33532 21456 33584
rect 21508 33572 21514 33584
rect 22465 33575 22523 33581
rect 22465 33572 22477 33575
rect 21508 33544 22477 33572
rect 21508 33532 21514 33544
rect 22465 33541 22477 33544
rect 22511 33572 22523 33575
rect 23474 33572 23480 33584
rect 22511 33544 23480 33572
rect 22511 33541 22523 33544
rect 22465 33535 22523 33541
rect 23474 33532 23480 33544
rect 23532 33532 23538 33584
rect 18322 33464 18328 33516
rect 18380 33464 18386 33516
rect 21266 33464 21272 33516
rect 21324 33504 21330 33516
rect 21324 33476 22324 33504
rect 21324 33464 21330 33476
rect 19794 33436 19800 33448
rect 17052 33408 19800 33436
rect 19794 33396 19800 33408
rect 19852 33396 19858 33448
rect 20070 33396 20076 33448
rect 20128 33396 20134 33448
rect 21177 33439 21235 33445
rect 21177 33405 21189 33439
rect 21223 33436 21235 33439
rect 22186 33436 22192 33448
rect 21223 33408 22192 33436
rect 21223 33405 21235 33408
rect 21177 33399 21235 33405
rect 22186 33396 22192 33408
rect 22244 33396 22250 33448
rect 19812 33368 19840 33396
rect 20162 33368 20168 33380
rect 19812 33340 20168 33368
rect 20162 33328 20168 33340
rect 20220 33328 20226 33380
rect 20990 33328 20996 33380
rect 21048 33368 21054 33380
rect 21545 33371 21603 33377
rect 21545 33368 21557 33371
rect 21048 33340 21557 33368
rect 21048 33328 21054 33340
rect 21545 33337 21557 33340
rect 21591 33337 21603 33371
rect 22296 33368 22324 33476
rect 24854 33464 24860 33516
rect 24912 33464 24918 33516
rect 22557 33439 22615 33445
rect 22557 33405 22569 33439
rect 22603 33405 22615 33439
rect 22557 33399 22615 33405
rect 22572 33368 22600 33399
rect 23382 33396 23388 33448
rect 23440 33436 23446 33448
rect 23477 33439 23535 33445
rect 23477 33436 23489 33439
rect 23440 33408 23489 33436
rect 23440 33396 23446 33408
rect 23477 33405 23489 33408
rect 23523 33405 23535 33439
rect 23477 33399 23535 33405
rect 23750 33396 23756 33448
rect 23808 33396 23814 33448
rect 22296 33340 22600 33368
rect 21545 33331 21603 33337
rect 1581 33303 1639 33309
rect 1581 33269 1593 33303
rect 1627 33300 1639 33303
rect 3418 33300 3424 33312
rect 1627 33272 3424 33300
rect 1627 33269 1639 33272
rect 1581 33263 1639 33269
rect 3418 33260 3424 33272
rect 3476 33260 3482 33312
rect 7834 33260 7840 33312
rect 7892 33300 7898 33312
rect 8205 33303 8263 33309
rect 8205 33300 8217 33303
rect 7892 33272 8217 33300
rect 7892 33260 7898 33272
rect 8205 33269 8217 33272
rect 8251 33269 8263 33303
rect 8205 33263 8263 33269
rect 12526 33260 12532 33312
rect 12584 33260 12590 33312
rect 13630 33260 13636 33312
rect 13688 33300 13694 33312
rect 15746 33300 15752 33312
rect 13688 33272 15752 33300
rect 13688 33260 13694 33272
rect 15746 33260 15752 33272
rect 15804 33260 15810 33312
rect 16022 33260 16028 33312
rect 16080 33300 16086 33312
rect 16574 33300 16580 33312
rect 16080 33272 16580 33300
rect 16080 33260 16086 33272
rect 16574 33260 16580 33272
rect 16632 33260 16638 33312
rect 21634 33260 21640 33312
rect 21692 33300 21698 33312
rect 22005 33303 22063 33309
rect 22005 33300 22017 33303
rect 21692 33272 22017 33300
rect 21692 33260 21698 33272
rect 22005 33269 22017 33272
rect 22051 33269 22063 33303
rect 22005 33263 22063 33269
rect 1104 33210 25852 33232
rect 1104 33158 2950 33210
rect 3002 33158 3014 33210
rect 3066 33158 3078 33210
rect 3130 33158 3142 33210
rect 3194 33158 3206 33210
rect 3258 33158 12950 33210
rect 13002 33158 13014 33210
rect 13066 33158 13078 33210
rect 13130 33158 13142 33210
rect 13194 33158 13206 33210
rect 13258 33158 22950 33210
rect 23002 33158 23014 33210
rect 23066 33158 23078 33210
rect 23130 33158 23142 33210
rect 23194 33158 23206 33210
rect 23258 33158 25852 33210
rect 1104 33136 25852 33158
rect 7558 33056 7564 33108
rect 7616 33056 7622 33108
rect 9398 33056 9404 33108
rect 9456 33056 9462 33108
rect 10870 33056 10876 33108
rect 10928 33056 10934 33108
rect 11882 33056 11888 33108
rect 11940 33056 11946 33108
rect 15930 33056 15936 33108
rect 15988 33096 15994 33108
rect 16117 33099 16175 33105
rect 16117 33096 16129 33099
rect 15988 33068 16129 33096
rect 15988 33056 15994 33068
rect 16117 33065 16129 33068
rect 16163 33065 16175 33099
rect 16117 33059 16175 33065
rect 16574 33056 16580 33108
rect 16632 33056 16638 33108
rect 17034 33056 17040 33108
rect 17092 33096 17098 33108
rect 17678 33096 17684 33108
rect 17092 33068 17684 33096
rect 17092 33056 17098 33068
rect 17678 33056 17684 33068
rect 17736 33056 17742 33108
rect 19521 33099 19579 33105
rect 19521 33065 19533 33099
rect 19567 33096 19579 33099
rect 22462 33096 22468 33108
rect 19567 33068 22468 33096
rect 19567 33065 19579 33068
rect 19521 33059 19579 33065
rect 22462 33056 22468 33068
rect 22520 33056 22526 33108
rect 22646 33056 22652 33108
rect 22704 33096 22710 33108
rect 25133 33099 25191 33105
rect 25133 33096 25145 33099
rect 22704 33068 25145 33096
rect 22704 33056 22710 33068
rect 25133 33065 25145 33068
rect 25179 33065 25191 33099
rect 25133 33059 25191 33065
rect 7101 33031 7159 33037
rect 7101 32997 7113 33031
rect 7147 33028 7159 33031
rect 7650 33028 7656 33040
rect 7147 33000 7656 33028
rect 7147 32997 7159 33000
rect 7101 32991 7159 32997
rect 7650 32988 7656 33000
rect 7708 32988 7714 33040
rect 8478 32988 8484 33040
rect 8536 33028 8542 33040
rect 9950 33028 9956 33040
rect 8536 33000 9956 33028
rect 8536 32988 8542 33000
rect 9950 32988 9956 33000
rect 10008 32988 10014 33040
rect 5353 32963 5411 32969
rect 5353 32929 5365 32963
rect 5399 32960 5411 32963
rect 5626 32960 5632 32972
rect 5399 32932 5632 32960
rect 5399 32929 5411 32932
rect 5353 32923 5411 32929
rect 5626 32920 5632 32932
rect 5684 32960 5690 32972
rect 6270 32960 6276 32972
rect 5684 32932 6276 32960
rect 5684 32920 5690 32932
rect 6270 32920 6276 32932
rect 6328 32920 6334 32972
rect 6914 32960 6920 32972
rect 6748 32932 6920 32960
rect 6748 32878 6776 32932
rect 6914 32920 6920 32932
rect 6972 32920 6978 32972
rect 8205 32963 8263 32969
rect 8205 32929 8217 32963
rect 8251 32960 8263 32963
rect 8294 32960 8300 32972
rect 8251 32932 8300 32960
rect 8251 32929 8263 32932
rect 8205 32923 8263 32929
rect 8220 32892 8248 32923
rect 8294 32920 8300 32932
rect 8352 32920 8358 32972
rect 8386 32920 8392 32972
rect 8444 32960 8450 32972
rect 10045 32963 10103 32969
rect 10045 32960 10057 32963
rect 8444 32932 10057 32960
rect 8444 32920 8450 32932
rect 10045 32929 10057 32932
rect 10091 32929 10103 32963
rect 10045 32923 10103 32929
rect 10597 32963 10655 32969
rect 10597 32929 10609 32963
rect 10643 32960 10655 32963
rect 11330 32960 11336 32972
rect 10643 32932 11336 32960
rect 10643 32929 10655 32932
rect 10597 32923 10655 32929
rect 6932 32864 8248 32892
rect 5629 32827 5687 32833
rect 5629 32793 5641 32827
rect 5675 32793 5687 32827
rect 5629 32787 5687 32793
rect 5644 32756 5672 32787
rect 6932 32756 6960 32864
rect 9766 32852 9772 32904
rect 9824 32852 9830 32904
rect 10060 32892 10088 32923
rect 11330 32920 11336 32932
rect 11388 32920 11394 32972
rect 11517 32963 11575 32969
rect 11517 32929 11529 32963
rect 11563 32960 11575 32963
rect 11900 32960 11928 33056
rect 14277 33031 14335 33037
rect 14277 32997 14289 33031
rect 14323 33028 14335 33031
rect 18690 33028 18696 33040
rect 14323 33000 18696 33028
rect 14323 32997 14335 33000
rect 14277 32991 14335 32997
rect 18690 32988 18696 33000
rect 18748 32988 18754 33040
rect 22830 33028 22836 33040
rect 20180 33000 22836 33028
rect 11563 32932 11928 32960
rect 11563 32929 11575 32932
rect 11517 32923 11575 32929
rect 14458 32920 14464 32972
rect 14516 32960 14522 32972
rect 14737 32963 14795 32969
rect 14737 32960 14749 32963
rect 14516 32932 14749 32960
rect 14516 32920 14522 32932
rect 14737 32929 14749 32932
rect 14783 32929 14795 32963
rect 14737 32923 14795 32929
rect 14826 32920 14832 32972
rect 14884 32920 14890 32972
rect 17034 32920 17040 32972
rect 17092 32920 17098 32972
rect 17218 32920 17224 32972
rect 17276 32960 17282 32972
rect 17402 32960 17408 32972
rect 17276 32932 17408 32960
rect 17276 32920 17282 32932
rect 17402 32920 17408 32932
rect 17460 32920 17466 32972
rect 20180 32969 20208 33000
rect 22830 32988 22836 33000
rect 22888 32988 22894 33040
rect 23014 32988 23020 33040
rect 23072 32988 23078 33040
rect 23658 32988 23664 33040
rect 23716 32988 23722 33040
rect 20165 32963 20223 32969
rect 20165 32929 20177 32963
rect 20211 32929 20223 32963
rect 20165 32923 20223 32929
rect 20714 32920 20720 32972
rect 20772 32960 20778 32972
rect 21361 32963 21419 32969
rect 21361 32960 21373 32963
rect 20772 32932 21373 32960
rect 20772 32920 20778 32932
rect 21361 32929 21373 32932
rect 21407 32960 21419 32963
rect 22557 32963 22615 32969
rect 22557 32960 22569 32963
rect 21407 32932 22569 32960
rect 21407 32929 21419 32932
rect 21361 32923 21419 32929
rect 22557 32929 22569 32932
rect 22603 32929 22615 32963
rect 22557 32923 22615 32929
rect 22646 32920 22652 32972
rect 22704 32960 22710 32972
rect 23385 32963 23443 32969
rect 23385 32960 23397 32963
rect 22704 32932 23397 32960
rect 22704 32920 22710 32932
rect 23385 32929 23397 32932
rect 23431 32929 23443 32963
rect 23385 32923 23443 32929
rect 11974 32892 11980 32904
rect 10060 32864 11980 32892
rect 11974 32852 11980 32864
rect 12032 32852 12038 32904
rect 14366 32852 14372 32904
rect 14424 32892 14430 32904
rect 15473 32895 15531 32901
rect 15473 32892 15485 32895
rect 14424 32864 15485 32892
rect 14424 32852 14430 32864
rect 15473 32861 15485 32864
rect 15519 32861 15531 32895
rect 15473 32855 15531 32861
rect 16298 32852 16304 32904
rect 16356 32892 16362 32904
rect 18785 32895 18843 32901
rect 18785 32892 18797 32895
rect 16356 32864 18797 32892
rect 16356 32852 16362 32864
rect 18785 32861 18797 32864
rect 18831 32892 18843 32895
rect 21269 32895 21327 32901
rect 18831 32864 20024 32892
rect 18831 32861 18843 32864
rect 18785 32855 18843 32861
rect 7742 32784 7748 32836
rect 7800 32824 7806 32836
rect 8021 32827 8079 32833
rect 8021 32824 8033 32827
rect 7800 32796 8033 32824
rect 7800 32784 7806 32796
rect 8021 32793 8033 32796
rect 8067 32793 8079 32827
rect 8021 32787 8079 32793
rect 8570 32784 8576 32836
rect 8628 32824 8634 32836
rect 12250 32824 12256 32836
rect 8628 32796 12256 32824
rect 8628 32784 8634 32796
rect 12250 32784 12256 32796
rect 12308 32824 12314 32836
rect 16666 32824 16672 32836
rect 12308 32796 16672 32824
rect 12308 32784 12314 32796
rect 16666 32784 16672 32796
rect 16724 32784 16730 32836
rect 19996 32833 20024 32864
rect 21269 32861 21281 32895
rect 21315 32892 21327 32895
rect 21450 32892 21456 32904
rect 21315 32864 21456 32892
rect 21315 32861 21327 32864
rect 21269 32855 21327 32861
rect 21450 32852 21456 32864
rect 21508 32892 21514 32904
rect 21726 32892 21732 32904
rect 21508 32864 21732 32892
rect 21508 32852 21514 32864
rect 21726 32852 21732 32864
rect 21784 32852 21790 32904
rect 21910 32852 21916 32904
rect 21968 32892 21974 32904
rect 22373 32895 22431 32901
rect 22373 32892 22385 32895
rect 21968 32864 22385 32892
rect 21968 32852 21974 32864
rect 22373 32861 22385 32864
rect 22419 32892 22431 32895
rect 23676 32892 23704 32988
rect 22419 32864 23704 32892
rect 24857 32895 24915 32901
rect 22419 32861 22431 32864
rect 22373 32855 22431 32861
rect 24857 32861 24869 32895
rect 24903 32892 24915 32895
rect 25314 32892 25320 32904
rect 24903 32864 25320 32892
rect 24903 32861 24915 32864
rect 24857 32855 24915 32861
rect 25314 32852 25320 32864
rect 25372 32852 25378 32904
rect 19981 32827 20039 32833
rect 16776 32796 19104 32824
rect 5644 32728 6960 32756
rect 7650 32716 7656 32768
rect 7708 32756 7714 32768
rect 7929 32759 7987 32765
rect 7929 32756 7941 32759
rect 7708 32728 7941 32756
rect 7708 32716 7714 32728
rect 7929 32725 7941 32728
rect 7975 32725 7987 32759
rect 7929 32719 7987 32725
rect 9766 32716 9772 32768
rect 9824 32756 9830 32768
rect 9861 32759 9919 32765
rect 9861 32756 9873 32759
rect 9824 32728 9873 32756
rect 9824 32716 9830 32728
rect 9861 32725 9873 32728
rect 9907 32725 9919 32759
rect 9861 32719 9919 32725
rect 10962 32716 10968 32768
rect 11020 32756 11026 32768
rect 11241 32759 11299 32765
rect 11241 32756 11253 32759
rect 11020 32728 11253 32756
rect 11020 32716 11026 32728
rect 11241 32725 11253 32728
rect 11287 32725 11299 32759
rect 11241 32719 11299 32725
rect 11330 32716 11336 32768
rect 11388 32756 11394 32768
rect 14274 32756 14280 32768
rect 11388 32728 14280 32756
rect 11388 32716 11394 32728
rect 14274 32716 14280 32728
rect 14332 32716 14338 32768
rect 14642 32716 14648 32768
rect 14700 32716 14706 32768
rect 14734 32716 14740 32768
rect 14792 32756 14798 32768
rect 16776 32756 16804 32796
rect 14792 32728 16804 32756
rect 14792 32716 14798 32728
rect 16942 32716 16948 32768
rect 17000 32716 17006 32768
rect 19076 32765 19104 32796
rect 19981 32793 19993 32827
rect 20027 32824 20039 32827
rect 21177 32827 21235 32833
rect 20027 32796 21128 32824
rect 20027 32793 20039 32796
rect 19981 32787 20039 32793
rect 19061 32759 19119 32765
rect 19061 32725 19073 32759
rect 19107 32756 19119 32759
rect 19889 32759 19947 32765
rect 19889 32756 19901 32759
rect 19107 32728 19901 32756
rect 19107 32725 19119 32728
rect 19061 32719 19119 32725
rect 19889 32725 19901 32728
rect 19935 32725 19947 32759
rect 19889 32719 19947 32725
rect 20809 32759 20867 32765
rect 20809 32725 20821 32759
rect 20855 32756 20867 32759
rect 20898 32756 20904 32768
rect 20855 32728 20904 32756
rect 20855 32725 20867 32728
rect 20809 32719 20867 32725
rect 20898 32716 20904 32728
rect 20956 32716 20962 32768
rect 21100 32756 21128 32796
rect 21177 32793 21189 32827
rect 21223 32824 21235 32827
rect 21358 32824 21364 32836
rect 21223 32796 21364 32824
rect 21223 32793 21235 32796
rect 21177 32787 21235 32793
rect 21358 32784 21364 32796
rect 21416 32784 21422 32836
rect 21910 32756 21916 32768
rect 21100 32728 21916 32756
rect 21910 32716 21916 32728
rect 21968 32716 21974 32768
rect 22005 32759 22063 32765
rect 22005 32725 22017 32759
rect 22051 32756 22063 32759
rect 22278 32756 22284 32768
rect 22051 32728 22284 32756
rect 22051 32725 22063 32728
rect 22005 32719 22063 32725
rect 22278 32716 22284 32728
rect 22336 32716 22342 32768
rect 22462 32716 22468 32768
rect 22520 32756 22526 32768
rect 22646 32756 22652 32768
rect 22520 32728 22652 32756
rect 22520 32716 22526 32728
rect 22646 32716 22652 32728
rect 22704 32716 22710 32768
rect 23198 32716 23204 32768
rect 23256 32716 23262 32768
rect 1104 32666 25852 32688
rect 1104 32614 7950 32666
rect 8002 32614 8014 32666
rect 8066 32614 8078 32666
rect 8130 32614 8142 32666
rect 8194 32614 8206 32666
rect 8258 32614 17950 32666
rect 18002 32614 18014 32666
rect 18066 32614 18078 32666
rect 18130 32614 18142 32666
rect 18194 32614 18206 32666
rect 18258 32614 25852 32666
rect 1104 32592 25852 32614
rect 4522 32512 4528 32564
rect 4580 32552 4586 32564
rect 4801 32555 4859 32561
rect 4801 32552 4813 32555
rect 4580 32524 4813 32552
rect 4580 32512 4586 32524
rect 4801 32521 4813 32524
rect 4847 32521 4859 32555
rect 4801 32515 4859 32521
rect 5169 32555 5227 32561
rect 5169 32521 5181 32555
rect 5215 32552 5227 32555
rect 5442 32552 5448 32564
rect 5215 32524 5448 32552
rect 5215 32521 5227 32524
rect 5169 32515 5227 32521
rect 4816 32484 4844 32515
rect 5442 32512 5448 32524
rect 5500 32512 5506 32564
rect 5534 32512 5540 32564
rect 5592 32512 5598 32564
rect 7009 32555 7067 32561
rect 7009 32521 7021 32555
rect 7055 32552 7067 32555
rect 7650 32552 7656 32564
rect 7055 32524 7656 32552
rect 7055 32521 7067 32524
rect 7009 32515 7067 32521
rect 7650 32512 7656 32524
rect 7708 32512 7714 32564
rect 9674 32552 9680 32564
rect 7760 32524 9680 32552
rect 5629 32487 5687 32493
rect 5629 32484 5641 32487
rect 4816 32456 5641 32484
rect 5552 32428 5580 32456
rect 5629 32453 5641 32456
rect 5675 32453 5687 32487
rect 7760 32484 7788 32524
rect 9674 32512 9680 32524
rect 9732 32512 9738 32564
rect 11238 32512 11244 32564
rect 11296 32552 11302 32564
rect 13725 32555 13783 32561
rect 13725 32552 13737 32555
rect 11296 32524 13737 32552
rect 11296 32512 11302 32524
rect 13725 32521 13737 32524
rect 13771 32521 13783 32555
rect 13725 32515 13783 32521
rect 14185 32555 14243 32561
rect 14185 32521 14197 32555
rect 14231 32552 14243 32555
rect 14231 32524 16068 32552
rect 14231 32521 14243 32524
rect 14185 32515 14243 32521
rect 5629 32447 5687 32453
rect 7668 32456 7788 32484
rect 5534 32376 5540 32428
rect 5592 32376 5598 32428
rect 6270 32376 6276 32428
rect 6328 32416 6334 32428
rect 7668 32425 7696 32456
rect 7834 32444 7840 32496
rect 7892 32484 7898 32496
rect 7929 32487 7987 32493
rect 7929 32484 7941 32487
rect 7892 32456 7941 32484
rect 7892 32444 7898 32456
rect 7929 32453 7941 32456
rect 7975 32453 7987 32487
rect 7929 32447 7987 32453
rect 8018 32444 8024 32496
rect 8076 32484 8082 32496
rect 8076 32456 8418 32484
rect 8076 32444 8082 32456
rect 9582 32444 9588 32496
rect 9640 32484 9646 32496
rect 13357 32487 13415 32493
rect 13357 32484 13369 32487
rect 9640 32456 13369 32484
rect 9640 32444 9646 32456
rect 13357 32453 13369 32456
rect 13403 32484 13415 32487
rect 13403 32456 14320 32484
rect 13403 32453 13415 32456
rect 13357 32447 13415 32453
rect 7653 32419 7711 32425
rect 7653 32416 7665 32419
rect 6328 32388 7665 32416
rect 6328 32376 6334 32388
rect 7653 32385 7665 32388
rect 7699 32385 7711 32419
rect 7653 32379 7711 32385
rect 9398 32376 9404 32428
rect 9456 32416 9462 32428
rect 9769 32419 9827 32425
rect 9769 32416 9781 32419
rect 9456 32388 9781 32416
rect 9456 32376 9462 32388
rect 9769 32385 9781 32388
rect 9815 32385 9827 32419
rect 9769 32379 9827 32385
rect 10226 32376 10232 32428
rect 10284 32416 10290 32428
rect 10686 32416 10692 32428
rect 10284 32388 10692 32416
rect 10284 32376 10290 32388
rect 10686 32376 10692 32388
rect 10744 32416 10750 32428
rect 14093 32419 14151 32425
rect 10744 32388 14044 32416
rect 10744 32376 10750 32388
rect 5813 32351 5871 32357
rect 5813 32317 5825 32351
rect 5859 32348 5871 32351
rect 6638 32348 6644 32360
rect 5859 32320 6644 32348
rect 5859 32317 5871 32320
rect 5813 32311 5871 32317
rect 6638 32308 6644 32320
rect 6696 32308 6702 32360
rect 6914 32308 6920 32360
rect 6972 32348 6978 32360
rect 8018 32348 8024 32360
rect 6972 32320 8024 32348
rect 6972 32308 6978 32320
rect 8018 32308 8024 32320
rect 8076 32308 8082 32360
rect 8294 32308 8300 32360
rect 8352 32348 8358 32360
rect 11701 32351 11759 32357
rect 11701 32348 11713 32351
rect 8352 32320 11713 32348
rect 8352 32308 8358 32320
rect 11701 32317 11713 32320
rect 11747 32317 11759 32351
rect 11701 32311 11759 32317
rect 12434 32308 12440 32360
rect 12492 32348 12498 32360
rect 12529 32351 12587 32357
rect 12529 32348 12541 32351
rect 12492 32320 12541 32348
rect 12492 32308 12498 32320
rect 12529 32317 12541 32320
rect 12575 32317 12587 32351
rect 12529 32311 12587 32317
rect 9401 32283 9459 32289
rect 9401 32249 9413 32283
rect 9447 32280 9459 32283
rect 10226 32280 10232 32292
rect 9447 32252 10232 32280
rect 9447 32249 9459 32252
rect 9401 32243 9459 32249
rect 10226 32240 10232 32252
rect 10284 32240 10290 32292
rect 14016 32280 14044 32388
rect 14093 32385 14105 32419
rect 14139 32416 14151 32419
rect 14182 32416 14188 32428
rect 14139 32388 14188 32416
rect 14139 32385 14151 32388
rect 14093 32379 14151 32385
rect 14182 32376 14188 32388
rect 14240 32376 14246 32428
rect 14292 32357 14320 32456
rect 15473 32419 15531 32425
rect 15473 32385 15485 32419
rect 15519 32416 15531 32419
rect 15930 32416 15936 32428
rect 15519 32388 15936 32416
rect 15519 32385 15531 32388
rect 15473 32379 15531 32385
rect 15930 32376 15936 32388
rect 15988 32376 15994 32428
rect 16040 32416 16068 32524
rect 16114 32512 16120 32564
rect 16172 32512 16178 32564
rect 17770 32512 17776 32564
rect 17828 32512 17834 32564
rect 19061 32555 19119 32561
rect 19061 32521 19073 32555
rect 19107 32552 19119 32555
rect 19426 32552 19432 32564
rect 19107 32524 19432 32552
rect 19107 32521 19119 32524
rect 19061 32515 19119 32521
rect 19426 32512 19432 32524
rect 19484 32552 19490 32564
rect 19702 32552 19708 32564
rect 19484 32524 19708 32552
rect 19484 32512 19490 32524
rect 19702 32512 19708 32524
rect 19760 32512 19766 32564
rect 20254 32512 20260 32564
rect 20312 32552 20318 32564
rect 20312 32524 23520 32552
rect 20312 32512 20318 32524
rect 16666 32444 16672 32496
rect 16724 32484 16730 32496
rect 16761 32487 16819 32493
rect 16761 32484 16773 32487
rect 16724 32456 16773 32484
rect 16724 32444 16730 32456
rect 16761 32453 16773 32456
rect 16807 32484 16819 32487
rect 17034 32484 17040 32496
rect 16807 32456 17040 32484
rect 16807 32453 16819 32456
rect 16761 32447 16819 32453
rect 17034 32444 17040 32456
rect 17092 32444 17098 32496
rect 17494 32444 17500 32496
rect 17552 32484 17558 32496
rect 17552 32456 19104 32484
rect 17552 32444 17558 32456
rect 18782 32416 18788 32428
rect 16040 32388 18788 32416
rect 18782 32376 18788 32388
rect 18840 32376 18846 32428
rect 18969 32419 19027 32425
rect 18969 32385 18981 32419
rect 19015 32385 19027 32419
rect 19076 32416 19104 32456
rect 19794 32444 19800 32496
rect 19852 32484 19858 32496
rect 20165 32487 20223 32493
rect 20165 32484 20177 32487
rect 19852 32456 20177 32484
rect 19852 32444 19858 32456
rect 20165 32453 20177 32456
rect 20211 32484 20223 32487
rect 20346 32484 20352 32496
rect 20211 32456 20352 32484
rect 20211 32453 20223 32456
rect 20165 32447 20223 32453
rect 20346 32444 20352 32456
rect 20404 32444 20410 32496
rect 21358 32444 21364 32496
rect 21416 32484 21422 32496
rect 21818 32484 21824 32496
rect 21416 32456 21824 32484
rect 21416 32444 21422 32456
rect 21818 32444 21824 32456
rect 21876 32484 21882 32496
rect 23198 32484 23204 32496
rect 21876 32456 23204 32484
rect 21876 32444 21882 32456
rect 23198 32444 23204 32456
rect 23256 32444 23262 32496
rect 21177 32419 21235 32425
rect 21177 32416 21189 32419
rect 19076 32388 21189 32416
rect 18969 32379 19027 32385
rect 21177 32385 21189 32388
rect 21223 32385 21235 32419
rect 21177 32379 21235 32385
rect 14277 32351 14335 32357
rect 14277 32317 14289 32351
rect 14323 32317 14335 32351
rect 14277 32311 14335 32317
rect 16574 32308 16580 32360
rect 16632 32348 16638 32360
rect 17865 32351 17923 32357
rect 17865 32348 17877 32351
rect 16632 32320 17877 32348
rect 16632 32308 16638 32320
rect 17865 32317 17877 32320
rect 17911 32317 17923 32351
rect 17865 32311 17923 32317
rect 17957 32351 18015 32357
rect 17957 32317 17969 32351
rect 18003 32317 18015 32351
rect 18984 32348 19012 32379
rect 22186 32376 22192 32428
rect 22244 32376 22250 32428
rect 22370 32376 22376 32428
rect 22428 32416 22434 32428
rect 23492 32425 23520 32524
rect 22833 32419 22891 32425
rect 22833 32416 22845 32419
rect 22428 32388 22845 32416
rect 22428 32376 22434 32388
rect 22833 32385 22845 32388
rect 22879 32385 22891 32419
rect 22833 32379 22891 32385
rect 23477 32419 23535 32425
rect 23477 32385 23489 32419
rect 23523 32385 23535 32419
rect 23477 32379 23535 32385
rect 24857 32419 24915 32425
rect 24857 32385 24869 32419
rect 24903 32416 24915 32419
rect 25317 32419 25375 32425
rect 25317 32416 25329 32419
rect 24903 32388 25329 32416
rect 24903 32385 24915 32388
rect 24857 32379 24915 32385
rect 25317 32385 25329 32388
rect 25363 32416 25375 32419
rect 25406 32416 25412 32428
rect 25363 32388 25412 32416
rect 25363 32385 25375 32388
rect 25317 32379 25375 32385
rect 25406 32376 25412 32388
rect 25464 32376 25470 32428
rect 17957 32311 18015 32317
rect 18432 32320 19012 32348
rect 15010 32280 15016 32292
rect 14016 32252 15016 32280
rect 15010 32240 15016 32252
rect 15068 32240 15074 32292
rect 16942 32280 16948 32292
rect 16408 32252 16948 32280
rect 8662 32172 8668 32224
rect 8720 32212 8726 32224
rect 9582 32212 9588 32224
rect 8720 32184 9588 32212
rect 8720 32172 8726 32184
rect 9582 32172 9588 32184
rect 9640 32172 9646 32224
rect 9858 32172 9864 32224
rect 9916 32212 9922 32224
rect 10873 32215 10931 32221
rect 10873 32212 10885 32215
rect 9916 32184 10885 32212
rect 9916 32172 9922 32184
rect 10873 32181 10885 32184
rect 10919 32181 10931 32215
rect 10873 32175 10931 32181
rect 13262 32172 13268 32224
rect 13320 32212 13326 32224
rect 13998 32212 14004 32224
rect 13320 32184 14004 32212
rect 13320 32172 13326 32184
rect 13998 32172 14004 32184
rect 14056 32212 14062 32224
rect 14182 32212 14188 32224
rect 14056 32184 14188 32212
rect 14056 32172 14062 32184
rect 14182 32172 14188 32184
rect 14240 32212 14246 32224
rect 14734 32212 14740 32224
rect 14240 32184 14740 32212
rect 14240 32172 14246 32184
rect 14734 32172 14740 32184
rect 14792 32172 14798 32224
rect 14826 32172 14832 32224
rect 14884 32212 14890 32224
rect 16408 32221 16436 32252
rect 16942 32240 16948 32252
rect 17000 32240 17006 32292
rect 17770 32240 17776 32292
rect 17828 32280 17834 32292
rect 17972 32280 18000 32311
rect 17828 32252 18000 32280
rect 17828 32240 17834 32252
rect 16393 32215 16451 32221
rect 16393 32212 16405 32215
rect 14884 32184 16405 32212
rect 14884 32172 14890 32184
rect 16393 32181 16405 32184
rect 16439 32181 16451 32215
rect 16393 32175 16451 32181
rect 16850 32172 16856 32224
rect 16908 32212 16914 32224
rect 17405 32215 17463 32221
rect 17405 32212 17417 32215
rect 16908 32184 17417 32212
rect 16908 32172 16914 32184
rect 17405 32181 17417 32184
rect 17451 32181 17463 32215
rect 17405 32175 17463 32181
rect 17678 32172 17684 32224
rect 17736 32212 17742 32224
rect 18432 32212 18460 32320
rect 18984 32280 19012 32320
rect 19242 32308 19248 32360
rect 19300 32308 19306 32360
rect 19334 32308 19340 32360
rect 19392 32348 19398 32360
rect 20257 32351 20315 32357
rect 20257 32348 20269 32351
rect 19392 32320 20269 32348
rect 19392 32308 19398 32320
rect 20257 32317 20269 32320
rect 20303 32317 20315 32351
rect 20257 32311 20315 32317
rect 20272 32280 20300 32311
rect 20438 32308 20444 32360
rect 20496 32308 20502 32360
rect 20714 32280 20720 32292
rect 18984 32252 19932 32280
rect 20272 32252 20720 32280
rect 17736 32184 18460 32212
rect 17736 32172 17742 32184
rect 18506 32172 18512 32224
rect 18564 32212 18570 32224
rect 18601 32215 18659 32221
rect 18601 32212 18613 32215
rect 18564 32184 18613 32212
rect 18564 32172 18570 32184
rect 18601 32181 18613 32184
rect 18647 32181 18659 32215
rect 18601 32175 18659 32181
rect 19518 32172 19524 32224
rect 19576 32212 19582 32224
rect 19797 32215 19855 32221
rect 19797 32212 19809 32215
rect 19576 32184 19809 32212
rect 19576 32172 19582 32184
rect 19797 32181 19809 32184
rect 19843 32181 19855 32215
rect 19904 32212 19932 32252
rect 20714 32240 20720 32252
rect 20772 32240 20778 32292
rect 21453 32283 21511 32289
rect 21453 32280 21465 32283
rect 20824 32252 21465 32280
rect 20824 32212 20852 32252
rect 21453 32249 21465 32252
rect 21499 32280 21511 32283
rect 25133 32283 25191 32289
rect 25133 32280 25145 32283
rect 21499 32252 25145 32280
rect 21499 32249 21511 32252
rect 21453 32243 21511 32249
rect 25133 32249 25145 32252
rect 25179 32249 25191 32283
rect 25133 32243 25191 32249
rect 19904 32184 20852 32212
rect 19797 32175 19855 32181
rect 20990 32172 20996 32224
rect 21048 32172 21054 32224
rect 21818 32172 21824 32224
rect 21876 32212 21882 32224
rect 22005 32215 22063 32221
rect 22005 32212 22017 32215
rect 21876 32184 22017 32212
rect 21876 32172 21882 32184
rect 22005 32181 22017 32184
rect 22051 32181 22063 32215
rect 22005 32175 22063 32181
rect 22462 32172 22468 32224
rect 22520 32212 22526 32224
rect 22649 32215 22707 32221
rect 22649 32212 22661 32215
rect 22520 32184 22661 32212
rect 22520 32172 22526 32184
rect 22649 32181 22661 32184
rect 22695 32181 22707 32215
rect 22649 32175 22707 32181
rect 22830 32172 22836 32224
rect 22888 32212 22894 32224
rect 23293 32215 23351 32221
rect 23293 32212 23305 32215
rect 22888 32184 23305 32212
rect 22888 32172 22894 32184
rect 23293 32181 23305 32184
rect 23339 32181 23351 32215
rect 23293 32175 23351 32181
rect 1104 32122 25852 32144
rect 1104 32070 2950 32122
rect 3002 32070 3014 32122
rect 3066 32070 3078 32122
rect 3130 32070 3142 32122
rect 3194 32070 3206 32122
rect 3258 32070 12950 32122
rect 13002 32070 13014 32122
rect 13066 32070 13078 32122
rect 13130 32070 13142 32122
rect 13194 32070 13206 32122
rect 13258 32070 22950 32122
rect 23002 32070 23014 32122
rect 23066 32070 23078 32122
rect 23130 32070 23142 32122
rect 23194 32070 23206 32122
rect 23258 32070 25852 32122
rect 1104 32048 25852 32070
rect 8021 32011 8079 32017
rect 8021 31977 8033 32011
rect 8067 32008 8079 32011
rect 8386 32008 8392 32020
rect 8067 31980 8392 32008
rect 8067 31977 8079 31980
rect 8021 31971 8079 31977
rect 8386 31968 8392 31980
rect 8444 31968 8450 32020
rect 8570 31968 8576 32020
rect 8628 31968 8634 32020
rect 9950 31968 9956 32020
rect 10008 32008 10014 32020
rect 11241 32011 11299 32017
rect 10008 31980 10916 32008
rect 10008 31968 10014 31980
rect 7834 31900 7840 31952
rect 7892 31940 7898 31952
rect 8588 31940 8616 31968
rect 7892 31912 8616 31940
rect 10888 31940 10916 31980
rect 11241 31977 11253 32011
rect 11287 32008 11299 32011
rect 11974 32008 11980 32020
rect 11287 31980 11980 32008
rect 11287 31977 11299 31980
rect 11241 31971 11299 31977
rect 11974 31968 11980 31980
rect 12032 31968 12038 32020
rect 12069 32011 12127 32017
rect 12069 31977 12081 32011
rect 12115 32008 12127 32011
rect 14642 32008 14648 32020
rect 12115 31980 14648 32008
rect 12115 31977 12127 31980
rect 12069 31971 12127 31977
rect 14642 31968 14648 31980
rect 14700 31968 14706 32020
rect 15930 31968 15936 32020
rect 15988 32008 15994 32020
rect 17037 32011 17095 32017
rect 17037 32008 17049 32011
rect 15988 31980 17049 32008
rect 15988 31968 15994 31980
rect 17037 31977 17049 31980
rect 17083 32008 17095 32011
rect 18598 32008 18604 32020
rect 17083 31980 18604 32008
rect 17083 31977 17095 31980
rect 17037 31971 17095 31977
rect 18598 31968 18604 31980
rect 18656 31968 18662 32020
rect 19242 31968 19248 32020
rect 19300 32008 19306 32020
rect 19429 32011 19487 32017
rect 19429 32008 19441 32011
rect 19300 31980 19441 32008
rect 19300 31968 19306 31980
rect 19429 31977 19441 31980
rect 19475 31977 19487 32011
rect 19429 31971 19487 31977
rect 20714 31968 20720 32020
rect 20772 32008 20778 32020
rect 20993 32011 21051 32017
rect 20993 32008 21005 32011
rect 20772 31980 21005 32008
rect 20772 31968 20778 31980
rect 20993 31977 21005 31980
rect 21039 32008 21051 32011
rect 21266 32008 21272 32020
rect 21039 31980 21272 32008
rect 21039 31977 21051 31980
rect 20993 31971 21051 31977
rect 21266 31968 21272 31980
rect 21324 31968 21330 32020
rect 23750 31968 23756 32020
rect 23808 32008 23814 32020
rect 24029 32011 24087 32017
rect 24029 32008 24041 32011
rect 23808 31980 24041 32008
rect 23808 31968 23814 31980
rect 24029 31977 24041 31980
rect 24075 31977 24087 32011
rect 24029 31971 24087 31977
rect 11701 31943 11759 31949
rect 11701 31940 11713 31943
rect 10888 31912 11713 31940
rect 7892 31900 7898 31912
rect 11701 31909 11713 31912
rect 11747 31940 11759 31943
rect 14090 31940 14096 31952
rect 11747 31912 14096 31940
rect 11747 31909 11759 31912
rect 11701 31903 11759 31909
rect 6270 31832 6276 31884
rect 6328 31832 6334 31884
rect 6549 31875 6607 31881
rect 6549 31841 6561 31875
rect 6595 31872 6607 31875
rect 7852 31872 7880 31900
rect 6595 31844 7880 31872
rect 6595 31841 6607 31844
rect 6549 31835 6607 31841
rect 8018 31832 8024 31884
rect 8076 31872 8082 31884
rect 8297 31875 8355 31881
rect 8297 31872 8309 31875
rect 8076 31844 8309 31872
rect 8076 31832 8082 31844
rect 8297 31841 8309 31844
rect 8343 31841 8355 31875
rect 8297 31835 8355 31841
rect 8036 31804 8064 31832
rect 7682 31776 8064 31804
rect 8312 31804 8340 31835
rect 9398 31832 9404 31884
rect 9456 31832 9462 31884
rect 9490 31832 9496 31884
rect 9548 31832 9554 31884
rect 9769 31875 9827 31881
rect 9769 31841 9781 31875
rect 9815 31872 9827 31875
rect 9858 31872 9864 31884
rect 9815 31844 9864 31872
rect 9815 31841 9827 31844
rect 9769 31835 9827 31841
rect 9858 31832 9864 31844
rect 9916 31832 9922 31884
rect 9416 31804 9444 31832
rect 8312 31776 9536 31804
rect 9508 31736 9536 31776
rect 9508 31708 9720 31736
rect 10994 31708 11652 31736
rect 9692 31668 9720 31708
rect 11072 31668 11100 31708
rect 11624 31680 11652 31708
rect 9692 31640 11100 31668
rect 11606 31628 11612 31680
rect 11664 31628 11670 31680
rect 12360 31668 12388 31912
rect 14090 31900 14096 31912
rect 14148 31900 14154 31952
rect 16942 31900 16948 31952
rect 17000 31940 17006 31952
rect 17497 31943 17555 31949
rect 17497 31940 17509 31943
rect 17000 31912 17509 31940
rect 17000 31900 17006 31912
rect 17497 31909 17509 31912
rect 17543 31909 17555 31943
rect 18693 31943 18751 31949
rect 18693 31940 18705 31943
rect 17497 31903 17555 31909
rect 17880 31912 18705 31940
rect 12713 31875 12771 31881
rect 12713 31841 12725 31875
rect 12759 31872 12771 31875
rect 12802 31872 12808 31884
rect 12759 31844 12808 31872
rect 12759 31841 12771 31844
rect 12713 31835 12771 31841
rect 12802 31832 12808 31844
rect 12860 31832 12866 31884
rect 13446 31832 13452 31884
rect 13504 31872 13510 31884
rect 17678 31872 17684 31884
rect 13504 31844 17684 31872
rect 13504 31832 13510 31844
rect 17678 31832 17684 31844
rect 17736 31832 17742 31884
rect 12434 31764 12440 31816
rect 12492 31764 12498 31816
rect 15286 31764 15292 31816
rect 15344 31764 15350 31816
rect 15562 31696 15568 31748
rect 15620 31696 15626 31748
rect 15654 31696 15660 31748
rect 15712 31736 15718 31748
rect 16022 31736 16028 31748
rect 15712 31708 16028 31736
rect 15712 31696 15718 31708
rect 16022 31696 16028 31708
rect 16080 31696 16086 31748
rect 12529 31671 12587 31677
rect 12529 31668 12541 31671
rect 12360 31640 12541 31668
rect 12529 31637 12541 31640
rect 12575 31637 12587 31671
rect 12529 31631 12587 31637
rect 15286 31628 15292 31680
rect 15344 31668 15350 31680
rect 16482 31668 16488 31680
rect 15344 31640 16488 31668
rect 15344 31628 15350 31640
rect 16482 31628 16488 31640
rect 16540 31628 16546 31680
rect 16574 31628 16580 31680
rect 16632 31668 16638 31680
rect 17880 31677 17908 31912
rect 18693 31909 18705 31912
rect 18739 31909 18751 31943
rect 18693 31903 18751 31909
rect 19610 31900 19616 31952
rect 19668 31940 19674 31952
rect 19797 31943 19855 31949
rect 19797 31940 19809 31943
rect 19668 31912 19809 31940
rect 19668 31900 19674 31912
rect 19797 31909 19809 31912
rect 19843 31909 19855 31943
rect 20809 31943 20867 31949
rect 20809 31940 20821 31943
rect 19797 31903 19855 31909
rect 20272 31912 20821 31940
rect 18046 31832 18052 31884
rect 18104 31832 18110 31884
rect 18598 31832 18604 31884
rect 18656 31872 18662 31884
rect 18877 31875 18935 31881
rect 18877 31872 18889 31875
rect 18656 31844 18889 31872
rect 18656 31832 18662 31844
rect 18877 31841 18889 31844
rect 18923 31841 18935 31875
rect 18877 31835 18935 31841
rect 19337 31875 19395 31881
rect 19337 31841 19349 31875
rect 19383 31872 19395 31875
rect 19426 31872 19432 31884
rect 19383 31844 19432 31872
rect 19383 31841 19395 31844
rect 19337 31835 19395 31841
rect 19426 31832 19432 31844
rect 19484 31832 19490 31884
rect 20272 31881 20300 31912
rect 20809 31909 20821 31912
rect 20855 31940 20867 31943
rect 21542 31940 21548 31952
rect 20855 31912 21548 31940
rect 20855 31909 20867 31912
rect 20809 31903 20867 31909
rect 21542 31900 21548 31912
rect 21600 31900 21606 31952
rect 22005 31943 22063 31949
rect 22005 31909 22017 31943
rect 22051 31940 22063 31943
rect 23290 31940 23296 31952
rect 22051 31912 23296 31940
rect 22051 31909 22063 31912
rect 22005 31903 22063 31909
rect 23290 31900 23296 31912
rect 23348 31900 23354 31952
rect 23474 31900 23480 31952
rect 23532 31940 23538 31952
rect 25133 31943 25191 31949
rect 25133 31940 25145 31943
rect 23532 31912 25145 31940
rect 23532 31900 23538 31912
rect 25133 31909 25145 31912
rect 25179 31909 25191 31943
rect 25133 31903 25191 31909
rect 20257 31875 20315 31881
rect 20257 31841 20269 31875
rect 20303 31841 20315 31875
rect 20257 31835 20315 31841
rect 20346 31832 20352 31884
rect 20404 31832 20410 31884
rect 20898 31832 20904 31884
rect 20956 31872 20962 31884
rect 22465 31875 22523 31881
rect 22465 31872 22477 31875
rect 20956 31844 22477 31872
rect 20956 31832 20962 31844
rect 22465 31841 22477 31844
rect 22511 31841 22523 31875
rect 22465 31835 22523 31841
rect 22557 31875 22615 31881
rect 22557 31841 22569 31875
rect 22603 31872 22615 31875
rect 23658 31872 23664 31884
rect 22603 31844 23664 31872
rect 22603 31841 22615 31844
rect 22557 31835 22615 31841
rect 23658 31832 23664 31844
rect 23716 31832 23722 31884
rect 17957 31807 18015 31813
rect 17957 31773 17969 31807
rect 18003 31804 18015 31807
rect 18616 31804 18644 31832
rect 18003 31776 18644 31804
rect 18003 31773 18015 31776
rect 17957 31767 18015 31773
rect 20162 31764 20168 31816
rect 20220 31764 20226 31816
rect 22646 31764 22652 31816
rect 22704 31804 22710 31816
rect 23385 31807 23443 31813
rect 23385 31804 23397 31807
rect 22704 31776 23397 31804
rect 22704 31764 22710 31776
rect 23385 31773 23397 31776
rect 23431 31773 23443 31807
rect 23385 31767 23443 31773
rect 24857 31807 24915 31813
rect 24857 31773 24869 31807
rect 24903 31804 24915 31807
rect 25314 31804 25320 31816
rect 24903 31776 25320 31804
rect 24903 31773 24915 31776
rect 24857 31767 24915 31773
rect 25314 31764 25320 31776
rect 25372 31764 25378 31816
rect 20990 31696 20996 31748
rect 21048 31736 21054 31748
rect 21266 31736 21272 31748
rect 21048 31708 21272 31736
rect 21048 31696 21054 31708
rect 21266 31696 21272 31708
rect 21324 31696 21330 31748
rect 22278 31696 22284 31748
rect 22336 31736 22342 31748
rect 22373 31739 22431 31745
rect 22373 31736 22385 31739
rect 22336 31708 22385 31736
rect 22336 31696 22342 31708
rect 22373 31705 22385 31708
rect 22419 31705 22431 31739
rect 22373 31699 22431 31705
rect 17865 31671 17923 31677
rect 17865 31668 17877 31671
rect 16632 31640 17877 31668
rect 16632 31628 16638 31640
rect 17865 31637 17877 31640
rect 17911 31637 17923 31671
rect 17865 31631 17923 31637
rect 18322 31628 18328 31680
rect 18380 31668 18386 31680
rect 18509 31671 18567 31677
rect 18509 31668 18521 31671
rect 18380 31640 18521 31668
rect 18380 31628 18386 31640
rect 18509 31637 18521 31640
rect 18555 31637 18567 31671
rect 18509 31631 18567 31637
rect 20254 31628 20260 31680
rect 20312 31668 20318 31680
rect 20438 31668 20444 31680
rect 20312 31640 20444 31668
rect 20312 31628 20318 31640
rect 20438 31628 20444 31640
rect 20496 31628 20502 31680
rect 1104 31578 25852 31600
rect 1104 31526 7950 31578
rect 8002 31526 8014 31578
rect 8066 31526 8078 31578
rect 8130 31526 8142 31578
rect 8194 31526 8206 31578
rect 8258 31526 17950 31578
rect 18002 31526 18014 31578
rect 18066 31526 18078 31578
rect 18130 31526 18142 31578
rect 18194 31526 18206 31578
rect 18258 31526 25852 31578
rect 1104 31504 25852 31526
rect 7285 31467 7343 31473
rect 7285 31433 7297 31467
rect 7331 31464 7343 31467
rect 7466 31464 7472 31476
rect 7331 31436 7472 31464
rect 7331 31433 7343 31436
rect 7285 31427 7343 31433
rect 7466 31424 7472 31436
rect 7524 31424 7530 31476
rect 13630 31464 13636 31476
rect 12912 31436 13636 31464
rect 11054 31396 11060 31408
rect 10902 31368 11060 31396
rect 11054 31356 11060 31368
rect 11112 31396 11118 31408
rect 11606 31396 11612 31408
rect 11112 31368 11612 31396
rect 11112 31356 11118 31368
rect 11606 31356 11612 31368
rect 11664 31356 11670 31408
rect 12802 31356 12808 31408
rect 12860 31396 12866 31408
rect 12912 31405 12940 31436
rect 13630 31424 13636 31436
rect 13688 31424 13694 31476
rect 15562 31424 15568 31476
rect 15620 31464 15626 31476
rect 16301 31467 16359 31473
rect 16301 31464 16313 31467
rect 15620 31436 16313 31464
rect 15620 31424 15626 31436
rect 16301 31433 16313 31436
rect 16347 31433 16359 31467
rect 16301 31427 16359 31433
rect 16390 31424 16396 31476
rect 16448 31464 16454 31476
rect 16853 31467 16911 31473
rect 16853 31464 16865 31467
rect 16448 31436 16865 31464
rect 16448 31424 16454 31436
rect 16853 31433 16865 31436
rect 16899 31433 16911 31467
rect 16853 31427 16911 31433
rect 17313 31467 17371 31473
rect 17313 31433 17325 31467
rect 17359 31464 17371 31467
rect 19794 31464 19800 31476
rect 17359 31436 19800 31464
rect 17359 31433 17371 31436
rect 17313 31427 17371 31433
rect 19794 31424 19800 31436
rect 19852 31424 19858 31476
rect 19978 31424 19984 31476
rect 20036 31424 20042 31476
rect 20162 31424 20168 31476
rect 20220 31464 20226 31476
rect 22186 31464 22192 31476
rect 20220 31436 22192 31464
rect 20220 31424 20226 31436
rect 22186 31424 22192 31436
rect 22244 31464 22250 31476
rect 22554 31464 22560 31476
rect 22244 31436 22560 31464
rect 22244 31424 22250 31436
rect 22554 31424 22560 31436
rect 22612 31424 22618 31476
rect 23842 31424 23848 31476
rect 23900 31464 23906 31476
rect 25133 31467 25191 31473
rect 25133 31464 25145 31467
rect 23900 31436 25145 31464
rect 23900 31424 23906 31436
rect 25133 31433 25145 31436
rect 25179 31433 25191 31467
rect 25133 31427 25191 31433
rect 12897 31399 12955 31405
rect 12897 31396 12909 31399
rect 12860 31368 12909 31396
rect 12860 31356 12866 31368
rect 12897 31365 12909 31368
rect 12943 31365 12955 31399
rect 12897 31359 12955 31365
rect 18601 31399 18659 31405
rect 18601 31365 18613 31399
rect 18647 31396 18659 31399
rect 19702 31396 19708 31408
rect 18647 31368 19708 31396
rect 18647 31365 18659 31368
rect 18601 31359 18659 31365
rect 19702 31356 19708 31368
rect 19760 31356 19766 31408
rect 19889 31399 19947 31405
rect 19889 31365 19901 31399
rect 19935 31396 19947 31399
rect 21634 31396 21640 31408
rect 19935 31368 21640 31396
rect 19935 31365 19947 31368
rect 19889 31359 19947 31365
rect 21634 31356 21640 31368
rect 21692 31356 21698 31408
rect 22094 31356 22100 31408
rect 22152 31396 22158 31408
rect 22373 31399 22431 31405
rect 22373 31396 22385 31399
rect 22152 31368 22385 31396
rect 22152 31356 22158 31368
rect 22373 31365 22385 31368
rect 22419 31365 22431 31399
rect 22373 31359 22431 31365
rect 3602 31288 3608 31340
rect 3660 31288 3666 31340
rect 7653 31331 7711 31337
rect 7653 31297 7665 31331
rect 7699 31328 7711 31331
rect 8481 31331 8539 31337
rect 8481 31328 8493 31331
rect 7699 31300 8493 31328
rect 7699 31297 7711 31300
rect 7653 31291 7711 31297
rect 8481 31297 8493 31300
rect 8527 31297 8539 31331
rect 8481 31291 8539 31297
rect 9398 31288 9404 31340
rect 9456 31288 9462 31340
rect 15657 31331 15715 31337
rect 14030 31314 14780 31328
rect 14016 31300 14780 31314
rect 3786 31220 3792 31272
rect 3844 31220 3850 31272
rect 4982 31220 4988 31272
rect 5040 31220 5046 31272
rect 6730 31220 6736 31272
rect 6788 31260 6794 31272
rect 6825 31263 6883 31269
rect 6825 31260 6837 31263
rect 6788 31232 6837 31260
rect 6788 31220 6794 31232
rect 6825 31229 6837 31232
rect 6871 31260 6883 31263
rect 7558 31260 7564 31272
rect 6871 31232 7564 31260
rect 6871 31229 6883 31232
rect 6825 31223 6883 31229
rect 7558 31220 7564 31232
rect 7616 31260 7622 31272
rect 7745 31263 7803 31269
rect 7745 31260 7757 31263
rect 7616 31232 7757 31260
rect 7616 31220 7622 31232
rect 7745 31229 7757 31232
rect 7791 31229 7803 31263
rect 7745 31223 7803 31229
rect 7926 31220 7932 31272
rect 7984 31220 7990 31272
rect 9677 31263 9735 31269
rect 9677 31229 9689 31263
rect 9723 31260 9735 31263
rect 10962 31260 10968 31272
rect 9723 31232 10968 31260
rect 9723 31229 9735 31232
rect 9677 31223 9735 31229
rect 10962 31220 10968 31232
rect 11020 31220 11026 31272
rect 12618 31220 12624 31272
rect 12676 31220 12682 31272
rect 7009 31195 7067 31201
rect 7009 31161 7021 31195
rect 7055 31192 7067 31195
rect 7190 31192 7196 31204
rect 7055 31164 7196 31192
rect 7055 31161 7067 31164
rect 7009 31155 7067 31161
rect 7190 31152 7196 31164
rect 7248 31192 7254 31204
rect 7944 31192 7972 31220
rect 7248 31164 7972 31192
rect 11149 31195 11207 31201
rect 7248 31152 7254 31164
rect 11149 31161 11161 31195
rect 11195 31192 11207 31195
rect 12434 31192 12440 31204
rect 11195 31164 12440 31192
rect 11195 31161 11207 31164
rect 11149 31155 11207 31161
rect 12434 31152 12440 31164
rect 12492 31152 12498 31204
rect 11606 31084 11612 31136
rect 11664 31124 11670 31136
rect 14016 31124 14044 31300
rect 14752 31269 14780 31300
rect 15657 31297 15669 31331
rect 15703 31328 15715 31331
rect 15703 31300 16344 31328
rect 15703 31297 15715 31300
rect 15657 31291 15715 31297
rect 16316 31272 16344 31300
rect 17126 31288 17132 31340
rect 17184 31328 17190 31340
rect 17221 31331 17279 31337
rect 17221 31328 17233 31331
rect 17184 31300 17233 31328
rect 17184 31288 17190 31300
rect 17221 31297 17233 31300
rect 17267 31297 17279 31331
rect 17221 31291 17279 31297
rect 18509 31331 18567 31337
rect 18509 31297 18521 31331
rect 18555 31328 18567 31331
rect 20438 31328 20444 31340
rect 18555 31300 20444 31328
rect 18555 31297 18567 31300
rect 18509 31291 18567 31297
rect 20438 31288 20444 31300
rect 20496 31288 20502 31340
rect 23842 31328 23848 31340
rect 23506 31300 23848 31328
rect 23842 31288 23848 31300
rect 23900 31288 23906 31340
rect 24486 31288 24492 31340
rect 24544 31288 24550 31340
rect 25314 31288 25320 31340
rect 25372 31288 25378 31340
rect 14737 31263 14795 31269
rect 14737 31229 14749 31263
rect 14783 31260 14795 31263
rect 15562 31260 15568 31272
rect 14783 31232 15568 31260
rect 14783 31229 14795 31232
rect 14737 31223 14795 31229
rect 15562 31220 15568 31232
rect 15620 31220 15626 31272
rect 16298 31220 16304 31272
rect 16356 31220 16362 31272
rect 17034 31220 17040 31272
rect 17092 31260 17098 31272
rect 17405 31263 17463 31269
rect 17405 31260 17417 31263
rect 17092 31232 17417 31260
rect 17092 31220 17098 31232
rect 17405 31229 17417 31232
rect 17451 31229 17463 31263
rect 17405 31223 17463 31229
rect 18693 31263 18751 31269
rect 18693 31229 18705 31263
rect 18739 31229 18751 31263
rect 18693 31223 18751 31229
rect 14918 31152 14924 31204
rect 14976 31192 14982 31204
rect 18141 31195 18199 31201
rect 18141 31192 18153 31195
rect 14976 31164 18153 31192
rect 14976 31152 14982 31164
rect 18141 31161 18153 31164
rect 18187 31161 18199 31195
rect 18141 31155 18199 31161
rect 11664 31096 14044 31124
rect 11664 31084 11670 31096
rect 14090 31084 14096 31136
rect 14148 31124 14154 31136
rect 14366 31124 14372 31136
rect 14148 31096 14372 31124
rect 14148 31084 14154 31096
rect 14366 31084 14372 31096
rect 14424 31084 14430 31136
rect 15010 31084 15016 31136
rect 15068 31124 15074 31136
rect 18708 31124 18736 31223
rect 20070 31220 20076 31272
rect 20128 31220 20134 31272
rect 22097 31263 22155 31269
rect 22097 31229 22109 31263
rect 22143 31260 22155 31263
rect 22143 31232 22232 31260
rect 22143 31229 22155 31232
rect 22097 31223 22155 31229
rect 15068 31096 18736 31124
rect 15068 31084 15074 31096
rect 19518 31084 19524 31136
rect 19576 31084 19582 31136
rect 22204 31124 22232 31232
rect 23382 31124 23388 31136
rect 22204 31096 23388 31124
rect 23382 31084 23388 31096
rect 23440 31084 23446 31136
rect 23658 31084 23664 31136
rect 23716 31124 23722 31136
rect 23845 31127 23903 31133
rect 23845 31124 23857 31127
rect 23716 31096 23857 31124
rect 23716 31084 23722 31096
rect 23845 31093 23857 31096
rect 23891 31093 23903 31127
rect 23845 31087 23903 31093
rect 24302 31084 24308 31136
rect 24360 31084 24366 31136
rect 24857 31127 24915 31133
rect 24857 31093 24869 31127
rect 24903 31124 24915 31127
rect 24946 31124 24952 31136
rect 24903 31096 24952 31124
rect 24903 31093 24915 31096
rect 24857 31087 24915 31093
rect 24946 31084 24952 31096
rect 25004 31084 25010 31136
rect 1104 31034 25852 31056
rect 1104 30982 2950 31034
rect 3002 30982 3014 31034
rect 3066 30982 3078 31034
rect 3130 30982 3142 31034
rect 3194 30982 3206 31034
rect 3258 30982 12950 31034
rect 13002 30982 13014 31034
rect 13066 30982 13078 31034
rect 13130 30982 13142 31034
rect 13194 30982 13206 31034
rect 13258 30982 22950 31034
rect 23002 30982 23014 31034
rect 23066 30982 23078 31034
rect 23130 30982 23142 31034
rect 23194 30982 23206 31034
rect 23258 30982 25852 31034
rect 1104 30960 25852 30982
rect 7282 30880 7288 30932
rect 7340 30920 7346 30932
rect 7745 30923 7803 30929
rect 7745 30920 7757 30923
rect 7340 30892 7757 30920
rect 7340 30880 7346 30892
rect 7745 30889 7757 30892
rect 7791 30889 7803 30923
rect 7745 30883 7803 30889
rect 8662 30880 8668 30932
rect 8720 30920 8726 30932
rect 8941 30923 8999 30929
rect 8941 30920 8953 30923
rect 8720 30892 8953 30920
rect 8720 30880 8726 30892
rect 8941 30889 8953 30892
rect 8987 30889 8999 30923
rect 8941 30883 8999 30889
rect 10502 30880 10508 30932
rect 10560 30920 10566 30932
rect 12529 30923 12587 30929
rect 12529 30920 12541 30923
rect 10560 30892 12541 30920
rect 10560 30880 10566 30892
rect 12529 30889 12541 30892
rect 12575 30889 12587 30923
rect 12529 30883 12587 30889
rect 15565 30923 15623 30929
rect 15565 30889 15577 30923
rect 15611 30920 15623 30923
rect 15746 30920 15752 30932
rect 15611 30892 15752 30920
rect 15611 30889 15623 30892
rect 15565 30883 15623 30889
rect 8389 30787 8447 30793
rect 8389 30753 8401 30787
rect 8435 30784 8447 30787
rect 8680 30784 8708 30880
rect 10870 30812 10876 30864
rect 10928 30852 10934 30864
rect 10928 30824 14872 30852
rect 10928 30812 10934 30824
rect 8435 30756 8708 30784
rect 8435 30753 8447 30756
rect 8389 30747 8447 30753
rect 11974 30744 11980 30796
rect 12032 30744 12038 30796
rect 14844 30793 14872 30824
rect 13081 30787 13139 30793
rect 13081 30753 13093 30787
rect 13127 30753 13139 30787
rect 13081 30747 13139 30753
rect 14829 30787 14887 30793
rect 14829 30753 14841 30787
rect 14875 30753 14887 30787
rect 14829 30747 14887 30753
rect 7926 30676 7932 30728
rect 7984 30716 7990 30728
rect 9677 30719 9735 30725
rect 7984 30688 8432 30716
rect 7984 30676 7990 30688
rect 8113 30651 8171 30657
rect 8113 30617 8125 30651
rect 8159 30648 8171 30651
rect 8294 30648 8300 30660
rect 8159 30620 8300 30648
rect 8159 30617 8171 30620
rect 8113 30611 8171 30617
rect 8294 30608 8300 30620
rect 8352 30608 8358 30660
rect 8404 30648 8432 30688
rect 9677 30685 9689 30719
rect 9723 30716 9735 30719
rect 12434 30716 12440 30728
rect 9723 30688 12440 30716
rect 9723 30685 9735 30688
rect 9677 30679 9735 30685
rect 12434 30676 12440 30688
rect 12492 30716 12498 30728
rect 12986 30716 12992 30728
rect 12492 30688 12992 30716
rect 12492 30676 12498 30688
rect 12986 30676 12992 30688
rect 13044 30676 13050 30728
rect 12253 30651 12311 30657
rect 12253 30648 12265 30651
rect 8404 30620 12265 30648
rect 12253 30617 12265 30620
rect 12299 30648 12311 30651
rect 13096 30648 13124 30747
rect 13998 30676 14004 30728
rect 14056 30716 14062 30728
rect 14274 30716 14280 30728
rect 14056 30688 14280 30716
rect 14056 30676 14062 30688
rect 14274 30676 14280 30688
rect 14332 30676 14338 30728
rect 14645 30719 14703 30725
rect 14645 30685 14657 30719
rect 14691 30716 14703 30719
rect 15580 30716 15608 30883
rect 15746 30880 15752 30892
rect 15804 30880 15810 30932
rect 15930 30880 15936 30932
rect 15988 30920 15994 30932
rect 19794 30920 19800 30932
rect 15988 30892 19800 30920
rect 15988 30880 15994 30892
rect 19794 30880 19800 30892
rect 19852 30880 19858 30932
rect 22738 30880 22744 30932
rect 22796 30920 22802 30932
rect 22833 30923 22891 30929
rect 22833 30920 22845 30923
rect 22796 30892 22845 30920
rect 22796 30880 22802 30892
rect 22833 30889 22845 30892
rect 22879 30889 22891 30923
rect 22833 30883 22891 30889
rect 24857 30923 24915 30929
rect 24857 30889 24869 30923
rect 24903 30920 24915 30923
rect 25314 30920 25320 30932
rect 24903 30892 25320 30920
rect 24903 30889 24915 30892
rect 24857 30883 24915 30889
rect 25314 30880 25320 30892
rect 25372 30880 25378 30932
rect 19429 30855 19487 30861
rect 16040 30824 17264 30852
rect 16040 30725 16068 30824
rect 16482 30744 16488 30796
rect 16540 30784 16546 30796
rect 17129 30787 17187 30793
rect 17129 30784 17141 30787
rect 16540 30756 17141 30784
rect 16540 30744 16546 30756
rect 17129 30753 17141 30756
rect 17175 30753 17187 30787
rect 17236 30784 17264 30824
rect 19429 30821 19441 30855
rect 19475 30852 19487 30855
rect 20714 30852 20720 30864
rect 19475 30824 20720 30852
rect 19475 30821 19487 30824
rect 19429 30815 19487 30821
rect 20714 30812 20720 30824
rect 20772 30812 20778 30864
rect 21821 30855 21879 30861
rect 21821 30821 21833 30855
rect 21867 30852 21879 30855
rect 22186 30852 22192 30864
rect 21867 30824 22192 30852
rect 21867 30821 21879 30824
rect 21821 30815 21879 30821
rect 22186 30812 22192 30824
rect 22244 30812 22250 30864
rect 22756 30852 22784 30880
rect 22296 30824 22784 30852
rect 17770 30784 17776 30796
rect 17236 30756 17776 30784
rect 17129 30747 17187 30753
rect 17770 30744 17776 30756
rect 17828 30784 17834 30796
rect 18877 30787 18935 30793
rect 18877 30784 18889 30787
rect 17828 30756 18889 30784
rect 17828 30744 17834 30756
rect 18877 30753 18889 30756
rect 18923 30753 18935 30787
rect 18877 30747 18935 30753
rect 20073 30787 20131 30793
rect 20073 30753 20085 30787
rect 20119 30784 20131 30787
rect 20162 30784 20168 30796
rect 20119 30756 20168 30784
rect 20119 30753 20131 30756
rect 20073 30747 20131 30753
rect 20162 30744 20168 30756
rect 20220 30744 20226 30796
rect 22296 30793 22324 30824
rect 22281 30787 22339 30793
rect 22281 30753 22293 30787
rect 22327 30753 22339 30787
rect 22281 30747 22339 30753
rect 22465 30787 22523 30793
rect 22465 30753 22477 30787
rect 22511 30784 22523 30787
rect 22738 30784 22744 30796
rect 22511 30756 22744 30784
rect 22511 30753 22523 30756
rect 22465 30747 22523 30753
rect 22738 30744 22744 30756
rect 22796 30744 22802 30796
rect 25130 30784 25136 30796
rect 22848 30756 25136 30784
rect 14691 30688 15608 30716
rect 16025 30719 16083 30725
rect 14691 30685 14703 30688
rect 14645 30679 14703 30685
rect 16025 30685 16037 30719
rect 16071 30685 16083 30719
rect 16025 30679 16083 30685
rect 19702 30676 19708 30728
rect 19760 30716 19766 30728
rect 22189 30719 22247 30725
rect 22189 30716 22201 30719
rect 19760 30688 22201 30716
rect 19760 30676 19766 30688
rect 22189 30685 22201 30688
rect 22235 30716 22247 30719
rect 22848 30716 22876 30756
rect 25130 30744 25136 30756
rect 25188 30744 25194 30796
rect 22235 30688 22876 30716
rect 22235 30685 22247 30688
rect 22189 30679 22247 30685
rect 23934 30676 23940 30728
rect 23992 30676 23998 30728
rect 25317 30719 25375 30725
rect 25317 30685 25329 30719
rect 25363 30716 25375 30719
rect 25498 30716 25504 30728
rect 25363 30688 25504 30716
rect 25363 30685 25375 30688
rect 25317 30679 25375 30685
rect 25498 30676 25504 30688
rect 25556 30676 25562 30728
rect 16206 30648 16212 30660
rect 12299 30620 13124 30648
rect 13740 30620 16212 30648
rect 12299 30617 12311 30620
rect 12253 30611 12311 30617
rect 5258 30540 5264 30592
rect 5316 30580 5322 30592
rect 7466 30580 7472 30592
rect 5316 30552 7472 30580
rect 5316 30540 5322 30552
rect 7466 30540 7472 30552
rect 7524 30580 7530 30592
rect 8205 30583 8263 30589
rect 8205 30580 8217 30583
rect 7524 30552 8217 30580
rect 7524 30540 7530 30552
rect 8205 30549 8217 30552
rect 8251 30549 8263 30583
rect 8205 30543 8263 30549
rect 9950 30540 9956 30592
rect 10008 30580 10014 30592
rect 10321 30583 10379 30589
rect 10321 30580 10333 30583
rect 10008 30552 10333 30580
rect 10008 30540 10014 30552
rect 10321 30549 10333 30552
rect 10367 30549 10379 30583
rect 10321 30543 10379 30549
rect 11974 30540 11980 30592
rect 12032 30580 12038 30592
rect 12897 30583 12955 30589
rect 12897 30580 12909 30583
rect 12032 30552 12909 30580
rect 12032 30540 12038 30552
rect 12897 30549 12909 30552
rect 12943 30549 12955 30583
rect 12897 30543 12955 30549
rect 12989 30583 13047 30589
rect 12989 30549 13001 30583
rect 13035 30580 13047 30583
rect 13740 30580 13768 30620
rect 16206 30608 16212 30620
rect 16264 30608 16270 30660
rect 17402 30608 17408 30660
rect 17460 30608 17466 30660
rect 18782 30648 18788 30660
rect 18630 30620 18788 30648
rect 13035 30552 13768 30580
rect 13035 30549 13047 30552
rect 12989 30543 13047 30549
rect 13998 30540 14004 30592
rect 14056 30580 14062 30592
rect 14277 30583 14335 30589
rect 14277 30580 14289 30583
rect 14056 30552 14289 30580
rect 14056 30540 14062 30552
rect 14277 30549 14289 30552
rect 14323 30549 14335 30583
rect 14277 30543 14335 30549
rect 14737 30583 14795 30589
rect 14737 30549 14749 30583
rect 14783 30580 14795 30583
rect 15378 30580 15384 30592
rect 14783 30552 15384 30580
rect 14783 30549 14795 30552
rect 14737 30543 14795 30549
rect 15378 30540 15384 30552
rect 15436 30540 15442 30592
rect 15562 30540 15568 30592
rect 15620 30580 15626 30592
rect 16669 30583 16727 30589
rect 16669 30580 16681 30583
rect 15620 30552 16681 30580
rect 15620 30540 15626 30552
rect 16669 30549 16681 30552
rect 16715 30549 16727 30583
rect 16669 30543 16727 30549
rect 18322 30540 18328 30592
rect 18380 30580 18386 30592
rect 18708 30580 18736 30620
rect 18782 30608 18788 30620
rect 18840 30608 18846 30660
rect 19797 30651 19855 30657
rect 19797 30617 19809 30651
rect 19843 30648 19855 30651
rect 20162 30648 20168 30660
rect 19843 30620 20168 30648
rect 19843 30617 19855 30620
rect 19797 30611 19855 30617
rect 20162 30608 20168 30620
rect 20220 30608 20226 30660
rect 18380 30552 18736 30580
rect 18380 30540 18386 30552
rect 19886 30540 19892 30592
rect 19944 30580 19950 30592
rect 20441 30583 20499 30589
rect 20441 30580 20453 30583
rect 19944 30552 20453 30580
rect 19944 30540 19950 30552
rect 20441 30549 20453 30552
rect 20487 30549 20499 30583
rect 20441 30543 20499 30549
rect 23753 30583 23811 30589
rect 23753 30549 23765 30583
rect 23799 30580 23811 30583
rect 24486 30580 24492 30592
rect 23799 30552 24492 30580
rect 23799 30549 23811 30552
rect 23753 30543 23811 30549
rect 24486 30540 24492 30552
rect 24544 30540 24550 30592
rect 25130 30540 25136 30592
rect 25188 30540 25194 30592
rect 1104 30490 25852 30512
rect 1104 30438 7950 30490
rect 8002 30438 8014 30490
rect 8066 30438 8078 30490
rect 8130 30438 8142 30490
rect 8194 30438 8206 30490
rect 8258 30438 17950 30490
rect 18002 30438 18014 30490
rect 18066 30438 18078 30490
rect 18130 30438 18142 30490
rect 18194 30438 18206 30490
rect 18258 30438 25852 30490
rect 1104 30416 25852 30438
rect 15654 30336 15660 30388
rect 15712 30376 15718 30388
rect 18322 30376 18328 30388
rect 15712 30348 16160 30376
rect 15712 30336 15718 30348
rect 10870 30308 10876 30320
rect 8864 30280 10876 30308
rect 8864 30249 8892 30280
rect 10870 30268 10876 30280
rect 10928 30268 10934 30320
rect 12618 30268 12624 30320
rect 12676 30308 12682 30320
rect 13722 30308 13728 30320
rect 12676 30280 13728 30308
rect 12676 30268 12682 30280
rect 13722 30268 13728 30280
rect 13780 30308 13786 30320
rect 16132 30308 16160 30348
rect 17696 30348 18328 30376
rect 16761 30311 16819 30317
rect 16761 30308 16773 30311
rect 13780 30280 14596 30308
rect 16054 30280 16773 30308
rect 13780 30268 13786 30280
rect 14568 30249 14596 30280
rect 16761 30277 16773 30280
rect 16807 30308 16819 30311
rect 17696 30308 17724 30348
rect 18322 30336 18328 30348
rect 18380 30336 18386 30388
rect 18690 30336 18696 30388
rect 18748 30376 18754 30388
rect 19426 30376 19432 30388
rect 18748 30348 19432 30376
rect 18748 30336 18754 30348
rect 19426 30336 19432 30348
rect 19484 30336 19490 30388
rect 19886 30336 19892 30388
rect 19944 30376 19950 30388
rect 21358 30376 21364 30388
rect 19944 30348 21364 30376
rect 19944 30336 19950 30348
rect 21358 30336 21364 30348
rect 21416 30336 21422 30388
rect 24946 30376 24952 30388
rect 24044 30348 24952 30376
rect 16807 30280 17724 30308
rect 16807 30277 16819 30280
rect 16761 30271 16819 30277
rect 18782 30268 18788 30320
rect 18840 30308 18846 30320
rect 18969 30311 19027 30317
rect 18969 30308 18981 30311
rect 18840 30280 18981 30308
rect 18840 30268 18846 30280
rect 18969 30277 18981 30280
rect 19015 30277 19027 30311
rect 18969 30271 19027 30277
rect 23658 30268 23664 30320
rect 23716 30268 23722 30320
rect 23934 30268 23940 30320
rect 23992 30308 23998 30320
rect 24044 30308 24072 30348
rect 24946 30336 24952 30348
rect 25004 30376 25010 30388
rect 25409 30379 25467 30385
rect 25409 30376 25421 30379
rect 25004 30348 25421 30376
rect 25004 30336 25010 30348
rect 25409 30345 25421 30348
rect 25455 30345 25467 30379
rect 25409 30339 25467 30345
rect 23992 30280 24150 30308
rect 23992 30268 23998 30280
rect 8849 30243 8907 30249
rect 8849 30209 8861 30243
rect 8895 30209 8907 30243
rect 8849 30203 8907 30209
rect 10781 30243 10839 30249
rect 10781 30209 10793 30243
rect 10827 30240 10839 30243
rect 11701 30243 11759 30249
rect 11701 30240 11713 30243
rect 10827 30212 11713 30240
rect 10827 30209 10839 30212
rect 10781 30203 10839 30209
rect 11701 30209 11713 30212
rect 11747 30209 11759 30243
rect 12897 30243 12955 30249
rect 12897 30240 12909 30243
rect 11701 30203 11759 30209
rect 12406 30212 12909 30240
rect 10137 30175 10195 30181
rect 10137 30141 10149 30175
rect 10183 30172 10195 30175
rect 10318 30172 10324 30184
rect 10183 30144 10324 30172
rect 10183 30141 10195 30144
rect 10137 30135 10195 30141
rect 10318 30132 10324 30144
rect 10376 30172 10382 30184
rect 10873 30175 10931 30181
rect 10873 30172 10885 30175
rect 10376 30144 10885 30172
rect 10376 30132 10382 30144
rect 10873 30141 10885 30144
rect 10919 30141 10931 30175
rect 10873 30135 10931 30141
rect 10962 30132 10968 30184
rect 11020 30132 11026 30184
rect 10413 30107 10471 30113
rect 10413 30073 10425 30107
rect 10459 30104 10471 30107
rect 12406 30104 12434 30212
rect 12897 30209 12909 30212
rect 12943 30209 12955 30243
rect 12897 30203 12955 30209
rect 14553 30243 14611 30249
rect 14553 30209 14565 30243
rect 14599 30209 14611 30243
rect 14553 30203 14611 30209
rect 17773 30243 17831 30249
rect 17773 30209 17785 30243
rect 17819 30209 17831 30243
rect 17773 30203 17831 30209
rect 12710 30132 12716 30184
rect 12768 30172 12774 30184
rect 12989 30175 13047 30181
rect 12989 30172 13001 30175
rect 12768 30144 13001 30172
rect 12768 30132 12774 30144
rect 12989 30141 13001 30144
rect 13035 30141 13047 30175
rect 12989 30135 13047 30141
rect 13078 30132 13084 30184
rect 13136 30132 13142 30184
rect 14829 30175 14887 30181
rect 14829 30141 14841 30175
rect 14875 30172 14887 30175
rect 15562 30172 15568 30184
rect 14875 30144 15568 30172
rect 14875 30141 14887 30144
rect 14829 30135 14887 30141
rect 15562 30132 15568 30144
rect 15620 30132 15626 30184
rect 17037 30107 17095 30113
rect 17037 30104 17049 30107
rect 10459 30076 12434 30104
rect 15856 30076 17049 30104
rect 10459 30073 10471 30076
rect 10413 30067 10471 30073
rect 8294 29996 8300 30048
rect 8352 30036 8358 30048
rect 9493 30039 9551 30045
rect 9493 30036 9505 30039
rect 8352 30008 9505 30036
rect 8352 29996 8358 30008
rect 9493 30005 9505 30008
rect 9539 30005 9551 30039
rect 9493 29999 9551 30005
rect 12529 30039 12587 30045
rect 12529 30005 12541 30039
rect 12575 30036 12587 30039
rect 12710 30036 12716 30048
rect 12575 30008 12716 30036
rect 12575 30005 12587 30008
rect 12529 29999 12587 30005
rect 12710 29996 12716 30008
rect 12768 29996 12774 30048
rect 14550 29996 14556 30048
rect 14608 30036 14614 30048
rect 15856 30036 15884 30076
rect 17037 30073 17049 30076
rect 17083 30104 17095 30107
rect 17788 30104 17816 30203
rect 19794 30200 19800 30252
rect 19852 30200 19858 30252
rect 23382 30200 23388 30252
rect 23440 30200 23446 30252
rect 17865 30175 17923 30181
rect 17865 30141 17877 30175
rect 17911 30141 17923 30175
rect 17865 30135 17923 30141
rect 18049 30175 18107 30181
rect 18049 30141 18061 30175
rect 18095 30172 18107 30175
rect 20898 30172 20904 30184
rect 18095 30144 20904 30172
rect 18095 30141 18107 30144
rect 18049 30135 18107 30141
rect 17083 30076 17816 30104
rect 17880 30104 17908 30135
rect 20898 30132 20904 30144
rect 20956 30132 20962 30184
rect 25406 30172 25412 30184
rect 22066 30144 25412 30172
rect 19337 30107 19395 30113
rect 17880 30076 18552 30104
rect 17083 30073 17095 30076
rect 17037 30067 17095 30073
rect 14608 30008 15884 30036
rect 14608 29996 14614 30008
rect 16298 29996 16304 30048
rect 16356 29996 16362 30048
rect 17405 30039 17463 30045
rect 17405 30005 17417 30039
rect 17451 30036 17463 30039
rect 18322 30036 18328 30048
rect 17451 30008 18328 30036
rect 17451 30005 17463 30008
rect 17405 29999 17463 30005
rect 18322 29996 18328 30008
rect 18380 29996 18386 30048
rect 18524 30045 18552 30076
rect 19337 30073 19349 30107
rect 19383 30104 19395 30107
rect 19794 30104 19800 30116
rect 19383 30076 19800 30104
rect 19383 30073 19395 30076
rect 19337 30067 19395 30073
rect 19794 30064 19800 30076
rect 19852 30104 19858 30116
rect 20162 30104 20168 30116
rect 19852 30076 20168 30104
rect 19852 30064 19858 30076
rect 20162 30064 20168 30076
rect 20220 30064 20226 30116
rect 18509 30039 18567 30045
rect 18509 30005 18521 30039
rect 18555 30036 18567 30039
rect 18690 30036 18696 30048
rect 18555 30008 18696 30036
rect 18555 30005 18567 30008
rect 18509 29999 18567 30005
rect 18690 29996 18696 30008
rect 18748 29996 18754 30048
rect 19613 30039 19671 30045
rect 19613 30005 19625 30039
rect 19659 30036 19671 30039
rect 22066 30036 22094 30144
rect 25406 30132 25412 30144
rect 25464 30132 25470 30184
rect 19659 30008 22094 30036
rect 19659 30005 19671 30008
rect 19613 29999 19671 30005
rect 22646 29996 22652 30048
rect 22704 30036 22710 30048
rect 23382 30036 23388 30048
rect 22704 30008 23388 30036
rect 22704 29996 22710 30008
rect 23382 29996 23388 30008
rect 23440 30036 23446 30048
rect 25133 30039 25191 30045
rect 25133 30036 25145 30039
rect 23440 30008 25145 30036
rect 23440 29996 23446 30008
rect 25133 30005 25145 30008
rect 25179 30005 25191 30039
rect 25133 29999 25191 30005
rect 1104 29946 25852 29968
rect 1104 29894 2950 29946
rect 3002 29894 3014 29946
rect 3066 29894 3078 29946
rect 3130 29894 3142 29946
rect 3194 29894 3206 29946
rect 3258 29894 12950 29946
rect 13002 29894 13014 29946
rect 13066 29894 13078 29946
rect 13130 29894 13142 29946
rect 13194 29894 13206 29946
rect 13258 29894 22950 29946
rect 23002 29894 23014 29946
rect 23066 29894 23078 29946
rect 23130 29894 23142 29946
rect 23194 29894 23206 29946
rect 23258 29894 25852 29946
rect 1104 29872 25852 29894
rect 15838 29792 15844 29844
rect 15896 29832 15902 29844
rect 15933 29835 15991 29841
rect 15933 29832 15945 29835
rect 15896 29804 15945 29832
rect 15896 29792 15902 29804
rect 15933 29801 15945 29804
rect 15979 29801 15991 29835
rect 15933 29795 15991 29801
rect 16206 29792 16212 29844
rect 16264 29832 16270 29844
rect 23934 29832 23940 29844
rect 16264 29804 23940 29832
rect 16264 29792 16270 29804
rect 23934 29792 23940 29804
rect 23992 29792 23998 29844
rect 15562 29724 15568 29776
rect 15620 29764 15626 29776
rect 16224 29764 16252 29792
rect 16390 29764 16396 29776
rect 15620 29736 16252 29764
rect 16316 29736 16396 29764
rect 15620 29724 15626 29736
rect 3878 29656 3884 29708
rect 3936 29696 3942 29708
rect 3973 29699 4031 29705
rect 3973 29696 3985 29699
rect 3936 29668 3985 29696
rect 3936 29656 3942 29668
rect 3973 29665 3985 29668
rect 4019 29665 4031 29699
rect 3973 29659 4031 29665
rect 9674 29656 9680 29708
rect 9732 29656 9738 29708
rect 9950 29656 9956 29708
rect 10008 29656 10014 29708
rect 10502 29656 10508 29708
rect 10560 29696 10566 29708
rect 12529 29699 12587 29705
rect 12529 29696 12541 29699
rect 10560 29668 12541 29696
rect 10560 29656 10566 29668
rect 12529 29665 12541 29668
rect 12575 29665 12587 29699
rect 12529 29659 12587 29665
rect 15654 29656 15660 29708
rect 15712 29696 15718 29708
rect 16316 29696 16344 29736
rect 16390 29724 16396 29736
rect 16448 29764 16454 29776
rect 19886 29764 19892 29776
rect 16448 29736 19892 29764
rect 16448 29724 16454 29736
rect 19886 29724 19892 29736
rect 19944 29724 19950 29776
rect 20070 29724 20076 29776
rect 20128 29764 20134 29776
rect 25133 29767 25191 29773
rect 25133 29764 25145 29767
rect 20128 29736 25145 29764
rect 20128 29724 20134 29736
rect 25133 29733 25145 29736
rect 25179 29733 25191 29767
rect 25133 29727 25191 29733
rect 15712 29668 16344 29696
rect 17681 29699 17739 29705
rect 15712 29656 15718 29668
rect 17681 29665 17693 29699
rect 17727 29696 17739 29699
rect 17770 29696 17776 29708
rect 17727 29668 17776 29696
rect 17727 29665 17739 29668
rect 17681 29659 17739 29665
rect 17770 29656 17776 29668
rect 17828 29656 17834 29708
rect 18322 29656 18328 29708
rect 18380 29696 18386 29708
rect 19981 29699 20039 29705
rect 19981 29696 19993 29699
rect 18380 29668 19993 29696
rect 18380 29656 18386 29668
rect 19981 29665 19993 29668
rect 20027 29665 20039 29699
rect 19981 29659 20039 29665
rect 20165 29699 20223 29705
rect 20165 29665 20177 29699
rect 20211 29696 20223 29699
rect 20898 29696 20904 29708
rect 20211 29668 20904 29696
rect 20211 29665 20223 29668
rect 20165 29659 20223 29665
rect 20898 29656 20904 29668
rect 20956 29656 20962 29708
rect 23290 29656 23296 29708
rect 23348 29656 23354 29708
rect 23382 29656 23388 29708
rect 23440 29656 23446 29708
rect 11054 29588 11060 29640
rect 11112 29588 11118 29640
rect 11885 29631 11943 29637
rect 11885 29628 11897 29631
rect 11440 29600 11897 29628
rect 3878 29520 3884 29572
rect 3936 29560 3942 29572
rect 4157 29563 4215 29569
rect 4157 29560 4169 29563
rect 3936 29532 4169 29560
rect 3936 29520 3942 29532
rect 4157 29529 4169 29532
rect 4203 29529 4215 29563
rect 4157 29523 4215 29529
rect 5813 29563 5871 29569
rect 5813 29529 5825 29563
rect 5859 29560 5871 29563
rect 6178 29560 6184 29572
rect 5859 29532 6184 29560
rect 5859 29529 5871 29532
rect 5813 29523 5871 29529
rect 6178 29520 6184 29532
rect 6236 29520 6242 29572
rect 11440 29504 11468 29600
rect 11885 29597 11897 29600
rect 11931 29597 11943 29631
rect 11885 29591 11943 29597
rect 16666 29588 16672 29640
rect 16724 29628 16730 29640
rect 17310 29628 17316 29640
rect 16724 29600 17316 29628
rect 16724 29588 16730 29600
rect 17310 29588 17316 29600
rect 17368 29588 17374 29640
rect 17494 29588 17500 29640
rect 17552 29628 17558 29640
rect 19889 29631 19947 29637
rect 17552 29600 18368 29628
rect 17552 29588 17558 29600
rect 14645 29563 14703 29569
rect 14645 29529 14657 29563
rect 14691 29560 14703 29563
rect 17405 29563 17463 29569
rect 14691 29532 16804 29560
rect 14691 29529 14703 29532
rect 14645 29523 14703 29529
rect 16776 29504 16804 29532
rect 17405 29529 17417 29563
rect 17451 29560 17463 29563
rect 18233 29563 18291 29569
rect 18233 29560 18245 29563
rect 17451 29532 18245 29560
rect 17451 29529 17463 29532
rect 17405 29523 17463 29529
rect 18233 29529 18245 29532
rect 18279 29529 18291 29563
rect 18340 29560 18368 29600
rect 19889 29597 19901 29631
rect 19935 29628 19947 29631
rect 20622 29628 20628 29640
rect 19935 29600 20628 29628
rect 19935 29597 19947 29600
rect 19889 29591 19947 29597
rect 20622 29588 20628 29600
rect 20680 29588 20686 29640
rect 22554 29588 22560 29640
rect 22612 29628 22618 29640
rect 23201 29631 23259 29637
rect 23201 29628 23213 29631
rect 22612 29600 23213 29628
rect 22612 29588 22618 29600
rect 23201 29597 23213 29600
rect 23247 29597 23259 29631
rect 23201 29591 23259 29597
rect 25314 29588 25320 29640
rect 25372 29588 25378 29640
rect 20254 29560 20260 29572
rect 18340 29532 20260 29560
rect 18233 29523 18291 29529
rect 20254 29520 20260 29532
rect 20312 29520 20318 29572
rect 24762 29560 24768 29572
rect 22848 29532 24768 29560
rect 7282 29452 7288 29504
rect 7340 29492 7346 29504
rect 7469 29495 7527 29501
rect 7469 29492 7481 29495
rect 7340 29464 7481 29492
rect 7340 29452 7346 29464
rect 7469 29461 7481 29464
rect 7515 29461 7527 29495
rect 7469 29455 7527 29461
rect 11422 29452 11428 29504
rect 11480 29452 11486 29504
rect 12250 29452 12256 29504
rect 12308 29492 12314 29504
rect 12897 29495 12955 29501
rect 12897 29492 12909 29495
rect 12308 29464 12909 29492
rect 12308 29452 12314 29464
rect 12897 29461 12909 29464
rect 12943 29492 12955 29495
rect 15286 29492 15292 29504
rect 12943 29464 15292 29492
rect 12943 29461 12955 29464
rect 12897 29455 12955 29461
rect 15286 29452 15292 29464
rect 15344 29452 15350 29504
rect 16758 29452 16764 29504
rect 16816 29452 16822 29504
rect 17034 29452 17040 29504
rect 17092 29452 17098 29504
rect 17494 29452 17500 29504
rect 17552 29452 17558 29504
rect 19521 29495 19579 29501
rect 19521 29461 19533 29495
rect 19567 29492 19579 29495
rect 19794 29492 19800 29504
rect 19567 29464 19800 29492
rect 19567 29461 19579 29464
rect 19521 29455 19579 29461
rect 19794 29452 19800 29464
rect 19852 29452 19858 29504
rect 22848 29501 22876 29532
rect 24762 29520 24768 29532
rect 24820 29520 24826 29572
rect 22833 29495 22891 29501
rect 22833 29461 22845 29495
rect 22879 29461 22891 29495
rect 22833 29455 22891 29461
rect 1104 29402 25852 29424
rect 1104 29350 7950 29402
rect 8002 29350 8014 29402
rect 8066 29350 8078 29402
rect 8130 29350 8142 29402
rect 8194 29350 8206 29402
rect 8258 29350 17950 29402
rect 18002 29350 18014 29402
rect 18066 29350 18078 29402
rect 18130 29350 18142 29402
rect 18194 29350 18206 29402
rect 18258 29350 25852 29402
rect 1104 29328 25852 29350
rect 3375 29291 3433 29297
rect 3375 29257 3387 29291
rect 3421 29288 3433 29291
rect 3786 29288 3792 29300
rect 3421 29260 3792 29288
rect 3421 29257 3433 29260
rect 3375 29251 3433 29257
rect 3786 29248 3792 29260
rect 3844 29248 3850 29300
rect 5074 29248 5080 29300
rect 5132 29288 5138 29300
rect 8938 29288 8944 29300
rect 5132 29260 8944 29288
rect 5132 29248 5138 29260
rect 8938 29248 8944 29260
rect 8996 29288 9002 29300
rect 9214 29288 9220 29300
rect 8996 29260 9220 29288
rect 8996 29248 9002 29260
rect 9214 29248 9220 29260
rect 9272 29248 9278 29300
rect 9766 29248 9772 29300
rect 9824 29248 9830 29300
rect 11054 29248 11060 29300
rect 11112 29288 11118 29300
rect 11517 29291 11575 29297
rect 11517 29288 11529 29291
rect 11112 29260 11529 29288
rect 11112 29248 11118 29260
rect 11517 29257 11529 29260
rect 11563 29257 11575 29291
rect 11517 29251 11575 29257
rect 13909 29291 13967 29297
rect 13909 29257 13921 29291
rect 13955 29288 13967 29291
rect 15194 29288 15200 29300
rect 13955 29260 15200 29288
rect 13955 29257 13967 29260
rect 13909 29251 13967 29257
rect 15194 29248 15200 29260
rect 15252 29248 15258 29300
rect 15933 29291 15991 29297
rect 15933 29257 15945 29291
rect 15979 29288 15991 29291
rect 16942 29288 16948 29300
rect 15979 29260 16948 29288
rect 15979 29257 15991 29260
rect 15933 29251 15991 29257
rect 16942 29248 16948 29260
rect 17000 29248 17006 29300
rect 17221 29291 17279 29297
rect 17221 29257 17233 29291
rect 17267 29288 17279 29291
rect 17310 29288 17316 29300
rect 17267 29260 17316 29288
rect 17267 29257 17279 29260
rect 17221 29251 17279 29257
rect 17310 29248 17316 29260
rect 17368 29248 17374 29300
rect 17494 29248 17500 29300
rect 17552 29288 17558 29300
rect 18049 29291 18107 29297
rect 18049 29288 18061 29291
rect 17552 29260 18061 29288
rect 17552 29248 17558 29260
rect 18049 29257 18061 29260
rect 18095 29257 18107 29291
rect 18049 29251 18107 29257
rect 18414 29248 18420 29300
rect 18472 29248 18478 29300
rect 18509 29291 18567 29297
rect 18509 29257 18521 29291
rect 18555 29288 18567 29291
rect 20070 29288 20076 29300
rect 18555 29260 20076 29288
rect 18555 29257 18567 29260
rect 18509 29251 18567 29257
rect 20070 29248 20076 29260
rect 20128 29248 20134 29300
rect 21818 29288 21824 29300
rect 20180 29260 21824 29288
rect 8570 29180 8576 29232
rect 8628 29220 8634 29232
rect 8628 29192 10824 29220
rect 8628 29180 8634 29192
rect 2222 29112 2228 29164
rect 2280 29152 2286 29164
rect 3272 29155 3330 29161
rect 3272 29152 3284 29155
rect 2280 29124 3284 29152
rect 2280 29112 2286 29124
rect 3272 29121 3284 29124
rect 3318 29121 3330 29155
rect 8662 29152 8668 29164
rect 8418 29124 8668 29152
rect 3272 29115 3330 29121
rect 8662 29112 8668 29124
rect 8720 29112 8726 29164
rect 9214 29112 9220 29164
rect 9272 29152 9278 29164
rect 10137 29155 10195 29161
rect 10137 29152 10149 29155
rect 9272 29124 10149 29152
rect 9272 29112 9278 29124
rect 10137 29121 10149 29124
rect 10183 29121 10195 29155
rect 10137 29115 10195 29121
rect 6454 29044 6460 29096
rect 6512 29084 6518 29096
rect 7009 29087 7067 29093
rect 7009 29084 7021 29087
rect 6512 29056 7021 29084
rect 6512 29044 6518 29056
rect 7009 29053 7021 29056
rect 7055 29053 7067 29087
rect 7009 29047 7067 29053
rect 10229 29087 10287 29093
rect 10229 29053 10241 29087
rect 10275 29053 10287 29087
rect 10229 29047 10287 29053
rect 10413 29087 10471 29093
rect 10413 29053 10425 29087
rect 10459 29084 10471 29087
rect 10686 29084 10692 29096
rect 10459 29056 10692 29084
rect 10459 29053 10471 29056
rect 10413 29047 10471 29053
rect 8754 28976 8760 29028
rect 8812 28976 8818 29028
rect 9493 29019 9551 29025
rect 9493 28985 9505 29019
rect 9539 29016 9551 29019
rect 9674 29016 9680 29028
rect 9539 28988 9680 29016
rect 9539 28985 9551 28988
rect 9493 28979 9551 28985
rect 9674 28976 9680 28988
rect 9732 29016 9738 29028
rect 10134 29016 10140 29028
rect 9732 28988 10140 29016
rect 9732 28976 9738 28988
rect 10134 28976 10140 28988
rect 10192 29016 10198 29028
rect 10244 29016 10272 29047
rect 10686 29044 10692 29056
rect 10744 29044 10750 29096
rect 10796 29084 10824 29192
rect 11330 29180 11336 29232
rect 11388 29220 11394 29232
rect 12250 29220 12256 29232
rect 11388 29192 12256 29220
rect 11388 29180 11394 29192
rect 12250 29180 12256 29192
rect 12308 29220 12314 29232
rect 12437 29223 12495 29229
rect 12437 29220 12449 29223
rect 12308 29192 12449 29220
rect 12308 29180 12314 29192
rect 12437 29189 12449 29192
rect 12483 29189 12495 29223
rect 12437 29183 12495 29189
rect 13081 29223 13139 29229
rect 13081 29189 13093 29223
rect 13127 29220 13139 29223
rect 15654 29220 15660 29232
rect 13127 29192 15660 29220
rect 13127 29189 13139 29192
rect 13081 29183 13139 29189
rect 12345 29155 12403 29161
rect 12345 29121 12357 29155
rect 12391 29152 12403 29155
rect 13096 29152 13124 29183
rect 15654 29180 15660 29192
rect 15712 29180 15718 29232
rect 15841 29223 15899 29229
rect 15841 29189 15853 29223
rect 15887 29220 15899 29223
rect 18432 29220 18460 29248
rect 20180 29220 20208 29260
rect 21818 29248 21824 29260
rect 21876 29248 21882 29300
rect 22002 29248 22008 29300
rect 22060 29288 22066 29300
rect 22373 29291 22431 29297
rect 22373 29288 22385 29291
rect 22060 29260 22385 29288
rect 22060 29248 22066 29260
rect 22373 29257 22385 29260
rect 22419 29257 22431 29291
rect 22373 29251 22431 29257
rect 23934 29248 23940 29300
rect 23992 29248 23998 29300
rect 25314 29248 25320 29300
rect 25372 29248 25378 29300
rect 25498 29248 25504 29300
rect 25556 29248 25562 29300
rect 15887 29192 18460 29220
rect 19306 29192 20208 29220
rect 15887 29189 15899 29192
rect 15841 29183 15899 29189
rect 12391 29124 13124 29152
rect 12391 29121 12403 29124
rect 12345 29115 12403 29121
rect 13354 29112 13360 29164
rect 13412 29152 13418 29164
rect 13817 29155 13875 29161
rect 13817 29152 13829 29155
rect 13412 29124 13829 29152
rect 13412 29112 13418 29124
rect 13817 29121 13829 29124
rect 13863 29121 13875 29155
rect 13817 29115 13875 29121
rect 17313 29155 17371 29161
rect 17313 29121 17325 29155
rect 17359 29152 17371 29155
rect 17678 29152 17684 29164
rect 17359 29124 17684 29152
rect 17359 29121 17371 29124
rect 17313 29115 17371 29121
rect 17678 29112 17684 29124
rect 17736 29112 17742 29164
rect 17954 29112 17960 29164
rect 18012 29152 18018 29164
rect 18417 29155 18475 29161
rect 18417 29152 18429 29155
rect 18012 29124 18429 29152
rect 18012 29112 18018 29124
rect 18417 29121 18429 29124
rect 18463 29121 18475 29155
rect 18417 29115 18475 29121
rect 12529 29087 12587 29093
rect 12529 29084 12541 29087
rect 10796 29056 12541 29084
rect 12529 29053 12541 29056
rect 12575 29053 12587 29087
rect 12529 29047 12587 29053
rect 14090 29044 14096 29096
rect 14148 29044 14154 29096
rect 14734 29044 14740 29096
rect 14792 29084 14798 29096
rect 16025 29087 16083 29093
rect 16025 29084 16037 29087
rect 14792 29056 16037 29084
rect 14792 29044 14798 29056
rect 16025 29053 16037 29056
rect 16071 29053 16083 29087
rect 16025 29047 16083 29053
rect 17402 29044 17408 29096
rect 17460 29044 17466 29096
rect 17586 29044 17592 29096
rect 17644 29084 17650 29096
rect 18601 29087 18659 29093
rect 18601 29084 18613 29087
rect 17644 29056 18613 29084
rect 17644 29044 17650 29056
rect 18601 29053 18613 29056
rect 18647 29084 18659 29087
rect 19306 29084 19334 29192
rect 20714 29180 20720 29232
rect 20772 29220 20778 29232
rect 22465 29223 22523 29229
rect 22465 29220 22477 29223
rect 20772 29192 22477 29220
rect 20772 29180 20778 29192
rect 22465 29189 22477 29192
rect 22511 29189 22523 29223
rect 22465 29183 22523 29189
rect 24578 29180 24584 29232
rect 24636 29220 24642 29232
rect 24673 29223 24731 29229
rect 24673 29220 24685 29223
rect 24636 29192 24685 29220
rect 24636 29180 24642 29192
rect 24673 29189 24685 29192
rect 24719 29189 24731 29223
rect 24673 29183 24731 29189
rect 19521 29155 19579 29161
rect 19521 29121 19533 29155
rect 19567 29152 19579 29155
rect 19794 29152 19800 29164
rect 19567 29124 19800 29152
rect 19567 29121 19579 29124
rect 19521 29115 19579 29121
rect 19794 29112 19800 29124
rect 19852 29152 19858 29164
rect 20165 29155 20223 29161
rect 20165 29152 20177 29155
rect 19852 29124 20177 29152
rect 19852 29112 19858 29124
rect 20165 29121 20177 29124
rect 20211 29121 20223 29155
rect 20806 29152 20812 29164
rect 20165 29115 20223 29121
rect 20272 29124 20812 29152
rect 20272 29096 20300 29124
rect 20806 29112 20812 29124
rect 20864 29112 20870 29164
rect 22738 29152 22744 29164
rect 21192 29124 22744 29152
rect 18647 29056 19334 29084
rect 18647 29053 18659 29056
rect 18601 29047 18659 29053
rect 20254 29044 20260 29096
rect 20312 29044 20318 29096
rect 20441 29087 20499 29093
rect 20441 29053 20453 29087
rect 20487 29084 20499 29087
rect 20530 29084 20536 29096
rect 20487 29056 20536 29084
rect 20487 29053 20499 29056
rect 20441 29047 20499 29053
rect 20530 29044 20536 29056
rect 20588 29084 20594 29096
rect 21192 29084 21220 29124
rect 22738 29112 22744 29124
rect 22796 29112 22802 29164
rect 23661 29155 23719 29161
rect 23661 29121 23673 29155
rect 23707 29152 23719 29155
rect 24118 29152 24124 29164
rect 23707 29124 24124 29152
rect 23707 29121 23719 29124
rect 23661 29115 23719 29121
rect 24118 29112 24124 29124
rect 24176 29112 24182 29164
rect 20588 29056 21220 29084
rect 20588 29044 20594 29056
rect 21266 29044 21272 29096
rect 21324 29044 21330 29096
rect 22462 29084 22468 29096
rect 21376 29056 22468 29084
rect 10192 28988 10272 29016
rect 10192 28976 10198 28988
rect 10778 28976 10784 29028
rect 10836 29016 10842 29028
rect 11977 29019 12035 29025
rect 11977 29016 11989 29019
rect 10836 28988 11989 29016
rect 10836 28976 10842 28988
rect 11977 28985 11989 28988
rect 12023 28985 12035 29019
rect 11977 28979 12035 28985
rect 12618 28976 12624 29028
rect 12676 29016 12682 29028
rect 13449 29019 13507 29025
rect 13449 29016 13461 29019
rect 12676 28988 13461 29016
rect 12676 28976 12682 28988
rect 13449 28985 13461 28988
rect 13495 28985 13507 29019
rect 13449 28979 13507 28985
rect 15470 28976 15476 29028
rect 15528 28976 15534 29028
rect 16853 29019 16911 29025
rect 16853 28985 16865 29019
rect 16899 29016 16911 29019
rect 18414 29016 18420 29028
rect 16899 28988 18420 29016
rect 16899 28985 16911 28988
rect 16853 28979 16911 28985
rect 18414 28976 18420 28988
rect 18472 28976 18478 29028
rect 19797 29019 19855 29025
rect 19797 28985 19809 29019
rect 19843 29016 19855 29019
rect 21376 29016 21404 29056
rect 22462 29044 22468 29056
rect 22520 29044 22526 29096
rect 22649 29087 22707 29093
rect 22649 29053 22661 29087
rect 22695 29084 22707 29087
rect 23290 29084 23296 29096
rect 22695 29056 23296 29084
rect 22695 29053 22707 29056
rect 22649 29047 22707 29053
rect 23290 29044 23296 29056
rect 23348 29044 23354 29096
rect 19843 28988 21404 29016
rect 19843 28985 19855 28988
rect 19797 28979 19855 28985
rect 21910 28976 21916 29028
rect 21968 29016 21974 29028
rect 22005 29019 22063 29025
rect 22005 29016 22017 29019
rect 21968 28988 22017 29016
rect 21968 28976 21974 28988
rect 22005 28985 22017 28988
rect 22051 28985 22063 29019
rect 22005 28979 22063 28985
rect 24857 29019 24915 29025
rect 24857 28985 24869 29019
rect 24903 29016 24915 29019
rect 25038 29016 25044 29028
rect 24903 28988 25044 29016
rect 24903 28985 24915 28988
rect 24857 28979 24915 28985
rect 25038 28976 25044 28988
rect 25096 28976 25102 29028
rect 7272 28951 7330 28957
rect 7272 28917 7284 28951
rect 7318 28948 7330 28951
rect 8294 28948 8300 28960
rect 7318 28920 8300 28948
rect 7318 28917 7330 28920
rect 7272 28911 7330 28917
rect 8294 28908 8300 28920
rect 8352 28908 8358 28960
rect 8662 28908 8668 28960
rect 8720 28948 8726 28960
rect 9125 28951 9183 28957
rect 9125 28948 9137 28951
rect 8720 28920 9137 28948
rect 8720 28908 8726 28920
rect 9125 28917 9137 28920
rect 9171 28948 9183 28951
rect 10962 28948 10968 28960
rect 9171 28920 10968 28948
rect 9171 28917 9183 28920
rect 9125 28911 9183 28917
rect 10962 28908 10968 28920
rect 11020 28908 11026 28960
rect 11606 28908 11612 28960
rect 11664 28948 11670 28960
rect 15010 28948 15016 28960
rect 11664 28920 15016 28948
rect 11664 28908 11670 28920
rect 15010 28908 15016 28920
rect 15068 28948 15074 28960
rect 17954 28948 17960 28960
rect 15068 28920 17960 28948
rect 15068 28908 15074 28920
rect 17954 28908 17960 28920
rect 18012 28908 18018 28960
rect 1104 28858 25852 28880
rect 1104 28806 2950 28858
rect 3002 28806 3014 28858
rect 3066 28806 3078 28858
rect 3130 28806 3142 28858
rect 3194 28806 3206 28858
rect 3258 28806 12950 28858
rect 13002 28806 13014 28858
rect 13066 28806 13078 28858
rect 13130 28806 13142 28858
rect 13194 28806 13206 28858
rect 13258 28806 22950 28858
rect 23002 28806 23014 28858
rect 23066 28806 23078 28858
rect 23130 28806 23142 28858
rect 23194 28806 23206 28858
rect 23258 28806 25852 28858
rect 1104 28784 25852 28806
rect 4062 28704 4068 28756
rect 4120 28744 4126 28756
rect 6365 28747 6423 28753
rect 6365 28744 6377 28747
rect 4120 28716 6377 28744
rect 4120 28704 4126 28716
rect 6365 28713 6377 28716
rect 6411 28744 6423 28747
rect 7650 28744 7656 28756
rect 6411 28716 7656 28744
rect 6411 28713 6423 28716
rect 6365 28707 6423 28713
rect 7650 28704 7656 28716
rect 7708 28704 7714 28756
rect 7742 28704 7748 28756
rect 7800 28744 7806 28756
rect 7837 28747 7895 28753
rect 7837 28744 7849 28747
rect 7800 28716 7849 28744
rect 7800 28704 7806 28716
rect 7837 28713 7849 28716
rect 7883 28713 7895 28747
rect 7837 28707 7895 28713
rect 7944 28716 10456 28744
rect 7944 28676 7972 28716
rect 7760 28648 7972 28676
rect 10428 28676 10456 28716
rect 10870 28704 10876 28756
rect 10928 28704 10934 28756
rect 11425 28747 11483 28753
rect 11425 28713 11437 28747
rect 11471 28744 11483 28747
rect 13354 28744 13360 28756
rect 11471 28716 13360 28744
rect 11471 28713 11483 28716
rect 11425 28707 11483 28713
rect 13354 28704 13360 28716
rect 13412 28704 13418 28756
rect 17954 28704 17960 28756
rect 18012 28704 18018 28756
rect 19150 28744 19156 28756
rect 18064 28716 19156 28744
rect 12621 28679 12679 28685
rect 10428 28648 12434 28676
rect 7760 28620 7788 28648
rect 1578 28568 1584 28620
rect 1636 28608 1642 28620
rect 3973 28611 4031 28617
rect 3973 28608 3985 28611
rect 1636 28580 3985 28608
rect 1636 28568 1642 28580
rect 3973 28577 3985 28580
rect 4019 28577 4031 28611
rect 3973 28571 4031 28577
rect 7742 28568 7748 28620
rect 7800 28568 7806 28620
rect 7834 28568 7840 28620
rect 7892 28608 7898 28620
rect 8389 28611 8447 28617
rect 8389 28608 8401 28611
rect 7892 28580 8401 28608
rect 7892 28568 7898 28580
rect 8389 28577 8401 28580
rect 8435 28577 8447 28611
rect 8389 28571 8447 28577
rect 12069 28611 12127 28617
rect 12069 28577 12081 28611
rect 12115 28577 12127 28611
rect 12406 28608 12434 28648
rect 12621 28645 12633 28679
rect 12667 28676 12679 28679
rect 13446 28676 13452 28688
rect 12667 28648 13452 28676
rect 12667 28645 12679 28648
rect 12621 28639 12679 28645
rect 13446 28636 13452 28648
rect 13504 28636 13510 28688
rect 13725 28679 13783 28685
rect 13725 28645 13737 28679
rect 13771 28676 13783 28679
rect 17586 28676 17592 28688
rect 13771 28648 17592 28676
rect 13771 28645 13783 28648
rect 13725 28639 13783 28645
rect 13173 28611 13231 28617
rect 13173 28608 13185 28611
rect 12406 28580 13185 28608
rect 12069 28571 12127 28577
rect 13173 28577 13185 28580
rect 13219 28577 13231 28611
rect 13173 28571 13231 28577
rect 6733 28543 6791 28549
rect 6733 28509 6745 28543
rect 6779 28540 6791 28543
rect 8754 28540 8760 28552
rect 6779 28512 8760 28540
rect 6779 28509 6791 28512
rect 6733 28503 6791 28509
rect 8754 28500 8760 28512
rect 8812 28500 8818 28552
rect 9122 28500 9128 28552
rect 9180 28500 9186 28552
rect 12084 28540 12112 28571
rect 12802 28540 12808 28552
rect 12084 28512 12808 28540
rect 12802 28500 12808 28512
rect 12860 28500 12866 28552
rect 12989 28543 13047 28549
rect 12989 28509 13001 28543
rect 13035 28540 13047 28543
rect 13740 28540 13768 28639
rect 17586 28636 17592 28648
rect 17644 28676 17650 28688
rect 18064 28676 18092 28716
rect 19150 28704 19156 28716
rect 19208 28704 19214 28756
rect 21085 28747 21143 28753
rect 21085 28713 21097 28747
rect 21131 28744 21143 28747
rect 22554 28744 22560 28756
rect 21131 28716 22560 28744
rect 21131 28713 21143 28716
rect 21085 28707 21143 28713
rect 22554 28704 22560 28716
rect 22612 28704 22618 28756
rect 17644 28648 18092 28676
rect 17644 28636 17650 28648
rect 18874 28636 18880 28688
rect 18932 28676 18938 28688
rect 23845 28679 23903 28685
rect 23845 28676 23857 28679
rect 18932 28648 23857 28676
rect 18932 28636 18938 28648
rect 23845 28645 23857 28648
rect 23891 28645 23903 28679
rect 23845 28639 23903 28645
rect 13814 28568 13820 28620
rect 13872 28608 13878 28620
rect 14829 28611 14887 28617
rect 14829 28608 14841 28611
rect 13872 28580 14841 28608
rect 13872 28568 13878 28580
rect 14829 28577 14841 28580
rect 14875 28577 14887 28611
rect 14829 28571 14887 28577
rect 16298 28568 16304 28620
rect 16356 28608 16362 28620
rect 16761 28611 16819 28617
rect 16761 28608 16773 28611
rect 16356 28580 16773 28608
rect 16356 28568 16362 28580
rect 16761 28577 16773 28580
rect 16807 28577 16819 28611
rect 16761 28571 16819 28577
rect 21729 28611 21787 28617
rect 21729 28577 21741 28611
rect 21775 28608 21787 28611
rect 23658 28608 23664 28620
rect 21775 28580 23664 28608
rect 21775 28577 21787 28580
rect 21729 28571 21787 28577
rect 23658 28568 23664 28580
rect 23716 28568 23722 28620
rect 13035 28512 13768 28540
rect 14645 28543 14703 28549
rect 13035 28509 13047 28512
rect 12989 28503 13047 28509
rect 14645 28509 14657 28543
rect 14691 28540 14703 28543
rect 15286 28540 15292 28552
rect 14691 28512 15292 28540
rect 14691 28509 14703 28512
rect 14645 28503 14703 28509
rect 15286 28500 15292 28512
rect 15344 28540 15350 28552
rect 15473 28543 15531 28549
rect 15473 28540 15485 28543
rect 15344 28512 15485 28540
rect 15344 28500 15350 28512
rect 15473 28509 15485 28512
rect 15519 28540 15531 28543
rect 16114 28540 16120 28552
rect 15519 28512 16120 28540
rect 15519 28509 15531 28512
rect 15473 28503 15531 28509
rect 16114 28500 16120 28512
rect 16172 28500 16178 28552
rect 16577 28543 16635 28549
rect 16577 28509 16589 28543
rect 16623 28540 16635 28543
rect 17034 28540 17040 28552
rect 16623 28512 17040 28540
rect 16623 28509 16635 28512
rect 16577 28503 16635 28509
rect 17034 28500 17040 28512
rect 17092 28500 17098 28552
rect 21266 28500 21272 28552
rect 21324 28540 21330 28552
rect 21453 28543 21511 28549
rect 21453 28540 21465 28543
rect 21324 28512 21465 28540
rect 21324 28500 21330 28512
rect 21453 28509 21465 28512
rect 21499 28509 21511 28543
rect 21453 28503 21511 28509
rect 24029 28543 24087 28549
rect 24029 28509 24041 28543
rect 24075 28509 24087 28543
rect 24029 28503 24087 28509
rect 3510 28432 3516 28484
rect 3568 28472 3574 28484
rect 4157 28475 4215 28481
rect 4157 28472 4169 28475
rect 3568 28444 4169 28472
rect 3568 28432 3574 28444
rect 4157 28441 4169 28444
rect 4203 28441 4215 28475
rect 4157 28435 4215 28441
rect 5718 28432 5724 28484
rect 5776 28472 5782 28484
rect 5813 28475 5871 28481
rect 5813 28472 5825 28475
rect 5776 28444 5825 28472
rect 5776 28432 5782 28444
rect 5813 28441 5825 28444
rect 5859 28441 5871 28475
rect 5813 28435 5871 28441
rect 7282 28432 7288 28484
rect 7340 28472 7346 28484
rect 8297 28475 8355 28481
rect 8297 28472 8309 28475
rect 7340 28444 8309 28472
rect 7340 28432 7346 28444
rect 8297 28441 8309 28444
rect 8343 28441 8355 28475
rect 8297 28435 8355 28441
rect 9398 28432 9404 28484
rect 9456 28432 9462 28484
rect 10962 28472 10968 28484
rect 10626 28444 10968 28472
rect 10962 28432 10968 28444
rect 11020 28432 11026 28484
rect 11793 28475 11851 28481
rect 11793 28441 11805 28475
rect 11839 28472 11851 28475
rect 12342 28472 12348 28484
rect 11839 28444 12348 28472
rect 11839 28441 11851 28444
rect 11793 28435 11851 28441
rect 12342 28432 12348 28444
rect 12400 28432 12406 28484
rect 13081 28475 13139 28481
rect 13081 28441 13093 28475
rect 13127 28472 13139 28475
rect 16482 28472 16488 28484
rect 13127 28444 16488 28472
rect 13127 28441 13139 28444
rect 13081 28435 13139 28441
rect 13740 28416 13768 28444
rect 16482 28432 16488 28444
rect 16540 28432 16546 28484
rect 16669 28475 16727 28481
rect 16669 28441 16681 28475
rect 16715 28472 16727 28475
rect 16850 28472 16856 28484
rect 16715 28444 16856 28472
rect 16715 28441 16727 28444
rect 16669 28435 16727 28441
rect 16850 28432 16856 28444
rect 16908 28432 16914 28484
rect 24044 28472 24072 28503
rect 24762 28500 24768 28552
rect 24820 28500 24826 28552
rect 25222 28472 25228 28484
rect 24044 28444 25228 28472
rect 25222 28432 25228 28444
rect 25280 28432 25286 28484
rect 6822 28364 6828 28416
rect 6880 28404 6886 28416
rect 7377 28407 7435 28413
rect 7377 28404 7389 28407
rect 6880 28376 7389 28404
rect 6880 28364 6886 28376
rect 7377 28373 7389 28376
rect 7423 28373 7435 28407
rect 7377 28367 7435 28373
rect 7650 28364 7656 28416
rect 7708 28404 7714 28416
rect 8205 28407 8263 28413
rect 8205 28404 8217 28407
rect 7708 28376 8217 28404
rect 7708 28364 7714 28376
rect 8205 28373 8217 28376
rect 8251 28404 8263 28407
rect 9582 28404 9588 28416
rect 8251 28376 9588 28404
rect 8251 28373 8263 28376
rect 8205 28367 8263 28373
rect 9582 28364 9588 28376
rect 9640 28364 9646 28416
rect 11054 28364 11060 28416
rect 11112 28404 11118 28416
rect 11885 28407 11943 28413
rect 11885 28404 11897 28407
rect 11112 28376 11897 28404
rect 11112 28364 11118 28376
rect 11885 28373 11897 28376
rect 11931 28373 11943 28407
rect 11885 28367 11943 28373
rect 13722 28364 13728 28416
rect 13780 28404 13786 28416
rect 13817 28407 13875 28413
rect 13817 28404 13829 28407
rect 13780 28376 13829 28404
rect 13780 28364 13786 28376
rect 13817 28373 13829 28376
rect 13863 28373 13875 28407
rect 13817 28367 13875 28373
rect 13906 28364 13912 28416
rect 13964 28404 13970 28416
rect 14277 28407 14335 28413
rect 14277 28404 14289 28407
rect 13964 28376 14289 28404
rect 13964 28364 13970 28376
rect 14277 28373 14289 28376
rect 14323 28373 14335 28407
rect 14277 28367 14335 28373
rect 14458 28364 14464 28416
rect 14516 28404 14522 28416
rect 14737 28407 14795 28413
rect 14737 28404 14749 28407
rect 14516 28376 14749 28404
rect 14516 28364 14522 28376
rect 14737 28373 14749 28376
rect 14783 28404 14795 28407
rect 15289 28407 15347 28413
rect 15289 28404 15301 28407
rect 14783 28376 15301 28404
rect 14783 28373 14795 28376
rect 14737 28367 14795 28373
rect 15289 28373 15301 28376
rect 15335 28373 15347 28407
rect 15289 28367 15347 28373
rect 16206 28364 16212 28416
rect 16264 28364 16270 28416
rect 17310 28364 17316 28416
rect 17368 28364 17374 28416
rect 17678 28364 17684 28416
rect 17736 28364 17742 28416
rect 20714 28364 20720 28416
rect 20772 28404 20778 28416
rect 21545 28407 21603 28413
rect 21545 28404 21557 28407
rect 20772 28376 21557 28404
rect 20772 28364 20778 28376
rect 21545 28373 21557 28376
rect 21591 28373 21603 28407
rect 21545 28367 21603 28373
rect 21818 28364 21824 28416
rect 21876 28404 21882 28416
rect 23750 28404 23756 28416
rect 21876 28376 23756 28404
rect 21876 28364 21882 28376
rect 23750 28364 23756 28376
rect 23808 28364 23814 28416
rect 24581 28407 24639 28413
rect 24581 28373 24593 28407
rect 24627 28404 24639 28407
rect 24762 28404 24768 28416
rect 24627 28376 24768 28404
rect 24627 28373 24639 28376
rect 24581 28367 24639 28373
rect 24762 28364 24768 28376
rect 24820 28364 24826 28416
rect 1104 28314 25852 28336
rect 1104 28262 7950 28314
rect 8002 28262 8014 28314
rect 8066 28262 8078 28314
rect 8130 28262 8142 28314
rect 8194 28262 8206 28314
rect 8258 28262 17950 28314
rect 18002 28262 18014 28314
rect 18066 28262 18078 28314
rect 18130 28262 18142 28314
rect 18194 28262 18206 28314
rect 18258 28262 25852 28314
rect 1104 28240 25852 28262
rect 8297 28203 8355 28209
rect 8297 28169 8309 28203
rect 8343 28200 8355 28203
rect 8570 28200 8576 28212
rect 8343 28172 8576 28200
rect 8343 28169 8355 28172
rect 8297 28163 8355 28169
rect 8570 28160 8576 28172
rect 8628 28160 8634 28212
rect 8662 28160 8668 28212
rect 8720 28160 8726 28212
rect 9398 28160 9404 28212
rect 9456 28200 9462 28212
rect 12345 28203 12403 28209
rect 12345 28200 12357 28203
rect 9456 28172 12357 28200
rect 9456 28160 9462 28172
rect 12345 28169 12357 28172
rect 12391 28169 12403 28203
rect 12345 28163 12403 28169
rect 13630 28160 13636 28212
rect 13688 28160 13694 28212
rect 14734 28160 14740 28212
rect 14792 28160 14798 28212
rect 15654 28160 15660 28212
rect 15712 28200 15718 28212
rect 17129 28203 17187 28209
rect 17129 28200 17141 28203
rect 15712 28172 17141 28200
rect 15712 28160 15718 28172
rect 17129 28169 17141 28172
rect 17175 28200 17187 28203
rect 17678 28200 17684 28212
rect 17175 28172 17684 28200
rect 17175 28169 17187 28172
rect 17129 28163 17187 28169
rect 17678 28160 17684 28172
rect 17736 28200 17742 28212
rect 17773 28203 17831 28209
rect 17773 28200 17785 28203
rect 17736 28172 17785 28200
rect 17736 28160 17742 28172
rect 17773 28169 17785 28172
rect 17819 28169 17831 28203
rect 21450 28200 21456 28212
rect 17773 28163 17831 28169
rect 18616 28172 21456 28200
rect 6822 28092 6828 28144
rect 6880 28092 6886 28144
rect 8680 28132 8708 28160
rect 10962 28132 10968 28144
rect 8050 28104 8708 28132
rect 10718 28104 10968 28132
rect 10962 28092 10968 28104
rect 11020 28092 11026 28144
rect 11422 28092 11428 28144
rect 11480 28132 11486 28144
rect 13648 28132 13676 28160
rect 11480 28104 13676 28132
rect 11480 28092 11486 28104
rect 11698 28024 11704 28076
rect 11756 28024 11762 28076
rect 2041 27999 2099 28005
rect 2041 27965 2053 27999
rect 2087 27965 2099 27999
rect 2041 27959 2099 27965
rect 2056 27928 2084 27959
rect 2222 27956 2228 28008
rect 2280 27956 2286 28008
rect 2774 27956 2780 28008
rect 2832 27956 2838 28008
rect 6454 27956 6460 28008
rect 6512 27996 6518 28008
rect 6549 27999 6607 28005
rect 6549 27996 6561 27999
rect 6512 27968 6561 27996
rect 6512 27956 6518 27968
rect 6549 27965 6561 27968
rect 6595 27965 6607 27999
rect 6549 27959 6607 27965
rect 9214 27956 9220 28008
rect 9272 27956 9278 28008
rect 9493 27999 9551 28005
rect 9493 27965 9505 27999
rect 9539 27996 9551 27999
rect 10502 27996 10508 28008
rect 9539 27968 10508 27996
rect 9539 27965 9551 27968
rect 9493 27959 9551 27965
rect 10502 27956 10508 27968
rect 10560 27956 10566 28008
rect 10965 27999 11023 28005
rect 10965 27965 10977 27999
rect 11011 27996 11023 27999
rect 11716 27996 11744 28024
rect 11011 27968 11744 27996
rect 11011 27965 11023 27968
rect 10965 27959 11023 27965
rect 12802 27956 12808 28008
rect 12860 27996 12866 28008
rect 12989 27999 13047 28005
rect 12989 27996 13001 27999
rect 12860 27968 13001 27996
rect 12860 27956 12866 27968
rect 12989 27965 13001 27968
rect 13035 27965 13047 27999
rect 12989 27959 13047 27965
rect 13265 27999 13323 28005
rect 13265 27965 13277 27999
rect 13311 27996 13323 27999
rect 13354 27996 13360 28008
rect 13311 27968 13360 27996
rect 13311 27965 13323 27968
rect 13265 27959 13323 27965
rect 13354 27956 13360 27968
rect 13412 27956 13418 28008
rect 4062 27928 4068 27940
rect 2056 27900 4068 27928
rect 4062 27888 4068 27900
rect 4120 27888 4126 27940
rect 11606 27928 11612 27940
rect 8496 27900 9352 27928
rect 5718 27820 5724 27872
rect 5776 27860 5782 27872
rect 8496 27860 8524 27900
rect 5776 27832 8524 27860
rect 9324 27860 9352 27900
rect 10980 27900 11612 27928
rect 10980 27860 11008 27900
rect 11606 27888 11612 27900
rect 11664 27888 11670 27940
rect 9324 27832 11008 27860
rect 5776 27820 5782 27832
rect 11054 27820 11060 27872
rect 11112 27860 11118 27872
rect 11241 27863 11299 27869
rect 11241 27860 11253 27863
rect 11112 27832 11253 27860
rect 11112 27820 11118 27832
rect 11241 27829 11253 27832
rect 11287 27829 11299 27863
rect 14384 27860 14412 28050
rect 15378 28024 15384 28076
rect 15436 28024 15442 28076
rect 18616 28073 18644 28172
rect 21450 28160 21456 28172
rect 21508 28160 21514 28212
rect 22112 28172 22692 28200
rect 21177 28135 21235 28141
rect 21177 28132 21189 28135
rect 20654 28104 21189 28132
rect 21177 28101 21189 28104
rect 21223 28132 21235 28135
rect 21634 28132 21640 28144
rect 21223 28104 21640 28132
rect 21223 28101 21235 28104
rect 21177 28095 21235 28101
rect 21634 28092 21640 28104
rect 21692 28132 21698 28144
rect 22112 28132 22140 28172
rect 21692 28104 22140 28132
rect 21692 28092 21698 28104
rect 18601 28067 18659 28073
rect 18601 28064 18613 28067
rect 17880 28036 18613 28064
rect 16114 27956 16120 28008
rect 16172 27996 16178 28008
rect 17880 28005 17908 28036
rect 18601 28033 18613 28036
rect 18647 28033 18659 28067
rect 20990 28064 20996 28076
rect 18601 28027 18659 28033
rect 20640 28036 20996 28064
rect 17865 27999 17923 28005
rect 17865 27996 17877 27999
rect 16172 27968 17877 27996
rect 16172 27956 16178 27968
rect 17865 27965 17877 27968
rect 17911 27965 17923 27999
rect 17865 27959 17923 27965
rect 18049 27999 18107 28005
rect 18049 27965 18061 27999
rect 18095 27965 18107 27999
rect 18049 27959 18107 27965
rect 14458 27888 14464 27940
rect 14516 27928 14522 27940
rect 17770 27928 17776 27940
rect 14516 27900 17776 27928
rect 14516 27888 14522 27900
rect 17770 27888 17776 27900
rect 17828 27928 17834 27940
rect 17954 27928 17960 27940
rect 17828 27900 17960 27928
rect 17828 27888 17834 27900
rect 17954 27888 17960 27900
rect 18012 27888 18018 27940
rect 18064 27928 18092 27959
rect 19150 27956 19156 28008
rect 19208 27956 19214 28008
rect 19429 27999 19487 28005
rect 19429 27965 19441 27999
rect 19475 27996 19487 27999
rect 19794 27996 19800 28008
rect 19475 27968 19800 27996
rect 19475 27965 19487 27968
rect 19429 27959 19487 27965
rect 19794 27956 19800 27968
rect 19852 27996 19858 28008
rect 20640 27996 20668 28036
rect 20990 28024 20996 28036
rect 21048 28024 21054 28076
rect 19852 27968 20668 27996
rect 19852 27956 19858 27968
rect 20898 27956 20904 28008
rect 20956 27956 20962 28008
rect 18509 27931 18567 27937
rect 18509 27928 18521 27931
rect 18064 27900 18521 27928
rect 18509 27897 18521 27900
rect 18555 27928 18567 27931
rect 18782 27928 18788 27940
rect 18555 27900 18788 27928
rect 18555 27897 18567 27900
rect 18509 27891 18567 27897
rect 18782 27888 18788 27900
rect 18840 27928 18846 27940
rect 18840 27900 19288 27928
rect 18840 27888 18846 27900
rect 19260 27872 19288 27900
rect 15105 27863 15163 27869
rect 15105 27860 15117 27863
rect 14384 27832 15117 27860
rect 11241 27823 11299 27829
rect 15105 27829 15117 27832
rect 15151 27860 15163 27863
rect 15930 27860 15936 27872
rect 15151 27832 15936 27860
rect 15151 27829 15163 27832
rect 15105 27823 15163 27829
rect 15930 27820 15936 27832
rect 15988 27820 15994 27872
rect 16022 27820 16028 27872
rect 16080 27820 16086 27872
rect 17405 27863 17463 27869
rect 17405 27829 17417 27863
rect 17451 27860 17463 27863
rect 18322 27860 18328 27872
rect 17451 27832 18328 27860
rect 17451 27829 17463 27832
rect 17405 27823 17463 27829
rect 18322 27820 18328 27832
rect 18380 27820 18386 27872
rect 19242 27820 19248 27872
rect 19300 27820 19306 27872
rect 21928 27860 21956 28104
rect 22186 28092 22192 28144
rect 22244 28132 22250 28144
rect 22554 28132 22560 28144
rect 22244 28104 22560 28132
rect 22244 28092 22250 28104
rect 22554 28092 22560 28104
rect 22612 28092 22618 28144
rect 22664 28132 22692 28172
rect 23750 28160 23756 28212
rect 23808 28160 23814 28212
rect 25222 28160 25228 28212
rect 25280 28160 25286 28212
rect 22664 28104 22770 28132
rect 24670 28092 24676 28144
rect 24728 28092 24734 28144
rect 22002 27956 22008 28008
rect 22060 27956 22066 28008
rect 22281 27999 22339 28005
rect 22281 27965 22293 27999
rect 22327 27996 22339 27999
rect 25130 27996 25136 28008
rect 22327 27968 25136 27996
rect 22327 27965 22339 27968
rect 22281 27959 22339 27965
rect 25130 27956 25136 27968
rect 25188 27956 25194 28008
rect 24857 27931 24915 27937
rect 24857 27897 24869 27931
rect 24903 27928 24915 27931
rect 25222 27928 25228 27940
rect 24903 27900 25228 27928
rect 24903 27897 24915 27900
rect 24857 27891 24915 27897
rect 25222 27888 25228 27900
rect 25280 27888 25286 27940
rect 22830 27860 22836 27872
rect 21928 27832 22836 27860
rect 22830 27820 22836 27832
rect 22888 27860 22894 27872
rect 23842 27860 23848 27872
rect 22888 27832 23848 27860
rect 22888 27820 22894 27832
rect 23842 27820 23848 27832
rect 23900 27860 23906 27872
rect 24121 27863 24179 27869
rect 24121 27860 24133 27863
rect 23900 27832 24133 27860
rect 23900 27820 23906 27832
rect 24121 27829 24133 27832
rect 24167 27829 24179 27863
rect 24121 27823 24179 27829
rect 1104 27770 25852 27792
rect 1104 27718 2950 27770
rect 3002 27718 3014 27770
rect 3066 27718 3078 27770
rect 3130 27718 3142 27770
rect 3194 27718 3206 27770
rect 3258 27718 12950 27770
rect 13002 27718 13014 27770
rect 13066 27718 13078 27770
rect 13130 27718 13142 27770
rect 13194 27718 13206 27770
rect 13258 27718 22950 27770
rect 23002 27718 23014 27770
rect 23066 27718 23078 27770
rect 23130 27718 23142 27770
rect 23194 27718 23206 27770
rect 23258 27718 25852 27770
rect 1104 27696 25852 27718
rect 7745 27659 7803 27665
rect 7745 27625 7757 27659
rect 7791 27656 7803 27659
rect 7834 27656 7840 27668
rect 7791 27628 7840 27656
rect 7791 27625 7803 27628
rect 7745 27619 7803 27625
rect 7834 27616 7840 27628
rect 7892 27616 7898 27668
rect 10962 27616 10968 27668
rect 11020 27656 11026 27668
rect 11057 27659 11115 27665
rect 11057 27656 11069 27659
rect 11020 27628 11069 27656
rect 11020 27616 11026 27628
rect 11057 27625 11069 27628
rect 11103 27625 11115 27659
rect 11057 27619 11115 27625
rect 15644 27659 15702 27665
rect 15644 27625 15656 27659
rect 15690 27656 15702 27659
rect 16022 27656 16028 27668
rect 15690 27628 16028 27656
rect 15690 27625 15702 27628
rect 15644 27619 15702 27625
rect 16022 27616 16028 27628
rect 16080 27616 16086 27668
rect 19150 27656 19156 27668
rect 17880 27628 19156 27656
rect 12989 27591 13047 27597
rect 12989 27557 13001 27591
rect 13035 27588 13047 27591
rect 14550 27588 14556 27600
rect 13035 27560 14556 27588
rect 13035 27557 13047 27560
rect 12989 27551 13047 27557
rect 14550 27548 14556 27560
rect 14608 27548 14614 27600
rect 8754 27480 8760 27532
rect 8812 27520 8818 27532
rect 11977 27523 12035 27529
rect 11977 27520 11989 27523
rect 8812 27492 11989 27520
rect 8812 27480 8818 27492
rect 11977 27489 11989 27492
rect 12023 27489 12035 27523
rect 11977 27483 12035 27489
rect 12066 27480 12072 27532
rect 12124 27520 12130 27532
rect 13541 27523 13599 27529
rect 13541 27520 13553 27523
rect 12124 27492 13553 27520
rect 12124 27480 12130 27492
rect 13541 27489 13553 27492
rect 13587 27489 13599 27523
rect 14090 27520 14096 27532
rect 13541 27483 13599 27489
rect 13648 27492 14096 27520
rect 3786 27412 3792 27464
rect 3844 27452 3850 27464
rect 4008 27455 4066 27461
rect 4008 27452 4020 27455
rect 3844 27424 4020 27452
rect 3844 27412 3850 27424
rect 4008 27421 4020 27424
rect 4054 27421 4066 27455
rect 4008 27415 4066 27421
rect 6641 27455 6699 27461
rect 6641 27421 6653 27455
rect 6687 27452 6699 27455
rect 8294 27452 8300 27464
rect 6687 27424 8300 27452
rect 6687 27421 6699 27424
rect 6641 27415 6699 27421
rect 8294 27412 8300 27424
rect 8352 27412 8358 27464
rect 11885 27455 11943 27461
rect 11885 27421 11897 27455
rect 11931 27452 11943 27455
rect 13648 27452 13676 27492
rect 14090 27480 14096 27492
rect 14148 27480 14154 27532
rect 15381 27523 15439 27529
rect 15381 27489 15393 27523
rect 15427 27520 15439 27523
rect 16390 27520 16396 27532
rect 15427 27492 16396 27520
rect 15427 27489 15439 27492
rect 15381 27483 15439 27489
rect 16390 27480 16396 27492
rect 16448 27520 16454 27532
rect 17880 27520 17908 27628
rect 19150 27616 19156 27628
rect 19208 27616 19214 27668
rect 22094 27616 22100 27668
rect 22152 27656 22158 27668
rect 22152 27628 22324 27656
rect 22152 27616 22158 27628
rect 17954 27548 17960 27600
rect 18012 27588 18018 27600
rect 18969 27591 19027 27597
rect 18969 27588 18981 27591
rect 18012 27560 18981 27588
rect 18012 27548 18018 27560
rect 18969 27557 18981 27560
rect 19015 27557 19027 27591
rect 18969 27551 19027 27557
rect 20625 27591 20683 27597
rect 20625 27557 20637 27591
rect 20671 27588 20683 27591
rect 22186 27588 22192 27600
rect 20671 27560 22192 27588
rect 20671 27557 20683 27560
rect 20625 27551 20683 27557
rect 18233 27523 18291 27529
rect 18233 27520 18245 27523
rect 16448 27492 17908 27520
rect 18064 27492 18245 27520
rect 16448 27480 16454 27492
rect 11931 27424 13676 27452
rect 11931 27421 11943 27424
rect 11885 27415 11943 27421
rect 13814 27412 13820 27464
rect 13872 27452 13878 27464
rect 14277 27455 14335 27461
rect 14277 27452 14289 27455
rect 13872 27424 14289 27452
rect 13872 27412 13878 27424
rect 14277 27421 14289 27424
rect 14323 27452 14335 27455
rect 14734 27452 14740 27464
rect 14323 27424 14740 27452
rect 14323 27421 14335 27424
rect 14277 27415 14335 27421
rect 14734 27412 14740 27424
rect 14792 27412 14798 27464
rect 17862 27412 17868 27464
rect 17920 27452 17926 27464
rect 18064 27452 18092 27492
rect 18233 27489 18245 27492
rect 18279 27489 18291 27523
rect 18233 27483 18291 27489
rect 17920 27424 18092 27452
rect 18141 27455 18199 27461
rect 17920 27412 17926 27424
rect 18141 27421 18153 27455
rect 18187 27452 18199 27455
rect 18414 27452 18420 27464
rect 18187 27424 18420 27452
rect 18187 27421 18199 27424
rect 18141 27415 18199 27421
rect 18414 27412 18420 27424
rect 18472 27412 18478 27464
rect 18984 27452 19012 27551
rect 22186 27548 22192 27560
rect 22244 27548 22250 27600
rect 19978 27480 19984 27532
rect 20036 27520 20042 27532
rect 20073 27523 20131 27529
rect 20073 27520 20085 27523
rect 20036 27492 20085 27520
rect 20036 27480 20042 27492
rect 20073 27489 20085 27492
rect 20119 27520 20131 27523
rect 20346 27520 20352 27532
rect 20119 27492 20352 27520
rect 20119 27489 20131 27492
rect 20073 27483 20131 27489
rect 20346 27480 20352 27492
rect 20404 27480 20410 27532
rect 21082 27480 21088 27532
rect 21140 27480 21146 27532
rect 21269 27523 21327 27529
rect 21269 27489 21281 27523
rect 21315 27520 21327 27523
rect 22296 27520 22324 27628
rect 22646 27520 22652 27532
rect 21315 27492 22652 27520
rect 21315 27489 21327 27492
rect 21269 27483 21327 27489
rect 22646 27480 22652 27492
rect 22704 27480 22710 27532
rect 23290 27480 23296 27532
rect 23348 27520 23354 27532
rect 24029 27523 24087 27529
rect 24029 27520 24041 27523
rect 23348 27492 24041 27520
rect 23348 27480 23354 27492
rect 24029 27489 24041 27492
rect 24075 27489 24087 27523
rect 24029 27483 24087 27489
rect 19797 27455 19855 27461
rect 19797 27452 19809 27455
rect 18984 27424 19809 27452
rect 19797 27421 19809 27424
rect 19843 27421 19855 27455
rect 19797 27415 19855 27421
rect 22002 27412 22008 27464
rect 22060 27452 22066 27464
rect 22281 27455 22339 27461
rect 22281 27452 22293 27455
rect 22060 27424 22293 27452
rect 22060 27412 22066 27424
rect 22281 27421 22293 27424
rect 22327 27421 22339 27455
rect 22281 27415 22339 27421
rect 3878 27344 3884 27396
rect 3936 27384 3942 27396
rect 4111 27387 4169 27393
rect 4111 27384 4123 27387
rect 3936 27356 4123 27384
rect 3936 27344 3942 27356
rect 4111 27353 4123 27356
rect 4157 27353 4169 27387
rect 4111 27347 4169 27353
rect 9122 27344 9128 27396
rect 9180 27384 9186 27396
rect 11793 27387 11851 27393
rect 11793 27384 11805 27387
rect 9180 27356 11805 27384
rect 9180 27344 9186 27356
rect 11793 27353 11805 27356
rect 11839 27353 11851 27387
rect 13449 27387 13507 27393
rect 13449 27384 13461 27387
rect 11793 27347 11851 27353
rect 12636 27356 13461 27384
rect 6730 27276 6736 27328
rect 6788 27316 6794 27328
rect 7285 27319 7343 27325
rect 7285 27316 7297 27319
rect 6788 27288 7297 27316
rect 6788 27276 6794 27288
rect 7285 27285 7297 27288
rect 7331 27285 7343 27319
rect 7285 27279 7343 27285
rect 9490 27276 9496 27328
rect 9548 27316 9554 27328
rect 9585 27319 9643 27325
rect 9585 27316 9597 27319
rect 9548 27288 9597 27316
rect 9548 27276 9554 27288
rect 9585 27285 9597 27288
rect 9631 27285 9643 27319
rect 9585 27279 9643 27285
rect 11425 27319 11483 27325
rect 11425 27285 11437 27319
rect 11471 27316 11483 27319
rect 12250 27316 12256 27328
rect 11471 27288 12256 27316
rect 11471 27285 11483 27288
rect 11425 27279 11483 27285
rect 12250 27276 12256 27288
rect 12308 27276 12314 27328
rect 12434 27276 12440 27328
rect 12492 27316 12498 27328
rect 12636 27325 12664 27356
rect 13449 27353 13461 27356
rect 13495 27384 13507 27387
rect 14458 27384 14464 27396
rect 13495 27356 14464 27384
rect 13495 27353 13507 27356
rect 13449 27347 13507 27353
rect 14458 27344 14464 27356
rect 14516 27344 14522 27396
rect 15930 27344 15936 27396
rect 15988 27384 15994 27396
rect 18049 27387 18107 27393
rect 15988 27356 16146 27384
rect 16960 27356 17816 27384
rect 15988 27344 15994 27356
rect 12621 27319 12679 27325
rect 12621 27316 12633 27319
rect 12492 27288 12633 27316
rect 12492 27276 12498 27288
rect 12621 27285 12633 27288
rect 12667 27285 12679 27319
rect 12621 27279 12679 27285
rect 13262 27276 13268 27328
rect 13320 27316 13326 27328
rect 13357 27319 13415 27325
rect 13357 27316 13369 27319
rect 13320 27288 13369 27316
rect 13320 27276 13326 27288
rect 13357 27285 13369 27288
rect 13403 27285 13415 27319
rect 13357 27279 13415 27285
rect 13538 27276 13544 27328
rect 13596 27316 13602 27328
rect 14921 27319 14979 27325
rect 14921 27316 14933 27319
rect 13596 27288 14933 27316
rect 13596 27276 13602 27288
rect 14921 27285 14933 27288
rect 14967 27285 14979 27319
rect 16040 27316 16068 27356
rect 16960 27316 16988 27356
rect 16040 27288 16988 27316
rect 17129 27319 17187 27325
rect 14921 27279 14979 27285
rect 17129 27285 17141 27319
rect 17175 27316 17187 27319
rect 17310 27316 17316 27328
rect 17175 27288 17316 27316
rect 17175 27285 17187 27288
rect 17129 27279 17187 27285
rect 17310 27276 17316 27288
rect 17368 27276 17374 27328
rect 17678 27276 17684 27328
rect 17736 27276 17742 27328
rect 17788 27316 17816 27356
rect 18049 27353 18061 27387
rect 18095 27384 18107 27387
rect 19334 27384 19340 27396
rect 18095 27356 19340 27384
rect 18095 27353 18107 27356
rect 18049 27347 18107 27353
rect 19334 27344 19340 27356
rect 19392 27344 19398 27396
rect 22557 27387 22615 27393
rect 22557 27353 22569 27387
rect 22603 27384 22615 27387
rect 22646 27384 22652 27396
rect 22603 27356 22652 27384
rect 22603 27353 22615 27356
rect 22557 27347 22615 27353
rect 22646 27344 22652 27356
rect 22704 27344 22710 27396
rect 22830 27344 22836 27396
rect 22888 27384 22894 27396
rect 24673 27387 24731 27393
rect 22888 27356 23046 27384
rect 22888 27344 22894 27356
rect 24673 27353 24685 27387
rect 24719 27353 24731 27387
rect 24673 27347 24731 27353
rect 24857 27387 24915 27393
rect 24857 27353 24869 27387
rect 24903 27384 24915 27387
rect 25314 27384 25320 27396
rect 24903 27356 25320 27384
rect 24903 27353 24915 27356
rect 24857 27347 24915 27353
rect 18693 27319 18751 27325
rect 18693 27316 18705 27319
rect 17788 27288 18705 27316
rect 18693 27285 18705 27288
rect 18739 27285 18751 27319
rect 18693 27279 18751 27285
rect 19429 27319 19487 27325
rect 19429 27285 19441 27319
rect 19475 27316 19487 27319
rect 19702 27316 19708 27328
rect 19475 27288 19708 27316
rect 19475 27285 19487 27288
rect 19429 27279 19487 27285
rect 19702 27276 19708 27288
rect 19760 27276 19766 27328
rect 19889 27319 19947 27325
rect 19889 27285 19901 27319
rect 19935 27316 19947 27319
rect 20438 27316 20444 27328
rect 19935 27288 20444 27316
rect 19935 27285 19947 27288
rect 19889 27279 19947 27285
rect 20438 27276 20444 27288
rect 20496 27276 20502 27328
rect 20622 27276 20628 27328
rect 20680 27316 20686 27328
rect 20993 27319 21051 27325
rect 20993 27316 21005 27319
rect 20680 27288 21005 27316
rect 20680 27276 20686 27288
rect 20993 27285 21005 27288
rect 21039 27285 21051 27319
rect 20993 27279 21051 27285
rect 22370 27276 22376 27328
rect 22428 27316 22434 27328
rect 24688 27316 24716 27347
rect 25314 27344 25320 27356
rect 25372 27344 25378 27396
rect 22428 27288 24716 27316
rect 22428 27276 22434 27288
rect 1104 27226 25852 27248
rect 1104 27174 7950 27226
rect 8002 27174 8014 27226
rect 8066 27174 8078 27226
rect 8130 27174 8142 27226
rect 8194 27174 8206 27226
rect 8258 27174 17950 27226
rect 18002 27174 18014 27226
rect 18066 27174 18078 27226
rect 18130 27174 18142 27226
rect 18194 27174 18206 27226
rect 18258 27174 25852 27226
rect 1104 27152 25852 27174
rect 7834 27112 7840 27124
rect 6840 27084 7840 27112
rect 6840 27053 6868 27084
rect 7834 27072 7840 27084
rect 7892 27112 7898 27124
rect 8570 27112 8576 27124
rect 7892 27084 8576 27112
rect 7892 27072 7898 27084
rect 8570 27072 8576 27084
rect 8628 27072 8634 27124
rect 8662 27072 8668 27124
rect 8720 27072 8726 27124
rect 9122 27072 9128 27124
rect 9180 27072 9186 27124
rect 9490 27072 9496 27124
rect 9548 27072 9554 27124
rect 15013 27115 15071 27121
rect 15013 27081 15025 27115
rect 15059 27112 15071 27115
rect 15102 27112 15108 27124
rect 15059 27084 15108 27112
rect 15059 27081 15071 27084
rect 15013 27075 15071 27081
rect 15102 27072 15108 27084
rect 15160 27112 15166 27124
rect 15378 27112 15384 27124
rect 15160 27084 15384 27112
rect 15160 27072 15166 27084
rect 15378 27072 15384 27084
rect 15436 27072 15442 27124
rect 16298 27072 16304 27124
rect 16356 27112 16362 27124
rect 17770 27112 17776 27124
rect 16356 27084 17776 27112
rect 16356 27072 16362 27084
rect 17770 27072 17776 27084
rect 17828 27072 17834 27124
rect 18509 27115 18567 27121
rect 18509 27081 18521 27115
rect 18555 27112 18567 27115
rect 18874 27112 18880 27124
rect 18555 27084 18880 27112
rect 18555 27081 18567 27084
rect 18509 27075 18567 27081
rect 18874 27072 18880 27084
rect 18932 27072 18938 27124
rect 20438 27072 20444 27124
rect 20496 27072 20502 27124
rect 22646 27072 22652 27124
rect 22704 27112 22710 27124
rect 23753 27115 23811 27121
rect 23753 27112 23765 27115
rect 22704 27084 23765 27112
rect 22704 27072 22710 27084
rect 23753 27081 23765 27084
rect 23799 27081 23811 27115
rect 23753 27075 23811 27081
rect 6825 27047 6883 27053
rect 6825 27013 6837 27047
rect 6871 27013 6883 27047
rect 8680 27044 8708 27072
rect 8050 27016 8708 27044
rect 10689 27047 10747 27053
rect 6825 27007 6883 27013
rect 10689 27013 10701 27047
rect 10735 27044 10747 27047
rect 11146 27044 11152 27056
rect 10735 27016 11152 27044
rect 10735 27013 10747 27016
rect 10689 27007 10747 27013
rect 11146 27004 11152 27016
rect 11204 27004 11210 27056
rect 13538 27004 13544 27056
rect 13596 27004 13602 27056
rect 17310 27004 17316 27056
rect 17368 27044 17374 27056
rect 19794 27044 19800 27056
rect 17368 27016 19800 27044
rect 17368 27004 17374 27016
rect 3418 26936 3424 26988
rect 3476 26936 3482 26988
rect 10962 26936 10968 26988
rect 11020 26976 11026 26988
rect 11701 26979 11759 26985
rect 11701 26976 11713 26979
rect 11020 26948 11713 26976
rect 11020 26936 11026 26948
rect 11701 26945 11713 26948
rect 11747 26976 11759 26979
rect 12066 26976 12072 26988
rect 11747 26948 12072 26976
rect 11747 26945 11759 26948
rect 11701 26939 11759 26945
rect 12066 26936 12072 26948
rect 12124 26936 12130 26988
rect 12802 26936 12808 26988
rect 12860 26976 12866 26988
rect 13265 26979 13323 26985
rect 13265 26976 13277 26979
rect 12860 26948 13277 26976
rect 12860 26936 12866 26948
rect 13265 26945 13277 26948
rect 13311 26945 13323 26979
rect 13265 26939 13323 26945
rect 14568 26948 14674 26976
rect 3602 26868 3608 26920
rect 3660 26868 3666 26920
rect 5166 26868 5172 26920
rect 5224 26868 5230 26920
rect 6454 26868 6460 26920
rect 6512 26908 6518 26920
rect 6549 26911 6607 26917
rect 6549 26908 6561 26911
rect 6512 26880 6561 26908
rect 6512 26868 6518 26880
rect 6549 26877 6561 26880
rect 6595 26877 6607 26911
rect 6549 26871 6607 26877
rect 8570 26868 8576 26920
rect 8628 26908 8634 26920
rect 8757 26911 8815 26917
rect 8757 26908 8769 26911
rect 8628 26880 8769 26908
rect 8628 26868 8634 26880
rect 8757 26877 8769 26880
rect 8803 26908 8815 26911
rect 8846 26908 8852 26920
rect 8803 26880 8852 26908
rect 8803 26877 8815 26880
rect 8757 26871 8815 26877
rect 8846 26868 8852 26880
rect 8904 26908 8910 26920
rect 9585 26911 9643 26917
rect 9585 26908 9597 26911
rect 8904 26880 9597 26908
rect 8904 26868 8910 26880
rect 9585 26877 9597 26880
rect 9631 26877 9643 26911
rect 9585 26871 9643 26877
rect 9769 26911 9827 26917
rect 9769 26877 9781 26911
rect 9815 26908 9827 26911
rect 10870 26908 10876 26920
rect 9815 26880 10876 26908
rect 9815 26877 9827 26880
rect 9769 26871 9827 26877
rect 10870 26868 10876 26880
rect 10928 26868 10934 26920
rect 8294 26800 8300 26852
rect 8352 26840 8358 26852
rect 10686 26840 10692 26852
rect 8352 26812 10692 26840
rect 8352 26800 8358 26812
rect 10686 26800 10692 26812
rect 10744 26800 10750 26852
rect 10042 26732 10048 26784
rect 10100 26772 10106 26784
rect 10781 26775 10839 26781
rect 10781 26772 10793 26775
rect 10100 26744 10793 26772
rect 10100 26732 10106 26744
rect 10781 26741 10793 26744
rect 10827 26741 10839 26775
rect 10781 26735 10839 26741
rect 11238 26732 11244 26784
rect 11296 26772 11302 26784
rect 12345 26775 12403 26781
rect 12345 26772 12357 26775
rect 11296 26744 12357 26772
rect 11296 26732 11302 26744
rect 12345 26741 12357 26744
rect 12391 26741 12403 26775
rect 12345 26735 12403 26741
rect 13262 26732 13268 26784
rect 13320 26772 13326 26784
rect 14090 26772 14096 26784
rect 13320 26744 14096 26772
rect 13320 26732 13326 26744
rect 14090 26732 14096 26744
rect 14148 26732 14154 26784
rect 14568 26772 14596 26948
rect 17218 26936 17224 26988
rect 17276 26936 17282 26988
rect 17954 26936 17960 26988
rect 18012 26976 18018 26988
rect 18417 26979 18475 26985
rect 18417 26976 18429 26979
rect 18012 26948 18429 26976
rect 18012 26936 18018 26948
rect 18417 26945 18429 26948
rect 18463 26945 18475 26979
rect 18417 26939 18475 26945
rect 16114 26868 16120 26920
rect 16172 26908 16178 26920
rect 17310 26908 17316 26920
rect 16172 26880 17316 26908
rect 16172 26868 16178 26880
rect 17310 26868 17316 26880
rect 17368 26868 17374 26920
rect 18708 26917 18736 27016
rect 19794 27004 19800 27016
rect 19852 27004 19858 27056
rect 22830 27004 22836 27056
rect 22888 27004 22894 27056
rect 24302 27004 24308 27056
rect 24360 27044 24366 27056
rect 24673 27047 24731 27053
rect 24673 27044 24685 27047
rect 24360 27016 24685 27044
rect 24360 27004 24366 27016
rect 24673 27013 24685 27016
rect 24719 27013 24731 27047
rect 24673 27007 24731 27013
rect 19426 26936 19432 26988
rect 19484 26936 19490 26988
rect 20809 26979 20867 26985
rect 20809 26945 20821 26979
rect 20855 26976 20867 26979
rect 20898 26976 20904 26988
rect 20855 26948 20904 26976
rect 20855 26945 20867 26948
rect 20809 26939 20867 26945
rect 20898 26936 20904 26948
rect 20956 26936 20962 26988
rect 17405 26911 17463 26917
rect 17405 26877 17417 26911
rect 17451 26877 17463 26911
rect 17405 26871 17463 26877
rect 18693 26911 18751 26917
rect 18693 26877 18705 26911
rect 18739 26877 18751 26911
rect 18693 26871 18751 26877
rect 14642 26800 14648 26852
rect 14700 26840 14706 26852
rect 17420 26840 17448 26871
rect 19794 26868 19800 26920
rect 19852 26908 19858 26920
rect 19889 26911 19947 26917
rect 19889 26908 19901 26911
rect 19852 26880 19901 26908
rect 19852 26868 19858 26880
rect 19889 26877 19901 26880
rect 19935 26877 19947 26911
rect 19889 26871 19947 26877
rect 22002 26868 22008 26920
rect 22060 26868 22066 26920
rect 22278 26868 22284 26920
rect 22336 26868 22342 26920
rect 22830 26868 22836 26920
rect 22888 26908 22894 26920
rect 24121 26911 24179 26917
rect 24121 26908 24133 26911
rect 22888 26880 24133 26908
rect 22888 26868 22894 26880
rect 24121 26877 24133 26880
rect 24167 26908 24179 26911
rect 25133 26911 25191 26917
rect 25133 26908 25145 26911
rect 24167 26880 25145 26908
rect 24167 26877 24179 26880
rect 24121 26871 24179 26877
rect 25133 26877 25145 26880
rect 25179 26877 25191 26911
rect 25133 26871 25191 26877
rect 14700 26812 17448 26840
rect 19245 26843 19303 26849
rect 14700 26800 14706 26812
rect 19245 26809 19257 26843
rect 19291 26840 19303 26843
rect 21266 26840 21272 26852
rect 19291 26812 21272 26840
rect 19291 26809 19303 26812
rect 19245 26803 19303 26809
rect 21266 26800 21272 26812
rect 21324 26800 21330 26852
rect 22020 26840 22048 26868
rect 24857 26843 24915 26849
rect 22020 26812 22094 26840
rect 15381 26775 15439 26781
rect 15381 26772 15393 26775
rect 14568 26744 15393 26772
rect 15381 26741 15393 26744
rect 15427 26772 15439 26775
rect 15930 26772 15936 26784
rect 15427 26744 15936 26772
rect 15427 26741 15439 26744
rect 15381 26735 15439 26741
rect 15930 26732 15936 26744
rect 15988 26732 15994 26784
rect 16114 26732 16120 26784
rect 16172 26772 16178 26784
rect 16393 26775 16451 26781
rect 16393 26772 16405 26775
rect 16172 26744 16405 26772
rect 16172 26732 16178 26744
rect 16393 26741 16405 26744
rect 16439 26741 16451 26775
rect 16393 26735 16451 26741
rect 16850 26732 16856 26784
rect 16908 26732 16914 26784
rect 18046 26732 18052 26784
rect 18104 26732 18110 26784
rect 20714 26732 20720 26784
rect 20772 26772 20778 26784
rect 21453 26775 21511 26781
rect 21453 26772 21465 26775
rect 20772 26744 21465 26772
rect 20772 26732 20778 26744
rect 21453 26741 21465 26744
rect 21499 26741 21511 26775
rect 22066 26772 22094 26812
rect 24857 26809 24869 26843
rect 24903 26840 24915 26843
rect 24946 26840 24952 26852
rect 24903 26812 24952 26840
rect 24903 26809 24915 26812
rect 24857 26803 24915 26809
rect 24946 26800 24952 26812
rect 25004 26800 25010 26852
rect 22830 26772 22836 26784
rect 22066 26744 22836 26772
rect 21453 26735 21511 26741
rect 22830 26732 22836 26744
rect 22888 26732 22894 26784
rect 1104 26682 25852 26704
rect 1104 26630 2950 26682
rect 3002 26630 3014 26682
rect 3066 26630 3078 26682
rect 3130 26630 3142 26682
rect 3194 26630 3206 26682
rect 3258 26630 12950 26682
rect 13002 26630 13014 26682
rect 13066 26630 13078 26682
rect 13130 26630 13142 26682
rect 13194 26630 13206 26682
rect 13258 26630 22950 26682
rect 23002 26630 23014 26682
rect 23066 26630 23078 26682
rect 23130 26630 23142 26682
rect 23194 26630 23206 26682
rect 23258 26630 25852 26682
rect 1104 26608 25852 26630
rect 3605 26571 3663 26577
rect 3605 26537 3617 26571
rect 3651 26568 3663 26571
rect 3694 26568 3700 26580
rect 3651 26540 3700 26568
rect 3651 26537 3663 26540
rect 3605 26531 3663 26537
rect 3694 26528 3700 26540
rect 3752 26528 3758 26580
rect 4249 26571 4307 26577
rect 4249 26537 4261 26571
rect 4295 26568 4307 26571
rect 4798 26568 4804 26580
rect 4295 26540 4804 26568
rect 4295 26537 4307 26540
rect 4249 26531 4307 26537
rect 4798 26528 4804 26540
rect 4856 26528 4862 26580
rect 6178 26528 6184 26580
rect 6236 26568 6242 26580
rect 6822 26568 6828 26580
rect 6236 26540 6828 26568
rect 6236 26528 6242 26540
rect 6822 26528 6828 26540
rect 6880 26528 6886 26580
rect 7742 26528 7748 26580
rect 7800 26568 7806 26580
rect 8205 26571 8263 26577
rect 8205 26568 8217 26571
rect 7800 26540 8217 26568
rect 7800 26528 7806 26540
rect 8205 26537 8217 26540
rect 8251 26537 8263 26571
rect 8205 26531 8263 26537
rect 8573 26571 8631 26577
rect 8573 26537 8585 26571
rect 8619 26568 8631 26571
rect 8662 26568 8668 26580
rect 8619 26540 8668 26568
rect 8619 26537 8631 26540
rect 8573 26531 8631 26537
rect 8662 26528 8668 26540
rect 8720 26528 8726 26580
rect 10226 26528 10232 26580
rect 10284 26568 10290 26580
rect 10413 26571 10471 26577
rect 10413 26568 10425 26571
rect 10284 26540 10425 26568
rect 10284 26528 10290 26540
rect 10413 26537 10425 26540
rect 10459 26537 10471 26571
rect 10413 26531 10471 26537
rect 12989 26571 13047 26577
rect 12989 26537 13001 26571
rect 13035 26568 13047 26571
rect 14826 26568 14832 26580
rect 13035 26540 14832 26568
rect 13035 26537 13047 26540
rect 12989 26531 13047 26537
rect 2222 26392 2228 26444
rect 2280 26432 2286 26444
rect 4433 26435 4491 26441
rect 4433 26432 4445 26435
rect 2280 26404 4445 26432
rect 2280 26392 2286 26404
rect 4433 26401 4445 26404
rect 4479 26401 4491 26435
rect 4433 26395 4491 26401
rect 6730 26392 6736 26444
rect 6788 26392 6794 26444
rect 6822 26392 6828 26444
rect 6880 26432 6886 26444
rect 10428 26432 10456 26531
rect 14826 26528 14832 26540
rect 14884 26528 14890 26580
rect 17218 26528 17224 26580
rect 17276 26568 17282 26580
rect 17681 26571 17739 26577
rect 17681 26568 17693 26571
rect 17276 26540 17693 26568
rect 17276 26528 17282 26540
rect 17681 26537 17693 26540
rect 17727 26537 17739 26571
rect 17681 26531 17739 26537
rect 10781 26503 10839 26509
rect 10781 26469 10793 26503
rect 10827 26500 10839 26503
rect 11790 26500 11796 26512
rect 10827 26472 11796 26500
rect 10827 26469 10839 26472
rect 10781 26463 10839 26469
rect 11790 26460 11796 26472
rect 11848 26460 11854 26512
rect 14921 26503 14979 26509
rect 14921 26500 14933 26503
rect 13464 26472 14933 26500
rect 11241 26435 11299 26441
rect 11241 26432 11253 26435
rect 6880 26404 10364 26432
rect 10428 26404 11253 26432
rect 6880 26392 6886 26404
rect 3694 26324 3700 26376
rect 3752 26364 3758 26376
rect 3973 26367 4031 26373
rect 3973 26364 3985 26367
rect 3752 26336 3985 26364
rect 3752 26324 3758 26336
rect 3973 26333 3985 26336
rect 4019 26333 4031 26367
rect 3973 26327 4031 26333
rect 6454 26324 6460 26376
rect 6512 26324 6518 26376
rect 8662 26364 8668 26376
rect 7866 26336 8668 26364
rect 8662 26324 8668 26336
rect 8720 26324 8726 26376
rect 9306 26324 9312 26376
rect 9364 26364 9370 26376
rect 9401 26367 9459 26373
rect 9401 26364 9413 26367
rect 9364 26336 9413 26364
rect 9364 26324 9370 26336
rect 9401 26333 9413 26336
rect 9447 26333 9459 26367
rect 10336 26364 10364 26404
rect 11241 26401 11253 26404
rect 11287 26401 11299 26435
rect 11241 26395 11299 26401
rect 11422 26392 11428 26444
rect 11480 26392 11486 26444
rect 12342 26392 12348 26444
rect 12400 26392 12406 26444
rect 13464 26441 13492 26472
rect 14921 26469 14933 26472
rect 14967 26469 14979 26503
rect 17696 26500 17724 26531
rect 17954 26528 17960 26580
rect 18012 26568 18018 26580
rect 18598 26568 18604 26580
rect 18012 26540 18604 26568
rect 18012 26528 18018 26540
rect 18598 26528 18604 26540
rect 18656 26528 18662 26580
rect 18690 26528 18696 26580
rect 18748 26568 18754 26580
rect 20533 26571 20591 26577
rect 20533 26568 20545 26571
rect 18748 26540 20545 26568
rect 18748 26528 18754 26540
rect 20533 26537 20545 26540
rect 20579 26568 20591 26571
rect 20622 26568 20628 26580
rect 20579 26540 20628 26568
rect 20579 26537 20591 26540
rect 20533 26531 20591 26537
rect 20622 26528 20628 26540
rect 20680 26528 20686 26580
rect 20806 26528 20812 26580
rect 20864 26528 20870 26580
rect 22094 26528 22100 26580
rect 22152 26568 22158 26580
rect 23937 26571 23995 26577
rect 23937 26568 23949 26571
rect 22152 26540 23949 26568
rect 22152 26528 22158 26540
rect 23937 26537 23949 26540
rect 23983 26537 23995 26571
rect 23937 26531 23995 26537
rect 25130 26528 25136 26580
rect 25188 26568 25194 26580
rect 25225 26571 25283 26577
rect 25225 26568 25237 26571
rect 25188 26540 25237 26568
rect 25188 26528 25194 26540
rect 25225 26537 25237 26540
rect 25271 26537 25283 26571
rect 25225 26531 25283 26537
rect 20993 26503 21051 26509
rect 20993 26500 21005 26503
rect 14921 26463 14979 26469
rect 15488 26472 16436 26500
rect 17696 26472 21005 26500
rect 13449 26435 13507 26441
rect 13449 26401 13461 26435
rect 13495 26401 13507 26435
rect 13449 26395 13507 26401
rect 13633 26435 13691 26441
rect 13633 26401 13645 26435
rect 13679 26432 13691 26435
rect 13814 26432 13820 26444
rect 13679 26404 13820 26432
rect 13679 26401 13691 26404
rect 13633 26395 13691 26401
rect 13814 26392 13820 26404
rect 13872 26392 13878 26444
rect 14090 26392 14096 26444
rect 14148 26432 14154 26444
rect 14185 26435 14243 26441
rect 14185 26432 14197 26435
rect 14148 26404 14197 26432
rect 14148 26392 14154 26404
rect 14185 26401 14197 26404
rect 14231 26432 14243 26435
rect 15488 26432 15516 26472
rect 14231 26404 15516 26432
rect 15565 26435 15623 26441
rect 14231 26401 14243 26404
rect 14185 26395 14243 26401
rect 15565 26401 15577 26435
rect 15611 26432 15623 26435
rect 16298 26432 16304 26444
rect 15611 26404 16304 26432
rect 15611 26401 15623 26404
rect 15565 26395 15623 26401
rect 10336 26336 12434 26364
rect 9401 26327 9459 26333
rect 5166 26256 5172 26308
rect 5224 26296 5230 26308
rect 11054 26296 11060 26308
rect 5224 26268 7144 26296
rect 5224 26256 5230 26268
rect 7116 26228 7144 26268
rect 8036 26268 11060 26296
rect 8036 26228 8064 26268
rect 11054 26256 11060 26268
rect 11112 26296 11118 26308
rect 12066 26296 12072 26308
rect 11112 26268 12072 26296
rect 11112 26256 11118 26268
rect 12066 26256 12072 26268
rect 12124 26256 12130 26308
rect 12406 26296 12434 26336
rect 13354 26324 13360 26376
rect 13412 26364 13418 26376
rect 13538 26364 13544 26376
rect 13412 26336 13544 26364
rect 13412 26324 13418 26336
rect 13538 26324 13544 26336
rect 13596 26364 13602 26376
rect 15580 26364 15608 26395
rect 16298 26392 16304 26404
rect 16356 26392 16362 26444
rect 13596 26336 15608 26364
rect 13596 26324 13602 26336
rect 16114 26324 16120 26376
rect 16172 26324 16178 26376
rect 16408 26364 16436 26472
rect 20993 26469 21005 26472
rect 21039 26469 21051 26503
rect 20993 26463 21051 26469
rect 21269 26503 21327 26509
rect 21269 26469 21281 26503
rect 21315 26500 21327 26503
rect 21542 26500 21548 26512
rect 21315 26472 21548 26500
rect 21315 26469 21327 26472
rect 21269 26463 21327 26469
rect 16666 26392 16672 26444
rect 16724 26392 16730 26444
rect 18046 26392 18052 26444
rect 18104 26432 18110 26444
rect 19889 26435 19947 26441
rect 19889 26432 19901 26435
rect 18104 26404 19901 26432
rect 18104 26392 18110 26404
rect 19889 26401 19901 26404
rect 19935 26401 19947 26435
rect 19889 26395 19947 26401
rect 20073 26435 20131 26441
rect 20073 26401 20085 26435
rect 20119 26432 20131 26435
rect 20898 26432 20904 26444
rect 20119 26404 20904 26432
rect 20119 26401 20131 26404
rect 20073 26395 20131 26401
rect 20898 26392 20904 26404
rect 20956 26392 20962 26444
rect 21008 26432 21036 26463
rect 21542 26460 21548 26472
rect 21600 26460 21606 26512
rect 21729 26435 21787 26441
rect 21729 26432 21741 26435
rect 21008 26404 21741 26432
rect 21729 26401 21741 26404
rect 21775 26401 21787 26435
rect 21729 26395 21787 26401
rect 16684 26364 16712 26392
rect 19150 26364 19156 26376
rect 16408 26336 19156 26364
rect 19150 26324 19156 26336
rect 19208 26324 19214 26376
rect 19794 26324 19800 26376
rect 19852 26324 19858 26376
rect 20438 26324 20444 26376
rect 20496 26324 20502 26376
rect 20806 26324 20812 26376
rect 20864 26364 20870 26376
rect 21637 26367 21695 26373
rect 21637 26364 21649 26367
rect 20864 26336 21649 26364
rect 20864 26324 20870 26336
rect 21637 26333 21649 26336
rect 21683 26333 21695 26367
rect 21637 26327 21695 26333
rect 14645 26299 14703 26305
rect 14645 26296 14657 26299
rect 12406 26268 14657 26296
rect 14645 26265 14657 26268
rect 14691 26296 14703 26299
rect 15289 26299 15347 26305
rect 15289 26296 15301 26299
rect 14691 26268 15301 26296
rect 14691 26265 14703 26268
rect 14645 26259 14703 26265
rect 15289 26265 15301 26268
rect 15335 26265 15347 26299
rect 15289 26259 15347 26265
rect 15381 26299 15439 26305
rect 15381 26265 15393 26299
rect 15427 26296 15439 26299
rect 15562 26296 15568 26308
rect 15427 26268 15568 26296
rect 15427 26265 15439 26268
rect 15381 26259 15439 26265
rect 7116 26200 8064 26228
rect 9766 26188 9772 26240
rect 9824 26228 9830 26240
rect 10045 26231 10103 26237
rect 10045 26228 10057 26231
rect 9824 26200 10057 26228
rect 9824 26188 9830 26200
rect 10045 26197 10057 26200
rect 10091 26197 10103 26231
rect 10045 26191 10103 26197
rect 11146 26188 11152 26240
rect 11204 26188 11210 26240
rect 13354 26188 13360 26240
rect 13412 26188 13418 26240
rect 15304 26228 15332 26259
rect 15562 26256 15568 26268
rect 15620 26256 15626 26308
rect 16666 26296 16672 26308
rect 15672 26268 16672 26296
rect 15672 26228 15700 26268
rect 16666 26256 16672 26268
rect 16724 26296 16730 26308
rect 18690 26296 18696 26308
rect 16724 26268 18696 26296
rect 16724 26256 16730 26268
rect 18690 26256 18696 26268
rect 18748 26256 18754 26308
rect 20456 26296 20484 26324
rect 19812 26268 20484 26296
rect 21744 26296 21772 26395
rect 21818 26392 21824 26444
rect 21876 26392 21882 26444
rect 22462 26392 22468 26444
rect 22520 26432 22526 26444
rect 22925 26435 22983 26441
rect 22925 26432 22937 26435
rect 22520 26404 22937 26432
rect 22520 26392 22526 26404
rect 22925 26401 22937 26404
rect 22971 26401 22983 26435
rect 22925 26395 22983 26401
rect 23109 26435 23167 26441
rect 23109 26401 23121 26435
rect 23155 26432 23167 26435
rect 24026 26432 24032 26444
rect 23155 26404 24032 26432
rect 23155 26401 23167 26404
rect 23109 26395 23167 26401
rect 24026 26392 24032 26404
rect 24084 26392 24090 26444
rect 22738 26324 22744 26376
rect 22796 26364 22802 26376
rect 23845 26367 23903 26373
rect 23845 26364 23857 26367
rect 22796 26336 23857 26364
rect 22796 26324 22802 26336
rect 23845 26333 23857 26336
rect 23891 26333 23903 26367
rect 23845 26327 23903 26333
rect 24578 26324 24584 26376
rect 24636 26324 24642 26376
rect 22370 26296 22376 26308
rect 21744 26268 22376 26296
rect 19812 26240 19840 26268
rect 22370 26256 22376 26268
rect 22428 26256 22434 26308
rect 22554 26256 22560 26308
rect 22612 26296 22618 26308
rect 22833 26299 22891 26305
rect 22833 26296 22845 26299
rect 22612 26268 22845 26296
rect 22612 26256 22618 26268
rect 22833 26265 22845 26268
rect 22879 26265 22891 26299
rect 22833 26259 22891 26265
rect 15304 26200 15700 26228
rect 16758 26188 16764 26240
rect 16816 26188 16822 26240
rect 19426 26188 19432 26240
rect 19484 26188 19490 26240
rect 19794 26188 19800 26240
rect 19852 26188 19858 26240
rect 22462 26188 22468 26240
rect 22520 26188 22526 26240
rect 1104 26138 25852 26160
rect 1104 26086 7950 26138
rect 8002 26086 8014 26138
rect 8066 26086 8078 26138
rect 8130 26086 8142 26138
rect 8194 26086 8206 26138
rect 8258 26086 17950 26138
rect 18002 26086 18014 26138
rect 18066 26086 18078 26138
rect 18130 26086 18142 26138
rect 18194 26086 18206 26138
rect 18258 26086 25852 26138
rect 1104 26064 25852 26086
rect 3510 26033 3516 26036
rect 3467 26027 3516 26033
rect 3467 25993 3479 26027
rect 3513 25993 3516 26027
rect 3467 25987 3516 25993
rect 3510 25984 3516 25987
rect 3568 25984 3574 26036
rect 8478 25984 8484 26036
rect 8536 26024 8542 26036
rect 8662 26024 8668 26036
rect 8536 25996 8668 26024
rect 8536 25984 8542 25996
rect 8662 25984 8668 25996
rect 8720 26024 8726 26036
rect 9493 26027 9551 26033
rect 9493 26024 9505 26027
rect 8720 25996 9505 26024
rect 8720 25984 8726 25996
rect 7742 25916 7748 25968
rect 7800 25916 7806 25968
rect 9048 25956 9076 25996
rect 9493 25993 9505 25996
rect 9539 25993 9551 26027
rect 9493 25987 9551 25993
rect 10597 26027 10655 26033
rect 10597 25993 10609 26027
rect 10643 26024 10655 26027
rect 10778 26024 10784 26036
rect 10643 25996 10784 26024
rect 10643 25993 10655 25996
rect 10597 25987 10655 25993
rect 8970 25928 9076 25956
rect 9508 25956 9536 25987
rect 10778 25984 10784 25996
rect 10836 25984 10842 26036
rect 11146 25984 11152 26036
rect 11204 26024 11210 26036
rect 11701 26027 11759 26033
rect 11701 26024 11713 26027
rect 11204 25996 11713 26024
rect 11204 25984 11210 25996
rect 11701 25993 11713 25996
rect 11747 25993 11759 26027
rect 11701 25987 11759 25993
rect 11790 25984 11796 26036
rect 11848 26024 11854 26036
rect 12989 26027 13047 26033
rect 12989 26024 13001 26027
rect 11848 25996 13001 26024
rect 11848 25984 11854 25996
rect 12989 25993 13001 25996
rect 13035 25993 13047 26027
rect 12989 25987 13047 25993
rect 13081 26027 13139 26033
rect 13081 25993 13093 26027
rect 13127 26024 13139 26027
rect 13906 26024 13912 26036
rect 13127 25996 13912 26024
rect 13127 25993 13139 25996
rect 13081 25987 13139 25993
rect 13906 25984 13912 25996
rect 13964 25984 13970 26036
rect 16758 26024 16764 26036
rect 14568 25996 16764 26024
rect 9508 25928 11192 25956
rect 11164 25900 11192 25928
rect 12066 25916 12072 25968
rect 12124 25956 12130 25968
rect 14568 25965 14596 25996
rect 16758 25984 16764 25996
rect 16816 25984 16822 26036
rect 18322 25984 18328 26036
rect 18380 25984 18386 26036
rect 19610 25984 19616 26036
rect 19668 25984 19674 26036
rect 19702 25984 19708 26036
rect 19760 25984 19766 26036
rect 22186 25984 22192 26036
rect 22244 26024 22250 26036
rect 22557 26027 22615 26033
rect 22557 26024 22569 26027
rect 22244 25996 22569 26024
rect 22244 25984 22250 25996
rect 22557 25993 22569 25996
rect 22603 25993 22615 26027
rect 22557 25987 22615 25993
rect 12161 25959 12219 25965
rect 12161 25956 12173 25959
rect 12124 25928 12173 25956
rect 12124 25916 12130 25928
rect 12161 25925 12173 25928
rect 12207 25925 12219 25959
rect 12161 25919 12219 25925
rect 14553 25959 14611 25965
rect 14553 25925 14565 25959
rect 14599 25925 14611 25959
rect 14553 25919 14611 25925
rect 16298 25916 16304 25968
rect 16356 25916 16362 25968
rect 18233 25959 18291 25965
rect 18233 25925 18245 25959
rect 18279 25956 18291 25959
rect 18414 25956 18420 25968
rect 18279 25928 18420 25956
rect 18279 25925 18291 25928
rect 18233 25919 18291 25925
rect 18414 25916 18420 25928
rect 18472 25916 18478 25968
rect 23382 25956 23388 25968
rect 21468 25928 23388 25956
rect 2682 25848 2688 25900
rect 2740 25888 2746 25900
rect 3364 25891 3422 25897
rect 3364 25888 3376 25891
rect 2740 25860 3376 25888
rect 2740 25848 2746 25860
rect 3364 25857 3376 25860
rect 3410 25857 3422 25891
rect 3364 25851 3422 25857
rect 3694 25848 3700 25900
rect 3752 25888 3758 25900
rect 3973 25891 4031 25897
rect 3973 25888 3985 25891
rect 3752 25860 3985 25888
rect 3752 25848 3758 25860
rect 3973 25857 3985 25860
rect 4019 25857 4031 25891
rect 3973 25851 4031 25857
rect 6546 25848 6552 25900
rect 6604 25888 6610 25900
rect 7469 25891 7527 25897
rect 7469 25888 7481 25891
rect 6604 25860 7481 25888
rect 6604 25848 6610 25860
rect 7469 25857 7481 25860
rect 7515 25857 7527 25891
rect 7469 25851 7527 25857
rect 10502 25848 10508 25900
rect 10560 25848 10566 25900
rect 11146 25848 11152 25900
rect 11204 25848 11210 25900
rect 11698 25848 11704 25900
rect 11756 25888 11762 25900
rect 15930 25888 15936 25900
rect 11756 25860 13216 25888
rect 15686 25860 15936 25888
rect 11756 25848 11762 25860
rect 3053 25823 3111 25829
rect 3053 25789 3065 25823
rect 3099 25820 3111 25823
rect 3712 25820 3740 25848
rect 3099 25792 3740 25820
rect 3099 25789 3111 25792
rect 3053 25783 3111 25789
rect 6822 25780 6828 25832
rect 6880 25780 6886 25832
rect 10686 25780 10692 25832
rect 10744 25780 10750 25832
rect 13188 25829 13216 25860
rect 15930 25848 15936 25860
rect 15988 25888 15994 25900
rect 16574 25888 16580 25900
rect 15988 25860 16580 25888
rect 15988 25848 15994 25860
rect 16574 25848 16580 25860
rect 16632 25848 16638 25900
rect 19150 25848 19156 25900
rect 19208 25888 19214 25900
rect 19610 25888 19616 25900
rect 19208 25860 19616 25888
rect 19208 25848 19214 25860
rect 19610 25848 19616 25860
rect 19668 25848 19674 25900
rect 21468 25897 21496 25928
rect 23382 25916 23388 25928
rect 23440 25916 23446 25968
rect 20993 25891 21051 25897
rect 20993 25857 21005 25891
rect 21039 25888 21051 25891
rect 21453 25891 21511 25897
rect 21453 25888 21465 25891
rect 21039 25860 21465 25888
rect 21039 25857 21051 25860
rect 20993 25851 21051 25857
rect 21453 25857 21465 25860
rect 21499 25857 21511 25891
rect 21453 25851 21511 25857
rect 22465 25891 22523 25897
rect 22465 25857 22477 25891
rect 22511 25888 22523 25891
rect 23293 25891 23351 25897
rect 23293 25888 23305 25891
rect 22511 25860 23305 25888
rect 22511 25857 22523 25860
rect 22465 25851 22523 25857
rect 23293 25857 23305 25860
rect 23339 25857 23351 25891
rect 23293 25851 23351 25857
rect 24118 25848 24124 25900
rect 24176 25848 24182 25900
rect 13173 25823 13231 25829
rect 13173 25789 13185 25823
rect 13219 25789 13231 25823
rect 13173 25783 13231 25789
rect 14277 25823 14335 25829
rect 14277 25789 14289 25823
rect 14323 25820 14335 25823
rect 18509 25823 18567 25829
rect 14323 25792 14412 25820
rect 14323 25789 14335 25792
rect 14277 25783 14335 25789
rect 3786 25712 3792 25764
rect 3844 25752 3850 25764
rect 4433 25755 4491 25761
rect 4433 25752 4445 25755
rect 3844 25724 4445 25752
rect 3844 25712 3850 25724
rect 4433 25721 4445 25724
rect 4479 25721 4491 25755
rect 4433 25715 4491 25721
rect 4249 25687 4307 25693
rect 4249 25653 4261 25687
rect 4295 25684 4307 25687
rect 4338 25684 4344 25696
rect 4295 25656 4344 25684
rect 4295 25653 4307 25656
rect 4249 25647 4307 25653
rect 4338 25644 4344 25656
rect 4396 25644 4402 25696
rect 9217 25687 9275 25693
rect 9217 25653 9229 25687
rect 9263 25684 9275 25687
rect 9306 25684 9312 25696
rect 9263 25656 9312 25684
rect 9263 25653 9275 25656
rect 9217 25647 9275 25653
rect 9306 25644 9312 25656
rect 9364 25644 9370 25696
rect 10137 25687 10195 25693
rect 10137 25653 10149 25687
rect 10183 25684 10195 25687
rect 10686 25684 10692 25696
rect 10183 25656 10692 25684
rect 10183 25653 10195 25656
rect 10137 25647 10195 25653
rect 10686 25644 10692 25656
rect 10744 25644 10750 25696
rect 11146 25644 11152 25696
rect 11204 25684 11210 25696
rect 11241 25687 11299 25693
rect 11241 25684 11253 25687
rect 11204 25656 11253 25684
rect 11204 25644 11210 25656
rect 11241 25653 11253 25656
rect 11287 25684 11299 25687
rect 12342 25684 12348 25696
rect 11287 25656 12348 25684
rect 11287 25653 11299 25656
rect 11241 25647 11299 25653
rect 12342 25644 12348 25656
rect 12400 25644 12406 25696
rect 12621 25687 12679 25693
rect 12621 25653 12633 25687
rect 12667 25684 12679 25687
rect 14090 25684 14096 25696
rect 12667 25656 14096 25684
rect 12667 25653 12679 25656
rect 12621 25647 12679 25653
rect 14090 25644 14096 25656
rect 14148 25644 14154 25696
rect 14384 25684 14412 25792
rect 18509 25789 18521 25823
rect 18555 25820 18567 25823
rect 18874 25820 18880 25832
rect 18555 25792 18880 25820
rect 18555 25789 18567 25792
rect 18509 25783 18567 25789
rect 18874 25780 18880 25792
rect 18932 25780 18938 25832
rect 19889 25823 19947 25829
rect 19889 25789 19901 25823
rect 19935 25820 19947 25823
rect 20622 25820 20628 25832
rect 19935 25792 20628 25820
rect 19935 25789 19947 25792
rect 19889 25783 19947 25789
rect 20622 25780 20628 25792
rect 20680 25780 20686 25832
rect 22741 25823 22799 25829
rect 22741 25789 22753 25823
rect 22787 25820 22799 25823
rect 23198 25820 23204 25832
rect 22787 25792 23204 25820
rect 22787 25789 22799 25792
rect 22741 25783 22799 25789
rect 23198 25780 23204 25792
rect 23256 25780 23262 25832
rect 25130 25780 25136 25832
rect 25188 25780 25194 25832
rect 17126 25712 17132 25764
rect 17184 25752 17190 25764
rect 21269 25755 21327 25761
rect 21269 25752 21281 25755
rect 17184 25724 21281 25752
rect 17184 25712 17190 25724
rect 21269 25721 21281 25724
rect 21315 25721 21327 25755
rect 21269 25715 21327 25721
rect 16390 25684 16396 25696
rect 14384 25656 16396 25684
rect 16390 25644 16396 25656
rect 16448 25644 16454 25696
rect 16574 25644 16580 25696
rect 16632 25684 16638 25696
rect 16669 25687 16727 25693
rect 16669 25684 16681 25687
rect 16632 25656 16681 25684
rect 16632 25644 16638 25656
rect 16669 25653 16681 25656
rect 16715 25653 16727 25687
rect 16669 25647 16727 25653
rect 17770 25644 17776 25696
rect 17828 25684 17834 25696
rect 17865 25687 17923 25693
rect 17865 25684 17877 25687
rect 17828 25656 17877 25684
rect 17828 25644 17834 25656
rect 17865 25653 17877 25656
rect 17911 25653 17923 25687
rect 17865 25647 17923 25653
rect 19242 25644 19248 25696
rect 19300 25644 19306 25696
rect 22097 25687 22155 25693
rect 22097 25653 22109 25687
rect 22143 25684 22155 25687
rect 22370 25684 22376 25696
rect 22143 25656 22376 25684
rect 22143 25653 22155 25656
rect 22097 25647 22155 25653
rect 22370 25644 22376 25656
rect 22428 25644 22434 25696
rect 1104 25594 25852 25616
rect 1104 25542 2950 25594
rect 3002 25542 3014 25594
rect 3066 25542 3078 25594
rect 3130 25542 3142 25594
rect 3194 25542 3206 25594
rect 3258 25542 12950 25594
rect 13002 25542 13014 25594
rect 13066 25542 13078 25594
rect 13130 25542 13142 25594
rect 13194 25542 13206 25594
rect 13258 25542 22950 25594
rect 23002 25542 23014 25594
rect 23066 25542 23078 25594
rect 23130 25542 23142 25594
rect 23194 25542 23206 25594
rect 23258 25542 25852 25594
rect 1104 25520 25852 25542
rect 4062 25440 4068 25492
rect 4120 25440 4126 25492
rect 7469 25483 7527 25489
rect 7469 25449 7481 25483
rect 7515 25480 7527 25483
rect 10502 25480 10508 25492
rect 7515 25452 10508 25480
rect 7515 25449 7527 25452
rect 7469 25443 7527 25449
rect 10502 25440 10508 25452
rect 10560 25440 10566 25492
rect 10594 25440 10600 25492
rect 10652 25480 10658 25492
rect 10962 25480 10968 25492
rect 10652 25452 10968 25480
rect 10652 25440 10658 25452
rect 10962 25440 10968 25452
rect 11020 25440 11026 25492
rect 12161 25483 12219 25489
rect 12161 25449 12173 25483
rect 12207 25480 12219 25483
rect 13354 25480 13360 25492
rect 12207 25452 13360 25480
rect 12207 25449 12219 25452
rect 12161 25443 12219 25449
rect 13354 25440 13360 25452
rect 13412 25440 13418 25492
rect 14090 25440 14096 25492
rect 14148 25480 14154 25492
rect 18414 25480 18420 25492
rect 14148 25452 18420 25480
rect 14148 25440 14154 25452
rect 18414 25440 18420 25452
rect 18472 25440 18478 25492
rect 22278 25440 22284 25492
rect 22336 25480 22342 25492
rect 23201 25483 23259 25489
rect 23201 25480 23213 25483
rect 22336 25452 23213 25480
rect 22336 25440 22342 25452
rect 23201 25449 23213 25452
rect 23247 25449 23259 25483
rect 23201 25443 23259 25449
rect 7834 25372 7840 25424
rect 7892 25412 7898 25424
rect 11146 25412 11152 25424
rect 7892 25384 8064 25412
rect 7892 25372 7898 25384
rect 4890 25304 4896 25356
rect 4948 25344 4954 25356
rect 7101 25347 7159 25353
rect 7101 25344 7113 25347
rect 4948 25316 7113 25344
rect 4948 25304 4954 25316
rect 7101 25313 7113 25316
rect 7147 25344 7159 25347
rect 7466 25344 7472 25356
rect 7147 25316 7472 25344
rect 7147 25313 7159 25316
rect 7101 25307 7159 25313
rect 7466 25304 7472 25316
rect 7524 25344 7530 25356
rect 8036 25353 8064 25384
rect 10612 25384 11152 25412
rect 7929 25347 7987 25353
rect 7929 25344 7941 25347
rect 7524 25316 7941 25344
rect 7524 25304 7530 25316
rect 7929 25313 7941 25316
rect 7975 25313 7987 25347
rect 7929 25307 7987 25313
rect 8021 25347 8079 25353
rect 8021 25313 8033 25347
rect 8067 25313 8079 25347
rect 8021 25307 8079 25313
rect 9214 25304 9220 25356
rect 9272 25344 9278 25356
rect 9858 25344 9864 25356
rect 9272 25316 9864 25344
rect 9272 25304 9278 25316
rect 9858 25304 9864 25316
rect 9916 25304 9922 25356
rect 4249 25279 4307 25285
rect 4249 25245 4261 25279
rect 4295 25245 4307 25279
rect 4249 25239 4307 25245
rect 4264 25208 4292 25239
rect 4798 25236 4804 25288
rect 4856 25236 4862 25288
rect 4982 25236 4988 25288
rect 5040 25276 5046 25288
rect 5040 25248 6776 25276
rect 5040 25236 5046 25248
rect 6454 25208 6460 25220
rect 4264 25180 6460 25208
rect 6454 25168 6460 25180
rect 6512 25168 6518 25220
rect 4246 25100 4252 25152
rect 4304 25140 4310 25152
rect 5445 25143 5503 25149
rect 5445 25140 5457 25143
rect 4304 25112 5457 25140
rect 4304 25100 4310 25112
rect 5445 25109 5457 25112
rect 5491 25109 5503 25143
rect 6748 25140 6776 25248
rect 6822 25236 6828 25288
rect 6880 25276 6886 25288
rect 7837 25279 7895 25285
rect 7837 25276 7849 25279
rect 6880 25248 7849 25276
rect 6880 25236 6886 25248
rect 7837 25245 7849 25248
rect 7883 25245 7895 25279
rect 10612 25262 10640 25384
rect 11146 25372 11152 25384
rect 11204 25372 11210 25424
rect 12434 25372 12440 25424
rect 12492 25412 12498 25424
rect 13262 25412 13268 25424
rect 12492 25384 13268 25412
rect 12492 25372 12498 25384
rect 13262 25372 13268 25384
rect 13320 25372 13326 25424
rect 21726 25372 21732 25424
rect 21784 25412 21790 25424
rect 23566 25412 23572 25424
rect 21784 25384 23572 25412
rect 21784 25372 21790 25384
rect 23566 25372 23572 25384
rect 23624 25372 23630 25424
rect 12526 25304 12532 25356
rect 12584 25344 12590 25356
rect 12621 25347 12679 25353
rect 12621 25344 12633 25347
rect 12584 25316 12633 25344
rect 12584 25304 12590 25316
rect 12621 25313 12633 25316
rect 12667 25313 12679 25347
rect 12621 25307 12679 25313
rect 12805 25347 12863 25353
rect 12805 25313 12817 25347
rect 12851 25344 12863 25347
rect 13538 25344 13544 25356
rect 12851 25316 13544 25344
rect 12851 25313 12863 25316
rect 12805 25307 12863 25313
rect 13538 25304 13544 25316
rect 13596 25304 13602 25356
rect 15102 25304 15108 25356
rect 15160 25304 15166 25356
rect 17126 25304 17132 25356
rect 17184 25344 17190 25356
rect 17221 25347 17279 25353
rect 17221 25344 17233 25347
rect 17184 25316 17233 25344
rect 17184 25304 17190 25316
rect 17221 25313 17233 25316
rect 17267 25313 17279 25347
rect 17221 25307 17279 25313
rect 17405 25347 17463 25353
rect 17405 25313 17417 25347
rect 17451 25344 17463 25347
rect 17494 25344 17500 25356
rect 17451 25316 17500 25344
rect 17451 25313 17463 25316
rect 17405 25307 17463 25313
rect 17494 25304 17500 25316
rect 17552 25304 17558 25356
rect 20625 25347 20683 25353
rect 20625 25313 20637 25347
rect 20671 25344 20683 25347
rect 20714 25344 20720 25356
rect 20671 25316 20720 25344
rect 20671 25313 20683 25316
rect 20625 25307 20683 25313
rect 20714 25304 20720 25316
rect 20772 25304 20778 25356
rect 21358 25304 21364 25356
rect 21416 25344 21422 25356
rect 21416 25316 23888 25344
rect 21416 25304 21422 25316
rect 13906 25276 13912 25288
rect 7837 25239 7895 25245
rect 10796 25248 13912 25276
rect 9493 25211 9551 25217
rect 9493 25177 9505 25211
rect 9539 25208 9551 25211
rect 9766 25208 9772 25220
rect 9539 25180 9772 25208
rect 9539 25177 9551 25180
rect 9493 25171 9551 25177
rect 9766 25168 9772 25180
rect 9824 25168 9830 25220
rect 10796 25140 10824 25248
rect 13906 25236 13912 25248
rect 13964 25276 13970 25288
rect 13964 25248 14780 25276
rect 13964 25236 13970 25248
rect 11517 25211 11575 25217
rect 11517 25177 11529 25211
rect 11563 25208 11575 25211
rect 12529 25211 12587 25217
rect 12529 25208 12541 25211
rect 11563 25180 12541 25208
rect 11563 25177 11575 25180
rect 11517 25171 11575 25177
rect 12529 25177 12541 25180
rect 12575 25177 12587 25211
rect 12529 25171 12587 25177
rect 13538 25168 13544 25220
rect 13596 25208 13602 25220
rect 13722 25208 13728 25220
rect 13596 25180 13728 25208
rect 13596 25168 13602 25180
rect 13722 25168 13728 25180
rect 13780 25168 13786 25220
rect 14752 25208 14780 25248
rect 14826 25236 14832 25288
rect 14884 25276 14890 25288
rect 14921 25279 14979 25285
rect 14921 25276 14933 25279
rect 14884 25248 14933 25276
rect 14884 25236 14890 25248
rect 14921 25245 14933 25248
rect 14967 25245 14979 25279
rect 14921 25239 14979 25245
rect 15013 25279 15071 25285
rect 15013 25245 15025 25279
rect 15059 25276 15071 25279
rect 15470 25276 15476 25288
rect 15059 25248 15476 25276
rect 15059 25245 15071 25248
rect 15013 25239 15071 25245
rect 15470 25236 15476 25248
rect 15528 25236 15534 25288
rect 19702 25236 19708 25288
rect 19760 25276 19766 25288
rect 23860 25285 23888 25316
rect 20349 25279 20407 25285
rect 20349 25276 20361 25279
rect 19760 25248 20361 25276
rect 19760 25236 19766 25248
rect 20349 25245 20361 25248
rect 20395 25245 20407 25279
rect 22557 25279 22615 25285
rect 22557 25276 22569 25279
rect 20349 25239 20407 25245
rect 22112 25248 22569 25276
rect 16485 25211 16543 25217
rect 16485 25208 16497 25211
rect 14752 25180 16497 25208
rect 16485 25177 16497 25180
rect 16531 25208 16543 25211
rect 17129 25211 17187 25217
rect 17129 25208 17141 25211
rect 16531 25180 17141 25208
rect 16531 25177 16543 25180
rect 16485 25171 16543 25177
rect 17129 25177 17141 25180
rect 17175 25208 17187 25211
rect 18598 25208 18604 25220
rect 17175 25180 18604 25208
rect 17175 25177 17187 25180
rect 17129 25171 17187 25177
rect 18598 25168 18604 25180
rect 18656 25168 18662 25220
rect 21634 25168 21640 25220
rect 21692 25168 21698 25220
rect 22112 25152 22140 25248
rect 22557 25245 22569 25248
rect 22603 25245 22615 25279
rect 22557 25239 22615 25245
rect 23845 25279 23903 25285
rect 23845 25245 23857 25279
rect 23891 25245 23903 25279
rect 23845 25239 23903 25245
rect 24486 25236 24492 25288
rect 24544 25276 24550 25288
rect 24857 25279 24915 25285
rect 24857 25276 24869 25279
rect 24544 25248 24869 25276
rect 24544 25236 24550 25248
rect 24857 25245 24869 25248
rect 24903 25245 24915 25279
rect 24857 25239 24915 25245
rect 6748 25112 10824 25140
rect 5445 25103 5503 25109
rect 12066 25100 12072 25152
rect 12124 25140 12130 25152
rect 12434 25140 12440 25152
rect 12124 25112 12440 25140
rect 12124 25100 12130 25112
rect 12434 25100 12440 25112
rect 12492 25100 12498 25152
rect 14553 25143 14611 25149
rect 14553 25109 14565 25143
rect 14599 25140 14611 25143
rect 14918 25140 14924 25152
rect 14599 25112 14924 25140
rect 14599 25109 14611 25112
rect 14553 25103 14611 25109
rect 14918 25100 14924 25112
rect 14976 25100 14982 25152
rect 16758 25100 16764 25152
rect 16816 25100 16822 25152
rect 17402 25100 17408 25152
rect 17460 25140 17466 25152
rect 17586 25140 17592 25152
rect 17460 25112 17592 25140
rect 17460 25100 17466 25112
rect 17586 25100 17592 25112
rect 17644 25100 17650 25152
rect 22094 25100 22100 25152
rect 22152 25100 22158 25152
rect 23934 25100 23940 25152
rect 23992 25100 23998 25152
rect 24670 25100 24676 25152
rect 24728 25100 24734 25152
rect 1104 25050 25852 25072
rect 1104 24998 7950 25050
rect 8002 24998 8014 25050
rect 8066 24998 8078 25050
rect 8130 24998 8142 25050
rect 8194 24998 8206 25050
rect 8258 24998 17950 25050
rect 18002 24998 18014 25050
rect 18066 24998 18078 25050
rect 18130 24998 18142 25050
rect 18194 24998 18206 25050
rect 18258 24998 25852 25050
rect 1104 24976 25852 24998
rect 7742 24896 7748 24948
rect 7800 24896 7806 24948
rect 9950 24896 9956 24948
rect 10008 24896 10014 24948
rect 11333 24939 11391 24945
rect 11333 24905 11345 24939
rect 11379 24936 11391 24939
rect 11422 24936 11428 24948
rect 11379 24908 11428 24936
rect 11379 24905 11391 24908
rect 11333 24899 11391 24905
rect 11422 24896 11428 24908
rect 11480 24936 11486 24948
rect 12066 24936 12072 24948
rect 11480 24908 12072 24936
rect 11480 24896 11486 24908
rect 12066 24896 12072 24908
rect 12124 24936 12130 24948
rect 12253 24939 12311 24945
rect 12253 24936 12265 24939
rect 12124 24908 12265 24936
rect 12124 24896 12130 24908
rect 12253 24905 12265 24908
rect 12299 24905 12311 24939
rect 12253 24899 12311 24905
rect 12710 24896 12716 24948
rect 12768 24936 12774 24948
rect 18322 24936 18328 24948
rect 12768 24908 18328 24936
rect 12768 24896 12774 24908
rect 18322 24896 18328 24908
rect 18380 24896 18386 24948
rect 19426 24896 19432 24948
rect 19484 24936 19490 24948
rect 19981 24939 20039 24945
rect 19981 24936 19993 24939
rect 19484 24908 19993 24936
rect 19484 24896 19490 24908
rect 19981 24905 19993 24908
rect 20027 24905 20039 24939
rect 19981 24899 20039 24905
rect 21634 24896 21640 24948
rect 21692 24936 21698 24948
rect 22005 24939 22063 24945
rect 22005 24936 22017 24939
rect 21692 24908 22017 24936
rect 21692 24896 21698 24908
rect 22005 24905 22017 24908
rect 22051 24936 22063 24939
rect 23658 24936 23664 24948
rect 22051 24908 23664 24936
rect 22051 24905 22063 24908
rect 22005 24899 22063 24905
rect 23658 24896 23664 24908
rect 23716 24936 23722 24948
rect 25041 24939 25099 24945
rect 25041 24936 25053 24939
rect 23716 24908 25053 24936
rect 23716 24896 23722 24908
rect 25041 24905 25053 24908
rect 25087 24936 25099 24939
rect 25130 24936 25136 24948
rect 25087 24908 25136 24936
rect 25087 24905 25099 24908
rect 25041 24899 25099 24905
rect 25130 24896 25136 24908
rect 25188 24896 25194 24948
rect 4246 24828 4252 24880
rect 4304 24828 4310 24880
rect 7760 24868 7788 24896
rect 7760 24840 8800 24868
rect 6549 24803 6607 24809
rect 5382 24772 6132 24800
rect 1673 24735 1731 24741
rect 1673 24701 1685 24735
rect 1719 24701 1731 24735
rect 1673 24695 1731 24701
rect 1857 24735 1915 24741
rect 1857 24701 1869 24735
rect 1903 24732 1915 24735
rect 1946 24732 1952 24744
rect 1903 24704 1952 24732
rect 1903 24701 1915 24704
rect 1857 24695 1915 24701
rect 1688 24664 1716 24695
rect 1946 24692 1952 24704
rect 2004 24692 2010 24744
rect 2866 24692 2872 24744
rect 2924 24692 2930 24744
rect 3970 24692 3976 24744
rect 4028 24692 4034 24744
rect 4338 24692 4344 24744
rect 4396 24732 4402 24744
rect 5721 24735 5779 24741
rect 5721 24732 5733 24735
rect 4396 24704 5733 24732
rect 4396 24692 4402 24704
rect 5721 24701 5733 24704
rect 5767 24701 5779 24735
rect 5721 24695 5779 24701
rect 3878 24664 3884 24676
rect 1688 24636 3884 24664
rect 3878 24624 3884 24636
rect 3936 24624 3942 24676
rect 6104 24608 6132 24772
rect 6549 24769 6561 24803
rect 6595 24800 6607 24803
rect 7742 24800 7748 24812
rect 6595 24772 7748 24800
rect 6595 24769 6607 24772
rect 6549 24763 6607 24769
rect 7742 24760 7748 24772
rect 7800 24760 7806 24812
rect 8662 24760 8668 24812
rect 8720 24760 8726 24812
rect 8772 24800 8800 24840
rect 9306 24828 9312 24880
rect 9364 24868 9370 24880
rect 12161 24871 12219 24877
rect 9364 24840 10824 24868
rect 9364 24828 9370 24840
rect 9861 24803 9919 24809
rect 8772 24772 8892 24800
rect 7558 24692 7564 24744
rect 7616 24732 7622 24744
rect 8021 24735 8079 24741
rect 8021 24732 8033 24735
rect 7616 24704 8033 24732
rect 7616 24692 7622 24704
rect 8021 24701 8033 24704
rect 8067 24732 8079 24735
rect 8754 24732 8760 24744
rect 8067 24704 8760 24732
rect 8067 24701 8079 24704
rect 8021 24695 8079 24701
rect 8754 24692 8760 24704
rect 8812 24692 8818 24744
rect 8864 24741 8892 24772
rect 9861 24769 9873 24803
rect 9907 24800 9919 24803
rect 10689 24803 10747 24809
rect 10689 24800 10701 24803
rect 9907 24772 10701 24800
rect 9907 24769 9919 24772
rect 9861 24763 9919 24769
rect 10689 24769 10701 24772
rect 10735 24769 10747 24803
rect 10796 24800 10824 24840
rect 12161 24837 12173 24871
rect 12207 24868 12219 24871
rect 12434 24868 12440 24880
rect 12207 24840 12440 24868
rect 12207 24837 12219 24840
rect 12161 24831 12219 24837
rect 12434 24828 12440 24840
rect 12492 24828 12498 24880
rect 13280 24840 13492 24868
rect 13280 24800 13308 24840
rect 10796 24772 13308 24800
rect 13357 24803 13415 24809
rect 10689 24763 10747 24769
rect 13357 24769 13369 24803
rect 13403 24769 13415 24803
rect 13464 24800 13492 24840
rect 17494 24828 17500 24880
rect 17552 24868 17558 24880
rect 17589 24871 17647 24877
rect 17589 24868 17601 24871
rect 17552 24840 17601 24868
rect 17552 24828 17558 24840
rect 17589 24837 17601 24840
rect 17635 24837 17647 24871
rect 17589 24831 17647 24837
rect 18046 24828 18052 24880
rect 18104 24828 18110 24880
rect 23290 24828 23296 24880
rect 23348 24828 23354 24880
rect 23676 24868 23704 24896
rect 23676 24840 23782 24868
rect 13464 24772 13584 24800
rect 13357 24763 13415 24769
rect 8849 24735 8907 24741
rect 8849 24701 8861 24735
rect 8895 24701 8907 24735
rect 8849 24695 8907 24701
rect 9398 24692 9404 24744
rect 9456 24732 9462 24744
rect 10045 24735 10103 24741
rect 10045 24732 10057 24735
rect 9456 24704 10057 24732
rect 9456 24692 9462 24704
rect 10045 24701 10057 24704
rect 10091 24701 10103 24735
rect 10045 24695 10103 24701
rect 10318 24692 10324 24744
rect 10376 24732 10382 24744
rect 12345 24735 12403 24741
rect 12345 24732 12357 24735
rect 10376 24704 12357 24732
rect 10376 24692 10382 24704
rect 12345 24701 12357 24704
rect 12391 24701 12403 24735
rect 12345 24695 12403 24701
rect 7650 24624 7656 24676
rect 7708 24664 7714 24676
rect 8297 24667 8355 24673
rect 7708 24636 8064 24664
rect 7708 24624 7714 24636
rect 1946 24556 1952 24608
rect 2004 24596 2010 24608
rect 3786 24596 3792 24608
rect 2004 24568 3792 24596
rect 2004 24556 2010 24568
rect 3786 24556 3792 24568
rect 3844 24556 3850 24608
rect 6086 24556 6092 24608
rect 6144 24556 6150 24608
rect 6822 24556 6828 24608
rect 6880 24596 6886 24608
rect 7193 24599 7251 24605
rect 7193 24596 7205 24599
rect 6880 24568 7205 24596
rect 6880 24556 6886 24568
rect 7193 24565 7205 24568
rect 7239 24565 7251 24599
rect 8036 24596 8064 24636
rect 8297 24633 8309 24667
rect 8343 24664 8355 24667
rect 13372 24664 13400 24763
rect 13446 24692 13452 24744
rect 13504 24692 13510 24744
rect 13556 24741 13584 24772
rect 15378 24760 15384 24812
rect 15436 24800 15442 24812
rect 15933 24803 15991 24809
rect 15933 24800 15945 24803
rect 15436 24772 15945 24800
rect 15436 24760 15442 24772
rect 15933 24769 15945 24772
rect 15979 24769 15991 24803
rect 15933 24763 15991 24769
rect 16025 24803 16083 24809
rect 16025 24769 16037 24803
rect 16071 24800 16083 24803
rect 16071 24772 16344 24800
rect 16071 24769 16083 24772
rect 16025 24763 16083 24769
rect 13541 24735 13599 24741
rect 13541 24701 13553 24735
rect 13587 24701 13599 24735
rect 13541 24695 13599 24701
rect 14921 24735 14979 24741
rect 14921 24701 14933 24735
rect 14967 24732 14979 24735
rect 15746 24732 15752 24744
rect 14967 24704 15752 24732
rect 14967 24701 14979 24704
rect 14921 24695 14979 24701
rect 15746 24692 15752 24704
rect 15804 24692 15810 24744
rect 16209 24735 16267 24741
rect 16209 24701 16221 24735
rect 16255 24701 16267 24735
rect 16316 24732 16344 24772
rect 16390 24760 16396 24812
rect 16448 24800 16454 24812
rect 17126 24800 17132 24812
rect 16448 24772 17132 24800
rect 16448 24760 16454 24772
rect 17126 24760 17132 24772
rect 17184 24800 17190 24812
rect 17313 24803 17371 24809
rect 17313 24800 17325 24803
rect 17184 24772 17325 24800
rect 17184 24760 17190 24772
rect 17313 24769 17325 24772
rect 17359 24769 17371 24803
rect 17313 24763 17371 24769
rect 19886 24760 19892 24812
rect 19944 24800 19950 24812
rect 20073 24803 20131 24809
rect 20073 24800 20085 24803
rect 19944 24772 20085 24800
rect 19944 24760 19950 24772
rect 20073 24769 20085 24772
rect 20119 24769 20131 24803
rect 20073 24763 20131 24769
rect 21913 24803 21971 24809
rect 21913 24769 21925 24803
rect 21959 24800 21971 24803
rect 22554 24800 22560 24812
rect 21959 24772 22560 24800
rect 21959 24769 21971 24772
rect 21913 24763 21971 24769
rect 22554 24760 22560 24772
rect 22612 24760 22618 24812
rect 16758 24732 16764 24744
rect 16316 24704 16764 24732
rect 16209 24695 16267 24701
rect 8343 24636 13400 24664
rect 16224 24664 16252 24695
rect 16758 24692 16764 24704
rect 16816 24692 16822 24744
rect 17954 24692 17960 24744
rect 18012 24732 18018 24744
rect 19061 24735 19119 24741
rect 19061 24732 19073 24735
rect 18012 24704 19073 24732
rect 18012 24692 18018 24704
rect 19061 24701 19073 24704
rect 19107 24701 19119 24735
rect 19061 24695 19119 24701
rect 20257 24735 20315 24741
rect 20257 24701 20269 24735
rect 20303 24732 20315 24735
rect 22094 24732 22100 24744
rect 20303 24704 22100 24732
rect 20303 24701 20315 24704
rect 20257 24695 20315 24701
rect 22094 24692 22100 24704
rect 22152 24692 22158 24744
rect 22830 24692 22836 24744
rect 22888 24732 22894 24744
rect 23017 24735 23075 24741
rect 23017 24732 23029 24735
rect 22888 24704 23029 24732
rect 22888 24692 22894 24704
rect 23017 24701 23029 24704
rect 23063 24701 23075 24735
rect 23017 24695 23075 24701
rect 16224 24636 17356 24664
rect 8343 24633 8355 24636
rect 8297 24627 8355 24633
rect 9493 24599 9551 24605
rect 9493 24596 9505 24599
rect 8036 24568 9505 24596
rect 7193 24559 7251 24565
rect 9493 24565 9505 24568
rect 9539 24565 9551 24599
rect 9493 24559 9551 24565
rect 10778 24556 10784 24608
rect 10836 24596 10842 24608
rect 11793 24599 11851 24605
rect 11793 24596 11805 24599
rect 10836 24568 11805 24596
rect 10836 24556 10842 24568
rect 11793 24565 11805 24568
rect 11839 24565 11851 24599
rect 11793 24559 11851 24565
rect 12989 24599 13047 24605
rect 12989 24565 13001 24599
rect 13035 24596 13047 24599
rect 15194 24596 15200 24608
rect 13035 24568 15200 24596
rect 13035 24565 13047 24568
rect 12989 24559 13047 24565
rect 15194 24556 15200 24568
rect 15252 24556 15258 24608
rect 15565 24599 15623 24605
rect 15565 24565 15577 24599
rect 15611 24596 15623 24599
rect 17218 24596 17224 24608
rect 15611 24568 17224 24596
rect 15611 24565 15623 24568
rect 15565 24559 15623 24565
rect 17218 24556 17224 24568
rect 17276 24556 17282 24608
rect 17328 24596 17356 24636
rect 18690 24624 18696 24676
rect 18748 24664 18754 24676
rect 19613 24667 19671 24673
rect 19613 24664 19625 24667
rect 18748 24636 19625 24664
rect 18748 24624 18754 24636
rect 19613 24633 19625 24636
rect 19659 24633 19671 24667
rect 19613 24627 19671 24633
rect 20346 24624 20352 24676
rect 20404 24664 20410 24676
rect 22373 24667 22431 24673
rect 22373 24664 22385 24667
rect 20404 24636 22385 24664
rect 20404 24624 20410 24636
rect 22373 24633 22385 24636
rect 22419 24633 22431 24667
rect 22373 24627 22431 24633
rect 17954 24596 17960 24608
rect 17328 24568 17960 24596
rect 17954 24556 17960 24568
rect 18012 24556 18018 24608
rect 23750 24556 23756 24608
rect 23808 24596 23814 24608
rect 24578 24596 24584 24608
rect 23808 24568 24584 24596
rect 23808 24556 23814 24568
rect 24578 24556 24584 24568
rect 24636 24596 24642 24608
rect 24765 24599 24823 24605
rect 24765 24596 24777 24599
rect 24636 24568 24777 24596
rect 24636 24556 24642 24568
rect 24765 24565 24777 24568
rect 24811 24565 24823 24599
rect 24765 24559 24823 24565
rect 1104 24506 25852 24528
rect 1104 24454 2950 24506
rect 3002 24454 3014 24506
rect 3066 24454 3078 24506
rect 3130 24454 3142 24506
rect 3194 24454 3206 24506
rect 3258 24454 12950 24506
rect 13002 24454 13014 24506
rect 13066 24454 13078 24506
rect 13130 24454 13142 24506
rect 13194 24454 13206 24506
rect 13258 24454 22950 24506
rect 23002 24454 23014 24506
rect 23066 24454 23078 24506
rect 23130 24454 23142 24506
rect 23194 24454 23206 24506
rect 23258 24454 25852 24506
rect 1104 24432 25852 24454
rect 4798 24352 4804 24404
rect 4856 24392 4862 24404
rect 5721 24395 5779 24401
rect 5721 24392 5733 24395
rect 4856 24364 5733 24392
rect 4856 24352 4862 24364
rect 5721 24361 5733 24364
rect 5767 24361 5779 24395
rect 5721 24355 5779 24361
rect 6454 24352 6460 24404
rect 6512 24352 6518 24404
rect 7466 24352 7472 24404
rect 7524 24392 7530 24404
rect 8570 24392 8576 24404
rect 7524 24364 8576 24392
rect 7524 24352 7530 24364
rect 8570 24352 8576 24364
rect 8628 24352 8634 24404
rect 9950 24352 9956 24404
rect 10008 24392 10014 24404
rect 10321 24395 10379 24401
rect 10321 24392 10333 24395
rect 10008 24364 10333 24392
rect 10008 24352 10014 24364
rect 10321 24361 10333 24364
rect 10367 24392 10379 24395
rect 11330 24392 11336 24404
rect 10367 24364 11336 24392
rect 10367 24361 10379 24364
rect 10321 24355 10379 24361
rect 11330 24352 11336 24364
rect 11388 24352 11394 24404
rect 12434 24352 12440 24404
rect 12492 24392 12498 24404
rect 12986 24392 12992 24404
rect 12492 24364 12992 24392
rect 12492 24352 12498 24364
rect 12986 24352 12992 24364
rect 13044 24352 13050 24404
rect 16114 24352 16120 24404
rect 16172 24392 16178 24404
rect 17405 24395 17463 24401
rect 17405 24392 17417 24395
rect 16172 24364 17417 24392
rect 16172 24352 16178 24364
rect 17405 24361 17417 24364
rect 17451 24361 17463 24395
rect 17405 24355 17463 24361
rect 25130 24352 25136 24404
rect 25188 24352 25194 24404
rect 6086 24284 6092 24336
rect 6144 24324 6150 24336
rect 8478 24324 8484 24336
rect 6144 24296 8484 24324
rect 6144 24284 6150 24296
rect 8478 24284 8484 24296
rect 8536 24284 8542 24336
rect 9582 24284 9588 24336
rect 9640 24324 9646 24336
rect 10505 24327 10563 24333
rect 10505 24324 10517 24327
rect 9640 24296 10517 24324
rect 9640 24284 9646 24296
rect 10505 24293 10517 24296
rect 10551 24293 10563 24327
rect 10505 24287 10563 24293
rect 12713 24327 12771 24333
rect 12713 24293 12725 24327
rect 12759 24324 12771 24327
rect 14090 24324 14096 24336
rect 12759 24296 14096 24324
rect 12759 24293 12771 24296
rect 12713 24287 12771 24293
rect 14090 24284 14096 24296
rect 14148 24284 14154 24336
rect 19981 24327 20039 24333
rect 19981 24293 19993 24327
rect 20027 24324 20039 24327
rect 23474 24324 23480 24336
rect 20027 24296 23480 24324
rect 20027 24293 20039 24296
rect 19981 24287 20039 24293
rect 23474 24284 23480 24296
rect 23532 24284 23538 24336
rect 2222 24148 2228 24200
rect 2280 24148 2286 24200
rect 3970 24148 3976 24200
rect 4028 24148 4034 24200
rect 6104 24188 6132 24284
rect 7098 24216 7104 24268
rect 7156 24216 7162 24268
rect 8662 24216 8668 24268
rect 8720 24256 8726 24268
rect 9125 24259 9183 24265
rect 9125 24256 9137 24259
rect 8720 24228 9137 24256
rect 8720 24216 8726 24228
rect 9125 24225 9137 24228
rect 9171 24225 9183 24259
rect 9125 24219 9183 24225
rect 9950 24216 9956 24268
rect 10008 24256 10014 24268
rect 10965 24259 11023 24265
rect 10965 24256 10977 24259
rect 10008 24228 10977 24256
rect 10008 24216 10014 24228
rect 10965 24225 10977 24228
rect 11011 24225 11023 24259
rect 10965 24219 11023 24225
rect 11238 24216 11244 24268
rect 11296 24216 11302 24268
rect 12434 24216 12440 24268
rect 12492 24256 12498 24268
rect 14921 24259 14979 24265
rect 14921 24256 14933 24259
rect 12492 24228 14933 24256
rect 12492 24216 12498 24228
rect 14921 24225 14933 24228
rect 14967 24225 14979 24259
rect 14921 24219 14979 24225
rect 15657 24259 15715 24265
rect 15657 24225 15669 24259
rect 15703 24256 15715 24259
rect 16390 24256 16396 24268
rect 15703 24228 16396 24256
rect 15703 24225 15715 24228
rect 15657 24219 15715 24225
rect 16390 24216 16396 24228
rect 16448 24216 16454 24268
rect 20346 24216 20352 24268
rect 20404 24256 20410 24268
rect 20441 24259 20499 24265
rect 20441 24256 20453 24259
rect 20404 24228 20453 24256
rect 20404 24216 20410 24228
rect 20441 24225 20453 24228
rect 20487 24225 20499 24259
rect 20441 24219 20499 24225
rect 20530 24216 20536 24268
rect 20588 24216 20594 24268
rect 21910 24216 21916 24268
rect 21968 24216 21974 24268
rect 22005 24259 22063 24265
rect 22005 24225 22017 24259
rect 22051 24256 22063 24259
rect 23750 24256 23756 24268
rect 22051 24228 23756 24256
rect 22051 24225 22063 24228
rect 22005 24219 22063 24225
rect 23750 24216 23756 24228
rect 23808 24216 23814 24268
rect 23845 24259 23903 24265
rect 23845 24225 23857 24259
rect 23891 24256 23903 24259
rect 24854 24256 24860 24268
rect 23891 24228 24860 24256
rect 23891 24225 23903 24228
rect 23845 24219 23903 24225
rect 24854 24216 24860 24228
rect 24912 24216 24918 24268
rect 5382 24160 6132 24188
rect 12342 24148 12348 24200
rect 12400 24188 12406 24200
rect 13173 24191 13231 24197
rect 13173 24188 13185 24191
rect 12400 24160 13185 24188
rect 12400 24148 12406 24160
rect 13173 24157 13185 24160
rect 13219 24157 13231 24191
rect 13173 24151 13231 24157
rect 14090 24148 14096 24200
rect 14148 24188 14154 24200
rect 14277 24191 14335 24197
rect 14277 24188 14289 24191
rect 14148 24160 14289 24188
rect 14148 24148 14154 24160
rect 14277 24157 14289 24160
rect 14323 24188 14335 24191
rect 14826 24188 14832 24200
rect 14323 24160 14832 24188
rect 14323 24157 14335 24160
rect 14277 24151 14335 24157
rect 14826 24148 14832 24160
rect 14884 24148 14890 24200
rect 17862 24148 17868 24200
rect 17920 24148 17926 24200
rect 19150 24148 19156 24200
rect 19208 24188 19214 24200
rect 19613 24191 19671 24197
rect 19613 24188 19625 24191
rect 19208 24160 19625 24188
rect 19208 24148 19214 24160
rect 19613 24157 19625 24160
rect 19659 24157 19671 24191
rect 19613 24151 19671 24157
rect 21821 24191 21879 24197
rect 21821 24157 21833 24191
rect 21867 24188 21879 24191
rect 22370 24188 22376 24200
rect 21867 24160 22376 24188
rect 21867 24157 21879 24160
rect 21821 24151 21879 24157
rect 4246 24080 4252 24132
rect 4304 24080 4310 24132
rect 9674 24080 9680 24132
rect 9732 24120 9738 24132
rect 10137 24123 10195 24129
rect 10137 24120 10149 24123
rect 9732 24092 10149 24120
rect 9732 24080 9738 24092
rect 10137 24089 10149 24092
rect 10183 24120 10195 24123
rect 10183 24092 10732 24120
rect 10183 24089 10195 24092
rect 10137 24083 10195 24089
rect 1854 24012 1860 24064
rect 1912 24052 1918 24064
rect 2041 24055 2099 24061
rect 2041 24052 2053 24055
rect 1912 24024 2053 24052
rect 1912 24012 1918 24024
rect 2041 24021 2053 24024
rect 2087 24021 2099 24055
rect 2041 24015 2099 24021
rect 6730 24012 6736 24064
rect 6788 24052 6794 24064
rect 6825 24055 6883 24061
rect 6825 24052 6837 24055
rect 6788 24024 6837 24052
rect 6788 24012 6794 24024
rect 6825 24021 6837 24024
rect 6871 24021 6883 24055
rect 6825 24015 6883 24021
rect 6917 24055 6975 24061
rect 6917 24021 6929 24055
rect 6963 24052 6975 24055
rect 9122 24052 9128 24064
rect 6963 24024 9128 24052
rect 6963 24021 6975 24024
rect 6917 24015 6975 24021
rect 9122 24012 9128 24024
rect 9180 24012 9186 24064
rect 10704 24052 10732 24092
rect 12986 24080 12992 24132
rect 13044 24080 13050 24132
rect 15933 24123 15991 24129
rect 15933 24089 15945 24123
rect 15979 24089 15991 24123
rect 15933 24083 15991 24089
rect 13354 24052 13360 24064
rect 10704 24024 13360 24052
rect 13354 24012 13360 24024
rect 13412 24012 13418 24064
rect 13446 24012 13452 24064
rect 13504 24052 13510 24064
rect 13722 24052 13728 24064
rect 13504 24024 13728 24052
rect 13504 24012 13510 24024
rect 13722 24012 13728 24024
rect 13780 24012 13786 24064
rect 15948 24052 15976 24083
rect 16574 24080 16580 24132
rect 16632 24080 16638 24132
rect 18509 24123 18567 24129
rect 18509 24120 18521 24123
rect 17236 24092 18521 24120
rect 17236 24052 17264 24092
rect 18509 24089 18521 24092
rect 18555 24089 18567 24123
rect 18509 24083 18567 24089
rect 15948 24024 17264 24052
rect 17862 24012 17868 24064
rect 17920 24052 17926 24064
rect 18046 24052 18052 24064
rect 17920 24024 18052 24052
rect 17920 24012 17926 24024
rect 18046 24012 18052 24024
rect 18104 24052 18110 24064
rect 18785 24055 18843 24061
rect 18785 24052 18797 24055
rect 18104 24024 18797 24052
rect 18104 24012 18110 24024
rect 18785 24021 18797 24024
rect 18831 24052 18843 24055
rect 19245 24055 19303 24061
rect 19245 24052 19257 24055
rect 18831 24024 19257 24052
rect 18831 24021 18843 24024
rect 18785 24015 18843 24021
rect 19245 24021 19257 24024
rect 19291 24021 19303 24055
rect 19628 24052 19656 24151
rect 22370 24148 22376 24160
rect 22428 24148 22434 24200
rect 22833 24191 22891 24197
rect 22833 24157 22845 24191
rect 22879 24157 22891 24191
rect 22833 24151 22891 24157
rect 19886 24080 19892 24132
rect 19944 24120 19950 24132
rect 22848 24120 22876 24151
rect 23566 24148 23572 24200
rect 23624 24188 23630 24200
rect 24673 24191 24731 24197
rect 24673 24188 24685 24191
rect 23624 24160 24685 24188
rect 23624 24148 23630 24160
rect 24673 24157 24685 24160
rect 24719 24157 24731 24191
rect 24673 24151 24731 24157
rect 25038 24120 25044 24132
rect 19944 24092 22094 24120
rect 22848 24092 25044 24120
rect 19944 24080 19950 24092
rect 20349 24055 20407 24061
rect 20349 24052 20361 24055
rect 19628 24024 20361 24052
rect 19245 24015 19303 24021
rect 20349 24021 20361 24024
rect 20395 24021 20407 24055
rect 20349 24015 20407 24021
rect 21453 24055 21511 24061
rect 21453 24021 21465 24055
rect 21499 24052 21511 24055
rect 21726 24052 21732 24064
rect 21499 24024 21732 24052
rect 21499 24021 21511 24024
rect 21453 24015 21511 24021
rect 21726 24012 21732 24024
rect 21784 24012 21790 24064
rect 22066 24052 22094 24092
rect 25038 24080 25044 24092
rect 25096 24080 25102 24132
rect 22646 24052 22652 24064
rect 22066 24024 22652 24052
rect 22646 24012 22652 24024
rect 22704 24012 22710 24064
rect 24394 24012 24400 24064
rect 24452 24052 24458 24064
rect 24765 24055 24823 24061
rect 24765 24052 24777 24055
rect 24452 24024 24777 24052
rect 24452 24012 24458 24024
rect 24765 24021 24777 24024
rect 24811 24021 24823 24055
rect 24765 24015 24823 24021
rect 1104 23962 25852 23984
rect 1104 23910 7950 23962
rect 8002 23910 8014 23962
rect 8066 23910 8078 23962
rect 8130 23910 8142 23962
rect 8194 23910 8206 23962
rect 8258 23910 17950 23962
rect 18002 23910 18014 23962
rect 18066 23910 18078 23962
rect 18130 23910 18142 23962
rect 18194 23910 18206 23962
rect 18258 23910 25852 23962
rect 1104 23888 25852 23910
rect 3602 23808 3608 23860
rect 3660 23848 3666 23860
rect 3835 23851 3893 23857
rect 3835 23848 3847 23851
rect 3660 23820 3847 23848
rect 3660 23808 3666 23820
rect 3835 23817 3847 23820
rect 3881 23817 3893 23851
rect 3835 23811 3893 23817
rect 4246 23808 4252 23860
rect 4304 23848 4310 23860
rect 5537 23851 5595 23857
rect 5537 23848 5549 23851
rect 4304 23820 5549 23848
rect 4304 23808 4310 23820
rect 5537 23817 5549 23820
rect 5583 23817 5595 23851
rect 5537 23811 5595 23817
rect 7098 23808 7104 23860
rect 7156 23848 7162 23860
rect 8297 23851 8355 23857
rect 8297 23848 8309 23851
rect 7156 23820 8309 23848
rect 7156 23808 7162 23820
rect 8297 23817 8309 23820
rect 8343 23817 8355 23851
rect 8297 23811 8355 23817
rect 8478 23808 8484 23860
rect 8536 23848 8542 23860
rect 8573 23851 8631 23857
rect 8573 23848 8585 23851
rect 8536 23820 8585 23848
rect 8536 23808 8542 23820
rect 8573 23817 8585 23820
rect 8619 23817 8631 23851
rect 8573 23811 8631 23817
rect 9582 23808 9588 23860
rect 9640 23808 9646 23860
rect 9674 23808 9680 23860
rect 9732 23808 9738 23860
rect 10873 23851 10931 23857
rect 10873 23848 10885 23851
rect 9784 23820 10885 23848
rect 6822 23740 6828 23792
rect 6880 23740 6886 23792
rect 8496 23780 8524 23808
rect 8050 23752 8524 23780
rect 9306 23740 9312 23792
rect 9364 23780 9370 23792
rect 9600 23780 9628 23808
rect 9784 23780 9812 23820
rect 10873 23817 10885 23820
rect 10919 23817 10931 23851
rect 10873 23811 10931 23817
rect 12529 23851 12587 23857
rect 12529 23817 12541 23851
rect 12575 23848 12587 23851
rect 13446 23848 13452 23860
rect 12575 23820 13452 23848
rect 12575 23817 12587 23820
rect 12529 23811 12587 23817
rect 13446 23808 13452 23820
rect 13504 23808 13510 23860
rect 13725 23851 13783 23857
rect 13725 23817 13737 23851
rect 13771 23848 13783 23851
rect 13998 23848 14004 23860
rect 13771 23820 14004 23848
rect 13771 23817 13783 23820
rect 13725 23811 13783 23817
rect 13998 23808 14004 23820
rect 14056 23848 14062 23860
rect 14369 23851 14427 23857
rect 14369 23848 14381 23851
rect 14056 23820 14381 23848
rect 14056 23808 14062 23820
rect 14369 23817 14381 23820
rect 14415 23848 14427 23851
rect 14458 23848 14464 23860
rect 14415 23820 14464 23848
rect 14415 23817 14427 23820
rect 14369 23811 14427 23817
rect 14458 23808 14464 23820
rect 14516 23808 14522 23860
rect 14645 23851 14703 23857
rect 14645 23817 14657 23851
rect 14691 23848 14703 23851
rect 14734 23848 14740 23860
rect 14691 23820 14740 23848
rect 14691 23817 14703 23820
rect 14645 23811 14703 23817
rect 13817 23783 13875 23789
rect 9364 23752 9812 23780
rect 11808 23752 12756 23780
rect 9364 23740 9370 23752
rect 2314 23672 2320 23724
rect 2372 23712 2378 23724
rect 3732 23715 3790 23721
rect 3732 23712 3744 23715
rect 2372 23684 3744 23712
rect 2372 23672 2378 23684
rect 3732 23681 3744 23684
rect 3778 23681 3790 23715
rect 3732 23675 3790 23681
rect 4893 23715 4951 23721
rect 4893 23681 4905 23715
rect 4939 23712 4951 23715
rect 5902 23712 5908 23724
rect 4939 23684 5908 23712
rect 4939 23681 4951 23684
rect 4893 23675 4951 23681
rect 5902 23672 5908 23684
rect 5960 23672 5966 23724
rect 9582 23672 9588 23724
rect 9640 23672 9646 23724
rect 10781 23715 10839 23721
rect 10781 23681 10793 23715
rect 10827 23712 10839 23715
rect 11698 23712 11704 23724
rect 10827 23684 11704 23712
rect 10827 23681 10839 23684
rect 10781 23675 10839 23681
rect 11698 23672 11704 23684
rect 11756 23672 11762 23724
rect 3970 23604 3976 23656
rect 4028 23644 4034 23656
rect 6546 23644 6552 23656
rect 4028 23616 6552 23644
rect 4028 23604 4034 23616
rect 6546 23604 6552 23616
rect 6604 23604 6610 23656
rect 7190 23604 7196 23656
rect 7248 23644 7254 23656
rect 7248 23616 9260 23644
rect 7248 23604 7254 23616
rect 6564 23508 6592 23604
rect 9232 23585 9260 23616
rect 9858 23604 9864 23656
rect 9916 23604 9922 23656
rect 10594 23604 10600 23656
rect 10652 23644 10658 23656
rect 10965 23647 11023 23653
rect 10965 23644 10977 23647
rect 10652 23616 10977 23644
rect 10652 23604 10658 23616
rect 10965 23613 10977 23616
rect 11011 23613 11023 23647
rect 10965 23607 11023 23613
rect 11054 23604 11060 23656
rect 11112 23644 11118 23656
rect 11808 23653 11836 23752
rect 12621 23715 12679 23721
rect 12621 23712 12633 23715
rect 12084 23684 12633 23712
rect 11793 23647 11851 23653
rect 11793 23644 11805 23647
rect 11112 23616 11805 23644
rect 11112 23604 11118 23616
rect 11793 23613 11805 23616
rect 11839 23613 11851 23647
rect 11793 23607 11851 23613
rect 9217 23579 9275 23585
rect 9217 23545 9229 23579
rect 9263 23545 9275 23579
rect 9217 23539 9275 23545
rect 10413 23579 10471 23585
rect 10413 23545 10425 23579
rect 10459 23576 10471 23579
rect 11974 23576 11980 23588
rect 10459 23548 11980 23576
rect 10459 23545 10471 23548
rect 10413 23539 10471 23545
rect 11974 23536 11980 23548
rect 12032 23536 12038 23588
rect 7834 23508 7840 23520
rect 6564 23480 7840 23508
rect 7834 23468 7840 23480
rect 7892 23468 7898 23520
rect 9030 23468 9036 23520
rect 9088 23508 9094 23520
rect 9766 23508 9772 23520
rect 9088 23480 9772 23508
rect 9088 23468 9094 23480
rect 9766 23468 9772 23480
rect 9824 23508 9830 23520
rect 11609 23511 11667 23517
rect 11609 23508 11621 23511
rect 9824 23480 11621 23508
rect 9824 23468 9830 23480
rect 11609 23477 11621 23480
rect 11655 23508 11667 23511
rect 12084 23508 12112 23684
rect 12621 23681 12633 23684
rect 12667 23681 12679 23715
rect 12621 23675 12679 23681
rect 12158 23604 12164 23656
rect 12216 23644 12222 23656
rect 12728 23653 12756 23752
rect 13817 23749 13829 23783
rect 13863 23780 13875 23783
rect 14660 23780 14688 23811
rect 14734 23808 14740 23820
rect 14792 23808 14798 23860
rect 15010 23808 15016 23860
rect 15068 23808 15074 23860
rect 15378 23808 15384 23860
rect 15436 23808 15442 23860
rect 15746 23808 15752 23860
rect 15804 23808 15810 23860
rect 17218 23808 17224 23860
rect 17276 23808 17282 23860
rect 17313 23851 17371 23857
rect 17313 23817 17325 23851
rect 17359 23848 17371 23851
rect 17678 23848 17684 23860
rect 17359 23820 17684 23848
rect 17359 23817 17371 23820
rect 17313 23811 17371 23817
rect 17678 23808 17684 23820
rect 17736 23808 17742 23860
rect 18049 23851 18107 23857
rect 18049 23817 18061 23851
rect 18095 23848 18107 23851
rect 19886 23848 19892 23860
rect 18095 23820 19892 23848
rect 18095 23817 18107 23820
rect 18049 23811 18107 23817
rect 19886 23808 19892 23820
rect 19944 23808 19950 23860
rect 20254 23808 20260 23860
rect 20312 23848 20318 23860
rect 20622 23848 20628 23860
rect 20312 23820 20628 23848
rect 20312 23808 20318 23820
rect 20622 23808 20628 23820
rect 20680 23848 20686 23860
rect 21453 23851 21511 23857
rect 21453 23848 21465 23851
rect 20680 23820 21465 23848
rect 20680 23808 20686 23820
rect 21453 23817 21465 23820
rect 21499 23817 21511 23851
rect 21453 23811 21511 23817
rect 21634 23808 21640 23860
rect 21692 23848 21698 23860
rect 21821 23851 21879 23857
rect 21821 23848 21833 23851
rect 21692 23820 21833 23848
rect 21692 23808 21698 23820
rect 21821 23817 21833 23820
rect 21867 23817 21879 23851
rect 21821 23811 21879 23817
rect 24026 23808 24032 23860
rect 24084 23848 24090 23860
rect 24578 23848 24584 23860
rect 24084 23820 24584 23848
rect 24084 23808 24090 23820
rect 24578 23808 24584 23820
rect 24636 23808 24642 23860
rect 13863 23752 14688 23780
rect 15028 23780 15056 23808
rect 15841 23783 15899 23789
rect 15841 23780 15853 23783
rect 15028 23752 15853 23780
rect 13863 23749 13875 23752
rect 13817 23743 13875 23749
rect 15841 23749 15853 23752
rect 15887 23780 15899 23783
rect 19150 23780 19156 23792
rect 15887 23752 19156 23780
rect 15887 23749 15899 23752
rect 15841 23743 15899 23749
rect 19150 23740 19156 23752
rect 19208 23740 19214 23792
rect 19978 23740 19984 23792
rect 20036 23740 20042 23792
rect 21652 23780 21680 23808
rect 21206 23752 21680 23780
rect 22738 23740 22744 23792
rect 22796 23780 22802 23792
rect 23109 23783 23167 23789
rect 23109 23780 23121 23783
rect 22796 23752 23121 23780
rect 22796 23740 22802 23752
rect 23109 23749 23121 23752
rect 23155 23749 23167 23783
rect 23109 23743 23167 23749
rect 23658 23740 23664 23792
rect 23716 23740 23722 23792
rect 25133 23783 25191 23789
rect 25133 23749 25145 23783
rect 25179 23780 25191 23783
rect 25406 23780 25412 23792
rect 25179 23752 25412 23780
rect 25179 23749 25191 23752
rect 25133 23743 25191 23749
rect 25406 23740 25412 23752
rect 25464 23740 25470 23792
rect 12986 23672 12992 23724
rect 13044 23712 13050 23724
rect 17310 23712 17316 23724
rect 13044 23684 17316 23712
rect 13044 23672 13050 23684
rect 17310 23672 17316 23684
rect 17368 23672 17374 23724
rect 18233 23715 18291 23721
rect 18233 23681 18245 23715
rect 18279 23712 18291 23715
rect 18322 23712 18328 23724
rect 18279 23684 18328 23712
rect 18279 23681 18291 23684
rect 18233 23675 18291 23681
rect 18322 23672 18328 23684
rect 18380 23672 18386 23724
rect 18598 23672 18604 23724
rect 18656 23712 18662 23724
rect 18782 23712 18788 23724
rect 18656 23684 18788 23712
rect 18656 23672 18662 23684
rect 18782 23672 18788 23684
rect 18840 23672 18846 23724
rect 22094 23672 22100 23724
rect 22152 23712 22158 23724
rect 22830 23712 22836 23724
rect 22152 23684 22836 23712
rect 22152 23672 22158 23684
rect 22830 23672 22836 23684
rect 22888 23672 22894 23724
rect 12713 23647 12771 23653
rect 12216 23616 12664 23644
rect 12216 23604 12222 23616
rect 12636 23576 12664 23616
rect 12713 23613 12725 23647
rect 12759 23613 12771 23647
rect 12713 23607 12771 23613
rect 13909 23647 13967 23653
rect 13909 23613 13921 23647
rect 13955 23613 13967 23647
rect 13909 23607 13967 23613
rect 16025 23647 16083 23653
rect 16025 23613 16037 23647
rect 16071 23613 16083 23647
rect 16025 23607 16083 23613
rect 13357 23579 13415 23585
rect 13357 23576 13369 23579
rect 12636 23548 13369 23576
rect 13357 23545 13369 23548
rect 13403 23545 13415 23579
rect 13357 23539 13415 23545
rect 13722 23536 13728 23588
rect 13780 23576 13786 23588
rect 13924 23576 13952 23607
rect 13780 23548 13952 23576
rect 16040 23576 16068 23607
rect 16114 23604 16120 23656
rect 16172 23644 16178 23656
rect 17405 23647 17463 23653
rect 17405 23644 17417 23647
rect 16172 23616 17417 23644
rect 16172 23604 16178 23616
rect 17405 23613 17417 23616
rect 17451 23613 17463 23647
rect 17405 23607 17463 23613
rect 17862 23604 17868 23656
rect 17920 23644 17926 23656
rect 18969 23647 19027 23653
rect 18969 23644 18981 23647
rect 17920 23616 18981 23644
rect 17920 23604 17926 23616
rect 18969 23613 18981 23616
rect 19015 23613 19027 23647
rect 18969 23607 19027 23613
rect 17494 23576 17500 23588
rect 16040 23548 17500 23576
rect 13780 23536 13786 23548
rect 17494 23536 17500 23548
rect 17552 23536 17558 23588
rect 11655 23480 12112 23508
rect 11655 23477 11667 23480
rect 11609 23471 11667 23477
rect 12158 23468 12164 23520
rect 12216 23468 12222 23520
rect 16850 23468 16856 23520
rect 16908 23468 16914 23520
rect 18984 23508 19012 23607
rect 19702 23604 19708 23656
rect 19760 23604 19766 23656
rect 20530 23604 20536 23656
rect 20588 23644 20594 23656
rect 22738 23644 22744 23656
rect 20588 23616 22744 23644
rect 20588 23604 20594 23616
rect 22738 23604 22744 23616
rect 22796 23604 22802 23656
rect 23658 23604 23664 23656
rect 23716 23644 23722 23656
rect 25317 23647 25375 23653
rect 25317 23644 25329 23647
rect 23716 23616 25329 23644
rect 23716 23604 23722 23616
rect 25317 23613 25329 23616
rect 25363 23613 25375 23647
rect 25317 23607 25375 23613
rect 19150 23508 19156 23520
rect 18984 23480 19156 23508
rect 19150 23468 19156 23480
rect 19208 23508 19214 23520
rect 20714 23508 20720 23520
rect 19208 23480 20720 23508
rect 19208 23468 19214 23480
rect 20714 23468 20720 23480
rect 20772 23468 20778 23520
rect 1104 23418 25852 23440
rect 1104 23366 2950 23418
rect 3002 23366 3014 23418
rect 3066 23366 3078 23418
rect 3130 23366 3142 23418
rect 3194 23366 3206 23418
rect 3258 23366 12950 23418
rect 13002 23366 13014 23418
rect 13066 23366 13078 23418
rect 13130 23366 13142 23418
rect 13194 23366 13206 23418
rect 13258 23366 22950 23418
rect 23002 23366 23014 23418
rect 23066 23366 23078 23418
rect 23130 23366 23142 23418
rect 23194 23366 23206 23418
rect 23258 23366 25852 23418
rect 1104 23344 25852 23366
rect 2774 23264 2780 23316
rect 2832 23304 2838 23316
rect 2832 23276 3004 23304
rect 2832 23264 2838 23276
rect 1581 23171 1639 23177
rect 1581 23137 1593 23171
rect 1627 23168 1639 23171
rect 2774 23168 2780 23180
rect 1627 23140 2780 23168
rect 1627 23137 1639 23140
rect 1581 23131 1639 23137
rect 2774 23128 2780 23140
rect 2832 23128 2838 23180
rect 2976 23177 3004 23276
rect 7742 23264 7748 23316
rect 7800 23304 7806 23316
rect 8021 23307 8079 23313
rect 8021 23304 8033 23307
rect 7800 23276 8033 23304
rect 7800 23264 7806 23276
rect 8021 23273 8033 23276
rect 8067 23273 8079 23307
rect 8021 23267 8079 23273
rect 8389 23307 8447 23313
rect 8389 23273 8401 23307
rect 8435 23304 8447 23307
rect 8478 23304 8484 23316
rect 8435 23276 8484 23304
rect 8435 23273 8447 23276
rect 8389 23267 8447 23273
rect 8478 23264 8484 23276
rect 8536 23264 8542 23316
rect 11514 23264 11520 23316
rect 11572 23304 11578 23316
rect 15838 23304 15844 23316
rect 11572 23276 15844 23304
rect 11572 23264 11578 23276
rect 15838 23264 15844 23276
rect 15896 23264 15902 23316
rect 18874 23264 18880 23316
rect 18932 23264 18938 23316
rect 20070 23264 20076 23316
rect 20128 23304 20134 23316
rect 21177 23307 21235 23313
rect 21177 23304 21189 23307
rect 20128 23276 21189 23304
rect 20128 23264 20134 23276
rect 21177 23273 21189 23276
rect 21223 23273 21235 23307
rect 21177 23267 21235 23273
rect 21545 23307 21603 23313
rect 21545 23273 21557 23307
rect 21591 23304 21603 23307
rect 21634 23304 21640 23316
rect 21591 23276 21640 23304
rect 21591 23273 21603 23276
rect 21545 23267 21603 23273
rect 11701 23239 11759 23245
rect 11701 23205 11713 23239
rect 11747 23236 11759 23239
rect 11790 23236 11796 23248
rect 11747 23208 11796 23236
rect 11747 23205 11759 23208
rect 11701 23199 11759 23205
rect 11790 23196 11796 23208
rect 11848 23196 11854 23248
rect 14277 23239 14335 23245
rect 14277 23205 14289 23239
rect 14323 23236 14335 23239
rect 17034 23236 17040 23248
rect 14323 23208 17040 23236
rect 14323 23205 14335 23208
rect 14277 23199 14335 23205
rect 17034 23196 17040 23208
rect 17092 23196 17098 23248
rect 2961 23171 3019 23177
rect 2961 23137 2973 23171
rect 3007 23137 3019 23171
rect 2961 23131 3019 23137
rect 6273 23171 6331 23177
rect 6273 23137 6285 23171
rect 6319 23168 6331 23171
rect 9950 23168 9956 23180
rect 6319 23140 9956 23168
rect 6319 23137 6331 23140
rect 6273 23131 6331 23137
rect 9950 23128 9956 23140
rect 10008 23168 10014 23180
rect 11057 23171 11115 23177
rect 11057 23168 11069 23171
rect 10008 23140 11069 23168
rect 10008 23128 10014 23140
rect 11057 23137 11069 23140
rect 11103 23168 11115 23171
rect 11977 23171 12035 23177
rect 11977 23168 11989 23171
rect 11103 23140 11989 23168
rect 11103 23137 11115 23140
rect 11057 23131 11115 23137
rect 11977 23137 11989 23140
rect 12023 23168 12035 23171
rect 12802 23168 12808 23180
rect 12023 23140 12808 23168
rect 12023 23137 12035 23140
rect 11977 23131 12035 23137
rect 12802 23128 12808 23140
rect 12860 23128 12866 23180
rect 14550 23128 14556 23180
rect 14608 23168 14614 23180
rect 14737 23171 14795 23177
rect 14737 23168 14749 23171
rect 14608 23140 14749 23168
rect 14608 23128 14614 23140
rect 14737 23137 14749 23140
rect 14783 23137 14795 23171
rect 14737 23131 14795 23137
rect 14826 23128 14832 23180
rect 14884 23128 14890 23180
rect 17126 23128 17132 23180
rect 17184 23128 17190 23180
rect 17405 23171 17463 23177
rect 17405 23137 17417 23171
rect 17451 23168 17463 23171
rect 19334 23168 19340 23180
rect 17451 23140 19340 23168
rect 17451 23137 17463 23140
rect 17405 23131 17463 23137
rect 19334 23128 19340 23140
rect 19392 23128 19398 23180
rect 19429 23171 19487 23177
rect 19429 23137 19441 23171
rect 19475 23168 19487 23171
rect 19702 23168 19708 23180
rect 19475 23140 19708 23168
rect 19475 23137 19487 23140
rect 19429 23131 19487 23137
rect 19702 23128 19708 23140
rect 19760 23168 19766 23180
rect 21082 23168 21088 23180
rect 19760 23140 21088 23168
rect 19760 23128 19766 23140
rect 21082 23128 21088 23140
rect 21140 23128 21146 23180
rect 4249 23103 4307 23109
rect 4249 23069 4261 23103
rect 4295 23100 4307 23103
rect 4338 23100 4344 23112
rect 4295 23072 4344 23100
rect 4295 23069 4307 23072
rect 4249 23063 4307 23069
rect 4338 23060 4344 23072
rect 4396 23060 4402 23112
rect 9582 23060 9588 23112
rect 9640 23060 9646 23112
rect 13386 23072 15424 23100
rect 1765 23035 1823 23041
rect 1765 23001 1777 23035
rect 1811 23032 1823 23035
rect 2038 23032 2044 23044
rect 1811 23004 2044 23032
rect 1811 23001 1823 23004
rect 1765 22995 1823 23001
rect 2038 22992 2044 23004
rect 2096 22992 2102 23044
rect 6549 23035 6607 23041
rect 6549 23001 6561 23035
rect 6595 23001 6607 23035
rect 8478 23032 8484 23044
rect 7774 23004 8484 23032
rect 6549 22995 6607 23001
rect 4430 22924 4436 22976
rect 4488 22964 4494 22976
rect 4893 22967 4951 22973
rect 4893 22964 4905 22967
rect 4488 22936 4905 22964
rect 4488 22924 4494 22936
rect 4893 22933 4905 22936
rect 4939 22933 4951 22967
rect 6564 22964 6592 22995
rect 8478 22992 8484 23004
rect 8536 23032 8542 23044
rect 8846 23032 8852 23044
rect 8536 23004 8852 23032
rect 8536 22992 8542 23004
rect 8846 22992 8852 23004
rect 8904 22992 8910 23044
rect 10226 22992 10232 23044
rect 10284 22992 10290 23044
rect 12253 23035 12311 23041
rect 12253 23001 12265 23035
rect 12299 23032 12311 23035
rect 12342 23032 12348 23044
rect 12299 23004 12348 23032
rect 12299 23001 12311 23004
rect 12253 22995 12311 23001
rect 12342 22992 12348 23004
rect 12400 22992 12406 23044
rect 14645 23035 14703 23041
rect 14645 23032 14657 23035
rect 13556 23004 14657 23032
rect 7558 22964 7564 22976
rect 6564 22936 7564 22964
rect 4893 22927 4951 22933
rect 7558 22924 7564 22936
rect 7616 22924 7622 22976
rect 10244 22964 10272 22992
rect 11425 22967 11483 22973
rect 11425 22964 11437 22967
rect 10244 22936 11437 22964
rect 11425 22933 11437 22936
rect 11471 22964 11483 22967
rect 11514 22964 11520 22976
rect 11471 22936 11520 22964
rect 11471 22933 11483 22936
rect 11425 22927 11483 22933
rect 11514 22924 11520 22936
rect 11572 22924 11578 22976
rect 11974 22924 11980 22976
rect 12032 22964 12038 22976
rect 13556 22964 13584 23004
rect 14645 23001 14657 23004
rect 14691 23001 14703 23035
rect 14645 22995 14703 23001
rect 15396 23032 15424 23072
rect 20806 23060 20812 23112
rect 20864 23100 20870 23112
rect 21560 23100 21588 23267
rect 21634 23264 21640 23276
rect 21692 23264 21698 23316
rect 24578 23264 24584 23316
rect 24636 23304 24642 23316
rect 24636 23276 25176 23304
rect 24636 23264 24642 23276
rect 23474 23196 23480 23248
rect 23532 23236 23538 23248
rect 23532 23208 25084 23236
rect 23532 23196 23538 23208
rect 25056 23177 25084 23208
rect 25148 23177 25176 23276
rect 22005 23171 22063 23177
rect 22005 23137 22017 23171
rect 22051 23168 22063 23171
rect 25041 23171 25099 23177
rect 22051 23140 24992 23168
rect 22051 23137 22063 23140
rect 22005 23131 22063 23137
rect 20864 23072 21588 23100
rect 22833 23103 22891 23109
rect 20864 23060 20870 23072
rect 22833 23069 22845 23103
rect 22879 23069 22891 23103
rect 22833 23063 22891 23069
rect 16574 23032 16580 23044
rect 15396 23004 16580 23032
rect 12032 22936 13584 22964
rect 13725 22967 13783 22973
rect 12032 22924 12038 22936
rect 13725 22933 13737 22967
rect 13771 22964 13783 22967
rect 13814 22964 13820 22976
rect 13771 22936 13820 22964
rect 13771 22933 13783 22936
rect 13725 22927 13783 22933
rect 13814 22924 13820 22936
rect 13872 22964 13878 22976
rect 14550 22964 14556 22976
rect 13872 22936 14556 22964
rect 13872 22924 13878 22936
rect 14550 22924 14556 22936
rect 14608 22924 14614 22976
rect 15396 22973 15424 23004
rect 16574 22992 16580 23004
rect 16632 23032 16638 23044
rect 17862 23032 17868 23044
rect 16632 23004 17868 23032
rect 16632 22992 16638 23004
rect 17862 22992 17868 23004
rect 17920 22992 17926 23044
rect 19705 23035 19763 23041
rect 19705 23001 19717 23035
rect 19751 23001 19763 23035
rect 22848 23032 22876 23063
rect 23842 23060 23848 23112
rect 23900 23060 23906 23112
rect 24964 23109 24992 23140
rect 25041 23137 25053 23171
rect 25087 23137 25099 23171
rect 25041 23131 25099 23137
rect 25133 23171 25191 23177
rect 25133 23137 25145 23171
rect 25179 23137 25191 23171
rect 25133 23131 25191 23137
rect 24949 23103 25007 23109
rect 24949 23069 24961 23103
rect 24995 23069 25007 23103
rect 24949 23063 25007 23069
rect 24670 23032 24676 23044
rect 22848 23004 24676 23032
rect 19705 22995 19763 23001
rect 15381 22967 15439 22973
rect 15381 22933 15393 22967
rect 15427 22964 15439 22967
rect 15562 22964 15568 22976
rect 15427 22936 15568 22964
rect 15427 22933 15439 22936
rect 15381 22927 15439 22933
rect 15562 22924 15568 22936
rect 15620 22924 15626 22976
rect 19720 22964 19748 22995
rect 24670 22992 24676 23004
rect 24728 22992 24734 23044
rect 20714 22964 20720 22976
rect 19720 22936 20720 22964
rect 20714 22924 20720 22936
rect 20772 22924 20778 22976
rect 23566 22924 23572 22976
rect 23624 22964 23630 22976
rect 24581 22967 24639 22973
rect 24581 22964 24593 22967
rect 23624 22936 24593 22964
rect 23624 22924 23630 22936
rect 24581 22933 24593 22936
rect 24627 22933 24639 22967
rect 24581 22927 24639 22933
rect 1104 22874 25852 22896
rect 1104 22822 7950 22874
rect 8002 22822 8014 22874
rect 8066 22822 8078 22874
rect 8130 22822 8142 22874
rect 8194 22822 8206 22874
rect 8258 22822 17950 22874
rect 18002 22822 18014 22874
rect 18066 22822 18078 22874
rect 18130 22822 18142 22874
rect 18194 22822 18206 22874
rect 18258 22822 25852 22874
rect 1104 22800 25852 22822
rect 2038 22720 2044 22772
rect 2096 22760 2102 22772
rect 2682 22760 2688 22772
rect 2096 22732 2688 22760
rect 2096 22720 2102 22732
rect 2682 22720 2688 22732
rect 2740 22760 2746 22772
rect 4801 22763 4859 22769
rect 4801 22760 4813 22763
rect 2740 22732 4813 22760
rect 2740 22720 2746 22732
rect 4801 22729 4813 22732
rect 4847 22729 4859 22763
rect 4801 22723 4859 22729
rect 7742 22720 7748 22772
rect 7800 22760 7806 22772
rect 8110 22760 8116 22772
rect 7800 22732 8116 22760
rect 7800 22720 7806 22732
rect 8110 22720 8116 22732
rect 8168 22720 8174 22772
rect 9766 22720 9772 22772
rect 9824 22760 9830 22772
rect 10137 22763 10195 22769
rect 10137 22760 10149 22763
rect 9824 22732 10149 22760
rect 9824 22720 9830 22732
rect 10137 22729 10149 22732
rect 10183 22760 10195 22763
rect 10781 22763 10839 22769
rect 10183 22732 10456 22760
rect 10183 22729 10195 22732
rect 10137 22723 10195 22729
rect 10428 22704 10456 22732
rect 10781 22729 10793 22763
rect 10827 22760 10839 22763
rect 11790 22760 11796 22772
rect 10827 22732 11796 22760
rect 10827 22729 10839 22732
rect 10781 22723 10839 22729
rect 11790 22720 11796 22732
rect 11848 22720 11854 22772
rect 12526 22720 12532 22772
rect 12584 22760 12590 22772
rect 13817 22763 13875 22769
rect 13817 22760 13829 22763
rect 12584 22732 13829 22760
rect 12584 22720 12590 22732
rect 13817 22729 13829 22732
rect 13863 22729 13875 22763
rect 13817 22723 13875 22729
rect 13906 22720 13912 22772
rect 13964 22720 13970 22772
rect 15838 22720 15844 22772
rect 15896 22760 15902 22772
rect 17681 22763 17739 22769
rect 17681 22760 17693 22763
rect 15896 22732 17693 22760
rect 15896 22720 15902 22732
rect 3694 22652 3700 22704
rect 3752 22692 3758 22704
rect 3973 22695 4031 22701
rect 3973 22692 3985 22695
rect 3752 22664 3985 22692
rect 3752 22652 3758 22664
rect 3973 22661 3985 22664
rect 4019 22661 4031 22695
rect 3973 22655 4031 22661
rect 8205 22695 8263 22701
rect 8205 22661 8217 22695
rect 8251 22692 8263 22695
rect 9401 22695 9459 22701
rect 9401 22692 9413 22695
rect 8251 22664 9413 22692
rect 8251 22661 8263 22664
rect 8205 22655 8263 22661
rect 9401 22661 9413 22664
rect 9447 22692 9459 22695
rect 10226 22692 10232 22704
rect 9447 22664 10232 22692
rect 9447 22661 9459 22664
rect 9401 22655 9459 22661
rect 3988 22624 4016 22655
rect 10226 22652 10232 22664
rect 10284 22652 10290 22704
rect 10410 22652 10416 22704
rect 10468 22692 10474 22704
rect 10873 22695 10931 22701
rect 10873 22692 10885 22695
rect 10468 22664 10885 22692
rect 10468 22652 10474 22664
rect 10873 22661 10885 22664
rect 10919 22661 10931 22695
rect 10873 22655 10931 22661
rect 11698 22652 11704 22704
rect 11756 22652 11762 22704
rect 12250 22652 12256 22704
rect 12308 22692 12314 22704
rect 12308 22664 16344 22692
rect 12308 22652 12314 22664
rect 4341 22627 4399 22633
rect 4341 22624 4353 22627
rect 3988 22596 4353 22624
rect 4341 22593 4353 22596
rect 4387 22624 4399 22627
rect 6362 22624 6368 22636
rect 4387 22596 6368 22624
rect 4387 22593 4399 22596
rect 4341 22587 4399 22593
rect 6362 22584 6368 22596
rect 6420 22584 6426 22636
rect 7098 22584 7104 22636
rect 7156 22584 7162 22636
rect 7834 22584 7840 22636
rect 7892 22624 7898 22636
rect 8941 22627 8999 22633
rect 8941 22624 8953 22627
rect 7892 22596 8953 22624
rect 7892 22584 7898 22596
rect 8941 22593 8953 22596
rect 8987 22593 8999 22627
rect 8941 22587 8999 22593
rect 10686 22584 10692 22636
rect 10744 22624 10750 22636
rect 12066 22624 12072 22636
rect 10744 22596 12072 22624
rect 10744 22584 10750 22596
rect 12066 22584 12072 22596
rect 12124 22584 12130 22636
rect 12618 22584 12624 22636
rect 12676 22624 12682 22636
rect 12989 22627 13047 22633
rect 12989 22624 13001 22627
rect 12676 22596 13001 22624
rect 12676 22584 12682 22596
rect 12989 22593 13001 22596
rect 13035 22593 13047 22627
rect 12989 22587 13047 22593
rect 14642 22584 14648 22636
rect 14700 22584 14706 22636
rect 16316 22633 16344 22664
rect 16301 22627 16359 22633
rect 16301 22593 16313 22627
rect 16347 22593 16359 22627
rect 17052 22624 17080 22732
rect 17681 22729 17693 22732
rect 17727 22729 17739 22763
rect 17681 22723 17739 22729
rect 24118 22720 24124 22772
rect 24176 22760 24182 22772
rect 24581 22763 24639 22769
rect 24581 22760 24593 22763
rect 24176 22732 24593 22760
rect 24176 22720 24182 22732
rect 24581 22729 24593 22732
rect 24627 22729 24639 22763
rect 24581 22723 24639 22729
rect 25130 22720 25136 22772
rect 25188 22720 25194 22772
rect 17126 22652 17132 22704
rect 17184 22692 17190 22704
rect 18322 22692 18328 22704
rect 17184 22664 18328 22692
rect 17184 22652 17190 22664
rect 18322 22652 18328 22664
rect 18380 22692 18386 22704
rect 18785 22695 18843 22701
rect 18785 22692 18797 22695
rect 18380 22664 18797 22692
rect 18380 22652 18386 22664
rect 18785 22661 18797 22664
rect 18831 22661 18843 22695
rect 25148 22692 25176 22720
rect 23598 22664 25176 22692
rect 18785 22655 18843 22661
rect 18049 22627 18107 22633
rect 18049 22624 18061 22627
rect 17052 22596 18061 22624
rect 16301 22587 16359 22593
rect 18049 22593 18061 22596
rect 18095 22593 18107 22627
rect 18049 22587 18107 22593
rect 10962 22516 10968 22568
rect 11020 22516 11026 22568
rect 14090 22516 14096 22568
rect 14148 22516 14154 22568
rect 17494 22516 17500 22568
rect 17552 22556 17558 22568
rect 18064 22556 18092 22587
rect 18874 22584 18880 22636
rect 18932 22624 18938 22636
rect 19429 22627 19487 22633
rect 19429 22624 19441 22627
rect 18932 22596 19441 22624
rect 18932 22584 18938 22596
rect 19429 22593 19441 22596
rect 19475 22593 19487 22627
rect 20530 22624 20536 22636
rect 19429 22587 19487 22593
rect 20272 22596 20536 22624
rect 20272 22556 20300 22596
rect 20530 22584 20536 22596
rect 20588 22624 20594 22636
rect 20588 22596 20633 22624
rect 20588 22584 20594 22596
rect 24762 22584 24768 22636
rect 24820 22584 24826 22636
rect 17552 22528 18000 22556
rect 18064 22528 20300 22556
rect 17552 22516 17558 22528
rect 9214 22448 9220 22500
rect 9272 22488 9278 22500
rect 11974 22488 11980 22500
rect 9272 22460 11980 22488
rect 9272 22448 9278 22460
rect 11974 22448 11980 22460
rect 12032 22448 12038 22500
rect 13449 22491 13507 22497
rect 13449 22457 13461 22491
rect 13495 22488 13507 22491
rect 17586 22488 17592 22500
rect 13495 22460 17592 22488
rect 13495 22457 13507 22460
rect 13449 22451 13507 22457
rect 17586 22448 17592 22460
rect 17644 22448 17650 22500
rect 17972 22488 18000 22528
rect 21082 22516 21088 22568
rect 21140 22556 21146 22568
rect 21269 22559 21327 22565
rect 21269 22556 21281 22559
rect 21140 22528 21281 22556
rect 21140 22516 21146 22528
rect 21269 22525 21281 22528
rect 21315 22556 21327 22559
rect 22094 22556 22100 22568
rect 21315 22528 22100 22556
rect 21315 22525 21327 22528
rect 21269 22519 21327 22525
rect 22094 22516 22100 22528
rect 22152 22516 22158 22568
rect 22373 22559 22431 22565
rect 22373 22525 22385 22559
rect 22419 22556 22431 22559
rect 24026 22556 24032 22568
rect 22419 22528 24032 22556
rect 22419 22525 22431 22528
rect 22373 22519 22431 22525
rect 24026 22516 24032 22528
rect 24084 22516 24090 22568
rect 24121 22559 24179 22565
rect 24121 22525 24133 22559
rect 24167 22525 24179 22559
rect 24121 22519 24179 22525
rect 17972 22460 22094 22488
rect 4617 22423 4675 22429
rect 4617 22389 4629 22423
rect 4663 22420 4675 22423
rect 5810 22420 5816 22432
rect 4663 22392 5816 22420
rect 4663 22389 4675 22392
rect 4617 22383 4675 22389
rect 5810 22380 5816 22392
rect 5868 22380 5874 22432
rect 7742 22380 7748 22432
rect 7800 22380 7806 22432
rect 10410 22380 10416 22432
rect 10468 22380 10474 22432
rect 12618 22380 12624 22432
rect 12676 22420 12682 22432
rect 12805 22423 12863 22429
rect 12805 22420 12817 22423
rect 12676 22392 12817 22420
rect 12676 22380 12682 22392
rect 12805 22389 12817 22392
rect 12851 22389 12863 22423
rect 12805 22383 12863 22389
rect 14550 22380 14556 22432
rect 14608 22420 14614 22432
rect 15289 22423 15347 22429
rect 15289 22420 15301 22423
rect 14608 22392 15301 22420
rect 14608 22380 14614 22392
rect 15289 22389 15301 22392
rect 15335 22389 15347 22423
rect 15289 22383 15347 22389
rect 16114 22380 16120 22432
rect 16172 22380 16178 22432
rect 20070 22380 20076 22432
rect 20128 22380 20134 22432
rect 22066 22420 22094 22460
rect 24136 22420 24164 22519
rect 22066 22392 24164 22420
rect 1104 22330 25852 22352
rect 1104 22278 2950 22330
rect 3002 22278 3014 22330
rect 3066 22278 3078 22330
rect 3130 22278 3142 22330
rect 3194 22278 3206 22330
rect 3258 22278 12950 22330
rect 13002 22278 13014 22330
rect 13066 22278 13078 22330
rect 13130 22278 13142 22330
rect 13194 22278 13206 22330
rect 13258 22278 22950 22330
rect 23002 22278 23014 22330
rect 23066 22278 23078 22330
rect 23130 22278 23142 22330
rect 23194 22278 23206 22330
rect 23258 22278 25852 22330
rect 1104 22256 25852 22278
rect 4420 22219 4478 22225
rect 4420 22185 4432 22219
rect 4466 22216 4478 22219
rect 5626 22216 5632 22228
rect 4466 22188 5632 22216
rect 4466 22185 4478 22188
rect 4420 22179 4478 22185
rect 5626 22176 5632 22188
rect 5684 22176 5690 22228
rect 14642 22216 14648 22228
rect 12406 22188 14648 22216
rect 8846 22148 8852 22160
rect 6886 22120 8852 22148
rect 3970 22040 3976 22092
rect 4028 22080 4034 22092
rect 4154 22080 4160 22092
rect 4028 22052 4160 22080
rect 4028 22040 4034 22052
rect 4154 22040 4160 22052
rect 4212 22040 4218 22092
rect 5902 22040 5908 22092
rect 5960 22040 5966 22092
rect 6886 22080 6914 22120
rect 8846 22108 8852 22120
rect 8904 22108 8910 22160
rect 12406 22148 12434 22188
rect 14642 22176 14648 22188
rect 14700 22216 14706 22228
rect 14700 22188 15148 22216
rect 14700 22176 14706 22188
rect 13814 22148 13820 22160
rect 11716 22120 12434 22148
rect 13096 22120 13820 22148
rect 11716 22092 11744 22120
rect 6104 22052 6914 22080
rect 1946 21972 1952 22024
rect 2004 22012 2010 22024
rect 2225 22015 2283 22021
rect 2225 22012 2237 22015
rect 2004 21984 2237 22012
rect 2004 21972 2010 21984
rect 2225 21981 2237 21984
rect 2271 21981 2283 22015
rect 2225 21975 2283 21981
rect 3326 21972 3332 22024
rect 3384 21972 3390 22024
rect 6104 21944 6132 22052
rect 8110 22040 8116 22092
rect 8168 22040 8174 22092
rect 9398 22040 9404 22092
rect 9456 22080 9462 22092
rect 9677 22083 9735 22089
rect 9677 22080 9689 22083
rect 9456 22052 9689 22080
rect 9456 22040 9462 22052
rect 9677 22049 9689 22052
rect 9723 22049 9735 22083
rect 9677 22043 9735 22049
rect 10686 22040 10692 22092
rect 10744 22080 10750 22092
rect 10781 22083 10839 22089
rect 10781 22080 10793 22083
rect 10744 22052 10793 22080
rect 10744 22040 10750 22052
rect 10781 22049 10793 22052
rect 10827 22080 10839 22083
rect 11609 22083 11667 22089
rect 11609 22080 11621 22083
rect 10827 22052 11621 22080
rect 10827 22049 10839 22052
rect 10781 22043 10839 22049
rect 11609 22049 11621 22052
rect 11655 22049 11667 22083
rect 11609 22043 11667 22049
rect 11698 22040 11704 22092
rect 11756 22040 11762 22092
rect 12526 22040 12532 22092
rect 12584 22080 12590 22092
rect 13096 22089 13124 22120
rect 13814 22108 13820 22120
rect 13872 22108 13878 22160
rect 14737 22151 14795 22157
rect 14737 22117 14749 22151
rect 14783 22117 14795 22151
rect 15120 22148 15148 22188
rect 20806 22176 20812 22228
rect 20864 22176 20870 22228
rect 22094 22176 22100 22228
rect 22152 22216 22158 22228
rect 23198 22216 23204 22228
rect 22152 22188 23204 22216
rect 22152 22176 22158 22188
rect 23198 22176 23204 22188
rect 23256 22176 23262 22228
rect 25130 22176 25136 22228
rect 25188 22176 25194 22228
rect 19978 22148 19984 22160
rect 15120 22120 15332 22148
rect 14737 22111 14795 22117
rect 13081 22083 13139 22089
rect 12584 22052 13032 22080
rect 12584 22040 12590 22052
rect 7650 21972 7656 22024
rect 7708 22012 7714 22024
rect 7929 22015 7987 22021
rect 7929 22012 7941 22015
rect 7708 21984 7941 22012
rect 7708 21972 7714 21984
rect 7929 21981 7941 21984
rect 7975 21981 7987 22015
rect 7929 21975 7987 21981
rect 8386 21972 8392 22024
rect 8444 22012 8450 22024
rect 8754 22012 8760 22024
rect 8444 21984 8760 22012
rect 8444 21972 8450 21984
rect 8754 21972 8760 21984
rect 8812 22012 8818 22024
rect 9493 22015 9551 22021
rect 9493 22012 9505 22015
rect 8812 21984 9505 22012
rect 8812 21972 8818 21984
rect 9493 21981 9505 21984
rect 9539 21981 9551 22015
rect 9493 21975 9551 21981
rect 12250 21972 12256 22024
rect 12308 22012 12314 22024
rect 12897 22015 12955 22021
rect 12897 22012 12909 22015
rect 12308 21984 12909 22012
rect 12308 21972 12314 21984
rect 12897 21981 12909 21984
rect 12943 21981 12955 22015
rect 13004 22012 13032 22052
rect 13081 22049 13093 22083
rect 13127 22080 13139 22083
rect 13541 22083 13599 22089
rect 13127 22052 13161 22080
rect 13127 22049 13139 22052
rect 13081 22043 13139 22049
rect 13541 22049 13553 22083
rect 13587 22080 13599 22083
rect 13906 22080 13912 22092
rect 13587 22052 13912 22080
rect 13587 22049 13599 22052
rect 13541 22043 13599 22049
rect 13906 22040 13912 22052
rect 13964 22040 13970 22092
rect 14182 22040 14188 22092
rect 14240 22040 14246 22092
rect 14752 22012 14780 22111
rect 15102 22040 15108 22092
rect 15160 22080 15166 22092
rect 15304 22089 15332 22120
rect 18064 22120 19984 22148
rect 15197 22083 15255 22089
rect 15197 22080 15209 22083
rect 15160 22052 15209 22080
rect 15160 22040 15166 22052
rect 15197 22049 15209 22052
rect 15243 22049 15255 22083
rect 15197 22043 15255 22049
rect 15289 22083 15347 22089
rect 15289 22049 15301 22083
rect 15335 22049 15347 22083
rect 15289 22043 15347 22049
rect 16482 22040 16488 22092
rect 16540 22040 16546 22092
rect 17770 22040 17776 22092
rect 17828 22080 17834 22092
rect 18064 22089 18092 22120
rect 19978 22108 19984 22120
rect 20036 22108 20042 22160
rect 17865 22083 17923 22089
rect 17865 22080 17877 22083
rect 17828 22052 17877 22080
rect 17828 22040 17834 22052
rect 17865 22049 17877 22052
rect 17911 22049 17923 22083
rect 17865 22043 17923 22049
rect 18049 22083 18107 22089
rect 18049 22049 18061 22083
rect 18095 22080 18107 22083
rect 18095 22052 18129 22080
rect 18095 22049 18107 22052
rect 18049 22043 18107 22049
rect 18598 22040 18604 22092
rect 18656 22040 18662 22092
rect 19334 22040 19340 22092
rect 19392 22080 19398 22092
rect 20073 22083 20131 22089
rect 20073 22080 20085 22083
rect 19392 22052 20085 22080
rect 19392 22040 19398 22052
rect 20073 22049 20085 22052
rect 20119 22049 20131 22083
rect 20073 22043 20131 22049
rect 22738 22040 22744 22092
rect 22796 22080 22802 22092
rect 22833 22083 22891 22089
rect 22833 22080 22845 22083
rect 22796 22052 22845 22080
rect 22796 22040 22802 22052
rect 22833 22049 22845 22052
rect 22879 22049 22891 22083
rect 22833 22043 22891 22049
rect 24026 22040 24032 22092
rect 24084 22040 24090 22092
rect 13004 21984 14780 22012
rect 12897 21975 12955 21981
rect 15010 21972 15016 22024
rect 15068 22012 15074 22024
rect 15068 21984 16528 22012
rect 15068 21972 15074 21984
rect 5658 21916 6132 21944
rect 6104 21888 6132 21916
rect 8021 21947 8079 21953
rect 8021 21913 8033 21947
rect 8067 21944 8079 21947
rect 16301 21947 16359 21953
rect 16301 21944 16313 21947
rect 8067 21916 9168 21944
rect 8067 21913 8079 21916
rect 8021 21907 8079 21913
rect 1762 21836 1768 21888
rect 1820 21876 1826 21888
rect 2041 21879 2099 21885
rect 2041 21876 2053 21879
rect 1820 21848 2053 21876
rect 1820 21836 1826 21848
rect 2041 21845 2053 21848
rect 2087 21845 2099 21879
rect 2041 21839 2099 21845
rect 2130 21836 2136 21888
rect 2188 21876 2194 21888
rect 3145 21879 3203 21885
rect 3145 21876 3157 21879
rect 2188 21848 3157 21876
rect 2188 21836 2194 21848
rect 3145 21845 3157 21848
rect 3191 21845 3203 21879
rect 3145 21839 3203 21845
rect 6086 21836 6092 21888
rect 6144 21876 6150 21888
rect 6181 21879 6239 21885
rect 6181 21876 6193 21879
rect 6144 21848 6193 21876
rect 6144 21836 6150 21848
rect 6181 21845 6193 21848
rect 6227 21845 6239 21879
rect 6181 21839 6239 21845
rect 6730 21836 6736 21888
rect 6788 21876 6794 21888
rect 7561 21879 7619 21885
rect 7561 21876 7573 21879
rect 6788 21848 7573 21876
rect 6788 21836 6794 21848
rect 7561 21845 7573 21848
rect 7607 21845 7619 21879
rect 7561 21839 7619 21845
rect 8386 21836 8392 21888
rect 8444 21876 8450 21888
rect 9140 21885 9168 21916
rect 12452 21916 16313 21944
rect 8665 21879 8723 21885
rect 8665 21876 8677 21879
rect 8444 21848 8677 21876
rect 8444 21836 8450 21848
rect 8665 21845 8677 21848
rect 8711 21845 8723 21879
rect 8665 21839 8723 21845
rect 9125 21879 9183 21885
rect 9125 21845 9137 21879
rect 9171 21845 9183 21879
rect 9125 21839 9183 21845
rect 9582 21836 9588 21888
rect 9640 21836 9646 21888
rect 11146 21836 11152 21888
rect 11204 21836 11210 21888
rect 11517 21879 11575 21885
rect 11517 21845 11529 21879
rect 11563 21876 11575 21879
rect 11606 21876 11612 21888
rect 11563 21848 11612 21876
rect 11563 21845 11575 21848
rect 11517 21839 11575 21845
rect 11606 21836 11612 21848
rect 11664 21836 11670 21888
rect 12452 21885 12480 21916
rect 16301 21913 16313 21916
rect 16347 21913 16359 21947
rect 16500 21944 16528 21984
rect 16574 21972 16580 22024
rect 16632 22012 16638 22024
rect 16758 22012 16764 22024
rect 16632 21984 16764 22012
rect 16632 21972 16638 21984
rect 16758 21972 16764 21984
rect 16816 21972 16822 22024
rect 18616 22012 18644 22040
rect 19429 22015 19487 22021
rect 19429 22012 19441 22015
rect 17880 21984 19441 22012
rect 17880 21944 17908 21984
rect 19429 21981 19441 21984
rect 19475 22012 19487 22015
rect 19475 21984 20484 22012
rect 19475 21981 19487 21984
rect 19429 21975 19487 21981
rect 16500 21916 17908 21944
rect 16301 21907 16359 21913
rect 12437 21879 12495 21885
rect 12437 21845 12449 21879
rect 12483 21845 12495 21879
rect 12437 21839 12495 21845
rect 12802 21836 12808 21888
rect 12860 21836 12866 21888
rect 14090 21836 14096 21888
rect 14148 21876 14154 21888
rect 14369 21879 14427 21885
rect 14369 21876 14381 21879
rect 14148 21848 14381 21876
rect 14148 21836 14154 21848
rect 14369 21845 14381 21848
rect 14415 21876 14427 21879
rect 15010 21876 15016 21888
rect 14415 21848 15016 21876
rect 14415 21845 14427 21848
rect 14369 21839 14427 21845
rect 15010 21836 15016 21848
rect 15068 21836 15074 21888
rect 15105 21879 15163 21885
rect 15105 21845 15117 21879
rect 15151 21876 15163 21879
rect 15654 21876 15660 21888
rect 15151 21848 15660 21876
rect 15151 21845 15163 21848
rect 15105 21839 15163 21845
rect 15654 21836 15660 21848
rect 15712 21836 15718 21888
rect 15930 21836 15936 21888
rect 15988 21836 15994 21888
rect 16393 21879 16451 21885
rect 16393 21845 16405 21879
rect 16439 21876 16451 21879
rect 16574 21876 16580 21888
rect 16439 21848 16580 21876
rect 16439 21845 16451 21848
rect 16393 21839 16451 21845
rect 16574 21836 16580 21848
rect 16632 21836 16638 21888
rect 16758 21836 16764 21888
rect 16816 21876 16822 21888
rect 17405 21879 17463 21885
rect 17405 21876 17417 21879
rect 16816 21848 17417 21876
rect 16816 21836 16822 21848
rect 17405 21845 17417 21848
rect 17451 21845 17463 21879
rect 17405 21839 17463 21845
rect 17494 21836 17500 21888
rect 17552 21876 17558 21888
rect 17773 21879 17831 21885
rect 17773 21876 17785 21879
rect 17552 21848 17785 21876
rect 17552 21836 17558 21848
rect 17773 21845 17785 21848
rect 17819 21845 17831 21879
rect 17773 21839 17831 21845
rect 17862 21836 17868 21888
rect 17920 21876 17926 21888
rect 20456 21885 20484 21984
rect 20806 21972 20812 22024
rect 20864 22012 20870 22024
rect 21082 22012 21088 22024
rect 20864 21984 21088 22012
rect 20864 21972 20870 21984
rect 21082 21972 21088 21984
rect 21140 21972 21146 22024
rect 23382 21972 23388 22024
rect 23440 21972 23446 22024
rect 20530 21904 20536 21956
rect 20588 21904 20594 21956
rect 21358 21904 21364 21956
rect 21416 21904 21422 21956
rect 21634 21904 21640 21956
rect 21692 21944 21698 21956
rect 24673 21947 24731 21953
rect 24673 21944 24685 21947
rect 21692 21916 21850 21944
rect 22664 21916 24685 21944
rect 21692 21904 21698 21916
rect 18601 21879 18659 21885
rect 18601 21876 18613 21879
rect 17920 21848 18613 21876
rect 17920 21836 17926 21848
rect 18601 21845 18613 21848
rect 18647 21845 18659 21879
rect 18601 21839 18659 21845
rect 20441 21879 20499 21885
rect 20441 21845 20453 21879
rect 20487 21876 20499 21879
rect 20898 21876 20904 21888
rect 20487 21848 20904 21876
rect 20487 21845 20499 21848
rect 20441 21839 20499 21845
rect 20898 21836 20904 21848
rect 20956 21836 20962 21888
rect 21266 21836 21272 21888
rect 21324 21876 21330 21888
rect 22664 21876 22692 21916
rect 24673 21913 24685 21916
rect 24719 21913 24731 21947
rect 24673 21907 24731 21913
rect 21324 21848 22692 21876
rect 21324 21836 21330 21848
rect 24118 21836 24124 21888
rect 24176 21876 24182 21888
rect 24765 21879 24823 21885
rect 24765 21876 24777 21879
rect 24176 21848 24777 21876
rect 24176 21836 24182 21848
rect 24765 21845 24777 21848
rect 24811 21845 24823 21879
rect 24765 21839 24823 21845
rect 1104 21786 25852 21808
rect 1104 21734 7950 21786
rect 8002 21734 8014 21786
rect 8066 21734 8078 21786
rect 8130 21734 8142 21786
rect 8194 21734 8206 21786
rect 8258 21734 17950 21786
rect 18002 21734 18014 21786
rect 18066 21734 18078 21786
rect 18130 21734 18142 21786
rect 18194 21734 18206 21786
rect 18258 21734 25852 21786
rect 1104 21712 25852 21734
rect 3326 21632 3332 21684
rect 3384 21672 3390 21684
rect 5169 21675 5227 21681
rect 5169 21672 5181 21675
rect 3384 21644 5181 21672
rect 3384 21632 3390 21644
rect 5169 21641 5181 21644
rect 5215 21641 5227 21675
rect 5169 21635 5227 21641
rect 5537 21675 5595 21681
rect 5537 21641 5549 21675
rect 5583 21672 5595 21675
rect 6641 21675 6699 21681
rect 6641 21672 6653 21675
rect 5583 21644 6653 21672
rect 5583 21641 5595 21644
rect 5537 21635 5595 21641
rect 6641 21641 6653 21644
rect 6687 21641 6699 21675
rect 6641 21635 6699 21641
rect 7009 21675 7067 21681
rect 7009 21641 7021 21675
rect 7055 21672 7067 21675
rect 7190 21672 7196 21684
rect 7055 21644 7196 21672
rect 7055 21641 7067 21644
rect 7009 21635 7067 21641
rect 7190 21632 7196 21644
rect 7248 21632 7254 21684
rect 10686 21672 10692 21684
rect 7668 21644 10692 21672
rect 2130 21604 2136 21616
rect 1872 21576 2136 21604
rect 1872 21545 1900 21576
rect 2130 21564 2136 21576
rect 2188 21564 2194 21616
rect 6270 21564 6276 21616
rect 6328 21604 6334 21616
rect 7668 21604 7696 21644
rect 10686 21632 10692 21644
rect 10744 21632 10750 21684
rect 10778 21632 10784 21684
rect 10836 21632 10842 21684
rect 11698 21672 11704 21684
rect 10888 21644 11704 21672
rect 6328 21576 7696 21604
rect 6328 21564 6334 21576
rect 7742 21564 7748 21616
rect 7800 21604 7806 21616
rect 8113 21607 8171 21613
rect 8113 21604 8125 21607
rect 7800 21576 8125 21604
rect 7800 21564 7806 21576
rect 8113 21573 8125 21576
rect 8159 21573 8171 21607
rect 8113 21567 8171 21573
rect 8846 21564 8852 21616
rect 8904 21564 8910 21616
rect 9861 21607 9919 21613
rect 9861 21573 9873 21607
rect 9907 21604 9919 21607
rect 10888 21604 10916 21644
rect 11698 21632 11704 21644
rect 11756 21632 11762 21684
rect 12802 21632 12808 21684
rect 12860 21672 12866 21684
rect 12897 21675 12955 21681
rect 12897 21672 12909 21675
rect 12860 21644 12909 21672
rect 12860 21632 12866 21644
rect 12897 21641 12909 21644
rect 12943 21641 12955 21675
rect 12897 21635 12955 21641
rect 14277 21675 14335 21681
rect 14277 21641 14289 21675
rect 14323 21641 14335 21675
rect 14277 21635 14335 21641
rect 14645 21675 14703 21681
rect 14645 21641 14657 21675
rect 14691 21672 14703 21675
rect 17129 21675 17187 21681
rect 14691 21644 15424 21672
rect 14691 21641 14703 21644
rect 14645 21635 14703 21641
rect 9907 21576 10916 21604
rect 9907 21573 9919 21576
rect 9861 21567 9919 21573
rect 10962 21564 10968 21616
rect 11020 21604 11026 21616
rect 11020 21576 12480 21604
rect 11020 21564 11026 21576
rect 1857 21539 1915 21545
rect 1857 21505 1869 21539
rect 1903 21505 1915 21539
rect 1857 21499 1915 21505
rect 5629 21539 5687 21545
rect 5629 21505 5641 21539
rect 5675 21536 5687 21539
rect 6914 21536 6920 21548
rect 5675 21508 6920 21536
rect 5675 21505 5687 21508
rect 5629 21499 5687 21505
rect 6914 21496 6920 21508
rect 6972 21496 6978 21548
rect 7834 21496 7840 21548
rect 7892 21496 7898 21548
rect 10873 21539 10931 21545
rect 10873 21505 10885 21539
rect 10919 21536 10931 21539
rect 12342 21536 12348 21548
rect 10919 21508 12348 21536
rect 10919 21505 10931 21508
rect 10873 21499 10931 21505
rect 12342 21496 12348 21508
rect 12400 21496 12406 21548
rect 12452 21536 12480 21576
rect 12710 21564 12716 21616
rect 12768 21604 12774 21616
rect 14292 21604 14320 21635
rect 15396 21613 15424 21644
rect 17129 21641 17141 21675
rect 17175 21672 17187 21675
rect 17494 21672 17500 21684
rect 17175 21644 17500 21672
rect 17175 21641 17187 21644
rect 17129 21635 17187 21641
rect 17494 21632 17500 21644
rect 17552 21632 17558 21684
rect 17586 21632 17592 21684
rect 17644 21632 17650 21684
rect 19978 21632 19984 21684
rect 20036 21672 20042 21684
rect 20073 21675 20131 21681
rect 20073 21672 20085 21675
rect 20036 21644 20085 21672
rect 20036 21632 20042 21644
rect 20073 21641 20085 21644
rect 20119 21641 20131 21675
rect 20073 21635 20131 21641
rect 12768 21576 14320 21604
rect 15381 21607 15439 21613
rect 12768 21564 12774 21576
rect 15381 21573 15393 21607
rect 15427 21604 15439 21607
rect 17862 21604 17868 21616
rect 15427 21576 17868 21604
rect 15427 21573 15439 21576
rect 15381 21567 15439 21573
rect 17862 21564 17868 21576
rect 17920 21564 17926 21616
rect 19150 21564 19156 21616
rect 19208 21564 19214 21616
rect 14090 21536 14096 21548
rect 12452 21508 14096 21536
rect 14090 21496 14096 21508
rect 14148 21536 14154 21548
rect 16117 21539 16175 21545
rect 14148 21508 14872 21536
rect 14148 21496 14154 21508
rect 2041 21471 2099 21477
rect 2041 21437 2053 21471
rect 2087 21468 2099 21471
rect 2314 21468 2320 21480
rect 2087 21440 2320 21468
rect 2087 21437 2099 21440
rect 2041 21431 2099 21437
rect 2314 21428 2320 21440
rect 2372 21428 2378 21480
rect 2866 21428 2872 21480
rect 2924 21428 2930 21480
rect 5813 21471 5871 21477
rect 5813 21437 5825 21471
rect 5859 21468 5871 21471
rect 5902 21468 5908 21480
rect 5859 21440 5908 21468
rect 5859 21437 5871 21440
rect 5813 21431 5871 21437
rect 5902 21428 5908 21440
rect 5960 21428 5966 21480
rect 7098 21428 7104 21480
rect 7156 21428 7162 21480
rect 7193 21471 7251 21477
rect 7193 21437 7205 21471
rect 7239 21437 7251 21471
rect 7193 21431 7251 21437
rect 7006 21360 7012 21412
rect 7064 21400 7070 21412
rect 7208 21400 7236 21431
rect 9950 21428 9956 21480
rect 10008 21468 10014 21480
rect 10965 21471 11023 21477
rect 10965 21468 10977 21471
rect 10008 21440 10977 21468
rect 10008 21428 10014 21440
rect 10965 21437 10977 21440
rect 11011 21437 11023 21471
rect 10965 21431 11023 21437
rect 11606 21428 11612 21480
rect 11664 21468 11670 21480
rect 12069 21471 12127 21477
rect 12069 21468 12081 21471
rect 11664 21440 12081 21468
rect 11664 21428 11670 21440
rect 12069 21437 12081 21440
rect 12115 21468 12127 21471
rect 13630 21468 13636 21480
rect 12115 21440 13636 21468
rect 12115 21437 12127 21440
rect 12069 21431 12127 21437
rect 13630 21428 13636 21440
rect 13688 21428 13694 21480
rect 13906 21428 13912 21480
rect 13964 21468 13970 21480
rect 14274 21468 14280 21480
rect 13964 21440 14280 21468
rect 13964 21428 13970 21440
rect 14274 21428 14280 21440
rect 14332 21468 14338 21480
rect 14844 21477 14872 21508
rect 16117 21505 16129 21539
rect 16163 21536 16175 21539
rect 17497 21539 17555 21545
rect 17497 21536 17509 21539
rect 16163 21508 17509 21536
rect 16163 21505 16175 21508
rect 16117 21499 16175 21505
rect 17497 21505 17509 21508
rect 17543 21505 17555 21539
rect 20088 21536 20116 21635
rect 20714 21632 20720 21684
rect 20772 21672 20778 21684
rect 21177 21675 21235 21681
rect 21177 21672 21189 21675
rect 20772 21644 21189 21672
rect 20772 21632 20778 21644
rect 21177 21641 21189 21644
rect 21223 21641 21235 21675
rect 21177 21635 21235 21641
rect 22462 21632 22468 21684
rect 22520 21632 22526 21684
rect 23382 21672 23388 21684
rect 23032 21644 23388 21672
rect 20533 21539 20591 21545
rect 20533 21536 20545 21539
rect 20088 21508 20545 21536
rect 17497 21499 17555 21505
rect 20533 21505 20545 21508
rect 20579 21505 20591 21539
rect 20533 21499 20591 21505
rect 22373 21539 22431 21545
rect 22373 21505 22385 21539
rect 22419 21536 22431 21539
rect 22419 21508 22600 21536
rect 22419 21505 22431 21508
rect 22373 21499 22431 21505
rect 14737 21471 14795 21477
rect 14737 21468 14749 21471
rect 14332 21440 14749 21468
rect 14332 21428 14338 21440
rect 14737 21437 14749 21440
rect 14783 21437 14795 21471
rect 14737 21431 14795 21437
rect 14829 21471 14887 21477
rect 14829 21437 14841 21471
rect 14875 21437 14887 21471
rect 14829 21431 14887 21437
rect 17773 21471 17831 21477
rect 17773 21437 17785 21471
rect 17819 21468 17831 21471
rect 18046 21468 18052 21480
rect 17819 21440 18052 21468
rect 17819 21437 17831 21440
rect 17773 21431 17831 21437
rect 18046 21428 18052 21440
rect 18104 21428 18110 21480
rect 18322 21428 18328 21480
rect 18380 21428 18386 21480
rect 18601 21471 18659 21477
rect 18601 21437 18613 21471
rect 18647 21468 18659 21471
rect 20070 21468 20076 21480
rect 18647 21440 20076 21468
rect 18647 21437 18659 21440
rect 18601 21431 18659 21437
rect 20070 21428 20076 21440
rect 20128 21428 20134 21480
rect 7064 21372 7236 21400
rect 7064 21360 7070 21372
rect 9490 21360 9496 21412
rect 9548 21400 9554 21412
rect 12250 21400 12256 21412
rect 9548 21372 12256 21400
rect 9548 21360 9554 21372
rect 12250 21360 12256 21372
rect 12308 21360 12314 21412
rect 13814 21360 13820 21412
rect 13872 21400 13878 21412
rect 18340 21400 18368 21428
rect 13872 21372 18368 21400
rect 13872 21360 13878 21372
rect 8478 21292 8484 21344
rect 8536 21332 8542 21344
rect 10413 21335 10471 21341
rect 10413 21332 10425 21335
rect 8536 21304 10425 21332
rect 8536 21292 8542 21304
rect 10413 21301 10425 21304
rect 10459 21301 10471 21335
rect 10413 21295 10471 21301
rect 13906 21292 13912 21344
rect 13964 21292 13970 21344
rect 14182 21292 14188 21344
rect 14240 21332 14246 21344
rect 15102 21332 15108 21344
rect 14240 21304 15108 21332
rect 14240 21292 14246 21304
rect 15102 21292 15108 21304
rect 15160 21292 15166 21344
rect 15654 21292 15660 21344
rect 15712 21332 15718 21344
rect 16574 21332 16580 21344
rect 15712 21304 16580 21332
rect 15712 21292 15718 21304
rect 16574 21292 16580 21304
rect 16632 21292 16638 21344
rect 16666 21292 16672 21344
rect 16724 21332 16730 21344
rect 16853 21335 16911 21341
rect 16853 21332 16865 21335
rect 16724 21304 16865 21332
rect 16724 21292 16730 21304
rect 16853 21301 16865 21304
rect 16899 21332 16911 21335
rect 17770 21332 17776 21344
rect 16899 21304 17776 21332
rect 16899 21301 16911 21304
rect 16853 21295 16911 21301
rect 17770 21292 17776 21304
rect 17828 21292 17834 21344
rect 17862 21292 17868 21344
rect 17920 21332 17926 21344
rect 19886 21332 19892 21344
rect 17920 21304 19892 21332
rect 17920 21292 17926 21304
rect 19886 21292 19892 21304
rect 19944 21292 19950 21344
rect 21818 21292 21824 21344
rect 21876 21332 21882 21344
rect 22005 21335 22063 21341
rect 22005 21332 22017 21335
rect 21876 21304 22017 21332
rect 21876 21292 21882 21304
rect 22005 21301 22017 21304
rect 22051 21301 22063 21335
rect 22572 21332 22600 21508
rect 22649 21471 22707 21477
rect 22649 21437 22661 21471
rect 22695 21468 22707 21471
rect 23032 21468 23060 21644
rect 23382 21632 23388 21644
rect 23440 21672 23446 21684
rect 24949 21675 25007 21681
rect 24949 21672 24961 21675
rect 23440 21644 24961 21672
rect 23440 21632 23446 21644
rect 24949 21641 24961 21644
rect 24995 21641 25007 21675
rect 24949 21635 25007 21641
rect 25130 21604 25136 21616
rect 24702 21576 25136 21604
rect 25130 21564 25136 21576
rect 25188 21604 25194 21616
rect 25225 21607 25283 21613
rect 25225 21604 25237 21607
rect 25188 21576 25237 21604
rect 25188 21564 25194 21576
rect 25225 21573 25237 21576
rect 25271 21573 25283 21607
rect 25225 21567 25283 21573
rect 23198 21496 23204 21548
rect 23256 21496 23262 21548
rect 22695 21440 23060 21468
rect 23477 21471 23535 21477
rect 22695 21437 22707 21440
rect 22649 21431 22707 21437
rect 23477 21437 23489 21471
rect 23523 21468 23535 21471
rect 24486 21468 24492 21480
rect 23523 21440 24492 21468
rect 23523 21437 23535 21440
rect 23477 21431 23535 21437
rect 24486 21428 24492 21440
rect 24544 21428 24550 21480
rect 23566 21332 23572 21344
rect 22572 21304 23572 21332
rect 22005 21295 22063 21301
rect 23566 21292 23572 21304
rect 23624 21292 23630 21344
rect 1104 21242 25852 21264
rect 1104 21190 2950 21242
rect 3002 21190 3014 21242
rect 3066 21190 3078 21242
rect 3130 21190 3142 21242
rect 3194 21190 3206 21242
rect 3258 21190 12950 21242
rect 13002 21190 13014 21242
rect 13066 21190 13078 21242
rect 13130 21190 13142 21242
rect 13194 21190 13206 21242
rect 13258 21190 22950 21242
rect 23002 21190 23014 21242
rect 23066 21190 23078 21242
rect 23130 21190 23142 21242
rect 23194 21190 23206 21242
rect 23258 21190 25852 21242
rect 1104 21168 25852 21190
rect 5626 21088 5632 21140
rect 5684 21128 5690 21140
rect 7009 21131 7067 21137
rect 7009 21128 7021 21131
rect 5684 21100 7021 21128
rect 5684 21088 5690 21100
rect 7009 21097 7021 21100
rect 7055 21097 7067 21131
rect 7009 21091 7067 21097
rect 7558 21088 7564 21140
rect 7616 21128 7622 21140
rect 8573 21131 8631 21137
rect 8573 21128 8585 21131
rect 7616 21100 8585 21128
rect 7616 21088 7622 21100
rect 8573 21097 8585 21100
rect 8619 21097 8631 21131
rect 8573 21091 8631 21097
rect 9122 21088 9128 21140
rect 9180 21088 9186 21140
rect 13630 21088 13636 21140
rect 13688 21128 13694 21140
rect 15838 21128 15844 21140
rect 13688 21100 15844 21128
rect 13688 21088 13694 21100
rect 15838 21088 15844 21100
rect 15896 21088 15902 21140
rect 16022 21088 16028 21140
rect 16080 21128 16086 21140
rect 16482 21128 16488 21140
rect 16080 21100 16488 21128
rect 16080 21088 16086 21100
rect 16482 21088 16488 21100
rect 16540 21088 16546 21140
rect 16574 21088 16580 21140
rect 16632 21128 16638 21140
rect 19794 21128 19800 21140
rect 16632 21100 19800 21128
rect 16632 21088 16638 21100
rect 19794 21088 19800 21100
rect 19852 21088 19858 21140
rect 21634 21088 21640 21140
rect 21692 21128 21698 21140
rect 21913 21131 21971 21137
rect 21913 21128 21925 21131
rect 21692 21100 21925 21128
rect 21692 21088 21698 21100
rect 21913 21097 21925 21100
rect 21959 21128 21971 21131
rect 22554 21128 22560 21140
rect 21959 21100 22560 21128
rect 21959 21097 21971 21100
rect 21913 21091 21971 21097
rect 22554 21088 22560 21100
rect 22612 21088 22618 21140
rect 9398 21020 9404 21072
rect 9456 21060 9462 21072
rect 17313 21063 17371 21069
rect 9456 21032 11836 21060
rect 9456 21020 9462 21032
rect 11808 21004 11836 21032
rect 17313 21029 17325 21063
rect 17359 21060 17371 21063
rect 19150 21060 19156 21072
rect 17359 21032 19156 21060
rect 17359 21029 17371 21032
rect 17313 21023 17371 21029
rect 19150 21020 19156 21032
rect 19208 21020 19214 21072
rect 1302 20952 1308 21004
rect 1360 20992 1366 21004
rect 2041 20995 2099 21001
rect 2041 20992 2053 20995
rect 1360 20964 2053 20992
rect 1360 20952 1366 20964
rect 2041 20961 2053 20964
rect 2087 20961 2099 20995
rect 2041 20955 2099 20961
rect 4154 20952 4160 21004
rect 4212 20952 4218 21004
rect 4430 20952 4436 21004
rect 4488 20952 4494 21004
rect 8202 20952 8208 21004
rect 8260 20992 8266 21004
rect 9677 20995 9735 21001
rect 9677 20992 9689 20995
rect 8260 20964 9689 20992
rect 8260 20952 8266 20964
rect 9677 20961 9689 20964
rect 9723 20961 9735 20995
rect 9677 20955 9735 20961
rect 11790 20952 11796 21004
rect 11848 20952 11854 21004
rect 14550 20952 14556 21004
rect 14608 20952 14614 21004
rect 15010 20952 15016 21004
rect 15068 20992 15074 21004
rect 15562 20992 15568 21004
rect 15068 20964 15568 20992
rect 15068 20952 15074 20964
rect 15562 20952 15568 20964
rect 15620 20992 15626 21004
rect 16945 20995 17003 21001
rect 16945 20992 16957 20995
rect 15620 20964 16957 20992
rect 15620 20952 15626 20964
rect 16945 20961 16957 20964
rect 16991 20961 17003 20995
rect 16945 20955 17003 20961
rect 17770 20952 17776 21004
rect 17828 20952 17834 21004
rect 17957 20995 18015 21001
rect 17957 20961 17969 20995
rect 18003 20961 18015 20995
rect 17957 20955 18015 20961
rect 1765 20927 1823 20933
rect 1765 20893 1777 20927
rect 1811 20924 1823 20927
rect 1854 20924 1860 20936
rect 1811 20896 1860 20924
rect 1811 20893 1823 20896
rect 1765 20887 1823 20893
rect 1854 20884 1860 20896
rect 1912 20884 1918 20936
rect 6365 20927 6423 20933
rect 6365 20893 6377 20927
rect 6411 20924 6423 20927
rect 7006 20924 7012 20936
rect 6411 20896 7012 20924
rect 6411 20893 6423 20896
rect 6365 20887 6423 20893
rect 7006 20884 7012 20896
rect 7064 20884 7070 20936
rect 7929 20927 7987 20933
rect 7929 20893 7941 20927
rect 7975 20924 7987 20927
rect 9398 20924 9404 20936
rect 7975 20896 9404 20924
rect 7975 20893 7987 20896
rect 7929 20887 7987 20893
rect 9398 20884 9404 20896
rect 9456 20884 9462 20936
rect 9585 20927 9643 20933
rect 9585 20893 9597 20927
rect 9631 20924 9643 20927
rect 11238 20924 11244 20936
rect 9631 20896 11244 20924
rect 9631 20893 9643 20896
rect 9585 20887 9643 20893
rect 11238 20884 11244 20896
rect 11296 20884 11302 20936
rect 11609 20927 11667 20933
rect 11609 20893 11621 20927
rect 11655 20924 11667 20927
rect 12158 20924 12164 20936
rect 11655 20896 12164 20924
rect 11655 20893 11667 20896
rect 11609 20887 11667 20893
rect 12158 20884 12164 20896
rect 12216 20884 12222 20936
rect 13814 20884 13820 20936
rect 13872 20924 13878 20936
rect 14277 20927 14335 20933
rect 14277 20924 14289 20927
rect 13872 20896 14289 20924
rect 13872 20884 13878 20896
rect 14277 20893 14289 20896
rect 14323 20893 14335 20927
rect 14277 20887 14335 20893
rect 16206 20884 16212 20936
rect 16264 20924 16270 20936
rect 16669 20927 16727 20933
rect 16669 20924 16681 20927
rect 16264 20896 16681 20924
rect 16264 20884 16270 20896
rect 16669 20893 16681 20896
rect 16715 20893 16727 20927
rect 16669 20887 16727 20893
rect 17678 20884 17684 20936
rect 17736 20884 17742 20936
rect 6086 20856 6092 20868
rect 5658 20828 6092 20856
rect 6086 20816 6092 20828
rect 6144 20816 6150 20868
rect 9493 20859 9551 20865
rect 9493 20825 9505 20859
rect 9539 20856 9551 20859
rect 9539 20828 11284 20856
rect 9539 20825 9551 20828
rect 9493 20819 9551 20825
rect 5902 20748 5908 20800
rect 5960 20748 5966 20800
rect 10226 20748 10232 20800
rect 10284 20748 10290 20800
rect 11256 20797 11284 20828
rect 13998 20816 14004 20868
rect 14056 20856 14062 20868
rect 15010 20856 15016 20868
rect 14056 20828 15016 20856
rect 14056 20816 14062 20828
rect 15010 20816 15016 20828
rect 15068 20816 15074 20868
rect 17972 20856 18000 20955
rect 18046 20952 18052 21004
rect 18104 20992 18110 21004
rect 18874 20992 18880 21004
rect 18104 20964 18880 20992
rect 18104 20952 18110 20964
rect 18874 20952 18880 20964
rect 18932 20952 18938 21004
rect 19889 20995 19947 21001
rect 19889 20961 19901 20995
rect 19935 20992 19947 20995
rect 20806 20992 20812 21004
rect 19935 20964 20812 20992
rect 19935 20961 19947 20964
rect 19889 20955 19947 20961
rect 20806 20952 20812 20964
rect 20864 20952 20870 21004
rect 23845 20995 23903 21001
rect 23845 20961 23857 20995
rect 23891 20992 23903 20995
rect 24854 20992 24860 21004
rect 23891 20964 24860 20992
rect 23891 20961 23903 20964
rect 23845 20955 23903 20961
rect 24854 20952 24860 20964
rect 24912 20952 24918 21004
rect 18414 20884 18420 20936
rect 18472 20924 18478 20936
rect 18693 20927 18751 20933
rect 18693 20924 18705 20927
rect 18472 20896 18705 20924
rect 18472 20884 18478 20896
rect 18693 20893 18705 20896
rect 18739 20893 18751 20927
rect 21634 20924 21640 20936
rect 21298 20896 21640 20924
rect 18693 20887 18751 20893
rect 21634 20884 21640 20896
rect 21692 20884 21698 20936
rect 22833 20927 22891 20933
rect 22833 20893 22845 20927
rect 22879 20924 22891 20927
rect 25222 20924 25228 20936
rect 22879 20896 25228 20924
rect 22879 20893 22891 20896
rect 22833 20887 22891 20893
rect 25222 20884 25228 20896
rect 25280 20884 25286 20936
rect 20165 20859 20223 20865
rect 20165 20856 20177 20859
rect 17972 20828 20177 20856
rect 20165 20825 20177 20828
rect 20211 20856 20223 20859
rect 20254 20856 20260 20868
rect 20211 20828 20260 20856
rect 20211 20825 20223 20828
rect 20165 20819 20223 20825
rect 20254 20816 20260 20828
rect 20312 20816 20318 20868
rect 11241 20791 11299 20797
rect 11241 20757 11253 20791
rect 11287 20757 11299 20791
rect 11241 20751 11299 20757
rect 11701 20791 11759 20797
rect 11701 20757 11713 20791
rect 11747 20788 11759 20791
rect 14274 20788 14280 20800
rect 11747 20760 14280 20788
rect 11747 20757 11759 20760
rect 11701 20751 11759 20757
rect 14274 20748 14280 20760
rect 14332 20748 14338 20800
rect 15838 20748 15844 20800
rect 15896 20788 15902 20800
rect 16485 20791 16543 20797
rect 16485 20788 16497 20791
rect 15896 20760 16497 20788
rect 15896 20748 15902 20760
rect 16485 20757 16497 20760
rect 16531 20757 16543 20791
rect 16485 20751 16543 20757
rect 18509 20791 18567 20797
rect 18509 20757 18521 20791
rect 18555 20788 18567 20791
rect 20438 20788 20444 20800
rect 18555 20760 20444 20788
rect 18555 20757 18567 20760
rect 18509 20751 18567 20757
rect 20438 20748 20444 20760
rect 20496 20748 20502 20800
rect 21634 20748 21640 20800
rect 21692 20748 21698 20800
rect 1104 20698 25852 20720
rect 1104 20646 7950 20698
rect 8002 20646 8014 20698
rect 8066 20646 8078 20698
rect 8130 20646 8142 20698
rect 8194 20646 8206 20698
rect 8258 20646 17950 20698
rect 18002 20646 18014 20698
rect 18066 20646 18078 20698
rect 18130 20646 18142 20698
rect 18194 20646 18206 20698
rect 18258 20646 25852 20698
rect 1104 20624 25852 20646
rect 2774 20544 2780 20596
rect 2832 20584 2838 20596
rect 3329 20587 3387 20593
rect 3329 20584 3341 20587
rect 2832 20556 3341 20584
rect 2832 20544 2838 20556
rect 3329 20553 3341 20556
rect 3375 20553 3387 20587
rect 3329 20547 3387 20553
rect 3878 20544 3884 20596
rect 3936 20584 3942 20596
rect 4157 20587 4215 20593
rect 4157 20584 4169 20587
rect 3936 20556 4169 20584
rect 3936 20544 3942 20556
rect 4157 20553 4169 20556
rect 4203 20553 4215 20587
rect 4157 20547 4215 20553
rect 7098 20544 7104 20596
rect 7156 20584 7162 20596
rect 8205 20587 8263 20593
rect 8205 20584 8217 20587
rect 7156 20556 8217 20584
rect 7156 20544 7162 20556
rect 8205 20553 8217 20556
rect 8251 20553 8263 20587
rect 8205 20547 8263 20553
rect 8573 20587 8631 20593
rect 8573 20553 8585 20587
rect 8619 20584 8631 20587
rect 8938 20584 8944 20596
rect 8619 20556 8944 20584
rect 8619 20553 8631 20556
rect 8573 20547 8631 20553
rect 8938 20544 8944 20556
rect 8996 20544 9002 20596
rect 9306 20544 9312 20596
rect 9364 20584 9370 20596
rect 9490 20584 9496 20596
rect 9364 20556 9496 20584
rect 9364 20544 9370 20556
rect 9490 20544 9496 20556
rect 9548 20544 9554 20596
rect 12161 20587 12219 20593
rect 12161 20553 12173 20587
rect 12207 20584 12219 20587
rect 12805 20587 12863 20593
rect 12805 20584 12817 20587
rect 12207 20556 12817 20584
rect 12207 20553 12219 20556
rect 12161 20547 12219 20553
rect 12805 20553 12817 20556
rect 12851 20584 12863 20587
rect 13538 20584 13544 20596
rect 12851 20556 13544 20584
rect 12851 20553 12863 20556
rect 12805 20547 12863 20553
rect 13538 20544 13544 20556
rect 13596 20544 13602 20596
rect 13722 20544 13728 20596
rect 13780 20584 13786 20596
rect 15013 20587 15071 20593
rect 15013 20584 15025 20587
rect 13780 20556 15025 20584
rect 13780 20544 13786 20556
rect 15013 20553 15025 20556
rect 15059 20553 15071 20587
rect 18233 20587 18291 20593
rect 18233 20584 18245 20587
rect 15013 20547 15071 20553
rect 17696 20556 18245 20584
rect 8956 20516 8984 20544
rect 9398 20516 9404 20528
rect 8956 20488 9404 20516
rect 9398 20476 9404 20488
rect 9456 20476 9462 20528
rect 13814 20516 13820 20528
rect 13280 20488 13820 20516
rect 3513 20451 3571 20457
rect 3513 20417 3525 20451
rect 3559 20448 3571 20451
rect 4246 20448 4252 20460
rect 3559 20420 4252 20448
rect 3559 20417 3571 20420
rect 3513 20411 3571 20417
rect 4246 20408 4252 20420
rect 4304 20408 4310 20460
rect 4341 20451 4399 20457
rect 4341 20417 4353 20451
rect 4387 20448 4399 20451
rect 6454 20448 6460 20460
rect 4387 20420 6460 20448
rect 4387 20417 4399 20420
rect 4341 20411 4399 20417
rect 6454 20408 6460 20420
rect 6512 20408 6518 20460
rect 7101 20451 7159 20457
rect 7101 20417 7113 20451
rect 7147 20417 7159 20451
rect 7101 20411 7159 20417
rect 8665 20451 8723 20457
rect 8665 20417 8677 20451
rect 8711 20448 8723 20451
rect 9214 20448 9220 20460
rect 8711 20420 9220 20448
rect 8711 20417 8723 20420
rect 8665 20411 8723 20417
rect 7116 20380 7144 20411
rect 9214 20408 9220 20420
rect 9272 20408 9278 20460
rect 13280 20457 13308 20488
rect 13814 20476 13820 20488
rect 13872 20476 13878 20528
rect 13998 20476 14004 20528
rect 14056 20476 14062 20528
rect 17696 20525 17724 20556
rect 18233 20553 18245 20556
rect 18279 20584 18291 20587
rect 19058 20584 19064 20596
rect 18279 20556 19064 20584
rect 18279 20553 18291 20556
rect 18233 20547 18291 20553
rect 19058 20544 19064 20556
rect 19116 20544 19122 20596
rect 19242 20544 19248 20596
rect 19300 20584 19306 20596
rect 19337 20587 19395 20593
rect 19337 20584 19349 20587
rect 19300 20556 19349 20584
rect 19300 20544 19306 20556
rect 19337 20553 19349 20556
rect 19383 20553 19395 20587
rect 19337 20547 19395 20553
rect 21269 20587 21327 20593
rect 21269 20553 21281 20587
rect 21315 20584 21327 20587
rect 21358 20584 21364 20596
rect 21315 20556 21364 20584
rect 21315 20553 21327 20556
rect 21269 20547 21327 20553
rect 21358 20544 21364 20556
rect 21416 20544 21422 20596
rect 17681 20519 17739 20525
rect 17681 20485 17693 20519
rect 17727 20485 17739 20519
rect 17681 20479 17739 20485
rect 23293 20519 23351 20525
rect 23293 20485 23305 20519
rect 23339 20516 23351 20519
rect 23382 20516 23388 20528
rect 23339 20488 23388 20516
rect 23339 20485 23351 20488
rect 23293 20479 23351 20485
rect 23382 20476 23388 20488
rect 23440 20476 23446 20528
rect 10965 20451 11023 20457
rect 10965 20417 10977 20451
rect 11011 20448 11023 20451
rect 12069 20451 12127 20457
rect 12069 20448 12081 20451
rect 11011 20420 12081 20448
rect 11011 20417 11023 20420
rect 10965 20411 11023 20417
rect 12069 20417 12081 20420
rect 12115 20417 12127 20451
rect 12069 20411 12127 20417
rect 13265 20451 13323 20457
rect 13265 20417 13277 20451
rect 13311 20417 13323 20451
rect 13265 20411 13323 20417
rect 15473 20451 15531 20457
rect 15473 20417 15485 20451
rect 15519 20448 15531 20451
rect 16022 20448 16028 20460
rect 15519 20420 16028 20448
rect 15519 20417 15531 20420
rect 15473 20411 15531 20417
rect 16022 20408 16028 20420
rect 16080 20408 16086 20460
rect 17037 20451 17095 20457
rect 17037 20417 17049 20451
rect 17083 20417 17095 20451
rect 17037 20411 17095 20417
rect 8849 20383 8907 20389
rect 8849 20380 8861 20383
rect 7116 20352 8861 20380
rect 8849 20349 8861 20352
rect 8895 20380 8907 20383
rect 9858 20380 9864 20392
rect 8895 20352 9864 20380
rect 8895 20349 8907 20352
rect 8849 20343 8907 20349
rect 9858 20340 9864 20352
rect 9916 20340 9922 20392
rect 12250 20340 12256 20392
rect 12308 20340 12314 20392
rect 13541 20383 13599 20389
rect 13541 20349 13553 20383
rect 13587 20380 13599 20383
rect 16117 20383 16175 20389
rect 16117 20380 16129 20383
rect 13587 20352 16129 20380
rect 13587 20349 13599 20352
rect 13541 20343 13599 20349
rect 16117 20349 16129 20352
rect 16163 20349 16175 20383
rect 17052 20380 17080 20411
rect 19150 20408 19156 20460
rect 19208 20448 19214 20460
rect 19245 20451 19303 20457
rect 19245 20448 19257 20451
rect 19208 20420 19257 20448
rect 19208 20408 19214 20420
rect 19245 20417 19257 20420
rect 19291 20417 19303 20451
rect 20625 20451 20683 20457
rect 20625 20448 20637 20451
rect 19245 20411 19303 20417
rect 19536 20420 20637 20448
rect 19536 20389 19564 20420
rect 20625 20417 20637 20420
rect 20671 20448 20683 20451
rect 21634 20448 21640 20460
rect 20671 20420 21640 20448
rect 20671 20417 20683 20420
rect 20625 20411 20683 20417
rect 21634 20408 21640 20420
rect 21692 20408 21698 20460
rect 22278 20408 22284 20460
rect 22336 20408 22342 20460
rect 24121 20451 24179 20457
rect 24121 20417 24133 20451
rect 24167 20448 24179 20451
rect 24946 20448 24952 20460
rect 24167 20420 24952 20448
rect 24167 20417 24179 20420
rect 24121 20411 24179 20417
rect 24946 20408 24952 20420
rect 25004 20408 25010 20460
rect 16117 20343 16175 20349
rect 16224 20352 17080 20380
rect 19521 20383 19579 20389
rect 9306 20272 9312 20324
rect 9364 20312 9370 20324
rect 11701 20315 11759 20321
rect 11701 20312 11713 20315
rect 9364 20284 11713 20312
rect 9364 20272 9370 20284
rect 11701 20281 11713 20284
rect 11747 20281 11759 20315
rect 16224 20312 16252 20352
rect 19521 20349 19533 20383
rect 19567 20349 19579 20383
rect 19521 20343 19579 20349
rect 23290 20340 23296 20392
rect 23348 20380 23354 20392
rect 24397 20383 24455 20389
rect 24397 20380 24409 20383
rect 23348 20352 24409 20380
rect 23348 20340 23354 20352
rect 24397 20349 24409 20352
rect 24443 20349 24455 20383
rect 24397 20343 24455 20349
rect 11701 20275 11759 20281
rect 12406 20284 12848 20312
rect 6086 20204 6092 20256
rect 6144 20244 6150 20256
rect 6730 20244 6736 20256
rect 6144 20216 6736 20244
rect 6144 20204 6150 20216
rect 6730 20204 6736 20216
rect 6788 20204 6794 20256
rect 7742 20204 7748 20256
rect 7800 20204 7806 20256
rect 12066 20204 12072 20256
rect 12124 20244 12130 20256
rect 12406 20244 12434 20284
rect 12124 20216 12434 20244
rect 12820 20244 12848 20284
rect 14752 20284 16252 20312
rect 16853 20315 16911 20321
rect 14752 20244 14780 20284
rect 16853 20281 16865 20315
rect 16899 20312 16911 20315
rect 22830 20312 22836 20324
rect 16899 20284 22836 20312
rect 16899 20281 16911 20284
rect 16853 20275 16911 20281
rect 22830 20272 22836 20284
rect 22888 20272 22894 20324
rect 12820 20216 14780 20244
rect 17773 20247 17831 20253
rect 12124 20204 12130 20216
rect 17773 20213 17785 20247
rect 17819 20244 17831 20247
rect 17862 20244 17868 20256
rect 17819 20216 17868 20244
rect 17819 20213 17831 20216
rect 17773 20207 17831 20213
rect 17862 20204 17868 20216
rect 17920 20204 17926 20256
rect 18046 20204 18052 20256
rect 18104 20244 18110 20256
rect 18877 20247 18935 20253
rect 18877 20244 18889 20247
rect 18104 20216 18889 20244
rect 18104 20204 18110 20216
rect 18877 20213 18889 20216
rect 18923 20213 18935 20247
rect 18877 20207 18935 20213
rect 1104 20154 25852 20176
rect 1104 20102 2950 20154
rect 3002 20102 3014 20154
rect 3066 20102 3078 20154
rect 3130 20102 3142 20154
rect 3194 20102 3206 20154
rect 3258 20102 12950 20154
rect 13002 20102 13014 20154
rect 13066 20102 13078 20154
rect 13130 20102 13142 20154
rect 13194 20102 13206 20154
rect 13258 20102 22950 20154
rect 23002 20102 23014 20154
rect 23066 20102 23078 20154
rect 23130 20102 23142 20154
rect 23194 20102 23206 20154
rect 23258 20102 25852 20154
rect 1104 20080 25852 20102
rect 6914 20000 6920 20052
rect 6972 20040 6978 20052
rect 7837 20043 7895 20049
rect 7837 20040 7849 20043
rect 6972 20012 7849 20040
rect 6972 20000 6978 20012
rect 7837 20009 7849 20012
rect 7883 20009 7895 20043
rect 7837 20003 7895 20009
rect 10134 20000 10140 20052
rect 10192 20040 10198 20052
rect 10597 20043 10655 20049
rect 10597 20040 10609 20043
rect 10192 20012 10609 20040
rect 10192 20000 10198 20012
rect 10597 20009 10609 20012
rect 10643 20040 10655 20043
rect 10870 20040 10876 20052
rect 10643 20012 10876 20040
rect 10643 20009 10655 20012
rect 10597 20003 10655 20009
rect 10870 20000 10876 20012
rect 10928 20000 10934 20052
rect 11238 20000 11244 20052
rect 11296 20000 11302 20052
rect 16574 20000 16580 20052
rect 16632 20040 16638 20052
rect 18046 20040 18052 20052
rect 16632 20012 18052 20040
rect 16632 20000 16638 20012
rect 18046 20000 18052 20012
rect 18104 20000 18110 20052
rect 18966 20000 18972 20052
rect 19024 20000 19030 20052
rect 6730 19932 6736 19984
rect 6788 19972 6794 19984
rect 7377 19975 7435 19981
rect 7377 19972 7389 19975
rect 6788 19944 7389 19972
rect 6788 19932 6794 19944
rect 7377 19941 7389 19944
rect 7423 19941 7435 19975
rect 7377 19935 7435 19941
rect 7558 19932 7564 19984
rect 7616 19972 7622 19984
rect 9125 19975 9183 19981
rect 9125 19972 9137 19975
rect 7616 19944 9137 19972
rect 7616 19932 7622 19944
rect 9125 19941 9137 19944
rect 9171 19941 9183 19975
rect 9125 19935 9183 19941
rect 10226 19932 10232 19984
rect 10284 19972 10290 19984
rect 10413 19975 10471 19981
rect 10413 19972 10425 19975
rect 10284 19944 10425 19972
rect 10284 19932 10290 19944
rect 10413 19941 10425 19944
rect 10459 19972 10471 19975
rect 13998 19972 14004 19984
rect 10459 19944 14004 19972
rect 10459 19941 10471 19944
rect 10413 19935 10471 19941
rect 13998 19932 14004 19944
rect 14056 19972 14062 19984
rect 15105 19975 15163 19981
rect 15105 19972 15117 19975
rect 14056 19944 15117 19972
rect 14056 19932 14062 19944
rect 15105 19941 15117 19944
rect 15151 19941 15163 19975
rect 15105 19935 15163 19941
rect 17957 19975 18015 19981
rect 17957 19941 17969 19975
rect 18003 19972 18015 19975
rect 19058 19972 19064 19984
rect 18003 19944 19064 19972
rect 18003 19941 18015 19944
rect 17957 19935 18015 19941
rect 19058 19932 19064 19944
rect 19116 19932 19122 19984
rect 4154 19864 4160 19916
rect 4212 19904 4218 19916
rect 5353 19907 5411 19913
rect 5353 19904 5365 19907
rect 4212 19876 5365 19904
rect 4212 19864 4218 19876
rect 5353 19873 5365 19876
rect 5399 19873 5411 19907
rect 5353 19867 5411 19873
rect 5629 19907 5687 19913
rect 5629 19873 5641 19907
rect 5675 19904 5687 19907
rect 7742 19904 7748 19916
rect 5675 19876 7748 19904
rect 5675 19873 5687 19876
rect 5629 19867 5687 19873
rect 7742 19864 7748 19876
rect 7800 19864 7806 19916
rect 8389 19907 8447 19913
rect 8389 19904 8401 19907
rect 7852 19876 8401 19904
rect 6730 19796 6736 19848
rect 6788 19796 6794 19848
rect 7006 19660 7012 19712
rect 7064 19700 7070 19712
rect 7101 19703 7159 19709
rect 7101 19700 7113 19703
rect 7064 19672 7113 19700
rect 7064 19660 7070 19672
rect 7101 19669 7113 19672
rect 7147 19700 7159 19703
rect 7852 19700 7880 19876
rect 8389 19873 8401 19876
rect 8435 19873 8447 19907
rect 8389 19867 8447 19873
rect 9398 19864 9404 19916
rect 9456 19904 9462 19916
rect 9677 19907 9735 19913
rect 9677 19904 9689 19907
rect 9456 19876 9689 19904
rect 9456 19864 9462 19876
rect 9677 19873 9689 19876
rect 9723 19873 9735 19907
rect 9677 19867 9735 19873
rect 11054 19864 11060 19916
rect 11112 19904 11118 19916
rect 11790 19904 11796 19916
rect 11112 19876 11796 19904
rect 11112 19864 11118 19876
rect 11790 19864 11796 19876
rect 11848 19864 11854 19916
rect 15194 19864 15200 19916
rect 15252 19904 15258 19916
rect 18966 19904 18972 19916
rect 15252 19876 17080 19904
rect 15252 19864 15258 19876
rect 8205 19839 8263 19845
rect 8205 19805 8217 19839
rect 8251 19836 8263 19839
rect 8478 19836 8484 19848
rect 8251 19808 8484 19836
rect 8251 19805 8263 19808
rect 8205 19799 8263 19805
rect 8478 19796 8484 19808
rect 8536 19796 8542 19848
rect 9490 19796 9496 19848
rect 9548 19796 9554 19848
rect 9585 19839 9643 19845
rect 9585 19805 9597 19839
rect 9631 19836 9643 19839
rect 10410 19836 10416 19848
rect 9631 19808 10416 19836
rect 9631 19805 9643 19808
rect 9585 19799 9643 19805
rect 10410 19796 10416 19808
rect 10468 19796 10474 19848
rect 12989 19839 13047 19845
rect 12989 19805 13001 19839
rect 13035 19836 13047 19839
rect 13722 19836 13728 19848
rect 13035 19808 13728 19836
rect 13035 19805 13047 19808
rect 12989 19799 13047 19805
rect 13722 19796 13728 19808
rect 13780 19796 13786 19848
rect 15841 19839 15899 19845
rect 15841 19805 15853 19839
rect 15887 19836 15899 19839
rect 16850 19836 16856 19848
rect 15887 19808 16856 19836
rect 15887 19805 15899 19808
rect 15841 19799 15899 19805
rect 16850 19796 16856 19808
rect 16908 19796 16914 19848
rect 17052 19845 17080 19876
rect 17788 19876 18972 19904
rect 17788 19845 17816 19876
rect 18966 19864 18972 19876
rect 19024 19864 19030 19916
rect 23845 19907 23903 19913
rect 23845 19873 23857 19907
rect 23891 19904 23903 19907
rect 24946 19904 24952 19916
rect 23891 19876 24952 19904
rect 23891 19873 23903 19876
rect 23845 19867 23903 19873
rect 24946 19864 24952 19876
rect 25004 19864 25010 19916
rect 17037 19839 17095 19845
rect 17037 19805 17049 19839
rect 17083 19805 17095 19839
rect 17037 19799 17095 19805
rect 17773 19839 17831 19845
rect 17773 19805 17785 19839
rect 17819 19805 17831 19839
rect 17773 19799 17831 19805
rect 18601 19839 18659 19845
rect 18601 19805 18613 19839
rect 18647 19836 18659 19839
rect 19518 19836 19524 19848
rect 18647 19808 19524 19836
rect 18647 19805 18659 19808
rect 18601 19799 18659 19805
rect 19518 19796 19524 19808
rect 19576 19796 19582 19848
rect 20438 19796 20444 19848
rect 20496 19796 20502 19848
rect 21450 19796 21456 19848
rect 21508 19836 21514 19848
rect 21545 19839 21603 19845
rect 21545 19836 21557 19839
rect 21508 19808 21557 19836
rect 21508 19796 21514 19808
rect 21545 19805 21557 19808
rect 21591 19805 21603 19839
rect 21545 19799 21603 19805
rect 22833 19839 22891 19845
rect 22833 19805 22845 19839
rect 22879 19836 22891 19839
rect 25314 19836 25320 19848
rect 22879 19808 25320 19836
rect 22879 19805 22891 19808
rect 22833 19799 22891 19805
rect 25314 19796 25320 19808
rect 25372 19796 25378 19848
rect 8297 19771 8355 19777
rect 8297 19737 8309 19771
rect 8343 19768 8355 19771
rect 11609 19771 11667 19777
rect 8343 19740 10364 19768
rect 8343 19737 8355 19740
rect 8297 19731 8355 19737
rect 10336 19712 10364 19740
rect 11609 19737 11621 19771
rect 11655 19768 11667 19771
rect 12802 19768 12808 19780
rect 11655 19740 12808 19768
rect 11655 19737 11667 19740
rect 11609 19731 11667 19737
rect 12802 19728 12808 19740
rect 12860 19728 12866 19780
rect 16022 19728 16028 19780
rect 16080 19728 16086 19780
rect 20254 19768 20260 19780
rect 16868 19740 20260 19768
rect 7147 19672 7880 19700
rect 7147 19669 7159 19672
rect 7101 19663 7159 19669
rect 10134 19660 10140 19712
rect 10192 19700 10198 19712
rect 10229 19703 10287 19709
rect 10229 19700 10241 19703
rect 10192 19672 10241 19700
rect 10192 19660 10198 19672
rect 10229 19669 10241 19672
rect 10275 19669 10287 19703
rect 10229 19663 10287 19669
rect 10318 19660 10324 19712
rect 10376 19660 10382 19712
rect 11701 19703 11759 19709
rect 11701 19669 11713 19703
rect 11747 19700 11759 19703
rect 12158 19700 12164 19712
rect 11747 19672 12164 19700
rect 11747 19669 11759 19672
rect 11701 19663 11759 19669
rect 12158 19660 12164 19672
rect 12216 19660 12222 19712
rect 13630 19660 13636 19712
rect 13688 19660 13694 19712
rect 16868 19709 16896 19740
rect 20254 19728 20260 19740
rect 20312 19728 20318 19780
rect 20625 19771 20683 19777
rect 20625 19737 20637 19771
rect 20671 19768 20683 19771
rect 22738 19768 22744 19780
rect 20671 19740 22744 19768
rect 20671 19737 20683 19740
rect 20625 19731 20683 19737
rect 22738 19728 22744 19740
rect 22796 19728 22802 19780
rect 24673 19771 24731 19777
rect 24673 19768 24685 19771
rect 22848 19740 24685 19768
rect 16853 19703 16911 19709
rect 16853 19669 16865 19703
rect 16899 19669 16911 19703
rect 16853 19663 16911 19669
rect 18417 19703 18475 19709
rect 18417 19669 18429 19703
rect 18463 19700 18475 19703
rect 18506 19700 18512 19712
rect 18463 19672 18512 19700
rect 18463 19669 18475 19672
rect 18417 19663 18475 19669
rect 18506 19660 18512 19672
rect 18564 19660 18570 19712
rect 22186 19660 22192 19712
rect 22244 19660 22250 19712
rect 22646 19660 22652 19712
rect 22704 19700 22710 19712
rect 22848 19700 22876 19740
rect 24673 19737 24685 19740
rect 24719 19737 24731 19771
rect 24673 19731 24731 19737
rect 22704 19672 22876 19700
rect 22704 19660 22710 19672
rect 24302 19660 24308 19712
rect 24360 19700 24366 19712
rect 24765 19703 24823 19709
rect 24765 19700 24777 19703
rect 24360 19672 24777 19700
rect 24360 19660 24366 19672
rect 24765 19669 24777 19672
rect 24811 19669 24823 19703
rect 24765 19663 24823 19669
rect 1104 19610 25852 19632
rect 1104 19558 7950 19610
rect 8002 19558 8014 19610
rect 8066 19558 8078 19610
rect 8130 19558 8142 19610
rect 8194 19558 8206 19610
rect 8258 19558 17950 19610
rect 18002 19558 18014 19610
rect 18066 19558 18078 19610
rect 18130 19558 18142 19610
rect 18194 19558 18206 19610
rect 18258 19558 25852 19610
rect 1104 19536 25852 19558
rect 9674 19456 9680 19508
rect 9732 19496 9738 19508
rect 10413 19499 10471 19505
rect 10413 19496 10425 19499
rect 9732 19468 10425 19496
rect 9732 19456 9738 19468
rect 10413 19465 10425 19468
rect 10459 19465 10471 19499
rect 10413 19459 10471 19465
rect 10502 19456 10508 19508
rect 10560 19496 10566 19508
rect 10870 19496 10876 19508
rect 10560 19468 10876 19496
rect 10560 19456 10566 19468
rect 10870 19456 10876 19468
rect 10928 19456 10934 19508
rect 12161 19499 12219 19505
rect 12161 19465 12173 19499
rect 12207 19496 12219 19499
rect 12710 19496 12716 19508
rect 12207 19468 12716 19496
rect 12207 19465 12219 19468
rect 12161 19459 12219 19465
rect 12710 19456 12716 19468
rect 12768 19456 12774 19508
rect 13265 19499 13323 19505
rect 13265 19465 13277 19499
rect 13311 19465 13323 19499
rect 21726 19496 21732 19508
rect 13265 19459 13323 19465
rect 19076 19468 21732 19496
rect 2038 19388 2044 19440
rect 2096 19428 2102 19440
rect 2133 19431 2191 19437
rect 2133 19428 2145 19431
rect 2096 19400 2145 19428
rect 2096 19388 2102 19400
rect 2133 19397 2145 19400
rect 2179 19397 2191 19431
rect 8662 19428 8668 19440
rect 2133 19391 2191 19397
rect 8128 19400 8668 19428
rect 8128 19369 8156 19400
rect 8662 19388 8668 19400
rect 8720 19388 8726 19440
rect 8846 19388 8852 19440
rect 8904 19388 8910 19440
rect 10781 19431 10839 19437
rect 10781 19397 10793 19431
rect 10827 19428 10839 19431
rect 10827 19400 12204 19428
rect 10827 19397 10839 19400
rect 10781 19391 10839 19397
rect 8113 19363 8171 19369
rect 8113 19329 8125 19363
rect 8159 19329 8171 19363
rect 8113 19323 8171 19329
rect 10134 19320 10140 19372
rect 10192 19360 10198 19372
rect 10870 19360 10876 19372
rect 10192 19332 10876 19360
rect 10192 19320 10198 19332
rect 10870 19320 10876 19332
rect 10928 19360 10934 19372
rect 10928 19332 11008 19360
rect 10928 19320 10934 19332
rect 10980 19301 11008 19332
rect 12066 19320 12072 19372
rect 12124 19320 12130 19372
rect 12176 19360 12204 19400
rect 12342 19388 12348 19440
rect 12400 19428 12406 19440
rect 13280 19428 13308 19459
rect 12400 19400 13308 19428
rect 13633 19431 13691 19437
rect 12400 19388 12406 19400
rect 13633 19397 13645 19431
rect 13679 19428 13691 19431
rect 13998 19428 14004 19440
rect 13679 19400 14004 19428
rect 13679 19397 13691 19400
rect 13633 19391 13691 19397
rect 13998 19388 14004 19400
rect 14056 19388 14062 19440
rect 19076 19428 19104 19468
rect 21726 19456 21732 19468
rect 21784 19456 21790 19508
rect 22002 19456 22008 19508
rect 22060 19496 22066 19508
rect 23753 19499 23811 19505
rect 23753 19496 23765 19499
rect 22060 19468 23765 19496
rect 22060 19456 22066 19468
rect 23753 19465 23765 19468
rect 23799 19465 23811 19499
rect 23753 19459 23811 19465
rect 18984 19400 19104 19428
rect 12618 19360 12624 19372
rect 12176 19332 12624 19360
rect 12618 19320 12624 19332
rect 12676 19320 12682 19372
rect 13740 19332 13952 19360
rect 13740 19304 13768 19332
rect 8389 19295 8447 19301
rect 8389 19261 8401 19295
rect 8435 19292 8447 19295
rect 10965 19295 11023 19301
rect 8435 19264 10272 19292
rect 8435 19261 8447 19264
rect 8389 19255 8447 19261
rect 10244 19236 10272 19264
rect 10965 19261 10977 19295
rect 11011 19261 11023 19295
rect 10965 19255 11023 19261
rect 11606 19252 11612 19304
rect 11664 19292 11670 19304
rect 12253 19295 12311 19301
rect 12253 19292 12265 19295
rect 11664 19264 12265 19292
rect 11664 19252 11670 19264
rect 12253 19261 12265 19264
rect 12299 19261 12311 19295
rect 12989 19295 13047 19301
rect 12253 19255 12311 19261
rect 12360 19264 12664 19292
rect 10226 19184 10232 19236
rect 10284 19224 10290 19236
rect 12360 19224 12388 19264
rect 10284 19196 12388 19224
rect 12636 19224 12664 19264
rect 12989 19261 13001 19295
rect 13035 19292 13047 19295
rect 13722 19292 13728 19304
rect 13035 19264 13728 19292
rect 13035 19261 13047 19264
rect 12989 19255 13047 19261
rect 13722 19252 13728 19264
rect 13780 19252 13786 19304
rect 13817 19295 13875 19301
rect 13817 19261 13829 19295
rect 13863 19261 13875 19295
rect 13924 19292 13952 19332
rect 17126 19320 17132 19372
rect 17184 19360 17190 19372
rect 17681 19363 17739 19369
rect 17681 19360 17693 19363
rect 17184 19332 17693 19360
rect 17184 19320 17190 19332
rect 17681 19329 17693 19332
rect 17727 19329 17739 19363
rect 17681 19323 17739 19329
rect 18325 19363 18383 19369
rect 18325 19329 18337 19363
rect 18371 19360 18383 19363
rect 18690 19360 18696 19372
rect 18371 19332 18696 19360
rect 18371 19329 18383 19332
rect 18325 19323 18383 19329
rect 18690 19320 18696 19332
rect 18748 19320 18754 19372
rect 18984 19369 19012 19400
rect 21174 19388 21180 19440
rect 21232 19428 21238 19440
rect 22554 19428 22560 19440
rect 21232 19400 22560 19428
rect 21232 19388 21238 19400
rect 22554 19388 22560 19400
rect 22612 19428 22618 19440
rect 22612 19400 22770 19428
rect 22612 19388 22618 19400
rect 18969 19363 19027 19369
rect 18969 19329 18981 19363
rect 19015 19329 19027 19363
rect 20378 19332 20760 19360
rect 18969 19323 19027 19329
rect 20732 19304 20760 19332
rect 15930 19292 15936 19304
rect 13924 19264 15936 19292
rect 13817 19255 13875 19261
rect 13446 19224 13452 19236
rect 12636 19196 13452 19224
rect 10284 19184 10290 19196
rect 13446 19184 13452 19196
rect 13504 19224 13510 19236
rect 13832 19224 13860 19255
rect 15930 19252 15936 19264
rect 15988 19252 15994 19304
rect 16022 19252 16028 19304
rect 16080 19292 16086 19304
rect 16942 19292 16948 19304
rect 16080 19264 16948 19292
rect 16080 19252 16086 19264
rect 16942 19252 16948 19264
rect 17000 19252 17006 19304
rect 19245 19295 19303 19301
rect 19245 19261 19257 19295
rect 19291 19292 19303 19295
rect 20622 19292 20628 19304
rect 19291 19264 20628 19292
rect 19291 19261 19303 19264
rect 19245 19255 19303 19261
rect 20622 19252 20628 19264
rect 20680 19252 20686 19304
rect 20714 19252 20720 19304
rect 20772 19292 20778 19304
rect 21174 19292 21180 19304
rect 20772 19264 21180 19292
rect 20772 19252 20778 19264
rect 21174 19252 21180 19264
rect 21232 19252 21238 19304
rect 21726 19252 21732 19304
rect 21784 19292 21790 19304
rect 22005 19295 22063 19301
rect 22005 19292 22017 19295
rect 21784 19264 22017 19292
rect 21784 19252 21790 19264
rect 22005 19261 22017 19264
rect 22051 19261 22063 19295
rect 22281 19295 22339 19301
rect 22281 19292 22293 19295
rect 22005 19255 22063 19261
rect 22112 19264 22293 19292
rect 14461 19227 14519 19233
rect 14461 19224 14473 19227
rect 13504 19196 13860 19224
rect 13924 19196 14473 19224
rect 13504 19184 13510 19196
rect 2222 19116 2228 19168
rect 2280 19116 2286 19168
rect 6362 19116 6368 19168
rect 6420 19156 6426 19168
rect 6822 19156 6828 19168
rect 6420 19128 6828 19156
rect 6420 19116 6426 19128
rect 6822 19116 6828 19128
rect 6880 19116 6886 19168
rect 7653 19159 7711 19165
rect 7653 19125 7665 19159
rect 7699 19156 7711 19159
rect 8570 19156 8576 19168
rect 7699 19128 8576 19156
rect 7699 19125 7711 19128
rect 7653 19119 7711 19125
rect 8570 19116 8576 19128
rect 8628 19116 8634 19168
rect 9858 19116 9864 19168
rect 9916 19116 9922 19168
rect 11698 19116 11704 19168
rect 11756 19116 11762 19168
rect 11974 19116 11980 19168
rect 12032 19156 12038 19168
rect 12713 19159 12771 19165
rect 12713 19156 12725 19159
rect 12032 19128 12725 19156
rect 12032 19116 12038 19128
rect 12713 19125 12725 19128
rect 12759 19125 12771 19159
rect 12713 19119 12771 19125
rect 13722 19116 13728 19168
rect 13780 19156 13786 19168
rect 13924 19156 13952 19196
rect 14461 19193 14473 19196
rect 14507 19193 14519 19227
rect 15010 19224 15016 19236
rect 14461 19187 14519 19193
rect 14660 19196 15016 19224
rect 13780 19128 13952 19156
rect 13780 19116 13786 19128
rect 13998 19116 14004 19168
rect 14056 19156 14062 19168
rect 14369 19159 14427 19165
rect 14369 19156 14381 19159
rect 14056 19128 14381 19156
rect 14056 19116 14062 19128
rect 14369 19125 14381 19128
rect 14415 19156 14427 19159
rect 14660 19156 14688 19196
rect 15010 19184 15016 19196
rect 15068 19184 15074 19236
rect 15102 19184 15108 19236
rect 15160 19224 15166 19236
rect 15160 19196 18184 19224
rect 15160 19184 15166 19196
rect 14415 19128 14688 19156
rect 14415 19125 14427 19128
rect 14369 19119 14427 19125
rect 14734 19116 14740 19168
rect 14792 19116 14798 19168
rect 17494 19116 17500 19168
rect 17552 19116 17558 19168
rect 18156 19165 18184 19196
rect 21910 19184 21916 19236
rect 21968 19224 21974 19236
rect 22112 19224 22140 19264
rect 22281 19261 22293 19264
rect 22327 19261 22339 19295
rect 22281 19255 22339 19261
rect 22646 19252 22652 19304
rect 22704 19292 22710 19304
rect 23566 19292 23572 19304
rect 22704 19264 23572 19292
rect 22704 19252 22710 19264
rect 23566 19252 23572 19264
rect 23624 19292 23630 19304
rect 24029 19295 24087 19301
rect 24029 19292 24041 19295
rect 23624 19264 24041 19292
rect 23624 19252 23630 19264
rect 24029 19261 24041 19264
rect 24075 19292 24087 19295
rect 24213 19295 24271 19301
rect 24213 19292 24225 19295
rect 24075 19264 24225 19292
rect 24075 19261 24087 19264
rect 24029 19255 24087 19261
rect 24213 19261 24225 19264
rect 24259 19261 24271 19295
rect 24213 19255 24271 19261
rect 21968 19196 22140 19224
rect 21968 19184 21974 19196
rect 18141 19159 18199 19165
rect 18141 19125 18153 19159
rect 18187 19156 18199 19159
rect 19242 19156 19248 19168
rect 18187 19128 19248 19156
rect 18187 19125 18199 19128
rect 18141 19119 18199 19125
rect 19242 19116 19248 19128
rect 19300 19116 19306 19168
rect 20717 19159 20775 19165
rect 20717 19125 20729 19159
rect 20763 19156 20775 19159
rect 20898 19156 20904 19168
rect 20763 19128 20904 19156
rect 20763 19125 20775 19128
rect 20717 19119 20775 19125
rect 20898 19116 20904 19128
rect 20956 19116 20962 19168
rect 1104 19066 25852 19088
rect 1104 19014 2950 19066
rect 3002 19014 3014 19066
rect 3066 19014 3078 19066
rect 3130 19014 3142 19066
rect 3194 19014 3206 19066
rect 3258 19014 12950 19066
rect 13002 19014 13014 19066
rect 13066 19014 13078 19066
rect 13130 19014 13142 19066
rect 13194 19014 13206 19066
rect 13258 19014 22950 19066
rect 23002 19014 23014 19066
rect 23066 19014 23078 19066
rect 23130 19014 23142 19066
rect 23194 19014 23206 19066
rect 23258 19014 25852 19066
rect 1104 18992 25852 19014
rect 7193 18955 7251 18961
rect 7193 18921 7205 18955
rect 7239 18952 7251 18955
rect 8570 18952 8576 18964
rect 7239 18924 8576 18952
rect 7239 18921 7251 18924
rect 7193 18915 7251 18921
rect 8570 18912 8576 18924
rect 8628 18912 8634 18964
rect 10873 18955 10931 18961
rect 10873 18921 10885 18955
rect 10919 18952 10931 18955
rect 11054 18952 11060 18964
rect 10919 18924 11060 18952
rect 10919 18921 10931 18924
rect 10873 18915 10931 18921
rect 11054 18912 11060 18924
rect 11112 18912 11118 18964
rect 12802 18912 12808 18964
rect 12860 18952 12866 18964
rect 12989 18955 13047 18961
rect 12989 18952 13001 18955
rect 12860 18924 13001 18952
rect 12860 18912 12866 18924
rect 12989 18921 13001 18924
rect 13035 18921 13047 18955
rect 12989 18915 13047 18921
rect 13538 18912 13544 18964
rect 13596 18912 13602 18964
rect 14274 18912 14280 18964
rect 14332 18912 14338 18964
rect 15930 18912 15936 18964
rect 15988 18952 15994 18964
rect 16485 18955 16543 18961
rect 16485 18952 16497 18955
rect 15988 18924 16497 18952
rect 15988 18912 15994 18924
rect 16485 18921 16497 18924
rect 16531 18921 16543 18955
rect 16485 18915 16543 18921
rect 16853 18955 16911 18961
rect 16853 18921 16865 18955
rect 16899 18952 16911 18955
rect 20346 18952 20352 18964
rect 16899 18924 20352 18952
rect 16899 18921 16911 18924
rect 16853 18915 16911 18921
rect 2314 18844 2320 18896
rect 2372 18884 2378 18896
rect 7377 18887 7435 18893
rect 7377 18884 7389 18887
rect 2372 18856 7389 18884
rect 2372 18844 2378 18856
rect 7377 18853 7389 18856
rect 7423 18853 7435 18887
rect 7377 18847 7435 18853
rect 10686 18844 10692 18896
rect 10744 18884 10750 18896
rect 11793 18887 11851 18893
rect 11793 18884 11805 18887
rect 10744 18856 11805 18884
rect 10744 18844 10750 18856
rect 11793 18853 11805 18856
rect 11839 18853 11851 18887
rect 13556 18884 13584 18912
rect 14366 18884 14372 18896
rect 13556 18856 14372 18884
rect 11793 18847 11851 18853
rect 14366 18844 14372 18856
rect 14424 18844 14430 18896
rect 1302 18776 1308 18828
rect 1360 18816 1366 18828
rect 2041 18819 2099 18825
rect 2041 18816 2053 18819
rect 1360 18788 2053 18816
rect 1360 18776 1366 18788
rect 2041 18785 2053 18788
rect 2087 18785 2099 18819
rect 2041 18779 2099 18785
rect 5902 18776 5908 18828
rect 5960 18816 5966 18828
rect 5960 18788 7972 18816
rect 5960 18776 5966 18788
rect 1762 18708 1768 18760
rect 1820 18708 1826 18760
rect 5813 18751 5871 18757
rect 5813 18717 5825 18751
rect 5859 18748 5871 18751
rect 6086 18748 6092 18760
rect 5859 18720 6092 18748
rect 5859 18717 5871 18720
rect 5813 18711 5871 18717
rect 6086 18708 6092 18720
rect 6144 18708 6150 18760
rect 6822 18708 6828 18760
rect 6880 18748 6886 18760
rect 7944 18757 7972 18788
rect 8662 18776 8668 18828
rect 8720 18816 8726 18828
rect 9125 18819 9183 18825
rect 9125 18816 9137 18819
rect 8720 18788 9137 18816
rect 8720 18776 8726 18788
rect 9125 18785 9137 18788
rect 9171 18816 9183 18819
rect 10962 18816 10968 18828
rect 9171 18788 10968 18816
rect 9171 18785 9183 18788
rect 9125 18779 9183 18785
rect 10962 18776 10968 18788
rect 11020 18776 11026 18828
rect 11882 18776 11888 18828
rect 11940 18816 11946 18828
rect 12250 18816 12256 18828
rect 11940 18788 12256 18816
rect 11940 18776 11946 18788
rect 12250 18776 12256 18788
rect 12308 18816 12314 18828
rect 12345 18819 12403 18825
rect 12345 18816 12357 18819
rect 12308 18788 12357 18816
rect 12308 18776 12314 18788
rect 12345 18785 12357 18788
rect 12391 18785 12403 18819
rect 12345 18779 12403 18785
rect 13449 18819 13507 18825
rect 13449 18785 13461 18819
rect 13495 18816 13507 18819
rect 13538 18816 13544 18828
rect 13495 18788 13544 18816
rect 13495 18785 13507 18788
rect 13449 18779 13507 18785
rect 13538 18776 13544 18788
rect 13596 18776 13602 18828
rect 13633 18819 13691 18825
rect 13633 18785 13645 18819
rect 13679 18816 13691 18819
rect 13722 18816 13728 18828
rect 13679 18788 13728 18816
rect 13679 18785 13691 18788
rect 13633 18779 13691 18785
rect 6917 18751 6975 18757
rect 6917 18748 6929 18751
rect 6880 18720 6929 18748
rect 6880 18708 6886 18720
rect 6917 18717 6929 18720
rect 6963 18717 6975 18751
rect 6917 18711 6975 18717
rect 7929 18751 7987 18757
rect 7929 18717 7941 18751
rect 7975 18717 7987 18751
rect 7929 18711 7987 18717
rect 8496 18720 9168 18748
rect 6730 18640 6736 18692
rect 6788 18680 6794 18692
rect 6788 18652 7328 18680
rect 6788 18640 6794 18652
rect 6457 18615 6515 18621
rect 6457 18581 6469 18615
rect 6503 18612 6515 18615
rect 6822 18612 6828 18624
rect 6503 18584 6828 18612
rect 6503 18581 6515 18584
rect 6457 18575 6515 18581
rect 6822 18572 6828 18584
rect 6880 18572 6886 18624
rect 7300 18612 7328 18652
rect 8496 18612 8524 18720
rect 9140 18680 9168 18720
rect 10870 18708 10876 18760
rect 10928 18748 10934 18760
rect 11425 18751 11483 18757
rect 11425 18748 11437 18751
rect 10928 18720 11437 18748
rect 10928 18708 10934 18720
rect 11425 18717 11437 18720
rect 11471 18748 11483 18751
rect 11974 18748 11980 18760
rect 11471 18720 11980 18748
rect 11471 18717 11483 18720
rect 11425 18711 11483 18717
rect 11974 18708 11980 18720
rect 12032 18748 12038 18760
rect 13648 18748 13676 18779
rect 13722 18776 13728 18788
rect 13780 18816 13786 18828
rect 14829 18819 14887 18825
rect 14829 18816 14841 18819
rect 13780 18788 14841 18816
rect 13780 18776 13786 18788
rect 14829 18785 14841 18788
rect 14875 18785 14887 18819
rect 14829 18779 14887 18785
rect 12032 18720 13676 18748
rect 14645 18751 14703 18757
rect 12032 18708 12038 18720
rect 14645 18717 14657 18751
rect 14691 18748 14703 18751
rect 15102 18748 15108 18760
rect 14691 18720 15108 18748
rect 14691 18717 14703 18720
rect 14645 18711 14703 18717
rect 15102 18708 15108 18720
rect 15160 18708 15166 18760
rect 16500 18748 16528 18915
rect 20346 18912 20352 18924
rect 20404 18912 20410 18964
rect 21358 18912 21364 18964
rect 21416 18952 21422 18964
rect 21910 18952 21916 18964
rect 21416 18924 21916 18952
rect 21416 18912 21422 18924
rect 21910 18912 21916 18924
rect 21968 18952 21974 18964
rect 24029 18955 24087 18961
rect 24029 18952 24041 18955
rect 21968 18924 24041 18952
rect 21968 18912 21974 18924
rect 24029 18921 24041 18924
rect 24075 18921 24087 18955
rect 24029 18915 24087 18921
rect 21085 18887 21143 18893
rect 21085 18853 21097 18887
rect 21131 18884 21143 18887
rect 22278 18884 22284 18896
rect 21131 18856 22284 18884
rect 21131 18853 21143 18856
rect 21085 18847 21143 18853
rect 22278 18844 22284 18856
rect 22336 18844 22342 18896
rect 16850 18776 16856 18828
rect 16908 18816 16914 18828
rect 17405 18819 17463 18825
rect 17405 18816 17417 18819
rect 16908 18788 17417 18816
rect 16908 18776 16914 18788
rect 17405 18785 17417 18788
rect 17451 18785 17463 18819
rect 17405 18779 17463 18785
rect 21542 18776 21548 18828
rect 21600 18776 21606 18828
rect 21637 18819 21695 18825
rect 21637 18785 21649 18819
rect 21683 18816 21695 18819
rect 22002 18816 22008 18828
rect 21683 18788 22008 18816
rect 21683 18785 21695 18788
rect 21637 18779 21695 18785
rect 22002 18776 22008 18788
rect 22060 18776 22066 18828
rect 22557 18819 22615 18825
rect 22557 18785 22569 18819
rect 22603 18816 22615 18819
rect 25225 18819 25283 18825
rect 25225 18816 25237 18819
rect 22603 18788 25237 18816
rect 22603 18785 22615 18788
rect 22557 18779 22615 18785
rect 25225 18785 25237 18788
rect 25271 18785 25283 18819
rect 25225 18779 25283 18785
rect 17221 18751 17279 18757
rect 17221 18748 17233 18751
rect 16500 18720 17233 18748
rect 17221 18717 17233 18720
rect 17267 18717 17279 18751
rect 17221 18711 17279 18717
rect 18598 18708 18604 18760
rect 18656 18748 18662 18760
rect 18693 18751 18751 18757
rect 18693 18748 18705 18751
rect 18656 18720 18705 18748
rect 18656 18708 18662 18720
rect 18693 18717 18705 18720
rect 18739 18748 18751 18751
rect 19337 18751 19395 18757
rect 19337 18748 19349 18751
rect 18739 18720 19349 18748
rect 18739 18717 18751 18720
rect 18693 18711 18751 18717
rect 19337 18717 19349 18720
rect 19383 18717 19395 18751
rect 19337 18711 19395 18717
rect 19797 18751 19855 18757
rect 19797 18717 19809 18751
rect 19843 18748 19855 18751
rect 20990 18748 20996 18760
rect 19843 18720 20996 18748
rect 19843 18717 19855 18720
rect 19797 18711 19855 18717
rect 20990 18708 20996 18720
rect 21048 18708 21054 18760
rect 21726 18708 21732 18760
rect 21784 18748 21790 18760
rect 22281 18751 22339 18757
rect 22281 18748 22293 18751
rect 21784 18720 22293 18748
rect 21784 18708 21790 18720
rect 22281 18717 22293 18720
rect 22327 18717 22339 18751
rect 22281 18711 22339 18717
rect 24578 18708 24584 18760
rect 24636 18708 24642 18760
rect 9401 18683 9459 18689
rect 9401 18680 9413 18683
rect 9140 18652 9413 18680
rect 9401 18649 9413 18652
rect 9447 18680 9459 18683
rect 12161 18683 12219 18689
rect 9447 18652 9812 18680
rect 10626 18652 11284 18680
rect 9447 18649 9459 18652
rect 9401 18643 9459 18649
rect 7300 18584 8524 18612
rect 8573 18615 8631 18621
rect 8573 18581 8585 18615
rect 8619 18612 8631 18615
rect 9674 18612 9680 18624
rect 8619 18584 9680 18612
rect 8619 18581 8631 18584
rect 8573 18575 8631 18581
rect 9674 18572 9680 18584
rect 9732 18572 9738 18624
rect 9784 18612 9812 18652
rect 11256 18624 11284 18652
rect 12161 18649 12173 18683
rect 12207 18680 12219 18683
rect 13998 18680 14004 18692
rect 12207 18652 14004 18680
rect 12207 18649 12219 18652
rect 12161 18643 12219 18649
rect 13998 18640 14004 18652
rect 14056 18640 14062 18692
rect 16022 18680 16028 18692
rect 14568 18652 16028 18680
rect 10134 18612 10140 18624
rect 9784 18584 10140 18612
rect 10134 18572 10140 18584
rect 10192 18572 10198 18624
rect 11238 18572 11244 18624
rect 11296 18572 11302 18624
rect 12253 18615 12311 18621
rect 12253 18581 12265 18615
rect 12299 18612 12311 18615
rect 12526 18612 12532 18624
rect 12299 18584 12532 18612
rect 12299 18581 12311 18584
rect 12253 18575 12311 18581
rect 12526 18572 12532 18584
rect 12584 18572 12590 18624
rect 13170 18572 13176 18624
rect 13228 18612 13234 18624
rect 13357 18615 13415 18621
rect 13357 18612 13369 18615
rect 13228 18584 13369 18612
rect 13228 18572 13234 18584
rect 13357 18581 13369 18584
rect 13403 18612 13415 18615
rect 14568 18612 14596 18652
rect 16022 18640 16028 18652
rect 16080 18640 16086 18692
rect 17313 18683 17371 18689
rect 17313 18649 17325 18683
rect 17359 18680 17371 18683
rect 17402 18680 17408 18692
rect 17359 18652 17408 18680
rect 17359 18649 17371 18652
rect 17313 18643 17371 18649
rect 17402 18640 17408 18652
rect 17460 18680 17466 18692
rect 17865 18683 17923 18689
rect 17865 18680 17877 18683
rect 17460 18652 17877 18680
rect 17460 18640 17466 18652
rect 17865 18649 17877 18652
rect 17911 18649 17923 18683
rect 17865 18643 17923 18649
rect 18877 18683 18935 18689
rect 18877 18649 18889 18683
rect 18923 18680 18935 18683
rect 18966 18680 18972 18692
rect 18923 18652 18972 18680
rect 18923 18649 18935 18652
rect 18877 18643 18935 18649
rect 18966 18640 18972 18652
rect 19024 18640 19030 18692
rect 19150 18640 19156 18692
rect 19208 18680 19214 18692
rect 21453 18683 21511 18689
rect 21453 18680 21465 18683
rect 19208 18652 21465 18680
rect 19208 18640 19214 18652
rect 21453 18649 21465 18652
rect 21499 18649 21511 18683
rect 21453 18643 21511 18649
rect 23566 18640 23572 18692
rect 23624 18640 23630 18692
rect 13403 18584 14596 18612
rect 13403 18581 13415 18584
rect 13357 18575 13415 18581
rect 14734 18572 14740 18624
rect 14792 18572 14798 18624
rect 15010 18572 15016 18624
rect 15068 18612 15074 18624
rect 17586 18612 17592 18624
rect 15068 18584 17592 18612
rect 15068 18572 15074 18584
rect 17586 18572 17592 18584
rect 17644 18612 17650 18624
rect 19518 18612 19524 18624
rect 17644 18584 19524 18612
rect 17644 18572 17650 18584
rect 19518 18572 19524 18584
rect 19576 18572 19582 18624
rect 19978 18572 19984 18624
rect 20036 18612 20042 18624
rect 20441 18615 20499 18621
rect 20441 18612 20453 18615
rect 20036 18584 20453 18612
rect 20036 18572 20042 18584
rect 20441 18581 20453 18584
rect 20487 18581 20499 18615
rect 20441 18575 20499 18581
rect 1104 18522 25852 18544
rect 1104 18470 7950 18522
rect 8002 18470 8014 18522
rect 8066 18470 8078 18522
rect 8130 18470 8142 18522
rect 8194 18470 8206 18522
rect 8258 18470 17950 18522
rect 18002 18470 18014 18522
rect 18066 18470 18078 18522
rect 18130 18470 18142 18522
rect 18194 18470 18206 18522
rect 18258 18470 25852 18522
rect 1104 18448 25852 18470
rect 4246 18368 4252 18420
rect 4304 18408 4310 18420
rect 5261 18411 5319 18417
rect 5261 18408 5273 18411
rect 4304 18380 5273 18408
rect 4304 18368 4310 18380
rect 5261 18377 5273 18380
rect 5307 18377 5319 18411
rect 5261 18371 5319 18377
rect 5629 18411 5687 18417
rect 5629 18377 5641 18411
rect 5675 18408 5687 18411
rect 7098 18408 7104 18420
rect 5675 18380 7104 18408
rect 5675 18377 5687 18380
rect 5629 18371 5687 18377
rect 7098 18368 7104 18380
rect 7156 18368 7162 18420
rect 9493 18411 9551 18417
rect 9493 18377 9505 18411
rect 9539 18408 9551 18411
rect 10042 18408 10048 18420
rect 9539 18380 10048 18408
rect 9539 18377 9551 18380
rect 9493 18371 9551 18377
rect 10042 18368 10048 18380
rect 10100 18368 10106 18420
rect 10318 18368 10324 18420
rect 10376 18408 10382 18420
rect 10413 18411 10471 18417
rect 10413 18408 10425 18411
rect 10376 18380 10425 18408
rect 10376 18368 10382 18380
rect 10413 18377 10425 18380
rect 10459 18377 10471 18411
rect 10413 18371 10471 18377
rect 10781 18411 10839 18417
rect 10781 18377 10793 18411
rect 10827 18408 10839 18411
rect 12805 18411 12863 18417
rect 12805 18408 12817 18411
rect 10827 18380 12817 18408
rect 10827 18377 10839 18380
rect 10781 18371 10839 18377
rect 12805 18377 12817 18380
rect 12851 18377 12863 18411
rect 12805 18371 12863 18377
rect 13170 18368 13176 18420
rect 13228 18368 13234 18420
rect 13265 18411 13323 18417
rect 13265 18377 13277 18411
rect 13311 18408 13323 18411
rect 13538 18408 13544 18420
rect 13311 18380 13544 18408
rect 13311 18377 13323 18380
rect 13265 18371 13323 18377
rect 6822 18300 6828 18352
rect 6880 18300 6886 18352
rect 6914 18300 6920 18352
rect 6972 18340 6978 18352
rect 8573 18343 8631 18349
rect 6972 18312 7314 18340
rect 6972 18300 6978 18312
rect 8573 18309 8585 18343
rect 8619 18340 8631 18343
rect 10226 18340 10232 18352
rect 8619 18312 10232 18340
rect 8619 18309 8631 18312
rect 8573 18303 8631 18309
rect 10226 18300 10232 18312
rect 10284 18300 10290 18352
rect 12342 18300 12348 18352
rect 12400 18340 12406 18352
rect 12529 18343 12587 18349
rect 12529 18340 12541 18343
rect 12400 18312 12541 18340
rect 12400 18300 12406 18312
rect 12529 18309 12541 18312
rect 12575 18340 12587 18343
rect 13280 18340 13308 18371
rect 13538 18368 13544 18380
rect 13596 18368 13602 18420
rect 13998 18368 14004 18420
rect 14056 18368 14062 18420
rect 14369 18411 14427 18417
rect 14369 18377 14381 18411
rect 14415 18408 14427 18411
rect 15105 18411 15163 18417
rect 15105 18408 15117 18411
rect 14415 18380 15117 18408
rect 14415 18377 14427 18380
rect 14369 18371 14427 18377
rect 15105 18377 15117 18380
rect 15151 18408 15163 18411
rect 18322 18408 18328 18420
rect 15151 18380 18328 18408
rect 15151 18377 15163 18380
rect 15105 18371 15163 18377
rect 18322 18368 18328 18380
rect 18380 18368 18386 18420
rect 19981 18411 20039 18417
rect 19981 18377 19993 18411
rect 20027 18408 20039 18411
rect 20714 18408 20720 18420
rect 20027 18380 20720 18408
rect 20027 18377 20039 18380
rect 19981 18371 20039 18377
rect 19996 18340 20024 18371
rect 20714 18368 20720 18380
rect 20772 18368 20778 18420
rect 12575 18312 13308 18340
rect 19366 18312 20024 18340
rect 20165 18343 20223 18349
rect 12575 18309 12587 18312
rect 12529 18303 12587 18309
rect 20165 18309 20177 18343
rect 20211 18340 20223 18343
rect 20441 18343 20499 18349
rect 20441 18340 20453 18343
rect 20211 18312 20453 18340
rect 20211 18309 20223 18312
rect 20165 18303 20223 18309
rect 20441 18309 20453 18312
rect 20487 18340 20499 18343
rect 20530 18340 20536 18352
rect 20487 18312 20536 18340
rect 20487 18309 20499 18312
rect 20441 18303 20499 18309
rect 20530 18300 20536 18312
rect 20588 18300 20594 18352
rect 9398 18232 9404 18284
rect 9456 18232 9462 18284
rect 10873 18275 10931 18281
rect 10873 18241 10885 18275
rect 10919 18272 10931 18275
rect 11974 18272 11980 18284
rect 10919 18244 11980 18272
rect 10919 18241 10931 18244
rect 10873 18235 10931 18241
rect 11974 18232 11980 18244
rect 12032 18232 12038 18284
rect 22281 18275 22339 18281
rect 22281 18241 22293 18275
rect 22327 18272 22339 18275
rect 23658 18272 23664 18284
rect 22327 18244 23664 18272
rect 22327 18241 22339 18244
rect 22281 18235 22339 18241
rect 23658 18232 23664 18244
rect 23716 18232 23722 18284
rect 24121 18275 24179 18281
rect 24121 18241 24133 18275
rect 24167 18272 24179 18275
rect 24394 18272 24400 18284
rect 24167 18244 24400 18272
rect 24167 18241 24179 18244
rect 24121 18235 24179 18241
rect 24394 18232 24400 18244
rect 24452 18232 24458 18284
rect 5721 18207 5779 18213
rect 5721 18173 5733 18207
rect 5767 18173 5779 18207
rect 5721 18167 5779 18173
rect 5905 18207 5963 18213
rect 5905 18173 5917 18207
rect 5951 18204 5963 18207
rect 6086 18204 6092 18216
rect 5951 18176 6092 18204
rect 5951 18173 5963 18176
rect 5905 18167 5963 18173
rect 5736 18068 5764 18167
rect 6086 18164 6092 18176
rect 6144 18164 6150 18216
rect 6546 18164 6552 18216
rect 6604 18164 6610 18216
rect 7374 18164 7380 18216
rect 7432 18204 7438 18216
rect 9030 18204 9036 18216
rect 7432 18176 9036 18204
rect 7432 18164 7438 18176
rect 9030 18164 9036 18176
rect 9088 18164 9094 18216
rect 9490 18164 9496 18216
rect 9548 18204 9554 18216
rect 9585 18207 9643 18213
rect 9585 18204 9597 18207
rect 9548 18176 9597 18204
rect 9548 18164 9554 18176
rect 9585 18173 9597 18176
rect 9631 18173 9643 18207
rect 9585 18167 9643 18173
rect 9600 18136 9628 18167
rect 9858 18164 9864 18216
rect 9916 18204 9922 18216
rect 10965 18207 11023 18213
rect 10965 18204 10977 18207
rect 9916 18176 10977 18204
rect 9916 18164 9922 18176
rect 10965 18173 10977 18176
rect 11011 18173 11023 18207
rect 10965 18167 11023 18173
rect 13446 18164 13452 18216
rect 13504 18164 13510 18216
rect 13814 18164 13820 18216
rect 13872 18204 13878 18216
rect 14461 18207 14519 18213
rect 14461 18204 14473 18207
rect 13872 18176 14473 18204
rect 13872 18164 13878 18176
rect 14461 18173 14473 18176
rect 14507 18173 14519 18207
rect 14461 18167 14519 18173
rect 14642 18164 14648 18216
rect 14700 18204 14706 18216
rect 15102 18204 15108 18216
rect 14700 18176 15108 18204
rect 14700 18164 14706 18176
rect 15102 18164 15108 18176
rect 15160 18164 15166 18216
rect 17865 18207 17923 18213
rect 17865 18173 17877 18207
rect 17911 18204 17923 18207
rect 17911 18176 18000 18204
rect 17911 18173 17923 18176
rect 17865 18167 17923 18173
rect 11606 18136 11612 18148
rect 9600 18108 11612 18136
rect 11606 18096 11612 18108
rect 11664 18096 11670 18148
rect 7466 18068 7472 18080
rect 5736 18040 7472 18068
rect 7466 18028 7472 18040
rect 7524 18028 7530 18080
rect 9030 18028 9036 18080
rect 9088 18028 9094 18080
rect 17972 18068 18000 18176
rect 18138 18164 18144 18216
rect 18196 18164 18202 18216
rect 21269 18207 21327 18213
rect 21269 18173 21281 18207
rect 21315 18204 21327 18207
rect 21726 18204 21732 18216
rect 21315 18176 21732 18204
rect 21315 18173 21327 18176
rect 21269 18167 21327 18173
rect 21726 18164 21732 18176
rect 21784 18164 21790 18216
rect 23293 18207 23351 18213
rect 23293 18173 23305 18207
rect 23339 18204 23351 18207
rect 23382 18204 23388 18216
rect 23339 18176 23388 18204
rect 23339 18173 23351 18176
rect 23293 18167 23351 18173
rect 23382 18164 23388 18176
rect 23440 18164 23446 18216
rect 24762 18164 24768 18216
rect 24820 18164 24826 18216
rect 19613 18139 19671 18145
rect 19613 18105 19625 18139
rect 19659 18136 19671 18139
rect 20990 18136 20996 18148
rect 19659 18108 20996 18136
rect 19659 18105 19671 18108
rect 19613 18099 19671 18105
rect 20990 18096 20996 18108
rect 21048 18096 21054 18148
rect 18690 18068 18696 18080
rect 17972 18040 18696 18068
rect 18690 18028 18696 18040
rect 18748 18028 18754 18080
rect 1104 17978 25852 18000
rect 1104 17926 2950 17978
rect 3002 17926 3014 17978
rect 3066 17926 3078 17978
rect 3130 17926 3142 17978
rect 3194 17926 3206 17978
rect 3258 17926 12950 17978
rect 13002 17926 13014 17978
rect 13066 17926 13078 17978
rect 13130 17926 13142 17978
rect 13194 17926 13206 17978
rect 13258 17926 22950 17978
rect 23002 17926 23014 17978
rect 23066 17926 23078 17978
rect 23130 17926 23142 17978
rect 23194 17926 23206 17978
rect 23258 17926 25852 17978
rect 1104 17904 25852 17926
rect 5534 17824 5540 17876
rect 5592 17864 5598 17876
rect 5810 17864 5816 17876
rect 5592 17836 5816 17864
rect 5592 17824 5598 17836
rect 5810 17824 5816 17836
rect 5868 17824 5874 17876
rect 6086 17824 6092 17876
rect 6144 17864 6150 17876
rect 6549 17867 6607 17873
rect 6549 17864 6561 17867
rect 6144 17836 6561 17864
rect 6144 17824 6150 17836
rect 6549 17833 6561 17836
rect 6595 17833 6607 17867
rect 6549 17827 6607 17833
rect 7098 17824 7104 17876
rect 7156 17824 7162 17876
rect 10413 17867 10471 17873
rect 10413 17833 10425 17867
rect 10459 17864 10471 17867
rect 11514 17864 11520 17876
rect 10459 17836 11520 17864
rect 10459 17833 10471 17836
rect 10413 17827 10471 17833
rect 7558 17688 7564 17740
rect 7616 17688 7622 17740
rect 7742 17688 7748 17740
rect 7800 17688 7806 17740
rect 8389 17731 8447 17737
rect 8389 17697 8401 17731
rect 8435 17728 8447 17731
rect 9398 17728 9404 17740
rect 8435 17700 9404 17728
rect 8435 17697 8447 17700
rect 8389 17691 8447 17697
rect 9398 17688 9404 17700
rect 9456 17688 9462 17740
rect 4798 17620 4804 17672
rect 4856 17620 4862 17672
rect 7469 17663 7527 17669
rect 7469 17629 7481 17663
rect 7515 17660 7527 17663
rect 9030 17660 9036 17672
rect 7515 17632 9036 17660
rect 7515 17629 7527 17632
rect 7469 17623 7527 17629
rect 9030 17620 9036 17632
rect 9088 17620 9094 17672
rect 9125 17663 9183 17669
rect 9125 17629 9137 17663
rect 9171 17660 9183 17663
rect 10428 17660 10456 17827
rect 11514 17824 11520 17836
rect 11572 17824 11578 17876
rect 17497 17867 17555 17873
rect 17497 17833 17509 17867
rect 17543 17864 17555 17867
rect 18138 17864 18144 17876
rect 17543 17836 18144 17864
rect 17543 17833 17555 17836
rect 17497 17827 17555 17833
rect 18138 17824 18144 17836
rect 18196 17824 18202 17876
rect 19337 17867 19395 17873
rect 19337 17833 19349 17867
rect 19383 17864 19395 17867
rect 20530 17864 20536 17876
rect 19383 17836 20536 17864
rect 19383 17833 19395 17836
rect 19337 17827 19395 17833
rect 11054 17688 11060 17740
rect 11112 17688 11118 17740
rect 11333 17731 11391 17737
rect 11333 17697 11345 17731
rect 11379 17728 11391 17731
rect 13630 17728 13636 17740
rect 11379 17700 13636 17728
rect 11379 17697 11391 17700
rect 11333 17691 11391 17697
rect 13630 17688 13636 17700
rect 13688 17688 13694 17740
rect 9171 17632 10456 17660
rect 9171 17629 9183 17632
rect 9125 17623 9183 17629
rect 14918 17620 14924 17672
rect 14976 17660 14982 17672
rect 15565 17663 15623 17669
rect 15565 17660 15577 17663
rect 14976 17632 15577 17660
rect 14976 17620 14982 17632
rect 15565 17629 15577 17632
rect 15611 17629 15623 17663
rect 15565 17623 15623 17629
rect 16209 17663 16267 17669
rect 16209 17629 16221 17663
rect 16255 17660 16267 17663
rect 16758 17660 16764 17672
rect 16255 17632 16764 17660
rect 16255 17629 16267 17632
rect 16209 17623 16267 17629
rect 16758 17620 16764 17632
rect 16816 17620 16822 17672
rect 16850 17620 16856 17672
rect 16908 17620 16914 17672
rect 17957 17663 18015 17669
rect 17957 17629 17969 17663
rect 18003 17660 18015 17663
rect 19352 17660 19380 17827
rect 20530 17824 20536 17836
rect 20588 17824 20594 17876
rect 21450 17824 21456 17876
rect 21508 17824 21514 17876
rect 23658 17824 23664 17876
rect 23716 17864 23722 17876
rect 24578 17864 24584 17876
rect 23716 17836 24584 17864
rect 23716 17824 23722 17836
rect 24578 17824 24584 17836
rect 24636 17824 24642 17876
rect 23566 17796 23572 17808
rect 23308 17768 23572 17796
rect 19702 17688 19708 17740
rect 19760 17728 19766 17740
rect 19760 17700 21772 17728
rect 19760 17688 19766 17700
rect 21744 17672 21772 17700
rect 22186 17688 22192 17740
rect 22244 17688 22250 17740
rect 18003 17632 19380 17660
rect 18003 17629 18015 17632
rect 17957 17623 18015 17629
rect 21726 17620 21732 17672
rect 21784 17660 21790 17672
rect 21913 17663 21971 17669
rect 21913 17660 21925 17663
rect 21784 17632 21925 17660
rect 21784 17620 21790 17632
rect 21913 17629 21925 17632
rect 21959 17629 21971 17663
rect 23308 17646 23336 17768
rect 23566 17756 23572 17768
rect 23624 17796 23630 17808
rect 23937 17799 23995 17805
rect 23937 17796 23949 17799
rect 23624 17768 23949 17796
rect 23624 17756 23630 17768
rect 23937 17765 23949 17768
rect 23983 17765 23995 17799
rect 23937 17759 23995 17765
rect 21913 17623 21971 17629
rect 5074 17552 5080 17604
rect 5132 17552 5138 17604
rect 6914 17592 6920 17604
rect 6302 17564 6920 17592
rect 6914 17552 6920 17564
rect 6972 17552 6978 17604
rect 9858 17552 9864 17604
rect 9916 17552 9922 17604
rect 9968 17564 10640 17592
rect 12558 17564 13216 17592
rect 9306 17484 9312 17536
rect 9364 17524 9370 17536
rect 9968 17524 9996 17564
rect 9364 17496 9996 17524
rect 9364 17484 9370 17496
rect 10502 17484 10508 17536
rect 10560 17484 10566 17536
rect 10612 17524 10640 17564
rect 13188 17533 13216 17564
rect 18690 17552 18696 17604
rect 18748 17552 18754 17604
rect 19978 17552 19984 17604
rect 20036 17552 20042 17604
rect 20714 17552 20720 17604
rect 20772 17552 20778 17604
rect 12805 17527 12863 17533
rect 12805 17524 12817 17527
rect 10612 17496 12817 17524
rect 12805 17493 12817 17496
rect 12851 17493 12863 17527
rect 12805 17487 12863 17493
rect 13173 17527 13231 17533
rect 13173 17493 13185 17527
rect 13219 17524 13231 17527
rect 13630 17524 13636 17536
rect 13219 17496 13636 17524
rect 13219 17493 13231 17496
rect 13173 17487 13231 17493
rect 13630 17484 13636 17496
rect 13688 17484 13694 17536
rect 13814 17484 13820 17536
rect 13872 17484 13878 17536
rect 15381 17527 15439 17533
rect 15381 17493 15393 17527
rect 15427 17524 15439 17527
rect 15470 17524 15476 17536
rect 15427 17496 15476 17524
rect 15427 17493 15439 17496
rect 15381 17487 15439 17493
rect 15470 17484 15476 17496
rect 15528 17484 15534 17536
rect 15562 17484 15568 17536
rect 15620 17524 15626 17536
rect 16301 17527 16359 17533
rect 16301 17524 16313 17527
rect 15620 17496 16313 17524
rect 15620 17484 15626 17496
rect 16301 17493 16313 17496
rect 16347 17493 16359 17527
rect 16301 17487 16359 17493
rect 1104 17434 25852 17456
rect 1104 17382 7950 17434
rect 8002 17382 8014 17434
rect 8066 17382 8078 17434
rect 8130 17382 8142 17434
rect 8194 17382 8206 17434
rect 8258 17382 17950 17434
rect 18002 17382 18014 17434
rect 18066 17382 18078 17434
rect 18130 17382 18142 17434
rect 18194 17382 18206 17434
rect 18258 17382 25852 17434
rect 1104 17360 25852 17382
rect 5074 17280 5080 17332
rect 5132 17320 5138 17332
rect 5997 17323 6055 17329
rect 5997 17320 6009 17323
rect 5132 17292 6009 17320
rect 5132 17280 5138 17292
rect 5997 17289 6009 17292
rect 6043 17289 6055 17323
rect 5997 17283 6055 17289
rect 6733 17323 6791 17329
rect 6733 17289 6745 17323
rect 6779 17320 6791 17323
rect 6914 17320 6920 17332
rect 6779 17292 6920 17320
rect 6779 17289 6791 17292
rect 6733 17283 6791 17289
rect 6914 17280 6920 17292
rect 6972 17280 6978 17332
rect 7466 17280 7472 17332
rect 7524 17280 7530 17332
rect 7837 17323 7895 17329
rect 7837 17289 7849 17323
rect 7883 17320 7895 17323
rect 7883 17292 9168 17320
rect 7883 17289 7895 17292
rect 7837 17283 7895 17289
rect 2225 17255 2283 17261
rect 2225 17221 2237 17255
rect 2271 17252 2283 17255
rect 2314 17252 2320 17264
rect 2271 17224 2320 17252
rect 2271 17221 2283 17224
rect 2225 17215 2283 17221
rect 2314 17212 2320 17224
rect 2372 17212 2378 17264
rect 7742 17252 7748 17264
rect 6886 17224 7748 17252
rect 5353 17187 5411 17193
rect 5353 17153 5365 17187
rect 5399 17184 5411 17187
rect 6886 17184 6914 17224
rect 7742 17212 7748 17224
rect 7800 17252 7806 17264
rect 9140 17252 9168 17292
rect 9214 17280 9220 17332
rect 9272 17320 9278 17332
rect 9861 17323 9919 17329
rect 9861 17320 9873 17323
rect 9272 17292 9873 17320
rect 9272 17280 9278 17292
rect 9861 17289 9873 17292
rect 9907 17289 9919 17323
rect 9861 17283 9919 17289
rect 10134 17280 10140 17332
rect 10192 17320 10198 17332
rect 10321 17323 10379 17329
rect 10321 17320 10333 17323
rect 10192 17292 10333 17320
rect 10192 17280 10198 17292
rect 10321 17289 10333 17292
rect 10367 17320 10379 17323
rect 10502 17320 10508 17332
rect 10367 17292 10508 17320
rect 10367 17289 10379 17292
rect 10321 17283 10379 17289
rect 10502 17280 10508 17292
rect 10560 17280 10566 17332
rect 11698 17320 11704 17332
rect 10612 17292 11704 17320
rect 10612 17252 10640 17292
rect 11698 17280 11704 17292
rect 11756 17280 11762 17332
rect 12066 17280 12072 17332
rect 12124 17320 12130 17332
rect 13081 17323 13139 17329
rect 13081 17320 13093 17323
rect 12124 17292 13093 17320
rect 12124 17280 12130 17292
rect 13081 17289 13093 17292
rect 13127 17289 13139 17323
rect 13081 17283 13139 17289
rect 15378 17280 15384 17332
rect 15436 17320 15442 17332
rect 15654 17320 15660 17332
rect 15436 17292 15660 17320
rect 15436 17280 15442 17292
rect 15654 17280 15660 17292
rect 15712 17280 15718 17332
rect 16025 17323 16083 17329
rect 16025 17289 16037 17323
rect 16071 17320 16083 17323
rect 16298 17320 16304 17332
rect 16071 17292 16304 17320
rect 16071 17289 16083 17292
rect 16025 17283 16083 17289
rect 16298 17280 16304 17292
rect 16356 17280 16362 17332
rect 19702 17320 19708 17332
rect 16960 17292 19708 17320
rect 7800 17224 7972 17252
rect 9140 17224 10640 17252
rect 7800 17212 7806 17224
rect 5399 17156 6914 17184
rect 7944 17184 7972 17224
rect 11054 17212 11060 17264
rect 11112 17252 11118 17264
rect 11790 17252 11796 17264
rect 11112 17224 11796 17252
rect 11112 17212 11118 17224
rect 11790 17212 11796 17224
rect 11848 17252 11854 17264
rect 12437 17255 12495 17261
rect 12437 17252 12449 17255
rect 11848 17224 12449 17252
rect 11848 17212 11854 17224
rect 12437 17221 12449 17224
rect 12483 17221 12495 17255
rect 12437 17215 12495 17221
rect 13449 17255 13507 17261
rect 13449 17221 13461 17255
rect 13495 17252 13507 17255
rect 15746 17252 15752 17264
rect 13495 17224 15752 17252
rect 13495 17221 13507 17224
rect 13449 17215 13507 17221
rect 15746 17212 15752 17224
rect 15804 17212 15810 17264
rect 16960 17252 16988 17292
rect 19702 17280 19708 17292
rect 19760 17280 19766 17332
rect 20622 17280 20628 17332
rect 20680 17320 20686 17332
rect 21269 17323 21327 17329
rect 21269 17320 21281 17323
rect 20680 17292 21281 17320
rect 20680 17280 20686 17292
rect 21269 17289 21281 17292
rect 21315 17289 21327 17323
rect 21269 17283 21327 17289
rect 16868 17224 16988 17252
rect 19521 17255 19579 17261
rect 9033 17187 9091 17193
rect 9033 17184 9045 17187
rect 7944 17156 8064 17184
rect 5399 17153 5411 17156
rect 5353 17147 5411 17153
rect 8036 17125 8064 17156
rect 8496 17156 9045 17184
rect 7929 17119 7987 17125
rect 7929 17116 7941 17119
rect 7852 17088 7941 17116
rect 7852 17060 7880 17088
rect 7929 17085 7941 17088
rect 7975 17085 7987 17119
rect 7929 17079 7987 17085
rect 8021 17119 8079 17125
rect 8021 17085 8033 17119
rect 8067 17085 8079 17119
rect 8021 17079 8079 17085
rect 5810 17008 5816 17060
rect 5868 17048 5874 17060
rect 5868 17020 6914 17048
rect 5868 17008 5874 17020
rect 1762 16940 1768 16992
rect 1820 16980 1826 16992
rect 2317 16983 2375 16989
rect 2317 16980 2329 16983
rect 1820 16952 2329 16980
rect 1820 16940 1826 16952
rect 2317 16949 2329 16952
rect 2363 16949 2375 16983
rect 2317 16943 2375 16949
rect 5902 16940 5908 16992
rect 5960 16980 5966 16992
rect 6546 16980 6552 16992
rect 5960 16952 6552 16980
rect 5960 16940 5966 16952
rect 6546 16940 6552 16952
rect 6604 16940 6610 16992
rect 6886 16980 6914 17020
rect 7834 17008 7840 17060
rect 7892 17008 7898 17060
rect 8496 16992 8524 17156
rect 9033 17153 9045 17156
rect 9079 17153 9091 17187
rect 9033 17147 9091 17153
rect 9122 17144 9128 17196
rect 9180 17144 9186 17196
rect 10229 17187 10287 17193
rect 10229 17153 10241 17187
rect 10275 17184 10287 17187
rect 10275 17156 10732 17184
rect 10275 17153 10287 17156
rect 10229 17147 10287 17153
rect 9306 17076 9312 17128
rect 9364 17076 9370 17128
rect 10318 17076 10324 17128
rect 10376 17116 10382 17128
rect 10413 17119 10471 17125
rect 10413 17116 10425 17119
rect 10376 17088 10425 17116
rect 10376 17076 10382 17088
rect 10413 17085 10425 17088
rect 10459 17085 10471 17119
rect 10413 17079 10471 17085
rect 8665 17051 8723 17057
rect 8665 17017 8677 17051
rect 8711 17048 8723 17051
rect 10502 17048 10508 17060
rect 8711 17020 10508 17048
rect 8711 17017 8723 17020
rect 8665 17011 8723 17017
rect 10502 17008 10508 17020
rect 10560 17008 10566 17060
rect 10704 17048 10732 17156
rect 11514 17144 11520 17196
rect 11572 17184 11578 17196
rect 11701 17187 11759 17193
rect 11701 17184 11713 17187
rect 11572 17156 11713 17184
rect 11572 17144 11578 17156
rect 11701 17153 11713 17156
rect 11747 17153 11759 17187
rect 14090 17184 14096 17196
rect 11701 17147 11759 17153
rect 12728 17156 14096 17184
rect 10778 17076 10784 17128
rect 10836 17116 10842 17128
rect 12728 17116 12756 17156
rect 10836 17088 12756 17116
rect 10836 17076 10842 17088
rect 12802 17076 12808 17128
rect 12860 17116 12866 17128
rect 13648 17125 13676 17156
rect 14090 17144 14096 17156
rect 14148 17144 14154 17196
rect 16868 17193 16896 17224
rect 19521 17221 19533 17255
rect 19567 17252 19579 17255
rect 19610 17252 19616 17264
rect 19567 17224 19616 17252
rect 19567 17221 19579 17224
rect 19521 17215 19579 17221
rect 19610 17212 19616 17224
rect 19668 17252 19674 17264
rect 20073 17255 20131 17261
rect 20073 17252 20085 17255
rect 19668 17224 20085 17252
rect 19668 17212 19674 17224
rect 20073 17221 20085 17224
rect 20119 17221 20131 17255
rect 20073 17215 20131 17221
rect 20714 17212 20720 17264
rect 20772 17252 20778 17264
rect 21545 17255 21603 17261
rect 21545 17252 21557 17255
rect 20772 17224 21557 17252
rect 20772 17212 20778 17224
rect 21545 17221 21557 17224
rect 21591 17252 21603 17255
rect 22186 17252 22192 17264
rect 21591 17224 22192 17252
rect 21591 17221 21603 17224
rect 21545 17215 21603 17221
rect 22186 17212 22192 17224
rect 22244 17212 22250 17264
rect 22830 17212 22836 17264
rect 22888 17252 22894 17264
rect 23201 17255 23259 17261
rect 23201 17252 23213 17255
rect 22888 17224 23213 17252
rect 22888 17212 22894 17224
rect 23201 17221 23213 17224
rect 23247 17221 23259 17255
rect 23201 17215 23259 17221
rect 15933 17187 15991 17193
rect 15933 17184 15945 17187
rect 15212 17156 15945 17184
rect 13541 17119 13599 17125
rect 13541 17116 13553 17119
rect 12860 17088 13553 17116
rect 12860 17076 12866 17088
rect 13541 17085 13553 17088
rect 13587 17085 13599 17119
rect 13541 17079 13599 17085
rect 13633 17119 13691 17125
rect 13633 17085 13645 17119
rect 13679 17116 13691 17119
rect 13679 17088 13713 17116
rect 13679 17085 13691 17088
rect 13633 17079 13691 17085
rect 10965 17051 11023 17057
rect 10965 17048 10977 17051
rect 10704 17020 10977 17048
rect 10965 17017 10977 17020
rect 11011 17048 11023 17051
rect 14274 17048 14280 17060
rect 11011 17020 12434 17048
rect 11011 17017 11023 17020
rect 10965 17011 11023 17017
rect 8478 16980 8484 16992
rect 6886 16952 8484 16980
rect 8478 16940 8484 16952
rect 8536 16940 8542 16992
rect 12406 16980 12434 17020
rect 13740 17020 14280 17048
rect 13740 16980 13768 17020
rect 14274 17008 14280 17020
rect 14332 17048 14338 17060
rect 14458 17048 14464 17060
rect 14332 17020 14464 17048
rect 14332 17008 14338 17020
rect 14458 17008 14464 17020
rect 14516 17008 14522 17060
rect 12406 16952 13768 16980
rect 13814 16940 13820 16992
rect 13872 16980 13878 16992
rect 15212 16989 15240 17156
rect 15933 17153 15945 17156
rect 15979 17153 15991 17187
rect 15933 17147 15991 17153
rect 16853 17187 16911 17193
rect 16853 17153 16865 17187
rect 16899 17153 16911 17187
rect 16853 17147 16911 17153
rect 18230 17144 18236 17196
rect 18288 17144 18294 17196
rect 19426 17144 19432 17196
rect 19484 17144 19490 17196
rect 20622 17144 20628 17196
rect 20680 17144 20686 17196
rect 22002 17144 22008 17196
rect 22060 17144 22066 17196
rect 23934 17144 23940 17196
rect 23992 17144 23998 17196
rect 15654 17076 15660 17128
rect 15712 17116 15718 17128
rect 16117 17119 16175 17125
rect 16117 17116 16129 17119
rect 15712 17088 16129 17116
rect 15712 17076 15718 17088
rect 16117 17085 16129 17088
rect 16163 17085 16175 17119
rect 16117 17079 16175 17085
rect 17129 17119 17187 17125
rect 17129 17085 17141 17119
rect 17175 17116 17187 17119
rect 18598 17116 18604 17128
rect 17175 17088 18604 17116
rect 17175 17085 17187 17088
rect 17129 17079 17187 17085
rect 18598 17076 18604 17088
rect 18656 17076 18662 17128
rect 19705 17119 19763 17125
rect 19705 17085 19717 17119
rect 19751 17116 19763 17119
rect 21450 17116 21456 17128
rect 19751 17088 21456 17116
rect 19751 17085 19763 17088
rect 19705 17079 19763 17085
rect 21450 17076 21456 17088
rect 21508 17076 21514 17128
rect 24670 17076 24676 17128
rect 24728 17076 24734 17128
rect 23382 17008 23388 17060
rect 23440 17008 23446 17060
rect 15197 16983 15255 16989
rect 15197 16980 15209 16983
rect 13872 16952 15209 16980
rect 13872 16940 13878 16952
rect 15197 16949 15209 16952
rect 15243 16949 15255 16983
rect 15197 16943 15255 16949
rect 15565 16983 15623 16989
rect 15565 16949 15577 16983
rect 15611 16980 15623 16983
rect 16482 16980 16488 16992
rect 15611 16952 16488 16980
rect 15611 16949 15623 16952
rect 15565 16943 15623 16949
rect 16482 16940 16488 16952
rect 16540 16940 16546 16992
rect 16850 16940 16856 16992
rect 16908 16980 16914 16992
rect 18601 16983 18659 16989
rect 18601 16980 18613 16983
rect 16908 16952 18613 16980
rect 16908 16940 16914 16952
rect 18601 16949 18613 16952
rect 18647 16949 18659 16983
rect 18601 16943 18659 16949
rect 19061 16983 19119 16989
rect 19061 16949 19073 16983
rect 19107 16980 19119 16983
rect 20438 16980 20444 16992
rect 19107 16952 20444 16980
rect 19107 16949 19119 16952
rect 19061 16943 19119 16949
rect 20438 16940 20444 16952
rect 20496 16940 20502 16992
rect 22002 16940 22008 16992
rect 22060 16980 22066 16992
rect 22649 16983 22707 16989
rect 22649 16980 22661 16983
rect 22060 16952 22661 16980
rect 22060 16940 22066 16952
rect 22649 16949 22661 16952
rect 22695 16949 22707 16983
rect 22649 16943 22707 16949
rect 1104 16890 25852 16912
rect 1104 16838 2950 16890
rect 3002 16838 3014 16890
rect 3066 16838 3078 16890
rect 3130 16838 3142 16890
rect 3194 16838 3206 16890
rect 3258 16838 12950 16890
rect 13002 16838 13014 16890
rect 13066 16838 13078 16890
rect 13130 16838 13142 16890
rect 13194 16838 13206 16890
rect 13258 16838 22950 16890
rect 23002 16838 23014 16890
rect 23066 16838 23078 16890
rect 23130 16838 23142 16890
rect 23194 16838 23206 16890
rect 23258 16838 25852 16890
rect 1104 16816 25852 16838
rect 6260 16779 6318 16785
rect 6260 16745 6272 16779
rect 6306 16776 6318 16779
rect 7926 16776 7932 16788
rect 6306 16748 7932 16776
rect 6306 16745 6318 16748
rect 6260 16739 6318 16745
rect 7926 16736 7932 16748
rect 7984 16736 7990 16788
rect 8478 16736 8484 16788
rect 8536 16736 8542 16788
rect 11514 16736 11520 16788
rect 11572 16776 11578 16788
rect 12713 16779 12771 16785
rect 12713 16776 12725 16779
rect 11572 16748 12725 16776
rect 11572 16736 11578 16748
rect 12713 16745 12725 16748
rect 12759 16745 12771 16779
rect 12713 16739 12771 16745
rect 12802 16736 12808 16788
rect 12860 16776 12866 16788
rect 12897 16779 12955 16785
rect 12897 16776 12909 16779
rect 12860 16748 12909 16776
rect 12860 16736 12866 16748
rect 12897 16745 12909 16748
rect 12943 16745 12955 16779
rect 12897 16739 12955 16745
rect 16298 16736 16304 16788
rect 16356 16776 16362 16788
rect 16393 16779 16451 16785
rect 16393 16776 16405 16779
rect 16356 16748 16405 16776
rect 16356 16736 16362 16748
rect 16393 16745 16405 16748
rect 16439 16745 16451 16779
rect 16393 16739 16451 16745
rect 19337 16779 19395 16785
rect 19337 16745 19349 16779
rect 19383 16776 19395 16779
rect 19426 16776 19432 16788
rect 19383 16748 19432 16776
rect 19383 16745 19395 16748
rect 19337 16739 19395 16745
rect 19426 16736 19432 16748
rect 19484 16736 19490 16788
rect 21177 16779 21235 16785
rect 21177 16745 21189 16779
rect 21223 16776 21235 16779
rect 23842 16776 23848 16788
rect 21223 16748 23848 16776
rect 21223 16745 21235 16748
rect 21177 16739 21235 16745
rect 23842 16736 23848 16748
rect 23900 16736 23906 16788
rect 9858 16708 9864 16720
rect 7668 16680 9864 16708
rect 4798 16600 4804 16652
rect 4856 16640 4862 16652
rect 5902 16640 5908 16652
rect 4856 16612 5908 16640
rect 4856 16600 4862 16612
rect 5902 16600 5908 16612
rect 5960 16640 5966 16652
rect 5997 16643 6055 16649
rect 5997 16640 6009 16643
rect 5960 16612 6009 16640
rect 5960 16600 5966 16612
rect 5997 16609 6009 16612
rect 6043 16609 6055 16643
rect 5997 16603 6055 16609
rect 6638 16600 6644 16652
rect 6696 16640 6702 16652
rect 7668 16640 7696 16680
rect 9858 16668 9864 16680
rect 9916 16668 9922 16720
rect 15194 16708 15200 16720
rect 13924 16680 15200 16708
rect 6696 16612 7696 16640
rect 6696 16600 6702 16612
rect 7742 16600 7748 16652
rect 7800 16600 7806 16652
rect 8938 16600 8944 16652
rect 8996 16640 9002 16652
rect 9582 16640 9588 16652
rect 8996 16612 9588 16640
rect 8996 16600 9002 16612
rect 9582 16600 9588 16612
rect 9640 16600 9646 16652
rect 9769 16643 9827 16649
rect 9769 16609 9781 16643
rect 9815 16640 9827 16643
rect 9950 16640 9956 16652
rect 9815 16612 9956 16640
rect 9815 16609 9827 16612
rect 9769 16603 9827 16609
rect 9950 16600 9956 16612
rect 10008 16640 10014 16652
rect 10873 16643 10931 16649
rect 10873 16640 10885 16643
rect 10008 16612 10885 16640
rect 10008 16600 10014 16612
rect 10873 16609 10885 16612
rect 10919 16609 10931 16643
rect 13924 16640 13952 16680
rect 15194 16668 15200 16680
rect 15252 16668 15258 16720
rect 18782 16708 18788 16720
rect 15580 16680 18788 16708
rect 10873 16603 10931 16609
rect 12406 16612 13952 16640
rect 14829 16643 14887 16649
rect 1765 16575 1823 16581
rect 1765 16541 1777 16575
rect 1811 16572 1823 16575
rect 2222 16572 2228 16584
rect 1811 16544 2228 16572
rect 1811 16541 1823 16544
rect 1765 16535 1823 16541
rect 2222 16532 2228 16544
rect 2280 16532 2286 16584
rect 9214 16532 9220 16584
rect 9272 16572 9278 16584
rect 9493 16575 9551 16581
rect 9493 16572 9505 16575
rect 9272 16544 9505 16572
rect 9272 16532 9278 16544
rect 9493 16541 9505 16544
rect 9539 16541 9551 16575
rect 9493 16535 9551 16541
rect 10686 16532 10692 16584
rect 10744 16532 10750 16584
rect 11514 16532 11520 16584
rect 11572 16532 11578 16584
rect 12066 16532 12072 16584
rect 12124 16572 12130 16584
rect 12406 16572 12434 16612
rect 14829 16609 14841 16643
rect 14875 16640 14887 16643
rect 14918 16640 14924 16652
rect 14875 16612 14924 16640
rect 14875 16609 14887 16612
rect 14829 16603 14887 16609
rect 14918 16600 14924 16612
rect 14976 16640 14982 16652
rect 15580 16649 15608 16680
rect 18782 16668 18788 16680
rect 18840 16668 18846 16720
rect 15565 16643 15623 16649
rect 15565 16640 15577 16643
rect 14976 16612 15577 16640
rect 14976 16600 14982 16612
rect 15565 16609 15577 16612
rect 15611 16609 15623 16643
rect 15565 16603 15623 16609
rect 15657 16643 15715 16649
rect 15657 16609 15669 16643
rect 15703 16609 15715 16643
rect 15657 16603 15715 16609
rect 12124 16544 12434 16572
rect 12124 16532 12130 16544
rect 15194 16532 15200 16584
rect 15252 16572 15258 16584
rect 15672 16572 15700 16603
rect 15746 16600 15752 16652
rect 15804 16640 15810 16652
rect 17586 16640 17592 16652
rect 15804 16612 17592 16640
rect 15804 16600 15810 16612
rect 17586 16600 17592 16612
rect 17644 16600 17650 16652
rect 18230 16640 18236 16652
rect 17880 16612 18236 16640
rect 16022 16572 16028 16584
rect 15252 16544 16028 16572
rect 15252 16532 15258 16544
rect 16022 16532 16028 16544
rect 16080 16532 16086 16584
rect 17770 16532 17776 16584
rect 17828 16572 17834 16584
rect 17880 16572 17908 16612
rect 18230 16600 18236 16612
rect 18288 16640 18294 16652
rect 18877 16643 18935 16649
rect 18877 16640 18889 16643
rect 18288 16612 18889 16640
rect 18288 16600 18294 16612
rect 18877 16609 18889 16612
rect 18923 16609 18935 16643
rect 18877 16603 18935 16609
rect 20533 16643 20591 16649
rect 20533 16609 20545 16643
rect 20579 16640 20591 16643
rect 20806 16640 20812 16652
rect 20579 16612 20812 16640
rect 20579 16609 20591 16612
rect 20533 16603 20591 16609
rect 20806 16600 20812 16612
rect 20864 16600 20870 16652
rect 20898 16600 20904 16652
rect 20956 16640 20962 16652
rect 21726 16640 21732 16652
rect 20956 16612 21732 16640
rect 20956 16600 20962 16612
rect 21726 16600 21732 16612
rect 21784 16600 21790 16652
rect 22002 16600 22008 16652
rect 22060 16600 22066 16652
rect 22462 16600 22468 16652
rect 22520 16640 22526 16652
rect 23753 16643 23811 16649
rect 23753 16640 23765 16643
rect 22520 16612 23765 16640
rect 22520 16600 22526 16612
rect 23753 16609 23765 16612
rect 23799 16609 23811 16643
rect 23753 16603 23811 16609
rect 17828 16544 17908 16572
rect 17957 16575 18015 16581
rect 17828 16532 17834 16544
rect 17957 16541 17969 16575
rect 18003 16572 18015 16575
rect 18322 16572 18328 16584
rect 18003 16544 18328 16572
rect 18003 16541 18015 16544
rect 17957 16535 18015 16541
rect 18322 16532 18328 16544
rect 18380 16532 18386 16584
rect 18598 16532 18604 16584
rect 18656 16532 18662 16584
rect 20254 16532 20260 16584
rect 20312 16572 20318 16584
rect 20349 16575 20407 16581
rect 20349 16572 20361 16575
rect 20312 16544 20361 16572
rect 20312 16532 20318 16544
rect 20349 16541 20361 16544
rect 20395 16541 20407 16575
rect 20349 16535 20407 16541
rect 1302 16464 1308 16516
rect 1360 16504 1366 16516
rect 2501 16507 2559 16513
rect 2501 16504 2513 16507
rect 1360 16476 2513 16504
rect 1360 16464 1366 16476
rect 2501 16473 2513 16476
rect 2547 16473 2559 16507
rect 7498 16476 7880 16504
rect 2501 16467 2559 16473
rect 6914 16396 6920 16448
rect 6972 16436 6978 16448
rect 7576 16436 7604 16476
rect 6972 16408 7604 16436
rect 7852 16436 7880 16476
rect 7926 16464 7932 16516
rect 7984 16504 7990 16516
rect 12161 16507 12219 16513
rect 12161 16504 12173 16507
rect 7984 16476 12173 16504
rect 7984 16464 7990 16476
rect 12161 16473 12173 16476
rect 12207 16473 12219 16507
rect 12161 16467 12219 16473
rect 14550 16464 14556 16516
rect 14608 16504 14614 16516
rect 19886 16504 19892 16516
rect 14608 16476 19892 16504
rect 14608 16464 14614 16476
rect 19886 16464 19892 16476
rect 19944 16464 19950 16516
rect 21082 16464 21088 16516
rect 21140 16464 21146 16516
rect 22646 16464 22652 16516
rect 22704 16464 22710 16516
rect 8113 16439 8171 16445
rect 8113 16436 8125 16439
rect 7852 16408 8125 16436
rect 6972 16396 6978 16408
rect 8113 16405 8125 16408
rect 8159 16436 8171 16439
rect 8478 16436 8484 16448
rect 8159 16408 8484 16436
rect 8159 16405 8171 16408
rect 8113 16399 8171 16405
rect 8478 16396 8484 16408
rect 8536 16436 8542 16448
rect 8665 16439 8723 16445
rect 8665 16436 8677 16439
rect 8536 16408 8677 16436
rect 8536 16396 8542 16408
rect 8665 16405 8677 16408
rect 8711 16405 8723 16439
rect 8665 16399 8723 16405
rect 9122 16396 9128 16448
rect 9180 16396 9186 16448
rect 9582 16396 9588 16448
rect 9640 16396 9646 16448
rect 10318 16396 10324 16448
rect 10376 16396 10382 16448
rect 10781 16439 10839 16445
rect 10781 16405 10793 16439
rect 10827 16436 10839 16439
rect 11054 16436 11060 16448
rect 10827 16408 11060 16436
rect 10827 16405 10839 16408
rect 10781 16399 10839 16405
rect 11054 16396 11060 16408
rect 11112 16396 11118 16448
rect 11238 16396 11244 16448
rect 11296 16436 11302 16448
rect 13630 16436 13636 16448
rect 11296 16408 13636 16436
rect 11296 16396 11302 16408
rect 13630 16396 13636 16408
rect 13688 16396 13694 16448
rect 15102 16396 15108 16448
rect 15160 16396 15166 16448
rect 15473 16439 15531 16445
rect 15473 16405 15485 16439
rect 15519 16436 15531 16439
rect 16114 16436 16120 16448
rect 15519 16408 16120 16436
rect 15519 16405 15531 16408
rect 15473 16399 15531 16405
rect 16114 16396 16120 16408
rect 16172 16436 16178 16448
rect 16209 16439 16267 16445
rect 16209 16436 16221 16439
rect 16172 16408 16221 16436
rect 16172 16396 16178 16408
rect 16209 16405 16221 16408
rect 16255 16436 16267 16439
rect 18414 16436 18420 16448
rect 16255 16408 18420 16436
rect 16255 16405 16267 16408
rect 16209 16399 16267 16405
rect 18414 16396 18420 16408
rect 18472 16396 18478 16448
rect 19518 16396 19524 16448
rect 19576 16436 19582 16448
rect 19613 16439 19671 16445
rect 19613 16436 19625 16439
rect 19576 16408 19625 16436
rect 19576 16396 19582 16408
rect 19613 16405 19625 16408
rect 19659 16405 19671 16439
rect 19613 16399 19671 16405
rect 20530 16396 20536 16448
rect 20588 16436 20594 16448
rect 23477 16439 23535 16445
rect 23477 16436 23489 16439
rect 20588 16408 23489 16436
rect 20588 16396 20594 16408
rect 23477 16405 23489 16408
rect 23523 16436 23535 16439
rect 24578 16436 24584 16448
rect 23523 16408 24584 16436
rect 23523 16405 23535 16408
rect 23477 16399 23535 16405
rect 24578 16396 24584 16408
rect 24636 16396 24642 16448
rect 1104 16346 25852 16368
rect 1104 16294 7950 16346
rect 8002 16294 8014 16346
rect 8066 16294 8078 16346
rect 8130 16294 8142 16346
rect 8194 16294 8206 16346
rect 8258 16294 17950 16346
rect 18002 16294 18014 16346
rect 18066 16294 18078 16346
rect 18130 16294 18142 16346
rect 18194 16294 18206 16346
rect 18258 16294 25852 16346
rect 1104 16272 25852 16294
rect 6362 16192 6368 16244
rect 6420 16232 6426 16244
rect 7009 16235 7067 16241
rect 7009 16232 7021 16235
rect 6420 16204 7021 16232
rect 6420 16192 6426 16204
rect 7009 16201 7021 16204
rect 7055 16201 7067 16235
rect 7009 16195 7067 16201
rect 7377 16235 7435 16241
rect 7377 16201 7389 16235
rect 7423 16232 7435 16235
rect 9122 16232 9128 16244
rect 7423 16204 9128 16232
rect 7423 16201 7435 16204
rect 7377 16195 7435 16201
rect 9122 16192 9128 16204
rect 9180 16192 9186 16244
rect 9582 16192 9588 16244
rect 9640 16192 9646 16244
rect 10045 16235 10103 16241
rect 10045 16201 10057 16235
rect 10091 16232 10103 16235
rect 11146 16232 11152 16244
rect 10091 16204 11152 16232
rect 10091 16201 10103 16204
rect 10045 16195 10103 16201
rect 11146 16192 11152 16204
rect 11204 16192 11210 16244
rect 11882 16232 11888 16244
rect 11808 16204 11888 16232
rect 7469 16167 7527 16173
rect 7469 16133 7481 16167
rect 7515 16164 7527 16167
rect 10318 16164 10324 16176
rect 7515 16136 10324 16164
rect 7515 16133 7527 16136
rect 7469 16127 7527 16133
rect 10318 16124 10324 16136
rect 10376 16124 10382 16176
rect 8202 16096 8208 16108
rect 7668 16068 8208 16096
rect 7668 16037 7696 16068
rect 8202 16056 8208 16068
rect 8260 16056 8266 16108
rect 9953 16099 10011 16105
rect 9953 16096 9965 16099
rect 9232 16068 9965 16096
rect 7653 16031 7711 16037
rect 7653 15997 7665 16031
rect 7699 15997 7711 16031
rect 7653 15991 7711 15997
rect 7742 15920 7748 15972
rect 7800 15960 7806 15972
rect 9232 15969 9260 16068
rect 9953 16065 9965 16068
rect 9999 16065 10011 16099
rect 11808 16096 11836 16204
rect 11882 16192 11888 16204
rect 11940 16232 11946 16244
rect 13538 16232 13544 16244
rect 11940 16204 13544 16232
rect 11940 16192 11946 16204
rect 13538 16192 13544 16204
rect 13596 16192 13602 16244
rect 16206 16192 16212 16244
rect 16264 16192 16270 16244
rect 16666 16192 16672 16244
rect 16724 16232 16730 16244
rect 17221 16235 17279 16241
rect 17221 16232 17233 16235
rect 16724 16204 17233 16232
rect 16724 16192 16730 16204
rect 17221 16201 17233 16204
rect 17267 16201 17279 16235
rect 17221 16195 17279 16201
rect 18782 16192 18788 16244
rect 18840 16192 18846 16244
rect 19150 16192 19156 16244
rect 19208 16192 19214 16244
rect 19518 16192 19524 16244
rect 19576 16192 19582 16244
rect 20346 16192 20352 16244
rect 20404 16232 20410 16244
rect 20809 16235 20867 16241
rect 20809 16232 20821 16235
rect 20404 16204 20821 16232
rect 20404 16192 20410 16204
rect 20809 16201 20821 16204
rect 20855 16201 20867 16235
rect 20809 16195 20867 16201
rect 22186 16192 22192 16244
rect 22244 16232 22250 16244
rect 22462 16232 22468 16244
rect 22244 16204 22468 16232
rect 22244 16192 22250 16204
rect 22462 16192 22468 16204
rect 22520 16232 22526 16244
rect 22646 16232 22652 16244
rect 22520 16204 22652 16232
rect 22520 16192 22526 16204
rect 22646 16192 22652 16204
rect 22704 16192 22710 16244
rect 12066 16124 12072 16176
rect 12124 16124 12130 16176
rect 15657 16167 15715 16173
rect 15657 16133 15669 16167
rect 15703 16164 15715 16167
rect 16224 16164 16252 16192
rect 15703 16136 16252 16164
rect 18800 16164 18828 16192
rect 19613 16167 19671 16173
rect 19613 16164 19625 16167
rect 18800 16136 19625 16164
rect 15703 16133 15715 16136
rect 15657 16127 15715 16133
rect 19613 16133 19625 16136
rect 19659 16133 19671 16167
rect 21358 16164 21364 16176
rect 19613 16127 19671 16133
rect 19812 16136 21364 16164
rect 13630 16096 13636 16108
rect 9953 16059 10011 16065
rect 10244 16068 11836 16096
rect 13202 16068 13636 16096
rect 9217 15963 9275 15969
rect 9217 15960 9229 15963
rect 7800 15932 9229 15960
rect 7800 15920 7806 15932
rect 9217 15929 9229 15932
rect 9263 15929 9275 15963
rect 9968 15960 9996 16059
rect 10244 16037 10272 16068
rect 13630 16056 13636 16068
rect 13688 16096 13694 16108
rect 13688 16068 14044 16096
rect 13688 16056 13694 16068
rect 10229 16031 10287 16037
rect 10229 15997 10241 16031
rect 10275 15997 10287 16031
rect 10229 15991 10287 15997
rect 10870 15988 10876 16040
rect 10928 16028 10934 16040
rect 11790 16028 11796 16040
rect 10928 16000 11796 16028
rect 10928 15988 10934 16000
rect 11790 15988 11796 16000
rect 11848 15988 11854 16040
rect 11698 15960 11704 15972
rect 9968 15932 11704 15960
rect 9217 15923 9275 15929
rect 11698 15920 11704 15932
rect 11756 15920 11762 15972
rect 8386 15852 8392 15904
rect 8444 15892 8450 15904
rect 8849 15895 8907 15901
rect 8849 15892 8861 15895
rect 8444 15864 8861 15892
rect 8444 15852 8450 15864
rect 8849 15861 8861 15864
rect 8895 15861 8907 15895
rect 8849 15855 8907 15861
rect 13538 15852 13544 15904
rect 13596 15852 13602 15904
rect 14016 15901 14044 16068
rect 19812 16037 19840 16136
rect 21358 16124 21364 16136
rect 21416 16124 21422 16176
rect 20717 16099 20775 16105
rect 20717 16065 20729 16099
rect 20763 16096 20775 16099
rect 21266 16096 21272 16108
rect 20763 16068 21272 16096
rect 20763 16065 20775 16068
rect 20717 16059 20775 16065
rect 21266 16056 21272 16068
rect 21324 16056 21330 16108
rect 22373 16099 22431 16105
rect 22373 16065 22385 16099
rect 22419 16096 22431 16099
rect 23201 16099 23259 16105
rect 23201 16096 23213 16099
rect 22419 16068 23213 16096
rect 22419 16065 22431 16068
rect 22373 16059 22431 16065
rect 23201 16065 23213 16068
rect 23247 16065 23259 16099
rect 23201 16059 23259 16065
rect 24118 16056 24124 16108
rect 24176 16056 24182 16108
rect 19797 16031 19855 16037
rect 19797 15997 19809 16031
rect 19843 15997 19855 16031
rect 19797 15991 19855 15997
rect 20990 15988 20996 16040
rect 21048 15988 21054 16040
rect 22465 16031 22523 16037
rect 22465 15997 22477 16031
rect 22511 15997 22523 16031
rect 22465 15991 22523 15997
rect 22649 16031 22707 16037
rect 22649 15997 22661 16031
rect 22695 16028 22707 16031
rect 23658 16028 23664 16040
rect 22695 16000 23664 16028
rect 22695 15997 22707 16000
rect 22649 15991 22707 15997
rect 15841 15963 15899 15969
rect 15841 15929 15853 15963
rect 15887 15960 15899 15963
rect 16298 15960 16304 15972
rect 15887 15932 16304 15960
rect 15887 15929 15899 15932
rect 15841 15923 15899 15929
rect 16298 15920 16304 15932
rect 16356 15920 16362 15972
rect 17402 15920 17408 15972
rect 17460 15960 17466 15972
rect 18601 15963 18659 15969
rect 18601 15960 18613 15963
rect 17460 15932 18613 15960
rect 17460 15920 17466 15932
rect 18601 15929 18613 15932
rect 18647 15929 18659 15963
rect 18601 15923 18659 15929
rect 20438 15920 20444 15972
rect 20496 15960 20502 15972
rect 22480 15960 22508 15991
rect 23658 15988 23664 16000
rect 23716 15988 23722 16040
rect 24762 15988 24768 16040
rect 24820 15988 24826 16040
rect 20496 15932 22508 15960
rect 20496 15920 20502 15932
rect 14001 15895 14059 15901
rect 14001 15861 14013 15895
rect 14047 15892 14059 15895
rect 17034 15892 17040 15904
rect 14047 15864 17040 15892
rect 14047 15861 14059 15864
rect 14001 15855 14059 15861
rect 17034 15852 17040 15864
rect 17092 15892 17098 15904
rect 17497 15895 17555 15901
rect 17497 15892 17509 15895
rect 17092 15864 17509 15892
rect 17092 15852 17098 15864
rect 17497 15861 17509 15864
rect 17543 15892 17555 15895
rect 17770 15892 17776 15904
rect 17543 15864 17776 15892
rect 17543 15861 17555 15864
rect 17497 15855 17555 15861
rect 17770 15852 17776 15864
rect 17828 15852 17834 15904
rect 17865 15895 17923 15901
rect 17865 15861 17877 15895
rect 17911 15892 17923 15895
rect 18230 15892 18236 15904
rect 17911 15864 18236 15892
rect 17911 15861 17923 15864
rect 17865 15855 17923 15861
rect 18230 15852 18236 15864
rect 18288 15852 18294 15904
rect 20349 15895 20407 15901
rect 20349 15861 20361 15895
rect 20395 15892 20407 15895
rect 21542 15892 21548 15904
rect 20395 15864 21548 15892
rect 20395 15861 20407 15864
rect 20349 15855 20407 15861
rect 21542 15852 21548 15864
rect 21600 15852 21606 15904
rect 22005 15895 22063 15901
rect 22005 15861 22017 15895
rect 22051 15892 22063 15895
rect 23474 15892 23480 15904
rect 22051 15864 23480 15892
rect 22051 15861 22063 15864
rect 22005 15855 22063 15861
rect 23474 15852 23480 15864
rect 23532 15852 23538 15904
rect 1104 15802 25852 15824
rect 1104 15750 2950 15802
rect 3002 15750 3014 15802
rect 3066 15750 3078 15802
rect 3130 15750 3142 15802
rect 3194 15750 3206 15802
rect 3258 15750 12950 15802
rect 13002 15750 13014 15802
rect 13066 15750 13078 15802
rect 13130 15750 13142 15802
rect 13194 15750 13206 15802
rect 13258 15750 22950 15802
rect 23002 15750 23014 15802
rect 23066 15750 23078 15802
rect 23130 15750 23142 15802
rect 23194 15750 23206 15802
rect 23258 15750 25852 15802
rect 1104 15728 25852 15750
rect 8202 15648 8208 15700
rect 8260 15688 8266 15700
rect 8481 15691 8539 15697
rect 8481 15688 8493 15691
rect 8260 15660 8493 15688
rect 8260 15648 8266 15660
rect 8481 15657 8493 15660
rect 8527 15657 8539 15691
rect 8481 15651 8539 15657
rect 10134 15648 10140 15700
rect 10192 15688 10198 15700
rect 10192 15660 11560 15688
rect 10192 15648 10198 15660
rect 11532 15620 11560 15660
rect 12158 15648 12164 15700
rect 12216 15688 12222 15700
rect 12989 15691 13047 15697
rect 12989 15688 13001 15691
rect 12216 15660 13001 15688
rect 12216 15648 12222 15660
rect 12989 15657 13001 15660
rect 13035 15657 13047 15691
rect 12989 15651 13047 15657
rect 15010 15648 15016 15700
rect 15068 15648 15074 15700
rect 15286 15648 15292 15700
rect 15344 15688 15350 15700
rect 17405 15691 17463 15697
rect 15344 15660 17356 15688
rect 15344 15648 15350 15660
rect 14090 15620 14096 15632
rect 11532 15592 14096 15620
rect 14090 15580 14096 15592
rect 14148 15580 14154 15632
rect 17328 15620 17356 15660
rect 17405 15657 17417 15691
rect 17451 15688 17463 15691
rect 18322 15688 18328 15700
rect 17451 15660 18328 15688
rect 17451 15657 17463 15660
rect 17405 15651 17463 15657
rect 18322 15648 18328 15660
rect 18380 15648 18386 15700
rect 18414 15648 18420 15700
rect 18472 15688 18478 15700
rect 20990 15688 20996 15700
rect 18472 15660 20996 15688
rect 18472 15648 18478 15660
rect 20990 15648 20996 15660
rect 21048 15648 21054 15700
rect 18969 15623 19027 15629
rect 18969 15620 18981 15623
rect 17328 15592 18981 15620
rect 7009 15555 7067 15561
rect 7009 15521 7021 15555
rect 7055 15552 7067 15555
rect 8570 15552 8576 15564
rect 7055 15524 8576 15552
rect 7055 15521 7067 15524
rect 7009 15515 7067 15521
rect 8570 15512 8576 15524
rect 8628 15512 8634 15564
rect 10229 15555 10287 15561
rect 10229 15521 10241 15555
rect 10275 15552 10287 15555
rect 10870 15552 10876 15564
rect 10275 15524 10876 15552
rect 10275 15521 10287 15524
rect 10229 15515 10287 15521
rect 10870 15512 10876 15524
rect 10928 15512 10934 15564
rect 12713 15555 12771 15561
rect 12713 15521 12725 15555
rect 12759 15552 12771 15555
rect 13541 15555 13599 15561
rect 13541 15552 13553 15555
rect 12759 15524 13553 15552
rect 12759 15521 12771 15524
rect 12713 15515 12771 15521
rect 13541 15521 13553 15524
rect 13587 15552 13599 15555
rect 13722 15552 13728 15564
rect 13587 15524 13728 15552
rect 13587 15521 13599 15524
rect 13541 15515 13599 15521
rect 13722 15512 13728 15524
rect 13780 15512 13786 15564
rect 18230 15552 18236 15564
rect 14384 15524 18236 15552
rect 6730 15444 6736 15496
rect 6788 15444 6794 15496
rect 9030 15444 9036 15496
rect 9088 15484 9094 15496
rect 9125 15487 9183 15493
rect 9125 15484 9137 15487
rect 9088 15456 9137 15484
rect 9088 15444 9094 15456
rect 9125 15453 9137 15456
rect 9171 15453 9183 15487
rect 9125 15447 9183 15453
rect 12529 15487 12587 15493
rect 12529 15453 12541 15487
rect 12575 15484 12587 15487
rect 13449 15487 13507 15493
rect 13449 15484 13461 15487
rect 12575 15456 13461 15484
rect 12575 15453 12587 15456
rect 12529 15447 12587 15453
rect 13449 15453 13461 15456
rect 13495 15484 13507 15487
rect 13630 15484 13636 15496
rect 13495 15456 13636 15484
rect 13495 15453 13507 15456
rect 13449 15447 13507 15453
rect 13630 15444 13636 15456
rect 13688 15484 13694 15496
rect 14384 15484 14412 15524
rect 18230 15512 18236 15524
rect 18288 15512 18294 15564
rect 18432 15561 18460 15592
rect 18969 15589 18981 15592
rect 19015 15589 19027 15623
rect 18969 15583 19027 15589
rect 19429 15623 19487 15629
rect 19429 15589 19441 15623
rect 19475 15620 19487 15623
rect 21174 15620 21180 15632
rect 19475 15592 21180 15620
rect 19475 15589 19487 15592
rect 19429 15583 19487 15589
rect 21174 15580 21180 15592
rect 21232 15580 21238 15632
rect 18417 15555 18475 15561
rect 18417 15521 18429 15555
rect 18463 15521 18475 15555
rect 18417 15515 18475 15521
rect 18601 15555 18659 15561
rect 18601 15521 18613 15555
rect 18647 15552 18659 15555
rect 18874 15552 18880 15564
rect 18647 15524 18880 15552
rect 18647 15521 18659 15524
rect 18601 15515 18659 15521
rect 18874 15512 18880 15524
rect 18932 15512 18938 15564
rect 19886 15512 19892 15564
rect 19944 15512 19950 15564
rect 20073 15555 20131 15561
rect 20073 15521 20085 15555
rect 20119 15552 20131 15555
rect 20530 15552 20536 15564
rect 20119 15524 20536 15552
rect 20119 15521 20131 15524
rect 20073 15515 20131 15521
rect 20530 15512 20536 15524
rect 20588 15512 20594 15564
rect 21266 15512 21272 15564
rect 21324 15512 21330 15564
rect 13688 15456 14412 15484
rect 14553 15487 14611 15493
rect 13688 15444 13694 15456
rect 14553 15453 14565 15487
rect 14599 15484 14611 15487
rect 15010 15484 15016 15496
rect 14599 15456 15016 15484
rect 14599 15453 14611 15456
rect 14553 15447 14611 15453
rect 15010 15444 15016 15456
rect 15068 15444 15074 15496
rect 15194 15444 15200 15496
rect 15252 15484 15258 15496
rect 15657 15487 15715 15493
rect 15657 15484 15669 15487
rect 15252 15456 15669 15484
rect 15252 15444 15258 15456
rect 15657 15453 15669 15456
rect 15703 15453 15715 15487
rect 15657 15447 15715 15453
rect 17034 15444 17040 15496
rect 17092 15444 17098 15496
rect 17402 15444 17408 15496
rect 17460 15484 17466 15496
rect 19797 15487 19855 15493
rect 19797 15484 19809 15487
rect 17460 15456 19809 15484
rect 17460 15444 17466 15456
rect 19797 15453 19809 15456
rect 19843 15453 19855 15487
rect 19797 15447 19855 15453
rect 20714 15444 20720 15496
rect 20772 15484 20778 15496
rect 20809 15487 20867 15493
rect 20809 15484 20821 15487
rect 20772 15456 20821 15484
rect 20772 15444 20778 15456
rect 20809 15453 20821 15456
rect 20855 15453 20867 15487
rect 20809 15447 20867 15453
rect 21634 15444 21640 15496
rect 21692 15484 21698 15496
rect 22097 15487 22155 15493
rect 22097 15484 22109 15487
rect 21692 15456 22109 15484
rect 21692 15444 21698 15456
rect 22097 15453 22109 15456
rect 22143 15453 22155 15487
rect 22097 15447 22155 15453
rect 22738 15444 22744 15496
rect 22796 15444 22802 15496
rect 24578 15444 24584 15496
rect 24636 15444 24642 15496
rect 8478 15416 8484 15428
rect 8234 15388 8484 15416
rect 7650 15308 7656 15360
rect 7708 15348 7714 15360
rect 8312 15348 8340 15388
rect 8478 15376 8484 15388
rect 8536 15376 8542 15428
rect 8754 15376 8760 15428
rect 8812 15416 8818 15428
rect 10134 15416 10140 15428
rect 8812 15388 10140 15416
rect 8812 15376 8818 15388
rect 10134 15376 10140 15388
rect 10192 15376 10198 15428
rect 10505 15419 10563 15425
rect 10505 15385 10517 15419
rect 10551 15416 10563 15419
rect 10778 15416 10784 15428
rect 10551 15388 10784 15416
rect 10551 15385 10563 15388
rect 10505 15379 10563 15385
rect 10778 15376 10784 15388
rect 10836 15376 10842 15428
rect 11238 15376 11244 15428
rect 11296 15376 11302 15428
rect 13262 15376 13268 15428
rect 13320 15416 13326 15428
rect 13357 15419 13415 15425
rect 13357 15416 13369 15419
rect 13320 15388 13369 15416
rect 13320 15376 13326 15388
rect 13357 15385 13369 15388
rect 13403 15416 13415 15419
rect 15562 15416 15568 15428
rect 13403 15388 15568 15416
rect 13403 15385 13415 15388
rect 13357 15379 13415 15385
rect 15562 15376 15568 15388
rect 15620 15416 15626 15428
rect 15838 15416 15844 15428
rect 15620 15388 15844 15416
rect 15620 15376 15626 15388
rect 15838 15376 15844 15388
rect 15896 15376 15902 15428
rect 15930 15376 15936 15428
rect 15988 15376 15994 15428
rect 20530 15416 20536 15428
rect 17972 15388 20536 15416
rect 7708 15320 8340 15348
rect 7708 15308 7714 15320
rect 9122 15308 9128 15360
rect 9180 15348 9186 15360
rect 9769 15351 9827 15357
rect 9769 15348 9781 15351
rect 9180 15320 9781 15348
rect 9180 15308 9186 15320
rect 9769 15317 9781 15320
rect 9815 15317 9827 15351
rect 9769 15311 9827 15317
rect 11514 15308 11520 15360
rect 11572 15348 11578 15360
rect 11977 15351 12035 15357
rect 11977 15348 11989 15351
rect 11572 15320 11989 15348
rect 11572 15308 11578 15320
rect 11977 15317 11989 15320
rect 12023 15348 12035 15351
rect 12342 15348 12348 15360
rect 12023 15320 12348 15348
rect 12023 15317 12035 15320
rect 11977 15311 12035 15317
rect 12342 15308 12348 15320
rect 12400 15308 12406 15360
rect 14642 15308 14648 15360
rect 14700 15308 14706 15360
rect 17972 15357 18000 15388
rect 20530 15376 20536 15388
rect 20588 15376 20594 15428
rect 23845 15419 23903 15425
rect 23845 15385 23857 15419
rect 23891 15416 23903 15419
rect 24946 15416 24952 15428
rect 23891 15388 24952 15416
rect 23891 15385 23903 15388
rect 23845 15379 23903 15385
rect 24946 15376 24952 15388
rect 25004 15376 25010 15428
rect 17957 15351 18015 15357
rect 17957 15317 17969 15351
rect 18003 15317 18015 15351
rect 17957 15311 18015 15317
rect 18230 15308 18236 15360
rect 18288 15348 18294 15360
rect 18325 15351 18383 15357
rect 18325 15348 18337 15351
rect 18288 15320 18337 15348
rect 18288 15308 18294 15320
rect 18325 15317 18337 15320
rect 18371 15317 18383 15351
rect 18325 15311 18383 15317
rect 20625 15351 20683 15357
rect 20625 15317 20637 15351
rect 20671 15348 20683 15351
rect 21082 15348 21088 15360
rect 20671 15320 21088 15348
rect 20671 15317 20683 15320
rect 20625 15311 20683 15317
rect 21082 15308 21088 15320
rect 21140 15308 21146 15360
rect 21358 15308 21364 15360
rect 21416 15348 21422 15360
rect 21913 15351 21971 15357
rect 21913 15348 21925 15351
rect 21416 15320 21925 15348
rect 21416 15308 21422 15320
rect 21913 15317 21925 15320
rect 21959 15317 21971 15351
rect 21913 15311 21971 15317
rect 22278 15308 22284 15360
rect 22336 15348 22342 15360
rect 25225 15351 25283 15357
rect 25225 15348 25237 15351
rect 22336 15320 25237 15348
rect 22336 15308 22342 15320
rect 25225 15317 25237 15320
rect 25271 15317 25283 15351
rect 25225 15311 25283 15317
rect 1104 15258 25852 15280
rect 1104 15206 7950 15258
rect 8002 15206 8014 15258
rect 8066 15206 8078 15258
rect 8130 15206 8142 15258
rect 8194 15206 8206 15258
rect 8258 15206 17950 15258
rect 18002 15206 18014 15258
rect 18066 15206 18078 15258
rect 18130 15206 18142 15258
rect 18194 15206 18206 15258
rect 18258 15206 25852 15258
rect 1104 15184 25852 15206
rect 7834 15104 7840 15156
rect 7892 15144 7898 15156
rect 11793 15147 11851 15153
rect 11793 15144 11805 15147
rect 7892 15116 11805 15144
rect 7892 15104 7898 15116
rect 11793 15113 11805 15116
rect 11839 15113 11851 15147
rect 11793 15107 11851 15113
rect 11974 15104 11980 15156
rect 12032 15144 12038 15156
rect 12989 15147 13047 15153
rect 12989 15144 13001 15147
rect 12032 15116 13001 15144
rect 12032 15104 12038 15116
rect 12989 15113 13001 15116
rect 13035 15113 13047 15147
rect 12989 15107 13047 15113
rect 13262 15104 13268 15156
rect 13320 15144 13326 15156
rect 13357 15147 13415 15153
rect 13357 15144 13369 15147
rect 13320 15116 13369 15144
rect 13320 15104 13326 15116
rect 13357 15113 13369 15116
rect 13403 15113 13415 15147
rect 13357 15107 13415 15113
rect 13722 15104 13728 15156
rect 13780 15144 13786 15156
rect 13998 15144 14004 15156
rect 13780 15116 14004 15144
rect 13780 15104 13786 15116
rect 13998 15104 14004 15116
rect 14056 15104 14062 15156
rect 14090 15104 14096 15156
rect 14148 15144 14154 15156
rect 14553 15147 14611 15153
rect 14553 15144 14565 15147
rect 14148 15116 14565 15144
rect 14148 15104 14154 15116
rect 14553 15113 14565 15116
rect 14599 15113 14611 15147
rect 14553 15107 14611 15113
rect 14645 15147 14703 15153
rect 14645 15113 14657 15147
rect 14691 15144 14703 15147
rect 15286 15144 15292 15156
rect 14691 15116 15292 15144
rect 14691 15113 14703 15116
rect 14645 15107 14703 15113
rect 15286 15104 15292 15116
rect 15344 15104 15350 15156
rect 15930 15104 15936 15156
rect 15988 15144 15994 15156
rect 16301 15147 16359 15153
rect 16301 15144 16313 15147
rect 15988 15116 16313 15144
rect 15988 15104 15994 15116
rect 16301 15113 16313 15116
rect 16347 15113 16359 15147
rect 16301 15107 16359 15113
rect 16482 15104 16488 15156
rect 16540 15144 16546 15156
rect 18049 15147 18107 15153
rect 18049 15144 18061 15147
rect 16540 15116 18061 15144
rect 16540 15104 16546 15116
rect 18049 15113 18061 15116
rect 18095 15113 18107 15147
rect 18049 15107 18107 15113
rect 20533 15147 20591 15153
rect 20533 15113 20545 15147
rect 20579 15144 20591 15147
rect 20622 15144 20628 15156
rect 20579 15116 20628 15144
rect 20579 15113 20591 15116
rect 20533 15107 20591 15113
rect 20622 15104 20628 15116
rect 20680 15104 20686 15156
rect 21450 15144 21456 15156
rect 21008 15116 21456 15144
rect 7650 15036 7656 15088
rect 7708 15076 7714 15088
rect 7745 15079 7803 15085
rect 7745 15076 7757 15079
rect 7708 15048 7757 15076
rect 7708 15036 7714 15048
rect 7745 15045 7757 15048
rect 7791 15045 7803 15079
rect 7745 15039 7803 15045
rect 8386 15036 8392 15088
rect 8444 15036 8450 15088
rect 10137 15079 10195 15085
rect 10137 15045 10149 15079
rect 10183 15076 10195 15079
rect 10778 15076 10784 15088
rect 10183 15048 10784 15076
rect 10183 15045 10195 15048
rect 10137 15039 10195 15045
rect 10778 15036 10784 15048
rect 10836 15036 10842 15088
rect 13446 15036 13452 15088
rect 13504 15076 13510 15088
rect 13504 15048 13584 15076
rect 13504 15036 13510 15048
rect 10505 15011 10563 15017
rect 10505 15008 10517 15011
rect 9522 14994 10517 15008
rect 9508 14980 10517 14994
rect 8113 14943 8171 14949
rect 8113 14909 8125 14943
rect 8159 14909 8171 14943
rect 8113 14903 8171 14909
rect 8128 14872 8156 14903
rect 8478 14900 8484 14952
rect 8536 14940 8542 14952
rect 9508 14940 9536 14980
rect 10505 14977 10517 14980
rect 10551 15008 10563 15011
rect 11238 15008 11244 15020
rect 10551 14980 11244 15008
rect 10551 14977 10563 14980
rect 10505 14971 10563 14977
rect 11238 14968 11244 14980
rect 11296 14968 11302 15020
rect 12161 15011 12219 15017
rect 12161 14977 12173 15011
rect 12207 15008 12219 15011
rect 12802 15008 12808 15020
rect 12207 14980 12808 15008
rect 12207 14977 12219 14980
rect 12161 14971 12219 14977
rect 12802 14968 12808 14980
rect 12860 14968 12866 15020
rect 8536 14912 9536 14940
rect 12253 14943 12311 14949
rect 8536 14900 8542 14912
rect 12253 14909 12265 14943
rect 12299 14909 12311 14943
rect 12253 14903 12311 14909
rect 8128 14844 8248 14872
rect 8220 14804 8248 14844
rect 8386 14804 8392 14816
rect 8220 14776 8392 14804
rect 8386 14764 8392 14776
rect 8444 14764 8450 14816
rect 12268 14804 12296 14903
rect 12342 14900 12348 14952
rect 12400 14900 12406 14952
rect 13556 14949 13584 15048
rect 16666 15036 16672 15088
rect 16724 15076 16730 15088
rect 16945 15079 17003 15085
rect 16945 15076 16957 15079
rect 16724 15048 16957 15076
rect 16724 15036 16730 15048
rect 16945 15045 16957 15048
rect 16991 15045 17003 15079
rect 21008 15076 21036 15116
rect 21450 15104 21456 15116
rect 21508 15104 21514 15156
rect 20286 15048 21036 15076
rect 16945 15039 17003 15045
rect 21082 15036 21088 15088
rect 21140 15076 21146 15088
rect 23293 15079 23351 15085
rect 23293 15076 23305 15079
rect 21140 15048 23305 15076
rect 21140 15036 21146 15048
rect 23293 15045 23305 15048
rect 23339 15045 23351 15079
rect 23293 15039 23351 15045
rect 14108 14980 14872 15008
rect 13449 14943 13507 14949
rect 13449 14909 13461 14943
rect 13495 14909 13507 14943
rect 13449 14903 13507 14909
rect 13541 14943 13599 14949
rect 13541 14909 13553 14943
rect 13587 14909 13599 14943
rect 13541 14903 13599 14909
rect 13464 14872 13492 14903
rect 13630 14872 13636 14884
rect 13464 14844 13636 14872
rect 13630 14832 13636 14844
rect 13688 14832 13694 14884
rect 14108 14804 14136 14980
rect 14734 14900 14740 14952
rect 14792 14900 14798 14952
rect 14844 14940 14872 14980
rect 15654 14968 15660 15020
rect 15712 14968 15718 15020
rect 17954 14968 17960 15020
rect 18012 14968 18018 15020
rect 21177 15011 21235 15017
rect 21177 14977 21189 15011
rect 21223 15008 21235 15011
rect 21818 15008 21824 15020
rect 21223 14980 21824 15008
rect 21223 14977 21235 14980
rect 21177 14971 21235 14977
rect 21818 14968 21824 14980
rect 21876 14968 21882 15020
rect 21910 14968 21916 15020
rect 21968 15008 21974 15020
rect 22557 15011 22615 15017
rect 22557 15008 22569 15011
rect 21968 14980 22569 15008
rect 21968 14968 21974 14980
rect 22557 14977 22569 14980
rect 22603 14977 22615 15011
rect 22557 14971 22615 14977
rect 24121 15011 24179 15017
rect 24121 14977 24133 15011
rect 24167 15008 24179 15011
rect 24302 15008 24308 15020
rect 24167 14980 24308 15008
rect 24167 14977 24179 14980
rect 24121 14971 24179 14977
rect 24302 14968 24308 14980
rect 24360 14968 24366 15020
rect 16114 14940 16120 14952
rect 14844 14912 16120 14940
rect 16114 14900 16120 14912
rect 16172 14900 16178 14952
rect 18230 14900 18236 14952
rect 18288 14900 18294 14952
rect 18322 14900 18328 14952
rect 18380 14940 18386 14952
rect 18690 14940 18696 14952
rect 18380 14912 18696 14940
rect 18380 14900 18386 14912
rect 18690 14900 18696 14912
rect 18748 14940 18754 14952
rect 18785 14943 18843 14949
rect 18785 14940 18797 14943
rect 18748 14912 18797 14940
rect 18748 14900 18754 14912
rect 18785 14909 18797 14912
rect 18831 14909 18843 14943
rect 18785 14903 18843 14909
rect 19061 14943 19119 14949
rect 19061 14909 19073 14943
rect 19107 14940 19119 14943
rect 19150 14940 19156 14952
rect 19107 14912 19156 14940
rect 19107 14909 19119 14912
rect 19061 14903 19119 14909
rect 19150 14900 19156 14912
rect 19208 14900 19214 14952
rect 19794 14900 19800 14952
rect 19852 14940 19858 14952
rect 22186 14940 22192 14952
rect 19852 14912 20116 14940
rect 19852 14900 19858 14912
rect 14185 14875 14243 14881
rect 14185 14841 14197 14875
rect 14231 14872 14243 14875
rect 16206 14872 16212 14884
rect 14231 14844 16212 14872
rect 14231 14841 14243 14844
rect 14185 14835 14243 14841
rect 16206 14832 16212 14844
rect 16264 14832 16270 14884
rect 20088 14872 20116 14912
rect 22066 14912 22192 14940
rect 22066 14872 22094 14912
rect 22186 14900 22192 14912
rect 22244 14900 22250 14952
rect 24670 14900 24676 14952
rect 24728 14900 24734 14952
rect 20088 14844 22094 14872
rect 22738 14832 22744 14884
rect 22796 14832 22802 14884
rect 23477 14875 23535 14881
rect 23477 14841 23489 14875
rect 23523 14872 23535 14875
rect 23934 14872 23940 14884
rect 23523 14844 23940 14872
rect 23523 14841 23535 14844
rect 23477 14835 23535 14841
rect 23934 14832 23940 14844
rect 23992 14832 23998 14884
rect 12268 14776 14136 14804
rect 16758 14764 16764 14816
rect 16816 14804 16822 14816
rect 17037 14807 17095 14813
rect 17037 14804 17049 14807
rect 16816 14776 17049 14804
rect 16816 14764 16822 14776
rect 17037 14773 17049 14776
rect 17083 14773 17095 14807
rect 17037 14767 17095 14773
rect 17589 14807 17647 14813
rect 17589 14773 17601 14807
rect 17635 14804 17647 14807
rect 19426 14804 19432 14816
rect 17635 14776 19432 14804
rect 17635 14773 17647 14776
rect 17589 14767 17647 14773
rect 19426 14764 19432 14776
rect 19484 14764 19490 14816
rect 19518 14764 19524 14816
rect 19576 14804 19582 14816
rect 20993 14807 21051 14813
rect 20993 14804 21005 14807
rect 19576 14776 21005 14804
rect 19576 14764 19582 14776
rect 20993 14773 21005 14776
rect 21039 14773 21051 14807
rect 20993 14767 21051 14773
rect 21450 14764 21456 14816
rect 21508 14804 21514 14816
rect 22646 14804 22652 14816
rect 21508 14776 22652 14804
rect 21508 14764 21514 14776
rect 22646 14764 22652 14776
rect 22704 14764 22710 14816
rect 1104 14714 25852 14736
rect 1104 14662 2950 14714
rect 3002 14662 3014 14714
rect 3066 14662 3078 14714
rect 3130 14662 3142 14714
rect 3194 14662 3206 14714
rect 3258 14662 12950 14714
rect 13002 14662 13014 14714
rect 13066 14662 13078 14714
rect 13130 14662 13142 14714
rect 13194 14662 13206 14714
rect 13258 14662 22950 14714
rect 23002 14662 23014 14714
rect 23066 14662 23078 14714
rect 23130 14662 23142 14714
rect 23194 14662 23206 14714
rect 23258 14662 25852 14714
rect 1104 14640 25852 14662
rect 8570 14560 8576 14612
rect 8628 14560 8634 14612
rect 11054 14560 11060 14612
rect 11112 14600 11118 14612
rect 12989 14603 13047 14609
rect 12989 14600 13001 14603
rect 11112 14572 13001 14600
rect 11112 14560 11118 14572
rect 12989 14569 13001 14572
rect 13035 14569 13047 14603
rect 12989 14563 13047 14569
rect 14826 14560 14832 14612
rect 14884 14560 14890 14612
rect 15654 14560 15660 14612
rect 15712 14600 15718 14612
rect 17037 14603 17095 14609
rect 17037 14600 17049 14603
rect 15712 14572 17049 14600
rect 15712 14560 15718 14572
rect 17037 14569 17049 14572
rect 17083 14569 17095 14603
rect 17037 14563 17095 14569
rect 17494 14560 17500 14612
rect 17552 14600 17558 14612
rect 21910 14600 21916 14612
rect 17552 14572 21916 14600
rect 17552 14560 17558 14572
rect 21910 14560 21916 14572
rect 21968 14560 21974 14612
rect 11790 14492 11796 14544
rect 11848 14532 11854 14544
rect 13814 14532 13820 14544
rect 11848 14504 13820 14532
rect 11848 14492 11854 14504
rect 13814 14492 13820 14504
rect 13872 14492 13878 14544
rect 19886 14492 19892 14544
rect 19944 14532 19950 14544
rect 20257 14535 20315 14541
rect 20257 14532 20269 14535
rect 19944 14504 20269 14532
rect 19944 14492 19950 14504
rect 20257 14501 20269 14504
rect 20303 14501 20315 14535
rect 20257 14495 20315 14501
rect 10045 14467 10103 14473
rect 10045 14433 10057 14467
rect 10091 14464 10103 14467
rect 10870 14464 10876 14476
rect 10091 14436 10876 14464
rect 10091 14433 10103 14436
rect 10045 14427 10103 14433
rect 10870 14424 10876 14436
rect 10928 14424 10934 14476
rect 11330 14424 11336 14476
rect 11388 14464 11394 14476
rect 12161 14467 12219 14473
rect 12161 14464 12173 14467
rect 11388 14436 12173 14464
rect 11388 14424 11394 14436
rect 7929 14399 7987 14405
rect 7929 14365 7941 14399
rect 7975 14396 7987 14399
rect 9950 14396 9956 14408
rect 7975 14368 9956 14396
rect 7975 14365 7987 14368
rect 7929 14359 7987 14365
rect 9950 14356 9956 14368
rect 10008 14356 10014 14408
rect 11440 14382 11468 14436
rect 12161 14433 12173 14436
rect 12207 14464 12219 14467
rect 12345 14467 12403 14473
rect 12345 14464 12357 14467
rect 12207 14436 12357 14464
rect 12207 14433 12219 14436
rect 12161 14427 12219 14433
rect 12345 14433 12357 14436
rect 12391 14433 12403 14467
rect 12345 14427 12403 14433
rect 13538 14424 13544 14476
rect 13596 14424 13602 14476
rect 17954 14424 17960 14476
rect 18012 14464 18018 14476
rect 19429 14467 19487 14473
rect 19429 14464 19441 14467
rect 18012 14436 19441 14464
rect 18012 14424 18018 14436
rect 19429 14433 19441 14436
rect 19475 14433 19487 14467
rect 19429 14427 19487 14433
rect 21269 14467 21327 14473
rect 21269 14433 21281 14467
rect 21315 14464 21327 14467
rect 22278 14464 22284 14476
rect 21315 14436 22284 14464
rect 21315 14433 21327 14436
rect 21269 14427 21327 14433
rect 22278 14424 22284 14436
rect 22336 14424 22342 14476
rect 13357 14399 13415 14405
rect 13357 14365 13369 14399
rect 13403 14396 13415 14399
rect 15102 14396 15108 14408
rect 13403 14368 15108 14396
rect 13403 14365 13415 14368
rect 13357 14359 13415 14365
rect 15102 14356 15108 14368
rect 15160 14356 15166 14408
rect 15194 14356 15200 14408
rect 15252 14396 15258 14408
rect 15289 14399 15347 14405
rect 15289 14396 15301 14399
rect 15252 14368 15301 14396
rect 15252 14356 15258 14368
rect 15289 14365 15301 14368
rect 15335 14365 15347 14399
rect 15289 14359 15347 14365
rect 17310 14356 17316 14408
rect 17368 14396 17374 14408
rect 17589 14399 17647 14405
rect 17589 14396 17601 14399
rect 17368 14368 17601 14396
rect 17368 14356 17374 14368
rect 17589 14365 17601 14368
rect 17635 14365 17647 14399
rect 17589 14359 17647 14365
rect 18414 14356 18420 14408
rect 18472 14396 18478 14408
rect 18877 14399 18935 14405
rect 18877 14396 18889 14399
rect 18472 14368 18889 14396
rect 18472 14356 18478 14368
rect 18877 14365 18889 14368
rect 18923 14365 18935 14399
rect 18877 14359 18935 14365
rect 20898 14356 20904 14408
rect 20956 14396 20962 14408
rect 20993 14399 21051 14405
rect 20993 14396 21005 14399
rect 20956 14368 21005 14396
rect 20956 14356 20962 14368
rect 20993 14365 21005 14368
rect 21039 14365 21051 14399
rect 20993 14359 21051 14365
rect 9674 14288 9680 14340
rect 9732 14328 9738 14340
rect 10321 14331 10379 14337
rect 10321 14328 10333 14331
rect 9732 14300 10333 14328
rect 9732 14288 9738 14300
rect 10321 14297 10333 14300
rect 10367 14297 10379 14331
rect 10321 14291 10379 14297
rect 12710 14288 12716 14340
rect 12768 14328 12774 14340
rect 13630 14328 13636 14340
rect 12768 14300 13636 14328
rect 12768 14288 12774 14300
rect 13630 14288 13636 14300
rect 13688 14288 13694 14340
rect 14369 14331 14427 14337
rect 14369 14297 14381 14331
rect 14415 14328 14427 14331
rect 14826 14328 14832 14340
rect 14415 14300 14832 14328
rect 14415 14297 14427 14300
rect 14369 14291 14427 14297
rect 14826 14288 14832 14300
rect 14884 14288 14890 14340
rect 15562 14288 15568 14340
rect 15620 14288 15626 14340
rect 17034 14328 17040 14340
rect 16790 14300 17040 14328
rect 17034 14288 17040 14300
rect 17092 14328 17098 14340
rect 17494 14328 17500 14340
rect 17092 14300 17500 14328
rect 17092 14288 17098 14300
rect 17494 14288 17500 14300
rect 17552 14288 17558 14340
rect 18601 14331 18659 14337
rect 18601 14297 18613 14331
rect 18647 14328 18659 14331
rect 18782 14328 18788 14340
rect 18647 14300 18788 14328
rect 18647 14297 18659 14300
rect 18601 14291 18659 14297
rect 18782 14288 18788 14300
rect 18840 14288 18846 14340
rect 22646 14328 22652 14340
rect 22494 14300 22652 14328
rect 22646 14288 22652 14300
rect 22704 14328 22710 14340
rect 23017 14331 23075 14337
rect 23017 14328 23029 14331
rect 22704 14300 23029 14328
rect 22704 14288 22710 14300
rect 23017 14297 23029 14300
rect 23063 14297 23075 14331
rect 23017 14291 23075 14297
rect 8662 14220 8668 14272
rect 8720 14260 8726 14272
rect 11606 14260 11612 14272
rect 8720 14232 11612 14260
rect 8720 14220 8726 14232
rect 11606 14220 11612 14232
rect 11664 14260 11670 14272
rect 11793 14263 11851 14269
rect 11793 14260 11805 14263
rect 11664 14232 11805 14260
rect 11664 14220 11670 14232
rect 11793 14229 11805 14232
rect 11839 14229 11851 14263
rect 11793 14223 11851 14229
rect 13446 14220 13452 14272
rect 13504 14220 13510 14272
rect 13814 14220 13820 14272
rect 13872 14260 13878 14272
rect 14461 14263 14519 14269
rect 14461 14260 14473 14263
rect 13872 14232 14473 14260
rect 13872 14220 13878 14232
rect 14461 14229 14473 14232
rect 14507 14229 14519 14263
rect 14461 14223 14519 14229
rect 17678 14220 17684 14272
rect 17736 14220 17742 14272
rect 22094 14220 22100 14272
rect 22152 14260 22158 14272
rect 22741 14263 22799 14269
rect 22741 14260 22753 14263
rect 22152 14232 22753 14260
rect 22152 14220 22158 14232
rect 22741 14229 22753 14232
rect 22787 14229 22799 14263
rect 22741 14223 22799 14229
rect 1104 14170 25852 14192
rect 1104 14118 7950 14170
rect 8002 14118 8014 14170
rect 8066 14118 8078 14170
rect 8130 14118 8142 14170
rect 8194 14118 8206 14170
rect 8258 14118 17950 14170
rect 18002 14118 18014 14170
rect 18066 14118 18078 14170
rect 18130 14118 18142 14170
rect 18194 14118 18206 14170
rect 18258 14118 25852 14170
rect 1104 14096 25852 14118
rect 9861 14059 9919 14065
rect 9861 14025 9873 14059
rect 9907 14056 9919 14059
rect 9950 14056 9956 14068
rect 9907 14028 9956 14056
rect 9907 14025 9919 14028
rect 9861 14019 9919 14025
rect 9950 14016 9956 14028
rect 10008 14016 10014 14068
rect 10229 14059 10287 14065
rect 10229 14025 10241 14059
rect 10275 14056 10287 14059
rect 11330 14056 11336 14068
rect 10275 14028 11336 14056
rect 10275 14025 10287 14028
rect 10229 14019 10287 14025
rect 10244 13988 10272 14019
rect 11330 14016 11336 14028
rect 11388 14016 11394 14068
rect 11698 14016 11704 14068
rect 11756 14056 11762 14068
rect 12069 14059 12127 14065
rect 12069 14056 12081 14059
rect 11756 14028 12081 14056
rect 11756 14016 11762 14028
rect 12069 14025 12081 14028
rect 12115 14025 12127 14059
rect 12069 14019 12127 14025
rect 12437 14059 12495 14065
rect 12437 14025 12449 14059
rect 12483 14025 12495 14059
rect 12437 14019 12495 14025
rect 9614 13960 10272 13988
rect 1762 13880 1768 13932
rect 1820 13880 1826 13932
rect 12084 13920 12112 14019
rect 12452 13988 12480 14019
rect 12526 14016 12532 14068
rect 12584 14056 12590 14068
rect 12894 14056 12900 14068
rect 12584 14028 12900 14056
rect 12584 14016 12590 14028
rect 12894 14016 12900 14028
rect 12952 14016 12958 14068
rect 13354 14016 13360 14068
rect 13412 14056 13418 14068
rect 13817 14059 13875 14065
rect 13817 14056 13829 14059
rect 13412 14028 13829 14056
rect 13412 14016 13418 14028
rect 13817 14025 13829 14028
rect 13863 14025 13875 14059
rect 13817 14019 13875 14025
rect 14918 14016 14924 14068
rect 14976 14016 14982 14068
rect 15562 14016 15568 14068
rect 15620 14056 15626 14068
rect 17497 14059 17555 14065
rect 17497 14056 17509 14059
rect 15620 14028 17509 14056
rect 15620 14016 15626 14028
rect 17497 14025 17509 14028
rect 17543 14025 17555 14059
rect 17497 14019 17555 14025
rect 19150 14016 19156 14068
rect 19208 14016 19214 14068
rect 20073 14059 20131 14065
rect 20073 14025 20085 14059
rect 20119 14056 20131 14059
rect 21910 14056 21916 14068
rect 20119 14028 21916 14056
rect 20119 14025 20131 14028
rect 20073 14019 20131 14025
rect 21910 14016 21916 14028
rect 21968 14016 21974 14068
rect 22830 14016 22836 14068
rect 22888 14056 22894 14068
rect 23017 14059 23075 14065
rect 23017 14056 23029 14059
rect 22888 14028 23029 14056
rect 22888 14016 22894 14028
rect 23017 14025 23029 14028
rect 23063 14025 23075 14059
rect 23017 14019 23075 14025
rect 15654 13988 15660 14000
rect 12452 13960 15660 13988
rect 15654 13948 15660 13960
rect 15712 13948 15718 14000
rect 17310 13948 17316 14000
rect 17368 13988 17374 14000
rect 17957 13991 18015 13997
rect 17957 13988 17969 13991
rect 17368 13960 17969 13988
rect 17368 13948 17374 13960
rect 17957 13957 17969 13960
rect 18003 13957 18015 13991
rect 17957 13951 18015 13957
rect 20530 13948 20536 14000
rect 20588 13948 20594 14000
rect 25130 13948 25136 14000
rect 25188 13948 25194 14000
rect 12805 13923 12863 13929
rect 12805 13920 12817 13923
rect 12084 13892 12817 13920
rect 12805 13889 12817 13892
rect 12851 13889 12863 13923
rect 12805 13883 12863 13889
rect 12894 13880 12900 13932
rect 12952 13920 12958 13932
rect 13449 13923 13507 13929
rect 13449 13920 13461 13923
rect 12952 13892 13461 13920
rect 12952 13880 12958 13892
rect 13449 13889 13461 13892
rect 13495 13889 13507 13923
rect 13449 13883 13507 13889
rect 14369 13923 14427 13929
rect 14369 13889 14381 13923
rect 14415 13920 14427 13923
rect 14918 13920 14924 13932
rect 14415 13892 14924 13920
rect 14415 13889 14427 13892
rect 14369 13883 14427 13889
rect 1302 13812 1308 13864
rect 1360 13852 1366 13864
rect 2041 13855 2099 13861
rect 2041 13852 2053 13855
rect 1360 13824 2053 13852
rect 1360 13812 1366 13824
rect 2041 13821 2053 13824
rect 2087 13821 2099 13855
rect 2041 13815 2099 13821
rect 5258 13812 5264 13864
rect 5316 13852 5322 13864
rect 6730 13852 6736 13864
rect 5316 13824 6736 13852
rect 5316 13812 5322 13824
rect 6730 13812 6736 13824
rect 6788 13852 6794 13864
rect 8113 13855 8171 13861
rect 8113 13852 8125 13855
rect 6788 13824 8125 13852
rect 6788 13812 6794 13824
rect 8113 13821 8125 13824
rect 8159 13852 8171 13855
rect 8389 13855 8447 13861
rect 8159 13824 8248 13852
rect 8159 13821 8171 13824
rect 8113 13815 8171 13821
rect 8220 13716 8248 13824
rect 8389 13821 8401 13855
rect 8435 13852 8447 13855
rect 8478 13852 8484 13864
rect 8435 13824 8484 13852
rect 8435 13821 8447 13824
rect 8389 13815 8447 13821
rect 8478 13812 8484 13824
rect 8536 13812 8542 13864
rect 12989 13855 13047 13861
rect 12989 13821 13001 13855
rect 13035 13821 13047 13855
rect 13464 13852 13492 13883
rect 14918 13880 14924 13892
rect 14976 13880 14982 13932
rect 16301 13923 16359 13929
rect 15488 13892 16252 13920
rect 14553 13855 14611 13861
rect 13464 13824 14504 13852
rect 12989 13815 13047 13821
rect 11698 13744 11704 13796
rect 11756 13784 11762 13796
rect 13004 13784 13032 13815
rect 11756 13756 13032 13784
rect 14476 13784 14504 13824
rect 14553 13821 14565 13855
rect 14599 13852 14611 13855
rect 14642 13852 14648 13864
rect 14599 13824 14648 13852
rect 14599 13821 14611 13824
rect 14553 13815 14611 13821
rect 14642 13812 14648 13824
rect 14700 13812 14706 13864
rect 15488 13852 15516 13892
rect 14752 13824 15516 13852
rect 14752 13784 14780 13824
rect 15562 13812 15568 13864
rect 15620 13852 15626 13864
rect 16224 13852 16252 13892
rect 16301 13889 16313 13923
rect 16347 13920 16359 13923
rect 16574 13920 16580 13932
rect 16347 13892 16580 13920
rect 16347 13889 16359 13892
rect 16301 13883 16359 13889
rect 16574 13880 16580 13892
rect 16632 13880 16638 13932
rect 16853 13923 16911 13929
rect 16853 13889 16865 13923
rect 16899 13920 16911 13923
rect 17034 13920 17040 13932
rect 16899 13892 17040 13920
rect 16899 13889 16911 13892
rect 16853 13883 16911 13889
rect 17034 13880 17040 13892
rect 17092 13880 17098 13932
rect 18509 13923 18567 13929
rect 18509 13889 18521 13923
rect 18555 13920 18567 13923
rect 18874 13920 18880 13932
rect 18555 13892 18880 13920
rect 18555 13889 18567 13892
rect 18509 13883 18567 13889
rect 18874 13880 18880 13892
rect 18932 13880 18938 13932
rect 20441 13923 20499 13929
rect 20441 13889 20453 13923
rect 20487 13920 20499 13923
rect 21269 13923 21327 13929
rect 21269 13920 21281 13923
rect 20487 13892 21281 13920
rect 20487 13889 20499 13892
rect 20441 13883 20499 13889
rect 21269 13889 21281 13892
rect 21315 13889 21327 13923
rect 21269 13883 21327 13889
rect 22554 13880 22560 13932
rect 22612 13920 22618 13932
rect 23201 13923 23259 13929
rect 23201 13920 23213 13923
rect 22612 13892 23213 13920
rect 22612 13880 22618 13892
rect 23201 13889 23213 13892
rect 23247 13889 23259 13923
rect 23201 13883 23259 13889
rect 23842 13880 23848 13932
rect 23900 13920 23906 13932
rect 23937 13923 23995 13929
rect 23937 13920 23949 13923
rect 23900 13892 23949 13920
rect 23900 13880 23906 13892
rect 23937 13889 23949 13892
rect 23983 13889 23995 13923
rect 23937 13883 23995 13889
rect 18138 13852 18144 13864
rect 15620 13824 16160 13852
rect 16224 13824 18144 13852
rect 15620 13812 15626 13824
rect 16132 13793 16160 13824
rect 18138 13812 18144 13824
rect 18196 13812 18202 13864
rect 19058 13812 19064 13864
rect 19116 13852 19122 13864
rect 19242 13852 19248 13864
rect 19116 13824 19248 13852
rect 19116 13812 19122 13824
rect 19242 13812 19248 13824
rect 19300 13812 19306 13864
rect 19426 13812 19432 13864
rect 19484 13852 19490 13864
rect 20254 13852 20260 13864
rect 19484 13824 20260 13852
rect 19484 13812 19490 13824
rect 20254 13812 20260 13824
rect 20312 13812 20318 13864
rect 20622 13812 20628 13864
rect 20680 13812 20686 13864
rect 14476 13756 14780 13784
rect 16117 13787 16175 13793
rect 11756 13744 11762 13756
rect 16117 13753 16129 13787
rect 16163 13753 16175 13787
rect 16117 13747 16175 13753
rect 8386 13716 8392 13728
rect 8220 13688 8392 13716
rect 8386 13676 8392 13688
rect 8444 13716 8450 13728
rect 8846 13716 8852 13728
rect 8444 13688 8852 13716
rect 8444 13676 8450 13688
rect 8846 13676 8852 13688
rect 8904 13676 8910 13728
rect 17494 13676 17500 13728
rect 17552 13716 17558 13728
rect 17773 13719 17831 13725
rect 17773 13716 17785 13719
rect 17552 13688 17785 13716
rect 17552 13676 17558 13688
rect 17773 13685 17785 13688
rect 17819 13685 17831 13719
rect 17773 13679 17831 13685
rect 1104 13626 25852 13648
rect 1104 13574 2950 13626
rect 3002 13574 3014 13626
rect 3066 13574 3078 13626
rect 3130 13574 3142 13626
rect 3194 13574 3206 13626
rect 3258 13574 12950 13626
rect 13002 13574 13014 13626
rect 13066 13574 13078 13626
rect 13130 13574 13142 13626
rect 13194 13574 13206 13626
rect 13258 13574 22950 13626
rect 23002 13574 23014 13626
rect 23066 13574 23078 13626
rect 23130 13574 23142 13626
rect 23194 13574 23206 13626
rect 23258 13574 25852 13626
rect 1104 13552 25852 13574
rect 8478 13472 8484 13524
rect 8536 13512 8542 13524
rect 12253 13515 12311 13521
rect 12253 13512 12265 13515
rect 8536 13484 12265 13512
rect 8536 13472 8542 13484
rect 12253 13481 12265 13484
rect 12299 13481 12311 13515
rect 12253 13475 12311 13481
rect 17681 13515 17739 13521
rect 17681 13481 17693 13515
rect 17727 13512 17739 13515
rect 19610 13512 19616 13524
rect 17727 13484 19616 13512
rect 17727 13481 17739 13484
rect 17681 13475 17739 13481
rect 19610 13472 19616 13484
rect 19668 13472 19674 13524
rect 16485 13447 16543 13453
rect 16485 13413 16497 13447
rect 16531 13444 16543 13447
rect 17770 13444 17776 13456
rect 16531 13416 17776 13444
rect 16531 13413 16543 13416
rect 16485 13407 16543 13413
rect 17770 13404 17776 13416
rect 17828 13404 17834 13456
rect 18785 13447 18843 13453
rect 18785 13444 18797 13447
rect 18156 13416 18797 13444
rect 18156 13388 18184 13416
rect 18785 13413 18797 13416
rect 18831 13413 18843 13447
rect 18785 13407 18843 13413
rect 20806 13404 20812 13456
rect 20864 13444 20870 13456
rect 20864 13416 22692 13444
rect 20864 13404 20870 13416
rect 10502 13336 10508 13388
rect 10560 13376 10566 13388
rect 10781 13379 10839 13385
rect 10781 13376 10793 13379
rect 10560 13348 10793 13376
rect 10560 13336 10566 13348
rect 10781 13345 10793 13348
rect 10827 13345 10839 13379
rect 10781 13339 10839 13345
rect 10962 13336 10968 13388
rect 11020 13336 11026 13388
rect 13538 13376 13544 13388
rect 11624 13348 13544 13376
rect 11624 13317 11652 13348
rect 13538 13336 13544 13348
rect 13596 13336 13602 13388
rect 13998 13336 14004 13388
rect 14056 13376 14062 13388
rect 14056 13348 16068 13376
rect 14056 13336 14062 13348
rect 11609 13311 11667 13317
rect 11609 13277 11621 13311
rect 11655 13277 11667 13311
rect 11609 13271 11667 13277
rect 14274 13268 14280 13320
rect 14332 13268 14338 13320
rect 15378 13268 15384 13320
rect 15436 13308 15442 13320
rect 15473 13311 15531 13317
rect 15473 13308 15485 13311
rect 15436 13280 15485 13308
rect 15436 13268 15442 13280
rect 15473 13277 15485 13280
rect 15519 13308 15531 13311
rect 15933 13311 15991 13317
rect 15933 13308 15945 13311
rect 15519 13280 15945 13308
rect 15519 13277 15531 13280
rect 15473 13271 15531 13277
rect 15933 13277 15945 13280
rect 15979 13277 15991 13311
rect 16040 13308 16068 13348
rect 16206 13336 16212 13388
rect 16264 13376 16270 13388
rect 16945 13379 17003 13385
rect 16945 13376 16957 13379
rect 16264 13348 16957 13376
rect 16264 13336 16270 13348
rect 16945 13345 16957 13348
rect 16991 13345 17003 13379
rect 16945 13339 17003 13345
rect 17034 13336 17040 13388
rect 17092 13336 17098 13388
rect 18138 13336 18144 13388
rect 18196 13336 18202 13388
rect 18325 13379 18383 13385
rect 18325 13345 18337 13379
rect 18371 13376 18383 13379
rect 18690 13376 18696 13388
rect 18371 13348 18696 13376
rect 18371 13345 18383 13348
rect 18325 13339 18383 13345
rect 18690 13336 18696 13348
rect 18748 13336 18754 13388
rect 19702 13336 19708 13388
rect 19760 13336 19766 13388
rect 19978 13336 19984 13388
rect 20036 13376 20042 13388
rect 20036 13348 20300 13376
rect 20036 13336 20042 13348
rect 19334 13308 19340 13320
rect 16040 13280 19340 13308
rect 15933 13271 15991 13277
rect 19334 13268 19340 13280
rect 19392 13268 19398 13320
rect 19521 13311 19579 13317
rect 19521 13277 19533 13311
rect 19567 13308 19579 13311
rect 19720 13308 19748 13336
rect 19886 13308 19892 13320
rect 19567 13280 19892 13308
rect 19567 13277 19579 13280
rect 19521 13271 19579 13277
rect 19886 13268 19892 13280
rect 19944 13268 19950 13320
rect 20272 13317 20300 13348
rect 20257 13311 20315 13317
rect 20257 13277 20269 13311
rect 20303 13308 20315 13311
rect 20717 13311 20775 13317
rect 20717 13308 20729 13311
rect 20303 13280 20729 13308
rect 20303 13277 20315 13280
rect 20257 13271 20315 13277
rect 20717 13277 20729 13280
rect 20763 13277 20775 13311
rect 20717 13271 20775 13277
rect 21085 13311 21143 13317
rect 21085 13277 21097 13311
rect 21131 13308 21143 13311
rect 22094 13308 22100 13320
rect 21131 13280 22100 13308
rect 21131 13277 21143 13280
rect 21085 13271 21143 13277
rect 22094 13268 22100 13280
rect 22152 13268 22158 13320
rect 22664 13317 22692 13416
rect 22649 13311 22707 13317
rect 22649 13277 22661 13311
rect 22695 13277 22707 13311
rect 22649 13271 22707 13277
rect 7098 13200 7104 13252
rect 7156 13240 7162 13252
rect 10689 13243 10747 13249
rect 10689 13240 10701 13243
rect 7156 13212 10701 13240
rect 7156 13200 7162 13212
rect 10689 13209 10701 13212
rect 10735 13209 10747 13243
rect 10689 13203 10747 13209
rect 13354 13200 13360 13252
rect 13412 13240 13418 13252
rect 13541 13243 13599 13249
rect 13541 13240 13553 13243
rect 13412 13212 13553 13240
rect 13412 13200 13418 13212
rect 13541 13209 13553 13212
rect 13587 13209 13599 13243
rect 13541 13203 13599 13209
rect 15657 13243 15715 13249
rect 15657 13209 15669 13243
rect 15703 13240 15715 13243
rect 16298 13240 16304 13252
rect 15703 13212 16304 13240
rect 15703 13209 15715 13212
rect 15657 13203 15715 13209
rect 16298 13200 16304 13212
rect 16356 13200 16362 13252
rect 18049 13243 18107 13249
rect 18049 13209 18061 13243
rect 18095 13240 18107 13243
rect 18414 13240 18420 13252
rect 18095 13212 18420 13240
rect 18095 13209 18107 13212
rect 18049 13203 18107 13209
rect 18414 13200 18420 13212
rect 18472 13200 18478 13252
rect 19705 13243 19763 13249
rect 19705 13209 19717 13243
rect 19751 13240 19763 13243
rect 19978 13240 19984 13252
rect 19751 13212 19984 13240
rect 19751 13209 19763 13212
rect 19705 13203 19763 13209
rect 19978 13200 19984 13212
rect 20036 13200 20042 13252
rect 20441 13243 20499 13249
rect 20441 13209 20453 13243
rect 20487 13240 20499 13243
rect 20530 13240 20536 13252
rect 20487 13212 20536 13240
rect 20487 13209 20499 13212
rect 20441 13203 20499 13209
rect 20530 13200 20536 13212
rect 20588 13200 20594 13252
rect 23845 13243 23903 13249
rect 23845 13209 23857 13243
rect 23891 13240 23903 13243
rect 24946 13240 24952 13252
rect 23891 13212 24952 13240
rect 23891 13209 23903 13212
rect 23845 13203 23903 13209
rect 24946 13200 24952 13212
rect 25004 13200 25010 13252
rect 10321 13175 10379 13181
rect 10321 13141 10333 13175
rect 10367 13172 10379 13175
rect 12342 13172 12348 13184
rect 10367 13144 12348 13172
rect 10367 13141 10379 13144
rect 10321 13135 10379 13141
rect 12342 13132 12348 13144
rect 12400 13132 12406 13184
rect 13630 13132 13636 13184
rect 13688 13132 13694 13184
rect 14918 13132 14924 13184
rect 14976 13132 14982 13184
rect 16850 13132 16856 13184
rect 16908 13132 16914 13184
rect 20806 13132 20812 13184
rect 20864 13172 20870 13184
rect 21729 13175 21787 13181
rect 21729 13172 21741 13175
rect 20864 13144 21741 13172
rect 20864 13132 20870 13144
rect 21729 13141 21741 13144
rect 21775 13141 21787 13175
rect 21729 13135 21787 13141
rect 1104 13082 25852 13104
rect 1104 13030 7950 13082
rect 8002 13030 8014 13082
rect 8066 13030 8078 13082
rect 8130 13030 8142 13082
rect 8194 13030 8206 13082
rect 8258 13030 17950 13082
rect 18002 13030 18014 13082
rect 18066 13030 18078 13082
rect 18130 13030 18142 13082
rect 18194 13030 18206 13082
rect 18258 13030 25852 13082
rect 1104 13008 25852 13030
rect 10597 12971 10655 12977
rect 10597 12937 10609 12971
rect 10643 12968 10655 12971
rect 10962 12968 10968 12980
rect 10643 12940 10968 12968
rect 10643 12937 10655 12940
rect 10597 12931 10655 12937
rect 10962 12928 10968 12940
rect 11020 12928 11026 12980
rect 12802 12928 12808 12980
rect 12860 12968 12866 12980
rect 13357 12971 13415 12977
rect 13357 12968 13369 12971
rect 12860 12940 13369 12968
rect 12860 12928 12866 12940
rect 13357 12937 13369 12940
rect 13403 12937 13415 12971
rect 13817 12971 13875 12977
rect 13817 12968 13829 12971
rect 13357 12931 13415 12937
rect 13648 12940 13829 12968
rect 9122 12860 9128 12912
rect 9180 12860 9186 12912
rect 13081 12903 13139 12909
rect 13081 12900 13093 12903
rect 12406 12872 13093 12900
rect 4982 12792 4988 12844
rect 5040 12832 5046 12844
rect 8754 12832 8760 12844
rect 5040 12804 8760 12832
rect 5040 12792 5046 12804
rect 8754 12792 8760 12804
rect 8812 12792 8818 12844
rect 10258 12804 10364 12832
rect 10336 12776 10364 12804
rect 11698 12792 11704 12844
rect 11756 12792 11762 12844
rect 8846 12724 8852 12776
rect 8904 12764 8910 12776
rect 9582 12764 9588 12776
rect 8904 12736 9588 12764
rect 8904 12724 8910 12736
rect 9582 12724 9588 12736
rect 9640 12724 9646 12776
rect 10318 12724 10324 12776
rect 10376 12764 10382 12776
rect 10873 12767 10931 12773
rect 10873 12764 10885 12767
rect 10376 12736 10885 12764
rect 10376 12724 10382 12736
rect 10873 12733 10885 12736
rect 10919 12733 10931 12767
rect 10873 12727 10931 12733
rect 11882 12656 11888 12708
rect 11940 12696 11946 12708
rect 12406 12696 12434 12872
rect 13081 12869 13093 12872
rect 13127 12900 13139 12903
rect 13648 12900 13676 12940
rect 13817 12937 13829 12940
rect 13863 12968 13875 12971
rect 13998 12968 14004 12980
rect 13863 12940 14004 12968
rect 13863 12937 13875 12940
rect 13817 12931 13875 12937
rect 13998 12928 14004 12940
rect 14056 12928 14062 12980
rect 15194 12968 15200 12980
rect 14568 12940 15200 12968
rect 13127 12872 13676 12900
rect 13127 12869 13139 12872
rect 13081 12863 13139 12869
rect 14568 12841 14596 12940
rect 15194 12928 15200 12940
rect 15252 12968 15258 12980
rect 18322 12968 18328 12980
rect 15252 12940 18328 12968
rect 15252 12928 15258 12940
rect 15286 12860 15292 12912
rect 15344 12860 15350 12912
rect 16850 12860 16856 12912
rect 16908 12900 16914 12912
rect 16945 12903 17003 12909
rect 16945 12900 16957 12903
rect 16908 12872 16957 12900
rect 16908 12860 16914 12872
rect 16945 12869 16957 12872
rect 16991 12869 17003 12903
rect 16945 12863 17003 12869
rect 17880 12841 17908 12940
rect 18322 12928 18328 12940
rect 18380 12928 18386 12980
rect 18874 12928 18880 12980
rect 18932 12968 18938 12980
rect 19613 12971 19671 12977
rect 19613 12968 19625 12971
rect 18932 12940 19625 12968
rect 18932 12928 18938 12940
rect 19613 12937 19625 12940
rect 19659 12937 19671 12971
rect 19613 12931 19671 12937
rect 19886 12928 19892 12980
rect 19944 12928 19950 12980
rect 21174 12928 21180 12980
rect 21232 12928 21238 12980
rect 20346 12900 20352 12912
rect 19366 12872 20352 12900
rect 20346 12860 20352 12872
rect 20404 12860 20410 12912
rect 21085 12903 21143 12909
rect 21085 12869 21097 12903
rect 21131 12900 21143 12903
rect 22741 12903 22799 12909
rect 22741 12900 22753 12903
rect 21131 12872 22753 12900
rect 21131 12869 21143 12872
rect 21085 12863 21143 12869
rect 22741 12869 22753 12872
rect 22787 12869 22799 12903
rect 22741 12863 22799 12869
rect 13725 12835 13783 12841
rect 13725 12801 13737 12835
rect 13771 12832 13783 12835
rect 14553 12835 14611 12841
rect 13771 12804 14504 12832
rect 13771 12801 13783 12804
rect 13725 12795 13783 12801
rect 13909 12767 13967 12773
rect 13909 12764 13921 12767
rect 13740 12736 13921 12764
rect 13740 12708 13768 12736
rect 13909 12733 13921 12736
rect 13955 12764 13967 12767
rect 14182 12764 14188 12776
rect 13955 12736 14188 12764
rect 13955 12733 13967 12736
rect 13909 12727 13967 12733
rect 14182 12724 14188 12736
rect 14240 12724 14246 12776
rect 11940 12668 12434 12696
rect 11940 12656 11946 12668
rect 13722 12656 13728 12708
rect 13780 12656 13786 12708
rect 12066 12588 12072 12640
rect 12124 12628 12130 12640
rect 12345 12631 12403 12637
rect 12345 12628 12357 12631
rect 12124 12600 12357 12628
rect 12124 12588 12130 12600
rect 12345 12597 12357 12600
rect 12391 12597 12403 12631
rect 14476 12628 14504 12804
rect 14553 12801 14565 12835
rect 14599 12801 14611 12835
rect 14553 12795 14611 12801
rect 17865 12835 17923 12841
rect 17865 12801 17877 12835
rect 17911 12801 17923 12835
rect 17865 12795 17923 12801
rect 22097 12835 22155 12841
rect 22097 12801 22109 12835
rect 22143 12832 22155 12835
rect 22186 12832 22192 12844
rect 22143 12804 22192 12832
rect 22143 12801 22155 12804
rect 22097 12795 22155 12801
rect 22186 12792 22192 12804
rect 22244 12832 22250 12844
rect 23201 12835 23259 12841
rect 23201 12832 23213 12835
rect 22244 12804 23213 12832
rect 22244 12792 22250 12804
rect 23201 12801 23213 12804
rect 23247 12801 23259 12835
rect 23201 12795 23259 12801
rect 23382 12792 23388 12844
rect 23440 12832 23446 12844
rect 23937 12835 23995 12841
rect 23937 12832 23949 12835
rect 23440 12804 23949 12832
rect 23440 12792 23446 12804
rect 23937 12801 23949 12804
rect 23983 12801 23995 12835
rect 23937 12795 23995 12801
rect 14829 12767 14887 12773
rect 14829 12733 14841 12767
rect 14875 12764 14887 12767
rect 15470 12764 15476 12776
rect 14875 12736 15476 12764
rect 14875 12733 14887 12736
rect 14829 12727 14887 12733
rect 15470 12724 15476 12736
rect 15528 12724 15534 12776
rect 16301 12767 16359 12773
rect 16301 12733 16313 12767
rect 16347 12764 16359 12767
rect 17034 12764 17040 12776
rect 16347 12736 17040 12764
rect 16347 12733 16359 12736
rect 16301 12727 16359 12733
rect 17034 12724 17040 12736
rect 17092 12724 17098 12776
rect 18141 12767 18199 12773
rect 18141 12733 18153 12767
rect 18187 12764 18199 12767
rect 20622 12764 20628 12776
rect 18187 12736 20628 12764
rect 18187 12733 18199 12736
rect 18141 12727 18199 12733
rect 20622 12724 20628 12736
rect 20680 12724 20686 12776
rect 21361 12767 21419 12773
rect 21361 12733 21373 12767
rect 21407 12764 21419 12767
rect 22002 12764 22008 12776
rect 21407 12736 22008 12764
rect 21407 12733 21419 12736
rect 21361 12727 21419 12733
rect 22002 12724 22008 12736
rect 22060 12724 22066 12776
rect 24762 12724 24768 12776
rect 24820 12724 24826 12776
rect 15194 12628 15200 12640
rect 14476 12600 15200 12628
rect 12345 12591 12403 12597
rect 15194 12588 15200 12600
rect 15252 12628 15258 12640
rect 15378 12628 15384 12640
rect 15252 12600 15384 12628
rect 15252 12588 15258 12600
rect 15378 12588 15384 12600
rect 15436 12588 15442 12640
rect 16114 12588 16120 12640
rect 16172 12628 16178 12640
rect 17494 12628 17500 12640
rect 16172 12600 17500 12628
rect 16172 12588 16178 12600
rect 17494 12588 17500 12600
rect 17552 12628 17558 12640
rect 20165 12631 20223 12637
rect 20165 12628 20177 12631
rect 17552 12600 20177 12628
rect 17552 12588 17558 12600
rect 20165 12597 20177 12600
rect 20211 12628 20223 12631
rect 20346 12628 20352 12640
rect 20211 12600 20352 12628
rect 20211 12597 20223 12600
rect 20165 12591 20223 12597
rect 20346 12588 20352 12600
rect 20404 12588 20410 12640
rect 20714 12588 20720 12640
rect 20772 12588 20778 12640
rect 22094 12588 22100 12640
rect 22152 12628 22158 12640
rect 22189 12631 22247 12637
rect 22189 12628 22201 12631
rect 22152 12600 22201 12628
rect 22152 12588 22158 12600
rect 22189 12597 22201 12600
rect 22235 12597 22247 12631
rect 22189 12591 22247 12597
rect 1104 12538 25852 12560
rect 1104 12486 2950 12538
rect 3002 12486 3014 12538
rect 3066 12486 3078 12538
rect 3130 12486 3142 12538
rect 3194 12486 3206 12538
rect 3258 12486 12950 12538
rect 13002 12486 13014 12538
rect 13066 12486 13078 12538
rect 13130 12486 13142 12538
rect 13194 12486 13206 12538
rect 13258 12486 22950 12538
rect 23002 12486 23014 12538
rect 23066 12486 23078 12538
rect 23130 12486 23142 12538
rect 23194 12486 23206 12538
rect 23258 12486 25852 12538
rect 1104 12464 25852 12486
rect 1854 12384 1860 12436
rect 1912 12424 1918 12436
rect 9490 12424 9496 12436
rect 1912 12396 9496 12424
rect 1912 12384 1918 12396
rect 9490 12384 9496 12396
rect 9548 12384 9554 12436
rect 11333 12427 11391 12433
rect 11333 12393 11345 12427
rect 11379 12424 11391 12427
rect 11698 12424 11704 12436
rect 11379 12396 11704 12424
rect 11379 12393 11391 12396
rect 11333 12387 11391 12393
rect 11698 12384 11704 12396
rect 11756 12384 11762 12436
rect 13446 12384 13452 12436
rect 13504 12424 13510 12436
rect 15197 12427 15255 12433
rect 15197 12424 15209 12427
rect 13504 12396 15209 12424
rect 13504 12384 13510 12396
rect 15197 12393 15209 12396
rect 15243 12393 15255 12427
rect 15197 12387 15255 12393
rect 16206 12384 16212 12436
rect 16264 12424 16270 12436
rect 16393 12427 16451 12433
rect 16393 12424 16405 12427
rect 16264 12396 16405 12424
rect 16264 12384 16270 12396
rect 16393 12393 16405 12396
rect 16439 12393 16451 12427
rect 21361 12427 21419 12433
rect 21361 12424 21373 12427
rect 16393 12387 16451 12393
rect 19168 12396 21373 12424
rect 14182 12316 14188 12368
rect 14240 12356 14246 12368
rect 14240 12328 15148 12356
rect 14240 12316 14246 12328
rect 9582 12248 9588 12300
rect 9640 12248 9646 12300
rect 10870 12248 10876 12300
rect 10928 12288 10934 12300
rect 10928 12260 11100 12288
rect 10928 12248 10934 12260
rect 11072 12220 11100 12260
rect 12066 12248 12072 12300
rect 12124 12248 12130 12300
rect 13541 12291 13599 12297
rect 13541 12257 13553 12291
rect 13587 12288 13599 12291
rect 14274 12288 14280 12300
rect 13587 12260 14280 12288
rect 13587 12257 13599 12260
rect 13541 12251 13599 12257
rect 14274 12248 14280 12260
rect 14332 12288 14338 12300
rect 15010 12288 15016 12300
rect 14332 12260 15016 12288
rect 14332 12248 14338 12260
rect 15010 12248 15016 12260
rect 15068 12248 15074 12300
rect 11790 12220 11796 12232
rect 11072 12192 11796 12220
rect 11790 12180 11796 12192
rect 11848 12180 11854 12232
rect 14366 12180 14372 12232
rect 14424 12220 14430 12232
rect 14829 12223 14887 12229
rect 14829 12220 14841 12223
rect 14424 12192 14841 12220
rect 14424 12180 14430 12192
rect 14829 12189 14841 12192
rect 14875 12189 14887 12223
rect 15120 12220 15148 12328
rect 15746 12316 15752 12368
rect 15804 12356 15810 12368
rect 18414 12356 18420 12368
rect 15804 12328 18420 12356
rect 15804 12316 15810 12328
rect 18414 12316 18420 12328
rect 18472 12316 18478 12368
rect 15841 12291 15899 12297
rect 15841 12257 15853 12291
rect 15887 12288 15899 12291
rect 16022 12288 16028 12300
rect 15887 12260 16028 12288
rect 15887 12257 15899 12260
rect 15841 12251 15899 12257
rect 16022 12248 16028 12260
rect 16080 12248 16086 12300
rect 16945 12291 17003 12297
rect 16945 12288 16957 12291
rect 16546 12260 16957 12288
rect 16546 12220 16574 12260
rect 16945 12257 16957 12260
rect 16991 12257 17003 12291
rect 16945 12251 17003 12257
rect 15120 12192 16574 12220
rect 18233 12223 18291 12229
rect 14829 12183 14887 12189
rect 18233 12189 18245 12223
rect 18279 12220 18291 12223
rect 18690 12220 18696 12232
rect 18279 12192 18696 12220
rect 18279 12189 18291 12192
rect 18233 12183 18291 12189
rect 18690 12180 18696 12192
rect 18748 12220 18754 12232
rect 19168 12220 19196 12396
rect 21361 12393 21373 12396
rect 21407 12393 21419 12427
rect 21361 12387 21419 12393
rect 22649 12359 22707 12365
rect 22649 12325 22661 12359
rect 22695 12356 22707 12359
rect 24854 12356 24860 12368
rect 22695 12328 24860 12356
rect 22695 12325 22707 12328
rect 22649 12319 22707 12325
rect 24854 12316 24860 12328
rect 24912 12316 24918 12368
rect 19613 12291 19671 12297
rect 19613 12257 19625 12291
rect 19659 12288 19671 12291
rect 20898 12288 20904 12300
rect 19659 12260 20904 12288
rect 19659 12257 19671 12260
rect 19613 12251 19671 12257
rect 20898 12248 20904 12260
rect 20956 12248 20962 12300
rect 21542 12248 21548 12300
rect 21600 12288 21606 12300
rect 21600 12260 22876 12288
rect 21600 12248 21606 12260
rect 18748 12192 19196 12220
rect 18748 12180 18754 12192
rect 21818 12180 21824 12232
rect 21876 12220 21882 12232
rect 22848 12229 22876 12260
rect 22005 12223 22063 12229
rect 22005 12220 22017 12223
rect 21876 12192 22017 12220
rect 21876 12180 21882 12192
rect 22005 12189 22017 12192
rect 22051 12189 22063 12223
rect 22005 12183 22063 12189
rect 22833 12223 22891 12229
rect 22833 12189 22845 12223
rect 22879 12189 22891 12223
rect 22833 12183 22891 12189
rect 23474 12180 23480 12232
rect 23532 12180 23538 12232
rect 9858 12112 9864 12164
rect 9916 12112 9922 12164
rect 10318 12152 10324 12164
rect 10244 12124 10324 12152
rect 2774 12044 2780 12096
rect 2832 12084 2838 12096
rect 5166 12084 5172 12096
rect 2832 12056 5172 12084
rect 2832 12044 2838 12056
rect 5166 12044 5172 12056
rect 5224 12044 5230 12096
rect 10244 12084 10272 12124
rect 10318 12112 10324 12124
rect 10376 12112 10382 12164
rect 15286 12152 15292 12164
rect 12452 12124 12558 12152
rect 13832 12124 15292 12152
rect 12452 12084 12480 12124
rect 13722 12084 13728 12096
rect 10244 12056 13728 12084
rect 13722 12044 13728 12056
rect 13780 12084 13786 12096
rect 13832 12093 13860 12124
rect 15286 12112 15292 12124
rect 15344 12152 15350 12164
rect 16206 12152 16212 12164
rect 15344 12124 16212 12152
rect 15344 12112 15350 12124
rect 16206 12112 16212 12124
rect 16264 12112 16270 12164
rect 16761 12155 16819 12161
rect 16761 12121 16773 12155
rect 16807 12152 16819 12155
rect 19518 12152 19524 12164
rect 16807 12124 19524 12152
rect 16807 12121 16819 12124
rect 16761 12115 16819 12121
rect 19518 12112 19524 12124
rect 19576 12152 19582 12164
rect 19794 12152 19800 12164
rect 19576 12124 19800 12152
rect 19576 12112 19582 12124
rect 19794 12112 19800 12124
rect 19852 12112 19858 12164
rect 19889 12155 19947 12161
rect 19889 12121 19901 12155
rect 19935 12121 19947 12155
rect 21174 12152 21180 12164
rect 21114 12124 21180 12152
rect 19889 12115 19947 12121
rect 13817 12087 13875 12093
rect 13817 12084 13829 12087
rect 13780 12056 13829 12084
rect 13780 12044 13786 12056
rect 13817 12053 13829 12056
rect 13863 12053 13875 12087
rect 13817 12047 13875 12053
rect 14274 12044 14280 12096
rect 14332 12084 14338 12096
rect 14461 12087 14519 12093
rect 14461 12084 14473 12087
rect 14332 12056 14473 12084
rect 14332 12044 14338 12056
rect 14461 12053 14473 12056
rect 14507 12053 14519 12087
rect 14461 12047 14519 12053
rect 15562 12044 15568 12096
rect 15620 12044 15626 12096
rect 15657 12087 15715 12093
rect 15657 12053 15669 12087
rect 15703 12084 15715 12087
rect 15746 12084 15752 12096
rect 15703 12056 15752 12084
rect 15703 12053 15715 12056
rect 15657 12047 15715 12053
rect 15746 12044 15752 12056
rect 15804 12044 15810 12096
rect 16850 12044 16856 12096
rect 16908 12084 16914 12096
rect 17402 12084 17408 12096
rect 16908 12056 17408 12084
rect 16908 12044 16914 12056
rect 17402 12044 17408 12056
rect 17460 12044 17466 12096
rect 17586 12044 17592 12096
rect 17644 12044 17650 12096
rect 18874 12044 18880 12096
rect 18932 12044 18938 12096
rect 19904 12084 19932 12115
rect 21174 12112 21180 12124
rect 21232 12152 21238 12164
rect 21232 12124 22416 12152
rect 21232 12112 21238 12124
rect 20806 12084 20812 12096
rect 19904 12056 20812 12084
rect 20806 12044 20812 12056
rect 20864 12044 20870 12096
rect 21821 12087 21879 12093
rect 21821 12053 21833 12087
rect 21867 12084 21879 12087
rect 22002 12084 22008 12096
rect 21867 12056 22008 12084
rect 21867 12053 21879 12056
rect 21821 12047 21879 12053
rect 22002 12044 22008 12056
rect 22060 12044 22066 12096
rect 22388 12093 22416 12124
rect 22373 12087 22431 12093
rect 22373 12053 22385 12087
rect 22419 12084 22431 12087
rect 22646 12084 22652 12096
rect 22419 12056 22652 12084
rect 22419 12053 22431 12056
rect 22373 12047 22431 12053
rect 22646 12044 22652 12056
rect 22704 12044 22710 12096
rect 23290 12044 23296 12096
rect 23348 12044 23354 12096
rect 1104 11994 25852 12016
rect 1104 11942 7950 11994
rect 8002 11942 8014 11994
rect 8066 11942 8078 11994
rect 8130 11942 8142 11994
rect 8194 11942 8206 11994
rect 8258 11942 17950 11994
rect 18002 11942 18014 11994
rect 18066 11942 18078 11994
rect 18130 11942 18142 11994
rect 18194 11942 18206 11994
rect 18258 11942 25852 11994
rect 1104 11920 25852 11942
rect 9858 11840 9864 11892
rect 9916 11880 9922 11892
rect 10873 11883 10931 11889
rect 10873 11880 10885 11883
rect 9916 11852 10885 11880
rect 9916 11840 9922 11852
rect 10873 11849 10885 11852
rect 10919 11849 10931 11883
rect 10873 11843 10931 11849
rect 14734 11840 14740 11892
rect 14792 11840 14798 11892
rect 15565 11883 15623 11889
rect 15565 11849 15577 11883
rect 15611 11880 15623 11883
rect 17586 11880 17592 11892
rect 15611 11852 17592 11880
rect 15611 11849 15623 11852
rect 15565 11843 15623 11849
rect 17586 11840 17592 11852
rect 17644 11840 17650 11892
rect 20622 11840 20628 11892
rect 20680 11880 20686 11892
rect 20809 11883 20867 11889
rect 20809 11880 20821 11883
rect 20680 11852 20821 11880
rect 20680 11840 20686 11852
rect 20809 11849 20821 11852
rect 20855 11849 20867 11883
rect 20809 11843 20867 11849
rect 21174 11840 21180 11892
rect 21232 11840 21238 11892
rect 5902 11772 5908 11824
rect 5960 11812 5966 11824
rect 10410 11812 10416 11824
rect 5960 11784 10416 11812
rect 5960 11772 5966 11784
rect 10410 11772 10416 11784
rect 10468 11772 10474 11824
rect 13722 11772 13728 11824
rect 13780 11772 13786 11824
rect 15654 11772 15660 11824
rect 15712 11772 15718 11824
rect 16206 11772 16212 11824
rect 16264 11772 16270 11824
rect 18322 11812 18328 11824
rect 17972 11784 18328 11812
rect 10229 11747 10287 11753
rect 10229 11713 10241 11747
rect 10275 11744 10287 11747
rect 10962 11744 10968 11756
rect 10275 11716 10968 11744
rect 10275 11713 10287 11716
rect 10229 11707 10287 11713
rect 10962 11704 10968 11716
rect 11020 11704 11026 11756
rect 11790 11704 11796 11756
rect 11848 11744 11854 11756
rect 12989 11747 13047 11753
rect 12989 11744 13001 11747
rect 11848 11716 13001 11744
rect 11848 11704 11854 11716
rect 12989 11713 13001 11716
rect 13035 11713 13047 11747
rect 12989 11707 13047 11713
rect 15010 11704 15016 11756
rect 15068 11744 15074 11756
rect 17972 11753 18000 11784
rect 18322 11772 18328 11784
rect 18380 11772 18386 11824
rect 20254 11772 20260 11824
rect 20312 11812 20318 11824
rect 21818 11812 21824 11824
rect 20312 11784 21824 11812
rect 20312 11772 20318 11784
rect 21818 11772 21824 11784
rect 21876 11772 21882 11824
rect 25130 11772 25136 11824
rect 25188 11772 25194 11824
rect 17957 11747 18015 11753
rect 15068 11716 15792 11744
rect 15068 11704 15074 11716
rect 10318 11636 10324 11688
rect 10376 11676 10382 11688
rect 11517 11679 11575 11685
rect 11517 11676 11529 11679
rect 10376 11648 11529 11676
rect 10376 11636 10382 11648
rect 11517 11645 11529 11648
rect 11563 11645 11575 11679
rect 11517 11639 11575 11645
rect 13265 11679 13323 11685
rect 13265 11645 13277 11679
rect 13311 11676 13323 11679
rect 14918 11676 14924 11688
rect 13311 11648 14924 11676
rect 13311 11645 13323 11648
rect 13265 11639 13323 11645
rect 14918 11636 14924 11648
rect 14976 11636 14982 11688
rect 15764 11685 15792 11716
rect 17957 11713 17969 11747
rect 18003 11713 18015 11747
rect 17957 11707 18015 11713
rect 15749 11679 15807 11685
rect 15749 11645 15761 11679
rect 15795 11645 15807 11679
rect 15749 11639 15807 11645
rect 18233 11679 18291 11685
rect 18233 11645 18245 11679
rect 18279 11676 18291 11679
rect 18874 11676 18880 11688
rect 18279 11648 18880 11676
rect 18279 11645 18291 11648
rect 18233 11639 18291 11645
rect 18874 11636 18880 11648
rect 18932 11636 18938 11688
rect 19352 11676 19380 11730
rect 19702 11704 19708 11756
rect 19760 11744 19766 11756
rect 20165 11747 20223 11753
rect 20165 11744 20177 11747
rect 19760 11716 20177 11744
rect 19760 11704 19766 11716
rect 20165 11713 20177 11716
rect 20211 11713 20223 11747
rect 20165 11707 20223 11713
rect 20346 11704 20352 11756
rect 20404 11744 20410 11756
rect 21174 11744 21180 11756
rect 20404 11716 21180 11744
rect 20404 11704 20410 11716
rect 21174 11704 21180 11716
rect 21232 11704 21238 11756
rect 22738 11704 22744 11756
rect 22796 11744 22802 11756
rect 23937 11747 23995 11753
rect 23937 11744 23949 11747
rect 22796 11716 23949 11744
rect 22796 11704 22802 11716
rect 23937 11713 23949 11716
rect 23983 11713 23995 11747
rect 23937 11707 23995 11713
rect 20364 11676 20392 11704
rect 19352 11648 20392 11676
rect 11606 11568 11612 11620
rect 11664 11608 11670 11620
rect 11790 11608 11796 11620
rect 11664 11580 11796 11608
rect 11664 11568 11670 11580
rect 11790 11568 11796 11580
rect 11848 11568 11854 11620
rect 15197 11611 15255 11617
rect 15197 11577 15209 11611
rect 15243 11608 15255 11611
rect 15243 11580 17540 11608
rect 15243 11577 15255 11580
rect 15197 11571 15255 11577
rect 11974 11500 11980 11552
rect 12032 11540 12038 11552
rect 16393 11543 16451 11549
rect 16393 11540 16405 11543
rect 12032 11512 16405 11540
rect 12032 11500 12038 11512
rect 16393 11509 16405 11512
rect 16439 11540 16451 11543
rect 16850 11540 16856 11552
rect 16439 11512 16856 11540
rect 16439 11509 16451 11512
rect 16393 11503 16451 11509
rect 16850 11500 16856 11512
rect 16908 11500 16914 11552
rect 17512 11540 17540 11580
rect 18322 11540 18328 11552
rect 17512 11512 18328 11540
rect 18322 11500 18328 11512
rect 18380 11500 18386 11552
rect 19702 11500 19708 11552
rect 19760 11500 19766 11552
rect 1104 11450 25852 11472
rect 1104 11398 2950 11450
rect 3002 11398 3014 11450
rect 3066 11398 3078 11450
rect 3130 11398 3142 11450
rect 3194 11398 3206 11450
rect 3258 11398 12950 11450
rect 13002 11398 13014 11450
rect 13066 11398 13078 11450
rect 13130 11398 13142 11450
rect 13194 11398 13206 11450
rect 13258 11398 22950 11450
rect 23002 11398 23014 11450
rect 23066 11398 23078 11450
rect 23130 11398 23142 11450
rect 23194 11398 23206 11450
rect 23258 11398 25852 11450
rect 1104 11376 25852 11398
rect 15470 11296 15476 11348
rect 15528 11296 15534 11348
rect 16669 11339 16727 11345
rect 16669 11305 16681 11339
rect 16715 11336 16727 11339
rect 21726 11336 21732 11348
rect 16715 11308 21732 11336
rect 16715 11305 16727 11308
rect 16669 11299 16727 11305
rect 21726 11296 21732 11308
rect 21784 11296 21790 11348
rect 16022 11228 16028 11280
rect 16080 11268 16086 11280
rect 17129 11271 17187 11277
rect 17129 11268 17141 11271
rect 16080 11240 17141 11268
rect 16080 11228 16086 11240
rect 17129 11237 17141 11240
rect 17175 11237 17187 11271
rect 17129 11231 17187 11237
rect 17770 11228 17776 11280
rect 17828 11268 17834 11280
rect 20165 11271 20223 11277
rect 17828 11240 19012 11268
rect 17828 11228 17834 11240
rect 12342 11160 12348 11212
rect 12400 11200 12406 11212
rect 12400 11172 16574 11200
rect 12400 11160 12406 11172
rect 14734 11092 14740 11144
rect 14792 11132 14798 11144
rect 14829 11135 14887 11141
rect 14829 11132 14841 11135
rect 14792 11104 14841 11132
rect 14792 11092 14798 11104
rect 14829 11101 14841 11104
rect 14875 11101 14887 11135
rect 14829 11095 14887 11101
rect 16022 11092 16028 11144
rect 16080 11092 16086 11144
rect 16546 11132 16574 11172
rect 18598 11160 18604 11212
rect 18656 11200 18662 11212
rect 18877 11203 18935 11209
rect 18877 11200 18889 11203
rect 18656 11172 18889 11200
rect 18656 11160 18662 11172
rect 18877 11169 18889 11172
rect 18923 11169 18935 11203
rect 18877 11163 18935 11169
rect 16853 11135 16911 11141
rect 16853 11132 16865 11135
rect 16546 11104 16865 11132
rect 16853 11101 16865 11104
rect 16899 11101 16911 11135
rect 16853 11095 16911 11101
rect 18417 11135 18475 11141
rect 18417 11101 18429 11135
rect 18463 11132 18475 11135
rect 18616 11132 18644 11160
rect 18463 11104 18644 11132
rect 18984 11132 19012 11240
rect 20165 11237 20177 11271
rect 20211 11237 20223 11271
rect 20165 11231 20223 11237
rect 21177 11271 21235 11277
rect 21177 11237 21189 11271
rect 21223 11268 21235 11271
rect 22186 11268 22192 11280
rect 21223 11240 22192 11268
rect 21223 11237 21235 11240
rect 21177 11231 21235 11237
rect 20180 11200 20208 11231
rect 22186 11228 22192 11240
rect 22244 11228 22250 11280
rect 23201 11271 23259 11277
rect 23201 11237 23213 11271
rect 23247 11268 23259 11271
rect 23382 11268 23388 11280
rect 23247 11240 23388 11268
rect 23247 11237 23259 11240
rect 23201 11231 23259 11237
rect 23382 11228 23388 11240
rect 23440 11228 23446 11280
rect 20180 11172 23428 11200
rect 20349 11135 20407 11141
rect 20349 11132 20361 11135
rect 18984 11104 20361 11132
rect 18463 11101 18475 11104
rect 18417 11095 18475 11101
rect 20349 11101 20361 11104
rect 20395 11101 20407 11135
rect 20349 11095 20407 11101
rect 21726 11092 21732 11144
rect 21784 11092 21790 11144
rect 23400 11141 23428 11172
rect 23385 11135 23443 11141
rect 23385 11101 23397 11135
rect 23431 11101 23443 11135
rect 23385 11095 23443 11101
rect 16209 11067 16267 11073
rect 16209 11033 16221 11067
rect 16255 11064 16267 11067
rect 16758 11064 16764 11076
rect 16255 11036 16764 11064
rect 16255 11033 16267 11036
rect 16209 11027 16267 11033
rect 16758 11024 16764 11036
rect 16816 11024 16822 11076
rect 18601 11067 18659 11073
rect 18601 11033 18613 11067
rect 18647 11064 18659 11067
rect 18690 11064 18696 11076
rect 18647 11036 18696 11064
rect 18647 11033 18659 11036
rect 18601 11027 18659 11033
rect 18690 11024 18696 11036
rect 18748 11024 18754 11076
rect 20993 11067 21051 11073
rect 20993 11033 21005 11067
rect 21039 11064 21051 11067
rect 21082 11064 21088 11076
rect 21039 11036 21088 11064
rect 21039 11033 21051 11036
rect 20993 11027 21051 11033
rect 21082 11024 21088 11036
rect 21140 11024 21146 11076
rect 21913 11067 21971 11073
rect 21913 11033 21925 11067
rect 21959 11064 21971 11067
rect 23842 11064 23848 11076
rect 21959 11036 23848 11064
rect 21959 11033 21971 11036
rect 21913 11027 21971 11033
rect 23842 11024 23848 11036
rect 23900 11024 23906 11076
rect 19518 10956 19524 11008
rect 19576 10956 19582 11008
rect 1104 10906 25852 10928
rect 1104 10854 7950 10906
rect 8002 10854 8014 10906
rect 8066 10854 8078 10906
rect 8130 10854 8142 10906
rect 8194 10854 8206 10906
rect 8258 10854 17950 10906
rect 18002 10854 18014 10906
rect 18066 10854 18078 10906
rect 18130 10854 18142 10906
rect 18194 10854 18206 10906
rect 18258 10854 25852 10906
rect 1104 10832 25852 10854
rect 19518 10752 19524 10804
rect 19576 10752 19582 10804
rect 19610 10752 19616 10804
rect 19668 10752 19674 10804
rect 21082 10752 21088 10804
rect 21140 10792 21146 10804
rect 21269 10795 21327 10801
rect 21269 10792 21281 10795
rect 21140 10764 21281 10792
rect 21140 10752 21146 10764
rect 21269 10761 21281 10764
rect 21315 10761 21327 10795
rect 21269 10755 21327 10761
rect 10042 10684 10048 10736
rect 10100 10724 10106 10736
rect 11977 10727 12035 10733
rect 11977 10724 11989 10727
rect 10100 10696 11989 10724
rect 10100 10684 10106 10696
rect 11977 10693 11989 10696
rect 12023 10724 12035 10727
rect 12437 10727 12495 10733
rect 12437 10724 12449 10727
rect 12023 10696 12449 10724
rect 12023 10693 12035 10696
rect 11977 10687 12035 10693
rect 12437 10693 12449 10696
rect 12483 10693 12495 10727
rect 12437 10687 12495 10693
rect 18322 10616 18328 10668
rect 18380 10656 18386 10668
rect 18509 10659 18567 10665
rect 18509 10656 18521 10659
rect 18380 10628 18521 10656
rect 18380 10616 18386 10628
rect 18509 10625 18521 10628
rect 18555 10625 18567 10659
rect 18509 10619 18567 10625
rect 20714 10616 20720 10668
rect 20772 10656 20778 10668
rect 22925 10659 22983 10665
rect 22925 10656 22937 10659
rect 20772 10628 22937 10656
rect 20772 10616 20778 10628
rect 22925 10625 22937 10628
rect 22971 10625 22983 10659
rect 22925 10619 22983 10625
rect 23934 10616 23940 10668
rect 23992 10616 23998 10668
rect 18782 10548 18788 10600
rect 18840 10588 18846 10600
rect 19150 10588 19156 10600
rect 18840 10560 19156 10588
rect 18840 10548 18846 10560
rect 19150 10548 19156 10560
rect 19208 10548 19214 10600
rect 19702 10548 19708 10600
rect 19760 10548 19766 10600
rect 24762 10548 24768 10600
rect 24820 10548 24826 10600
rect 12161 10523 12219 10529
rect 12161 10489 12173 10523
rect 12207 10520 12219 10523
rect 12526 10520 12532 10532
rect 12207 10492 12532 10520
rect 12207 10489 12219 10492
rect 12161 10483 12219 10489
rect 12526 10480 12532 10492
rect 12584 10480 12590 10532
rect 18325 10523 18383 10529
rect 18325 10489 18337 10523
rect 18371 10520 18383 10523
rect 20622 10520 20628 10532
rect 18371 10492 20628 10520
rect 18371 10489 18383 10492
rect 18325 10483 18383 10489
rect 20622 10480 20628 10492
rect 20680 10480 20686 10532
rect 19153 10455 19211 10461
rect 19153 10421 19165 10455
rect 19199 10452 19211 10455
rect 21174 10452 21180 10464
rect 19199 10424 21180 10452
rect 19199 10421 19211 10424
rect 19153 10415 19211 10421
rect 21174 10412 21180 10424
rect 21232 10412 21238 10464
rect 22554 10412 22560 10464
rect 22612 10452 22618 10464
rect 22741 10455 22799 10461
rect 22741 10452 22753 10455
rect 22612 10424 22753 10452
rect 22612 10412 22618 10424
rect 22741 10421 22753 10424
rect 22787 10421 22799 10455
rect 22741 10415 22799 10421
rect 1104 10362 25852 10384
rect 1104 10310 2950 10362
rect 3002 10310 3014 10362
rect 3066 10310 3078 10362
rect 3130 10310 3142 10362
rect 3194 10310 3206 10362
rect 3258 10310 12950 10362
rect 13002 10310 13014 10362
rect 13066 10310 13078 10362
rect 13130 10310 13142 10362
rect 13194 10310 13206 10362
rect 13258 10310 22950 10362
rect 23002 10310 23014 10362
rect 23066 10310 23078 10362
rect 23130 10310 23142 10362
rect 23194 10310 23206 10362
rect 23258 10310 25852 10362
rect 1104 10288 25852 10310
rect 12618 10004 12624 10056
rect 12676 10044 12682 10056
rect 14553 10047 14611 10053
rect 14553 10044 14565 10047
rect 12676 10016 14565 10044
rect 12676 10004 12682 10016
rect 14553 10013 14565 10016
rect 14599 10013 14611 10047
rect 14553 10007 14611 10013
rect 16853 10047 16911 10053
rect 16853 10013 16865 10047
rect 16899 10044 16911 10047
rect 18506 10044 18512 10056
rect 16899 10016 18512 10044
rect 16899 10013 16911 10016
rect 16853 10007 16911 10013
rect 18506 10004 18512 10016
rect 18564 10004 18570 10056
rect 21910 10004 21916 10056
rect 21968 10044 21974 10056
rect 22189 10047 22247 10053
rect 22189 10044 22201 10047
rect 21968 10016 22201 10044
rect 21968 10004 21974 10016
rect 22189 10013 22201 10016
rect 22235 10013 22247 10047
rect 22189 10007 22247 10013
rect 22646 10004 22652 10056
rect 22704 10004 22710 10056
rect 22830 10004 22836 10056
rect 22888 10044 22894 10056
rect 24857 10047 24915 10053
rect 24857 10044 24869 10047
rect 22888 10016 24869 10044
rect 22888 10004 22894 10016
rect 24857 10013 24869 10016
rect 24903 10013 24915 10047
rect 24857 10007 24915 10013
rect 14737 9979 14795 9985
rect 14737 9945 14749 9979
rect 14783 9976 14795 9979
rect 14826 9976 14832 9988
rect 14783 9948 14832 9976
rect 14783 9945 14795 9948
rect 14737 9939 14795 9945
rect 14826 9936 14832 9948
rect 14884 9936 14890 9988
rect 23845 9979 23903 9985
rect 23845 9945 23857 9979
rect 23891 9976 23903 9979
rect 24946 9976 24952 9988
rect 23891 9948 24952 9976
rect 23891 9945 23903 9948
rect 23845 9939 23903 9945
rect 24946 9936 24952 9948
rect 25004 9936 25010 9988
rect 16942 9868 16948 9920
rect 17000 9868 17006 9920
rect 21818 9868 21824 9920
rect 21876 9908 21882 9920
rect 22005 9911 22063 9917
rect 22005 9908 22017 9911
rect 21876 9880 22017 9908
rect 21876 9868 21882 9880
rect 22005 9877 22017 9880
rect 22051 9877 22063 9911
rect 22005 9871 22063 9877
rect 23566 9868 23572 9920
rect 23624 9908 23630 9920
rect 24673 9911 24731 9917
rect 24673 9908 24685 9911
rect 23624 9880 24685 9908
rect 23624 9868 23630 9880
rect 24673 9877 24685 9880
rect 24719 9877 24731 9911
rect 24673 9871 24731 9877
rect 1104 9818 25852 9840
rect 1104 9766 7950 9818
rect 8002 9766 8014 9818
rect 8066 9766 8078 9818
rect 8130 9766 8142 9818
rect 8194 9766 8206 9818
rect 8258 9766 17950 9818
rect 18002 9766 18014 9818
rect 18066 9766 18078 9818
rect 18130 9766 18142 9818
rect 18194 9766 18206 9818
rect 18258 9766 25852 9818
rect 1104 9744 25852 9766
rect 22465 9707 22523 9713
rect 22465 9673 22477 9707
rect 22511 9704 22523 9707
rect 22646 9704 22652 9716
rect 22511 9676 22652 9704
rect 22511 9673 22523 9676
rect 22465 9667 22523 9673
rect 22646 9664 22652 9676
rect 22704 9664 22710 9716
rect 10042 9596 10048 9648
rect 10100 9636 10106 9648
rect 14090 9636 14096 9648
rect 10100 9608 14096 9636
rect 10100 9596 10106 9608
rect 14090 9596 14096 9608
rect 14148 9596 14154 9648
rect 16945 9639 17003 9645
rect 16945 9605 16957 9639
rect 16991 9636 17003 9639
rect 17494 9636 17500 9648
rect 16991 9608 17500 9636
rect 16991 9605 17003 9608
rect 16945 9599 17003 9605
rect 17494 9596 17500 9608
rect 17552 9596 17558 9648
rect 18877 9639 18935 9645
rect 18877 9605 18889 9639
rect 18923 9636 18935 9639
rect 19058 9636 19064 9648
rect 18923 9608 19064 9636
rect 18923 9605 18935 9608
rect 18877 9599 18935 9605
rect 19058 9596 19064 9608
rect 19116 9596 19122 9648
rect 22002 9596 22008 9648
rect 22060 9636 22066 9648
rect 22060 9608 23428 9636
rect 22060 9596 22066 9608
rect 7650 9528 7656 9580
rect 7708 9568 7714 9580
rect 12434 9568 12440 9580
rect 7708 9540 12440 9568
rect 7708 9528 7714 9540
rect 12434 9528 12440 9540
rect 12492 9528 12498 9580
rect 20622 9528 20628 9580
rect 20680 9568 20686 9580
rect 23400 9577 23428 9608
rect 22649 9571 22707 9577
rect 22649 9568 22661 9571
rect 20680 9540 22661 9568
rect 20680 9528 20686 9540
rect 22649 9537 22661 9540
rect 22695 9537 22707 9571
rect 22649 9531 22707 9537
rect 23385 9571 23443 9577
rect 23385 9537 23397 9571
rect 23431 9537 23443 9571
rect 23385 9531 23443 9537
rect 23842 9528 23848 9580
rect 23900 9568 23906 9580
rect 23937 9571 23995 9577
rect 23937 9568 23949 9571
rect 23900 9540 23949 9568
rect 23900 9528 23906 9540
rect 23937 9537 23949 9540
rect 23983 9537 23995 9571
rect 23937 9531 23995 9537
rect 2866 9460 2872 9512
rect 2924 9500 2930 9512
rect 5718 9500 5724 9512
rect 2924 9472 5724 9500
rect 2924 9460 2930 9472
rect 5718 9460 5724 9472
rect 5776 9460 5782 9512
rect 7466 9460 7472 9512
rect 7524 9500 7530 9512
rect 7561 9503 7619 9509
rect 7561 9500 7573 9503
rect 7524 9472 7573 9500
rect 7524 9460 7530 9472
rect 7561 9469 7573 9472
rect 7607 9469 7619 9503
rect 7561 9463 7619 9469
rect 24670 9460 24676 9512
rect 24728 9460 24734 9512
rect 17129 9435 17187 9441
rect 17129 9401 17141 9435
rect 17175 9432 17187 9435
rect 17402 9432 17408 9444
rect 17175 9404 17408 9432
rect 17175 9401 17187 9404
rect 17129 9395 17187 9401
rect 17402 9392 17408 9404
rect 17460 9392 17466 9444
rect 19061 9435 19119 9441
rect 19061 9401 19073 9435
rect 19107 9432 19119 9435
rect 22830 9432 22836 9444
rect 19107 9404 22836 9432
rect 19107 9401 19119 9404
rect 19061 9395 19119 9401
rect 22830 9392 22836 9404
rect 22888 9392 22894 9444
rect 23201 9367 23259 9373
rect 23201 9333 23213 9367
rect 23247 9364 23259 9367
rect 23474 9364 23480 9376
rect 23247 9336 23480 9364
rect 23247 9333 23259 9336
rect 23201 9327 23259 9333
rect 23474 9324 23480 9336
rect 23532 9324 23538 9376
rect 1104 9274 25852 9296
rect 1104 9222 2950 9274
rect 3002 9222 3014 9274
rect 3066 9222 3078 9274
rect 3130 9222 3142 9274
rect 3194 9222 3206 9274
rect 3258 9222 12950 9274
rect 13002 9222 13014 9274
rect 13066 9222 13078 9274
rect 13130 9222 13142 9274
rect 13194 9222 13206 9274
rect 13258 9222 22950 9274
rect 23002 9222 23014 9274
rect 23066 9222 23078 9274
rect 23130 9222 23142 9274
rect 23194 9222 23206 9274
rect 23258 9222 25852 9274
rect 1104 9200 25852 9222
rect 7098 9120 7104 9172
rect 7156 9120 7162 9172
rect 7745 9027 7803 9033
rect 7745 8993 7757 9027
rect 7791 9024 7803 9027
rect 9030 9024 9036 9036
rect 7791 8996 9036 9024
rect 7791 8993 7803 8996
rect 7745 8987 7803 8993
rect 9030 8984 9036 8996
rect 9088 8984 9094 9036
rect 7466 8916 7472 8968
rect 7524 8916 7530 8968
rect 23290 8916 23296 8968
rect 23348 8956 23354 8968
rect 23845 8959 23903 8965
rect 23845 8956 23857 8959
rect 23348 8928 23857 8956
rect 23348 8916 23354 8928
rect 23845 8925 23857 8928
rect 23891 8925 23903 8959
rect 23845 8919 23903 8925
rect 24854 8916 24860 8968
rect 24912 8916 24918 8968
rect 7561 8891 7619 8897
rect 7561 8888 7573 8891
rect 6886 8860 7573 8888
rect 5626 8780 5632 8832
rect 5684 8820 5690 8832
rect 6886 8820 6914 8860
rect 7561 8857 7573 8860
rect 7607 8857 7619 8891
rect 7561 8851 7619 8857
rect 9490 8848 9496 8900
rect 9548 8888 9554 8900
rect 13906 8888 13912 8900
rect 9548 8860 13912 8888
rect 9548 8848 9554 8860
rect 13906 8848 13912 8860
rect 13964 8848 13970 8900
rect 23308 8860 24716 8888
rect 23308 8832 23336 8860
rect 5684 8792 6914 8820
rect 5684 8780 5690 8792
rect 23290 8780 23296 8832
rect 23348 8780 23354 8832
rect 23934 8780 23940 8832
rect 23992 8780 23998 8832
rect 24688 8829 24716 8860
rect 24673 8823 24731 8829
rect 24673 8789 24685 8823
rect 24719 8789 24731 8823
rect 24673 8783 24731 8789
rect 1104 8730 25852 8752
rect 1104 8678 7950 8730
rect 8002 8678 8014 8730
rect 8066 8678 8078 8730
rect 8130 8678 8142 8730
rect 8194 8678 8206 8730
rect 8258 8678 17950 8730
rect 18002 8678 18014 8730
rect 18066 8678 18078 8730
rect 18130 8678 18142 8730
rect 18194 8678 18206 8730
rect 18258 8678 25852 8730
rect 1104 8656 25852 8678
rect 5258 8616 5264 8628
rect 3988 8588 5264 8616
rect 3988 8489 4016 8588
rect 5258 8576 5264 8588
rect 5316 8576 5322 8628
rect 6365 8551 6423 8557
rect 6365 8548 6377 8551
rect 5474 8520 6377 8548
rect 6365 8517 6377 8520
rect 6411 8548 6423 8551
rect 10318 8548 10324 8560
rect 6411 8520 10324 8548
rect 6411 8517 6423 8520
rect 6365 8511 6423 8517
rect 10318 8508 10324 8520
rect 10376 8508 10382 8560
rect 17034 8508 17040 8560
rect 17092 8548 17098 8560
rect 18877 8551 18935 8557
rect 18877 8548 18889 8551
rect 17092 8520 18889 8548
rect 17092 8508 17098 8520
rect 18877 8517 18889 8520
rect 18923 8517 18935 8551
rect 18877 8511 18935 8517
rect 20809 8551 20867 8557
rect 20809 8517 20821 8551
rect 20855 8548 20867 8551
rect 21358 8548 21364 8560
rect 20855 8520 21364 8548
rect 20855 8517 20867 8520
rect 20809 8511 20867 8517
rect 21358 8508 21364 8520
rect 21416 8508 21422 8560
rect 25130 8508 25136 8560
rect 25188 8508 25194 8560
rect 3973 8483 4031 8489
rect 3973 8449 3985 8483
rect 4019 8449 4031 8483
rect 3973 8443 4031 8449
rect 5997 8483 6055 8489
rect 5997 8449 6009 8483
rect 6043 8480 6055 8483
rect 6822 8480 6828 8492
rect 6043 8452 6828 8480
rect 6043 8449 6055 8452
rect 5997 8443 6055 8449
rect 6822 8440 6828 8452
rect 6880 8440 6886 8492
rect 22281 8483 22339 8489
rect 22281 8449 22293 8483
rect 22327 8480 22339 8483
rect 22370 8480 22376 8492
rect 22327 8452 22376 8480
rect 22327 8449 22339 8452
rect 22281 8443 22339 8449
rect 22370 8440 22376 8452
rect 22428 8440 22434 8492
rect 23382 8440 23388 8492
rect 23440 8480 23446 8492
rect 23937 8483 23995 8489
rect 23937 8480 23949 8483
rect 23440 8452 23949 8480
rect 23440 8440 23446 8452
rect 23937 8449 23949 8452
rect 23983 8449 23995 8483
rect 23937 8443 23995 8449
rect 2774 8372 2780 8424
rect 2832 8412 2838 8424
rect 4249 8415 4307 8421
rect 4249 8412 4261 8415
rect 2832 8384 4261 8412
rect 2832 8372 2838 8384
rect 4249 8381 4261 8384
rect 4295 8381 4307 8415
rect 4249 8375 4307 8381
rect 22738 8372 22744 8424
rect 22796 8372 22802 8424
rect 19061 8347 19119 8353
rect 19061 8313 19073 8347
rect 19107 8344 19119 8347
rect 20438 8344 20444 8356
rect 19107 8316 20444 8344
rect 19107 8313 19119 8316
rect 19061 8307 19119 8313
rect 20438 8304 20444 8316
rect 20496 8304 20502 8356
rect 20993 8347 21051 8353
rect 20993 8313 21005 8347
rect 21039 8344 21051 8347
rect 21266 8344 21272 8356
rect 21039 8316 21272 8344
rect 21039 8313 21051 8316
rect 20993 8307 21051 8313
rect 21266 8304 21272 8316
rect 21324 8304 21330 8356
rect 1104 8186 25852 8208
rect 1104 8134 2950 8186
rect 3002 8134 3014 8186
rect 3066 8134 3078 8186
rect 3130 8134 3142 8186
rect 3194 8134 3206 8186
rect 3258 8134 12950 8186
rect 13002 8134 13014 8186
rect 13066 8134 13078 8186
rect 13130 8134 13142 8186
rect 13194 8134 13206 8186
rect 13258 8134 22950 8186
rect 23002 8134 23014 8186
rect 23066 8134 23078 8186
rect 23130 8134 23142 8186
rect 23194 8134 23206 8186
rect 23258 8134 25852 8186
rect 1104 8112 25852 8134
rect 23290 7896 23296 7948
rect 23348 7896 23354 7948
rect 19794 7828 19800 7880
rect 19852 7868 19858 7880
rect 20625 7871 20683 7877
rect 20625 7868 20637 7871
rect 19852 7840 20637 7868
rect 19852 7828 19858 7840
rect 20625 7837 20637 7840
rect 20671 7837 20683 7871
rect 20625 7831 20683 7837
rect 21174 7828 21180 7880
rect 21232 7868 21238 7880
rect 21637 7871 21695 7877
rect 21637 7868 21649 7871
rect 21232 7840 21649 7868
rect 21232 7828 21238 7840
rect 21637 7837 21649 7840
rect 21683 7837 21695 7871
rect 21637 7831 21695 7837
rect 22833 7871 22891 7877
rect 22833 7837 22845 7871
rect 22879 7868 22891 7871
rect 23566 7868 23572 7880
rect 22879 7840 23572 7868
rect 22879 7837 22891 7840
rect 22833 7831 22891 7837
rect 23566 7828 23572 7840
rect 23624 7828 23630 7880
rect 20254 7692 20260 7744
rect 20312 7732 20318 7744
rect 20441 7735 20499 7741
rect 20441 7732 20453 7735
rect 20312 7704 20453 7732
rect 20312 7692 20318 7704
rect 20441 7701 20453 7704
rect 20487 7701 20499 7735
rect 20441 7695 20499 7701
rect 21453 7735 21511 7741
rect 21453 7701 21465 7735
rect 21499 7732 21511 7735
rect 24670 7732 24676 7744
rect 21499 7704 24676 7732
rect 21499 7701 21511 7704
rect 21453 7695 21511 7701
rect 24670 7692 24676 7704
rect 24728 7692 24734 7744
rect 1104 7642 25852 7664
rect 1104 7590 7950 7642
rect 8002 7590 8014 7642
rect 8066 7590 8078 7642
rect 8130 7590 8142 7642
rect 8194 7590 8206 7642
rect 8258 7590 17950 7642
rect 18002 7590 18014 7642
rect 18066 7590 18078 7642
rect 18130 7590 18142 7642
rect 18194 7590 18206 7642
rect 18258 7590 25852 7642
rect 1104 7568 25852 7590
rect 15194 7420 15200 7472
rect 15252 7460 15258 7472
rect 18509 7463 18567 7469
rect 18509 7460 18521 7463
rect 15252 7432 18521 7460
rect 15252 7420 15258 7432
rect 18509 7429 18521 7432
rect 18555 7429 18567 7463
rect 18509 7423 18567 7429
rect 19429 7463 19487 7469
rect 19429 7429 19441 7463
rect 19475 7429 19487 7463
rect 19429 7423 19487 7429
rect 15838 7352 15844 7404
rect 15896 7392 15902 7404
rect 19444 7392 19472 7423
rect 20438 7420 20444 7472
rect 20496 7460 20502 7472
rect 20496 7432 22140 7460
rect 20496 7420 20502 7432
rect 15896 7364 19472 7392
rect 20257 7395 20315 7401
rect 15896 7352 15902 7364
rect 20257 7361 20269 7395
rect 20303 7392 20315 7395
rect 20714 7392 20720 7404
rect 20303 7364 20720 7392
rect 20303 7361 20315 7364
rect 20257 7355 20315 7361
rect 20714 7352 20720 7364
rect 20772 7352 20778 7404
rect 22112 7401 22140 7432
rect 25130 7420 25136 7472
rect 25188 7420 25194 7472
rect 22097 7395 22155 7401
rect 22097 7361 22109 7395
rect 22143 7361 22155 7395
rect 22097 7355 22155 7361
rect 23937 7395 23995 7401
rect 23937 7361 23949 7395
rect 23983 7361 23995 7395
rect 23937 7355 23995 7361
rect 16206 7284 16212 7336
rect 16264 7324 16270 7336
rect 21269 7327 21327 7333
rect 16264 7296 20300 7324
rect 16264 7284 16270 7296
rect 17678 7216 17684 7268
rect 17736 7256 17742 7268
rect 19613 7259 19671 7265
rect 19613 7256 19625 7259
rect 17736 7228 19625 7256
rect 17736 7216 17742 7228
rect 19613 7225 19625 7228
rect 19659 7225 19671 7259
rect 20272 7256 20300 7296
rect 21269 7293 21281 7327
rect 21315 7324 21327 7327
rect 21634 7324 21640 7336
rect 21315 7296 21640 7324
rect 21315 7293 21327 7296
rect 21269 7287 21327 7293
rect 21634 7284 21640 7296
rect 21692 7284 21698 7336
rect 22278 7284 22284 7336
rect 22336 7324 22342 7336
rect 22557 7327 22615 7333
rect 22557 7324 22569 7327
rect 22336 7296 22569 7324
rect 22336 7284 22342 7296
rect 22557 7293 22569 7296
rect 22603 7293 22615 7327
rect 22557 7287 22615 7293
rect 23952 7256 23980 7355
rect 20272 7228 23980 7256
rect 19613 7219 19671 7225
rect 18601 7191 18659 7197
rect 18601 7157 18613 7191
rect 18647 7188 18659 7191
rect 20622 7188 20628 7200
rect 18647 7160 20628 7188
rect 18647 7157 18659 7160
rect 18601 7151 18659 7157
rect 20622 7148 20628 7160
rect 20680 7148 20686 7200
rect 1104 7098 25852 7120
rect 1104 7046 2950 7098
rect 3002 7046 3014 7098
rect 3066 7046 3078 7098
rect 3130 7046 3142 7098
rect 3194 7046 3206 7098
rect 3258 7046 12950 7098
rect 13002 7046 13014 7098
rect 13066 7046 13078 7098
rect 13130 7046 13142 7098
rect 13194 7046 13206 7098
rect 13258 7046 22950 7098
rect 23002 7046 23014 7098
rect 23066 7046 23078 7098
rect 23130 7046 23142 7098
rect 23194 7046 23206 7098
rect 23258 7046 25852 7098
rect 1104 7024 25852 7046
rect 15562 6740 15568 6792
rect 15620 6780 15626 6792
rect 20257 6783 20315 6789
rect 20257 6780 20269 6783
rect 15620 6752 20269 6780
rect 15620 6740 15626 6752
rect 20257 6749 20269 6752
rect 20303 6749 20315 6783
rect 20257 6743 20315 6749
rect 20809 6783 20867 6789
rect 20809 6749 20821 6783
rect 20855 6749 20867 6783
rect 20809 6743 20867 6749
rect 22833 6783 22891 6789
rect 22833 6749 22845 6783
rect 22879 6780 22891 6783
rect 23382 6780 23388 6792
rect 22879 6752 23388 6780
rect 22879 6749 22891 6752
rect 22833 6743 22891 6749
rect 3050 6672 3056 6724
rect 3108 6712 3114 6724
rect 6086 6712 6092 6724
rect 3108 6684 6092 6712
rect 3108 6672 3114 6684
rect 6086 6672 6092 6684
rect 6144 6672 6150 6724
rect 20073 6647 20131 6653
rect 20073 6613 20085 6647
rect 20119 6644 20131 6647
rect 20824 6644 20852 6743
rect 23382 6740 23388 6752
rect 23440 6740 23446 6792
rect 22002 6672 22008 6724
rect 22060 6672 22066 6724
rect 23845 6715 23903 6721
rect 23845 6681 23857 6715
rect 23891 6712 23903 6715
rect 25774 6712 25780 6724
rect 23891 6684 25780 6712
rect 23891 6681 23903 6684
rect 23845 6675 23903 6681
rect 25774 6672 25780 6684
rect 25832 6672 25838 6724
rect 20119 6616 20852 6644
rect 20119 6613 20131 6616
rect 20073 6607 20131 6613
rect 1104 6554 25852 6576
rect 1104 6502 7950 6554
rect 8002 6502 8014 6554
rect 8066 6502 8078 6554
rect 8130 6502 8142 6554
rect 8194 6502 8206 6554
rect 8258 6502 17950 6554
rect 18002 6502 18014 6554
rect 18066 6502 18078 6554
rect 18130 6502 18142 6554
rect 18194 6502 18206 6554
rect 18258 6502 25852 6554
rect 1104 6480 25852 6502
rect 11790 6400 11796 6452
rect 11848 6440 11854 6452
rect 17957 6443 18015 6449
rect 17957 6440 17969 6443
rect 11848 6412 17969 6440
rect 11848 6400 11854 6412
rect 17957 6409 17969 6412
rect 18003 6409 18015 6443
rect 17957 6403 18015 6409
rect 5534 6264 5540 6316
rect 5592 6304 5598 6316
rect 9766 6304 9772 6316
rect 5592 6276 9772 6304
rect 5592 6264 5598 6276
rect 9766 6264 9772 6276
rect 9824 6264 9830 6316
rect 17972 6304 18000 6403
rect 18233 6307 18291 6313
rect 18233 6304 18245 6307
rect 17972 6276 18245 6304
rect 18233 6273 18245 6276
rect 18279 6273 18291 6307
rect 18233 6267 18291 6273
rect 20254 6264 20260 6316
rect 20312 6264 20318 6316
rect 22186 6264 22192 6316
rect 22244 6264 22250 6316
rect 23474 6264 23480 6316
rect 23532 6304 23538 6316
rect 23937 6307 23995 6313
rect 23937 6304 23949 6307
rect 23532 6276 23949 6304
rect 23532 6264 23538 6276
rect 23937 6273 23949 6276
rect 23983 6273 23995 6307
rect 23937 6267 23995 6273
rect 19245 6239 19303 6245
rect 19245 6205 19257 6239
rect 19291 6205 19303 6239
rect 19245 6199 19303 6205
rect 21269 6239 21327 6245
rect 21269 6205 21281 6239
rect 21315 6236 21327 6239
rect 21726 6236 21732 6248
rect 21315 6208 21732 6236
rect 21315 6205 21327 6208
rect 21269 6199 21327 6205
rect 19260 6168 19288 6199
rect 21726 6196 21732 6208
rect 21784 6196 21790 6248
rect 21910 6196 21916 6248
rect 21968 6236 21974 6248
rect 22465 6239 22523 6245
rect 22465 6236 22477 6239
rect 21968 6208 22477 6236
rect 21968 6196 21974 6208
rect 22465 6205 22477 6208
rect 22511 6205 22523 6239
rect 22465 6199 22523 6205
rect 24762 6196 24768 6248
rect 24820 6196 24826 6248
rect 22186 6168 22192 6180
rect 19260 6140 22192 6168
rect 22186 6128 22192 6140
rect 22244 6128 22250 6180
rect 1104 6010 25852 6032
rect 1104 5958 2950 6010
rect 3002 5958 3014 6010
rect 3066 5958 3078 6010
rect 3130 5958 3142 6010
rect 3194 5958 3206 6010
rect 3258 5958 12950 6010
rect 13002 5958 13014 6010
rect 13066 5958 13078 6010
rect 13130 5958 13142 6010
rect 13194 5958 13206 6010
rect 13258 5958 22950 6010
rect 23002 5958 23014 6010
rect 23066 5958 23078 6010
rect 23130 5958 23142 6010
rect 23194 5958 23206 6010
rect 23258 5958 25852 6010
rect 1104 5936 25852 5958
rect 20714 5856 20720 5908
rect 20772 5896 20778 5908
rect 24765 5899 24823 5905
rect 24765 5896 24777 5899
rect 20772 5868 24777 5896
rect 20772 5856 20778 5868
rect 24765 5865 24777 5868
rect 24811 5865 24823 5899
rect 24765 5859 24823 5865
rect 10594 5788 10600 5840
rect 10652 5828 10658 5840
rect 11882 5828 11888 5840
rect 10652 5800 11888 5828
rect 10652 5788 10658 5800
rect 11882 5788 11888 5800
rect 11940 5788 11946 5840
rect 20438 5720 20444 5772
rect 20496 5760 20502 5772
rect 20993 5763 21051 5769
rect 20993 5760 21005 5763
rect 20496 5732 21005 5760
rect 20496 5720 20502 5732
rect 20993 5729 21005 5732
rect 21039 5729 21051 5763
rect 20993 5723 21051 5729
rect 21542 5720 21548 5772
rect 21600 5760 21606 5772
rect 22833 5763 22891 5769
rect 22833 5760 22845 5763
rect 21600 5732 22845 5760
rect 21600 5720 21606 5732
rect 22833 5729 22845 5732
rect 22879 5729 22891 5763
rect 22833 5723 22891 5729
rect 9306 5652 9312 5704
rect 9364 5692 9370 5704
rect 13446 5692 13452 5704
rect 9364 5664 13452 5692
rect 9364 5652 9370 5664
rect 13446 5652 13452 5664
rect 13504 5652 13510 5704
rect 20530 5652 20536 5704
rect 20588 5652 20594 5704
rect 20622 5652 20628 5704
rect 20680 5692 20686 5704
rect 22373 5695 22431 5701
rect 22373 5692 22385 5695
rect 20680 5664 22385 5692
rect 20680 5652 20686 5664
rect 22373 5661 22385 5664
rect 22419 5661 22431 5695
rect 22373 5655 22431 5661
rect 2682 5584 2688 5636
rect 2740 5624 2746 5636
rect 9398 5624 9404 5636
rect 2740 5596 9404 5624
rect 2740 5584 2746 5596
rect 9398 5584 9404 5596
rect 9456 5584 9462 5636
rect 21818 5584 21824 5636
rect 21876 5624 21882 5636
rect 24673 5627 24731 5633
rect 24673 5624 24685 5627
rect 21876 5596 24685 5624
rect 21876 5584 21882 5596
rect 24673 5593 24685 5596
rect 24719 5593 24731 5627
rect 24673 5587 24731 5593
rect 5166 5516 5172 5568
rect 5224 5556 5230 5568
rect 6270 5556 6276 5568
rect 5224 5528 6276 5556
rect 5224 5516 5230 5528
rect 6270 5516 6276 5528
rect 6328 5516 6334 5568
rect 12618 5516 12624 5568
rect 12676 5556 12682 5568
rect 14550 5556 14556 5568
rect 12676 5528 14556 5556
rect 12676 5516 12682 5528
rect 14550 5516 14556 5528
rect 14608 5516 14614 5568
rect 1104 5466 25852 5488
rect 1104 5414 7950 5466
rect 8002 5414 8014 5466
rect 8066 5414 8078 5466
rect 8130 5414 8142 5466
rect 8194 5414 8206 5466
rect 8258 5414 17950 5466
rect 18002 5414 18014 5466
rect 18066 5414 18078 5466
rect 18130 5414 18142 5466
rect 18194 5414 18206 5466
rect 18258 5414 25852 5466
rect 1104 5392 25852 5414
rect 18785 5287 18843 5293
rect 18785 5253 18797 5287
rect 18831 5284 18843 5287
rect 19518 5284 19524 5296
rect 18831 5256 19524 5284
rect 18831 5253 18843 5256
rect 18785 5247 18843 5253
rect 19518 5244 19524 5256
rect 19576 5244 19582 5296
rect 17770 5176 17776 5228
rect 17828 5176 17834 5228
rect 19058 5176 19064 5228
rect 19116 5216 19122 5228
rect 19429 5219 19487 5225
rect 19429 5216 19441 5219
rect 19116 5188 19441 5216
rect 19116 5176 19122 5188
rect 19429 5185 19441 5188
rect 19475 5185 19487 5219
rect 19429 5179 19487 5185
rect 22094 5176 22100 5228
rect 22152 5176 22158 5228
rect 23934 5176 23940 5228
rect 23992 5176 23998 5228
rect 19334 5108 19340 5160
rect 19392 5148 19398 5160
rect 19889 5151 19947 5157
rect 19889 5148 19901 5151
rect 19392 5120 19901 5148
rect 19392 5108 19398 5120
rect 19889 5117 19901 5120
rect 19935 5117 19947 5151
rect 19889 5111 19947 5117
rect 22462 5108 22468 5160
rect 22520 5108 22526 5160
rect 24762 5108 24768 5160
rect 24820 5108 24826 5160
rect 1104 4922 25852 4944
rect 1104 4870 2950 4922
rect 3002 4870 3014 4922
rect 3066 4870 3078 4922
rect 3130 4870 3142 4922
rect 3194 4870 3206 4922
rect 3258 4870 12950 4922
rect 13002 4870 13014 4922
rect 13066 4870 13078 4922
rect 13130 4870 13142 4922
rect 13194 4870 13206 4922
rect 13258 4870 22950 4922
rect 23002 4870 23014 4922
rect 23066 4870 23078 4922
rect 23130 4870 23142 4922
rect 23194 4870 23206 4922
rect 23258 4870 25852 4922
rect 1104 4848 25852 4870
rect 22370 4768 22376 4820
rect 22428 4808 22434 4820
rect 24765 4811 24823 4817
rect 24765 4808 24777 4811
rect 22428 4780 24777 4808
rect 22428 4768 22434 4780
rect 24765 4777 24777 4780
rect 24811 4777 24823 4811
rect 24765 4771 24823 4777
rect 17770 4700 17776 4752
rect 17828 4740 17834 4752
rect 17828 4712 23520 4740
rect 17828 4700 17834 4712
rect 19886 4632 19892 4684
rect 19944 4632 19950 4684
rect 20714 4632 20720 4684
rect 20772 4672 20778 4684
rect 21729 4675 21787 4681
rect 21729 4672 21741 4675
rect 20772 4644 21741 4672
rect 20772 4632 20778 4644
rect 21729 4641 21741 4644
rect 21775 4641 21787 4675
rect 21729 4635 21787 4641
rect 22554 4632 22560 4684
rect 22612 4672 22618 4684
rect 23492 4681 23520 4712
rect 23201 4675 23259 4681
rect 23201 4672 23213 4675
rect 22612 4644 23213 4672
rect 22612 4632 22618 4644
rect 23201 4641 23213 4644
rect 23247 4641 23259 4675
rect 23201 4635 23259 4641
rect 23477 4675 23535 4681
rect 23477 4641 23489 4675
rect 23523 4641 23535 4675
rect 23477 4635 23535 4641
rect 17678 4564 17684 4616
rect 17736 4564 17742 4616
rect 18690 4564 18696 4616
rect 18748 4604 18754 4616
rect 19429 4607 19487 4613
rect 19429 4604 19441 4607
rect 18748 4576 19441 4604
rect 18748 4564 18754 4576
rect 19429 4573 19441 4576
rect 19475 4573 19487 4607
rect 19429 4567 19487 4573
rect 21266 4564 21272 4616
rect 21324 4564 21330 4616
rect 24670 4564 24676 4616
rect 24728 4564 24734 4616
rect 18601 4539 18659 4545
rect 18601 4505 18613 4539
rect 18647 4536 18659 4539
rect 20622 4536 20628 4548
rect 18647 4508 20628 4536
rect 18647 4505 18659 4508
rect 18601 4499 18659 4505
rect 20622 4496 20628 4508
rect 20680 4496 20686 4548
rect 1104 4378 25852 4400
rect 1104 4326 7950 4378
rect 8002 4326 8014 4378
rect 8066 4326 8078 4378
rect 8130 4326 8142 4378
rect 8194 4326 8206 4378
rect 8258 4326 17950 4378
rect 18002 4326 18014 4378
rect 18066 4326 18078 4378
rect 18130 4326 18142 4378
rect 18194 4326 18206 4378
rect 18258 4326 25852 4378
rect 1104 4304 25852 4326
rect 2590 4224 2596 4276
rect 2648 4264 2654 4276
rect 8294 4264 8300 4276
rect 2648 4236 8300 4264
rect 2648 4224 2654 4236
rect 8294 4224 8300 4236
rect 8352 4224 8358 4276
rect 15102 4156 15108 4208
rect 15160 4196 15166 4208
rect 16482 4196 16488 4208
rect 15160 4168 16488 4196
rect 15160 4156 15166 4168
rect 16482 4156 16488 4168
rect 16540 4156 16546 4208
rect 1765 4131 1823 4137
rect 1765 4128 1777 4131
rect 1504 4100 1777 4128
rect 1504 3924 1532 4100
rect 1765 4097 1777 4100
rect 1811 4097 1823 4131
rect 1765 4091 1823 4097
rect 11974 4088 11980 4140
rect 12032 4088 12038 4140
rect 13538 4088 13544 4140
rect 13596 4088 13602 4140
rect 16114 4088 16120 4140
rect 16172 4088 16178 4140
rect 16206 4088 16212 4140
rect 16264 4128 16270 4140
rect 16301 4131 16359 4137
rect 16301 4128 16313 4131
rect 16264 4100 16313 4128
rect 16264 4088 16270 4100
rect 16301 4097 16313 4100
rect 16347 4097 16359 4131
rect 16301 4091 16359 4097
rect 16666 4088 16672 4140
rect 16724 4128 16730 4140
rect 16853 4131 16911 4137
rect 16853 4128 16865 4131
rect 16724 4100 16865 4128
rect 16724 4088 16730 4100
rect 16853 4097 16865 4100
rect 16899 4097 16911 4131
rect 16853 4091 16911 4097
rect 18877 4131 18935 4137
rect 18877 4097 18889 4131
rect 18923 4128 18935 4131
rect 19242 4128 19248 4140
rect 18923 4100 19248 4128
rect 18923 4097 18935 4100
rect 18877 4091 18935 4097
rect 19242 4088 19248 4100
rect 19300 4088 19306 4140
rect 19978 4088 19984 4140
rect 20036 4128 20042 4140
rect 22005 4131 22063 4137
rect 22005 4128 22017 4131
rect 20036 4100 22017 4128
rect 20036 4088 20042 4100
rect 22005 4097 22017 4100
rect 22051 4097 22063 4131
rect 22005 4091 22063 4097
rect 22830 4088 22836 4140
rect 22888 4128 22894 4140
rect 23845 4131 23903 4137
rect 23845 4128 23857 4131
rect 22888 4100 23857 4128
rect 22888 4088 22894 4100
rect 23845 4097 23857 4100
rect 23891 4097 23903 4131
rect 23845 4091 23903 4097
rect 2866 4020 2872 4072
rect 2924 4060 2930 4072
rect 5074 4060 5080 4072
rect 2924 4032 5080 4060
rect 2924 4020 2930 4032
rect 5074 4020 5080 4032
rect 5132 4020 5138 4072
rect 11333 4063 11391 4069
rect 11333 4029 11345 4063
rect 11379 4060 11391 4063
rect 11606 4060 11612 4072
rect 11379 4032 11612 4060
rect 11379 4029 11391 4032
rect 11333 4023 11391 4029
rect 11606 4020 11612 4032
rect 11664 4060 11670 4072
rect 11701 4063 11759 4069
rect 11701 4060 11713 4063
rect 11664 4032 11713 4060
rect 11664 4020 11670 4032
rect 11701 4029 11713 4032
rect 11747 4029 11759 4063
rect 11701 4023 11759 4029
rect 13446 4020 13452 4072
rect 13504 4060 13510 4072
rect 14001 4063 14059 4069
rect 14001 4060 14013 4063
rect 13504 4032 14013 4060
rect 13504 4020 13510 4032
rect 14001 4029 14013 4032
rect 14047 4029 14059 4063
rect 14001 4023 14059 4029
rect 16390 4020 16396 4072
rect 16448 4060 16454 4072
rect 17313 4063 17371 4069
rect 17313 4060 17325 4063
rect 16448 4032 17325 4060
rect 16448 4020 16454 4032
rect 17313 4029 17325 4032
rect 17359 4029 17371 4063
rect 17313 4023 17371 4029
rect 17494 4020 17500 4072
rect 17552 4060 17558 4072
rect 19153 4063 19211 4069
rect 19153 4060 19165 4063
rect 17552 4032 19165 4060
rect 17552 4020 17558 4032
rect 19153 4029 19165 4032
rect 19199 4029 19211 4063
rect 19153 4023 19211 4029
rect 20070 4020 20076 4072
rect 20128 4060 20134 4072
rect 22465 4063 22523 4069
rect 22465 4060 22477 4063
rect 20128 4032 22477 4060
rect 20128 4020 20134 4032
rect 22465 4029 22477 4032
rect 22511 4029 22523 4063
rect 22465 4023 22523 4029
rect 24305 4063 24363 4069
rect 24305 4029 24317 4063
rect 24351 4029 24363 4063
rect 24305 4023 24363 4029
rect 1581 3995 1639 4001
rect 1581 3961 1593 3995
rect 1627 3992 1639 3995
rect 2774 3992 2780 4004
rect 1627 3964 2780 3992
rect 1627 3961 1639 3964
rect 1581 3955 1639 3961
rect 2774 3952 2780 3964
rect 2832 3952 2838 4004
rect 9030 3952 9036 4004
rect 9088 3992 9094 4004
rect 9953 3995 10011 4001
rect 9953 3992 9965 3995
rect 9088 3964 9965 3992
rect 9088 3952 9094 3964
rect 9953 3961 9965 3964
rect 9999 3961 10011 3995
rect 9953 3955 10011 3961
rect 21174 3952 21180 4004
rect 21232 3992 21238 4004
rect 24320 3992 24348 4023
rect 21232 3964 24348 3992
rect 21232 3952 21238 3964
rect 2041 3927 2099 3933
rect 2041 3924 2053 3927
rect 1504 3896 2053 3924
rect 2041 3893 2053 3896
rect 2087 3924 2099 3927
rect 2866 3924 2872 3936
rect 2087 3896 2872 3924
rect 2087 3893 2099 3896
rect 2041 3887 2099 3893
rect 2866 3884 2872 3896
rect 2924 3884 2930 3936
rect 6086 3884 6092 3936
rect 6144 3924 6150 3936
rect 6365 3927 6423 3933
rect 6365 3924 6377 3927
rect 6144 3896 6377 3924
rect 6144 3884 6150 3896
rect 6365 3893 6377 3896
rect 6411 3893 6423 3927
rect 6365 3887 6423 3893
rect 9398 3884 9404 3936
rect 9456 3924 9462 3936
rect 9493 3927 9551 3933
rect 9493 3924 9505 3927
rect 9456 3896 9505 3924
rect 9456 3884 9462 3896
rect 9493 3893 9505 3896
rect 9539 3893 9551 3927
rect 9493 3887 9551 3893
rect 9766 3884 9772 3936
rect 9824 3884 9830 3936
rect 10502 3884 10508 3936
rect 10560 3924 10566 3936
rect 11057 3927 11115 3933
rect 11057 3924 11069 3927
rect 10560 3896 11069 3924
rect 10560 3884 10566 3896
rect 11057 3893 11069 3896
rect 11103 3893 11115 3927
rect 11057 3887 11115 3893
rect 19518 3884 19524 3936
rect 19576 3924 19582 3936
rect 22094 3924 22100 3936
rect 19576 3896 22100 3924
rect 19576 3884 19582 3896
rect 22094 3884 22100 3896
rect 22152 3884 22158 3936
rect 1104 3834 25852 3856
rect 1104 3782 2950 3834
rect 3002 3782 3014 3834
rect 3066 3782 3078 3834
rect 3130 3782 3142 3834
rect 3194 3782 3206 3834
rect 3258 3782 12950 3834
rect 13002 3782 13014 3834
rect 13066 3782 13078 3834
rect 13130 3782 13142 3834
rect 13194 3782 13206 3834
rect 13258 3782 22950 3834
rect 23002 3782 23014 3834
rect 23066 3782 23078 3834
rect 23130 3782 23142 3834
rect 23194 3782 23206 3834
rect 23258 3782 25852 3834
rect 1104 3760 25852 3782
rect 5261 3723 5319 3729
rect 5261 3689 5273 3723
rect 5307 3720 5319 3723
rect 5534 3720 5540 3732
rect 5307 3692 5540 3720
rect 5307 3689 5319 3692
rect 5261 3683 5319 3689
rect 5534 3680 5540 3692
rect 5592 3680 5598 3732
rect 5994 3680 6000 3732
rect 6052 3720 6058 3732
rect 6733 3723 6791 3729
rect 6733 3720 6745 3723
rect 6052 3692 6745 3720
rect 6052 3680 6058 3692
rect 6733 3689 6745 3692
rect 6779 3689 6791 3723
rect 6733 3683 6791 3689
rect 7374 3680 7380 3732
rect 7432 3720 7438 3732
rect 8205 3723 8263 3729
rect 8205 3720 8217 3723
rect 7432 3692 8217 3720
rect 7432 3680 7438 3692
rect 8205 3689 8217 3692
rect 8251 3689 8263 3723
rect 8205 3683 8263 3689
rect 9309 3723 9367 3729
rect 9309 3689 9321 3723
rect 9355 3720 9367 3723
rect 9490 3720 9496 3732
rect 9355 3692 9496 3720
rect 9355 3689 9367 3692
rect 9309 3683 9367 3689
rect 9490 3680 9496 3692
rect 9548 3680 9554 3732
rect 10042 3680 10048 3732
rect 10100 3680 10106 3732
rect 1765 3655 1823 3661
rect 1765 3621 1777 3655
rect 1811 3652 1823 3655
rect 5626 3652 5632 3664
rect 1811 3624 5632 3652
rect 1811 3621 1823 3624
rect 1765 3615 1823 3621
rect 5626 3612 5632 3624
rect 5684 3612 5690 3664
rect 5905 3655 5963 3661
rect 5905 3621 5917 3655
rect 5951 3652 5963 3655
rect 16114 3652 16120 3664
rect 5951 3624 16120 3652
rect 5951 3621 5963 3624
rect 5905 3615 5963 3621
rect 16114 3612 16120 3624
rect 16172 3612 16178 3664
rect 19150 3612 19156 3664
rect 19208 3652 19214 3664
rect 19208 3624 21312 3652
rect 19208 3612 19214 3624
rect 7561 3587 7619 3593
rect 7561 3553 7573 3587
rect 7607 3584 7619 3587
rect 8294 3584 8300 3596
rect 7607 3556 8300 3584
rect 7607 3553 7619 3556
rect 7561 3547 7619 3553
rect 8294 3544 8300 3556
rect 8352 3544 8358 3596
rect 12710 3544 12716 3596
rect 12768 3584 12774 3596
rect 12805 3587 12863 3593
rect 12805 3584 12817 3587
rect 12768 3556 12817 3584
rect 12768 3544 12774 3556
rect 12805 3553 12817 3556
rect 12851 3553 12863 3587
rect 12805 3547 12863 3553
rect 14918 3544 14924 3596
rect 14976 3584 14982 3596
rect 15473 3587 15531 3593
rect 15473 3584 15485 3587
rect 14976 3556 15485 3584
rect 14976 3544 14982 3556
rect 15473 3553 15485 3556
rect 15519 3553 15531 3587
rect 15473 3547 15531 3553
rect 16022 3544 16028 3596
rect 16080 3584 16086 3596
rect 17313 3587 17371 3593
rect 17313 3584 17325 3587
rect 16080 3556 17325 3584
rect 16080 3544 16086 3556
rect 17313 3553 17325 3556
rect 17359 3553 17371 3587
rect 17313 3547 17371 3553
rect 17770 3544 17776 3596
rect 17828 3584 17834 3596
rect 19889 3587 19947 3593
rect 19889 3584 19901 3587
rect 17828 3556 19901 3584
rect 17828 3544 17834 3556
rect 19889 3553 19901 3556
rect 19935 3553 19947 3587
rect 19889 3547 19947 3553
rect 1670 3476 1676 3528
rect 1728 3516 1734 3528
rect 1949 3519 2007 3525
rect 1949 3516 1961 3519
rect 1728 3488 1961 3516
rect 1728 3476 1734 3488
rect 1949 3485 1961 3488
rect 1995 3516 2007 3519
rect 2409 3519 2467 3525
rect 2409 3516 2421 3519
rect 1995 3488 2421 3516
rect 1995 3485 2007 3488
rect 1949 3479 2007 3485
rect 2409 3485 2421 3488
rect 2455 3485 2467 3519
rect 5077 3519 5135 3525
rect 5077 3516 5089 3519
rect 2409 3479 2467 3485
rect 4908 3488 5089 3516
rect 3145 3451 3203 3457
rect 3145 3417 3157 3451
rect 3191 3448 3203 3451
rect 3326 3448 3332 3460
rect 3191 3420 3332 3448
rect 3191 3417 3203 3420
rect 3145 3411 3203 3417
rect 3326 3408 3332 3420
rect 3384 3408 3390 3460
rect 4908 3392 4936 3488
rect 5077 3485 5089 3488
rect 5123 3485 5135 3519
rect 5077 3479 5135 3485
rect 6086 3476 6092 3528
rect 6144 3476 6150 3528
rect 6454 3476 6460 3528
rect 6512 3516 6518 3528
rect 6549 3519 6607 3525
rect 6549 3516 6561 3519
rect 6512 3488 6561 3516
rect 6512 3476 6518 3488
rect 6549 3485 6561 3488
rect 6595 3485 6607 3519
rect 8021 3519 8079 3525
rect 8021 3516 8033 3519
rect 6549 3479 6607 3485
rect 7852 3488 8033 3516
rect 7852 3392 7880 3488
rect 8021 3485 8033 3488
rect 8067 3485 8079 3519
rect 8021 3479 8079 3485
rect 9125 3519 9183 3525
rect 9125 3485 9137 3519
rect 9171 3516 9183 3519
rect 9398 3516 9404 3528
rect 9171 3488 9404 3516
rect 9171 3485 9183 3488
rect 9125 3479 9183 3485
rect 9398 3476 9404 3488
rect 9456 3476 9462 3528
rect 9766 3476 9772 3528
rect 9824 3516 9830 3528
rect 9861 3519 9919 3525
rect 9861 3516 9873 3519
rect 9824 3488 9873 3516
rect 9824 3476 9830 3488
rect 9861 3485 9873 3488
rect 9907 3485 9919 3519
rect 9861 3479 9919 3485
rect 10505 3519 10563 3525
rect 10505 3485 10517 3519
rect 10551 3516 10563 3519
rect 10870 3516 10876 3528
rect 10551 3488 10876 3516
rect 10551 3485 10563 3488
rect 10505 3479 10563 3485
rect 10870 3476 10876 3488
rect 10928 3516 10934 3528
rect 10965 3519 11023 3525
rect 10965 3516 10977 3519
rect 10928 3488 10977 3516
rect 10928 3476 10934 3488
rect 10965 3485 10977 3488
rect 11011 3485 11023 3519
rect 10965 3479 11023 3485
rect 11241 3519 11299 3525
rect 11241 3485 11253 3519
rect 11287 3485 11299 3519
rect 11241 3479 11299 3485
rect 12529 3519 12587 3525
rect 12529 3485 12541 3519
rect 12575 3516 12587 3519
rect 13630 3516 13636 3528
rect 12575 3488 13636 3516
rect 12575 3485 12587 3488
rect 12529 3479 12587 3485
rect 11256 3448 11284 3479
rect 13630 3476 13636 3488
rect 13688 3476 13694 3528
rect 15102 3476 15108 3528
rect 15160 3476 15166 3528
rect 16298 3476 16304 3528
rect 16356 3516 16362 3528
rect 16853 3519 16911 3525
rect 16853 3516 16865 3519
rect 16356 3488 16865 3516
rect 16356 3476 16362 3488
rect 16853 3485 16865 3488
rect 16899 3485 16911 3519
rect 16853 3479 16911 3485
rect 17586 3476 17592 3528
rect 17644 3516 17650 3528
rect 21284 3525 21312 3624
rect 21729 3587 21787 3593
rect 21729 3553 21741 3587
rect 21775 3553 21787 3587
rect 21729 3547 21787 3553
rect 19429 3519 19487 3525
rect 19429 3516 19441 3519
rect 17644 3488 19441 3516
rect 17644 3476 17650 3488
rect 19429 3485 19441 3488
rect 19475 3485 19487 3519
rect 19429 3479 19487 3485
rect 21269 3519 21327 3525
rect 21269 3485 21281 3519
rect 21315 3485 21327 3519
rect 21269 3479 21327 3485
rect 14734 3448 14740 3460
rect 11256 3420 14740 3448
rect 14734 3408 14740 3420
rect 14792 3408 14798 3460
rect 18966 3408 18972 3460
rect 19024 3448 19030 3460
rect 21744 3448 21772 3547
rect 19024 3420 21772 3448
rect 19024 3408 19030 3420
rect 22186 3408 22192 3460
rect 22244 3448 22250 3460
rect 24946 3448 24952 3460
rect 22244 3420 24952 3448
rect 22244 3408 22250 3420
rect 24946 3408 24952 3420
rect 25004 3408 25010 3460
rect 2038 3340 2044 3392
rect 2096 3380 2102 3392
rect 2225 3383 2283 3389
rect 2225 3380 2237 3383
rect 2096 3352 2237 3380
rect 2096 3340 2102 3352
rect 2225 3349 2237 3352
rect 2271 3349 2283 3383
rect 2225 3343 2283 3349
rect 2774 3340 2780 3392
rect 2832 3380 2838 3392
rect 2869 3383 2927 3389
rect 2869 3380 2881 3383
rect 2832 3352 2881 3380
rect 2832 3340 2838 3352
rect 2869 3349 2881 3352
rect 2915 3349 2927 3383
rect 2869 3343 2927 3349
rect 3237 3383 3295 3389
rect 3237 3349 3249 3383
rect 3283 3380 3295 3383
rect 3510 3380 3516 3392
rect 3283 3352 3516 3380
rect 3283 3349 3295 3352
rect 3237 3343 3295 3349
rect 3510 3340 3516 3352
rect 3568 3340 3574 3392
rect 3605 3383 3663 3389
rect 3605 3349 3617 3383
rect 3651 3380 3663 3383
rect 3878 3380 3884 3392
rect 3651 3352 3884 3380
rect 3651 3349 3663 3352
rect 3605 3343 3663 3349
rect 3878 3340 3884 3352
rect 3936 3340 3942 3392
rect 4801 3383 4859 3389
rect 4801 3349 4813 3383
rect 4847 3380 4859 3383
rect 4890 3380 4896 3392
rect 4847 3352 4896 3380
rect 4847 3349 4859 3352
rect 4801 3343 4859 3349
rect 4890 3340 4896 3352
rect 4948 3340 4954 3392
rect 6822 3340 6828 3392
rect 6880 3380 6886 3392
rect 7193 3383 7251 3389
rect 7193 3380 7205 3383
rect 6880 3352 7205 3380
rect 6880 3340 6886 3352
rect 7193 3349 7205 3352
rect 7239 3349 7251 3383
rect 7193 3343 7251 3349
rect 7745 3383 7803 3389
rect 7745 3349 7757 3383
rect 7791 3380 7803 3383
rect 7834 3380 7840 3392
rect 7791 3352 7840 3380
rect 7791 3349 7803 3352
rect 7745 3343 7803 3349
rect 7834 3340 7840 3352
rect 7892 3340 7898 3392
rect 8662 3340 8668 3392
rect 8720 3340 8726 3392
rect 10689 3383 10747 3389
rect 10689 3349 10701 3383
rect 10735 3380 10747 3383
rect 11238 3380 11244 3392
rect 10735 3352 11244 3380
rect 10735 3349 10747 3352
rect 10689 3343 10747 3349
rect 11238 3340 11244 3352
rect 11296 3340 11302 3392
rect 22002 3340 22008 3392
rect 22060 3380 22066 3392
rect 22830 3380 22836 3392
rect 22060 3352 22836 3380
rect 22060 3340 22066 3352
rect 22830 3340 22836 3352
rect 22888 3340 22894 3392
rect 23566 3340 23572 3392
rect 23624 3380 23630 3392
rect 24118 3380 24124 3392
rect 23624 3352 24124 3380
rect 23624 3340 23630 3352
rect 24118 3340 24124 3352
rect 24176 3380 24182 3392
rect 25409 3383 25467 3389
rect 25409 3380 25421 3383
rect 24176 3352 25421 3380
rect 24176 3340 24182 3352
rect 25409 3349 25421 3352
rect 25455 3349 25467 3383
rect 25409 3343 25467 3349
rect 1104 3290 25852 3312
rect 1104 3238 7950 3290
rect 8002 3238 8014 3290
rect 8066 3238 8078 3290
rect 8130 3238 8142 3290
rect 8194 3238 8206 3290
rect 8258 3238 17950 3290
rect 18002 3238 18014 3290
rect 18066 3238 18078 3290
rect 18130 3238 18142 3290
rect 18194 3238 18206 3290
rect 18258 3238 25852 3290
rect 1104 3216 25852 3238
rect 2682 3136 2688 3188
rect 2740 3136 2746 3188
rect 5166 3136 5172 3188
rect 5224 3136 5230 3188
rect 5902 3136 5908 3188
rect 5960 3136 5966 3188
rect 7006 3136 7012 3188
rect 7064 3136 7070 3188
rect 7282 3136 7288 3188
rect 7340 3176 7346 3188
rect 7745 3179 7803 3185
rect 7745 3176 7757 3179
rect 7340 3148 7757 3176
rect 7340 3136 7346 3148
rect 7745 3145 7757 3148
rect 7791 3145 7803 3179
rect 7745 3139 7803 3145
rect 8478 3136 8484 3188
rect 8536 3136 8542 3188
rect 11882 3136 11888 3188
rect 11940 3136 11946 3188
rect 22646 3136 22652 3188
rect 22704 3176 22710 3188
rect 24857 3179 24915 3185
rect 24857 3176 24869 3179
rect 22704 3148 24869 3176
rect 22704 3136 22710 3148
rect 24857 3145 24869 3148
rect 24903 3145 24915 3179
rect 24857 3139 24915 3145
rect 23566 3068 23572 3120
rect 23624 3068 23630 3120
rect 1857 3043 1915 3049
rect 1857 3009 1869 3043
rect 1903 3040 1915 3043
rect 2038 3040 2044 3052
rect 1903 3012 2044 3040
rect 1903 3009 1915 3012
rect 1857 3003 1915 3009
rect 2038 3000 2044 3012
rect 2096 3000 2102 3052
rect 2501 3043 2559 3049
rect 2501 3009 2513 3043
rect 2547 3040 2559 3043
rect 2774 3040 2780 3052
rect 2547 3012 2780 3040
rect 2547 3009 2559 3012
rect 2501 3003 2559 3009
rect 2774 3000 2780 3012
rect 2832 3000 2838 3052
rect 4709 3043 4767 3049
rect 4709 3009 4721 3043
rect 4755 3040 4767 3043
rect 4985 3043 5043 3049
rect 4985 3040 4997 3043
rect 4755 3012 4997 3040
rect 4755 3009 4767 3012
rect 4709 3003 4767 3009
rect 4985 3009 4997 3012
rect 5031 3040 5043 3043
rect 5350 3040 5356 3052
rect 5031 3012 5356 3040
rect 5031 3009 5043 3012
rect 4985 3003 5043 3009
rect 5350 3000 5356 3012
rect 5408 3000 5414 3052
rect 5718 3000 5724 3052
rect 5776 3000 5782 3052
rect 6822 3000 6828 3052
rect 6880 3000 6886 3052
rect 7561 3043 7619 3049
rect 7561 3009 7573 3043
rect 7607 3040 7619 3043
rect 8202 3040 8208 3052
rect 7607 3012 8208 3040
rect 7607 3009 7619 3012
rect 7561 3003 7619 3009
rect 8202 3000 8208 3012
rect 8260 3000 8266 3052
rect 8297 3043 8355 3049
rect 8297 3009 8309 3043
rect 8343 3040 8355 3043
rect 8662 3040 8668 3052
rect 8343 3012 8668 3040
rect 8343 3009 8355 3012
rect 8297 3003 8355 3009
rect 8662 3000 8668 3012
rect 8720 3000 8726 3052
rect 9306 3000 9312 3052
rect 9364 3000 9370 3052
rect 10594 3000 10600 3052
rect 10652 3000 10658 3052
rect 11238 3000 11244 3052
rect 11296 3040 11302 3052
rect 11701 3043 11759 3049
rect 11701 3040 11713 3043
rect 11296 3012 11713 3040
rect 11296 3000 11302 3012
rect 11701 3009 11713 3012
rect 11747 3009 11759 3043
rect 11701 3003 11759 3009
rect 12618 3000 12624 3052
rect 12676 3000 12682 3052
rect 14274 3000 14280 3052
rect 14332 3000 14338 3052
rect 16758 3000 16764 3052
rect 16816 3040 16822 3052
rect 16853 3043 16911 3049
rect 16853 3040 16865 3043
rect 16816 3012 16865 3040
rect 16816 3000 16822 3012
rect 16853 3009 16865 3012
rect 16899 3009 16911 3043
rect 16853 3003 16911 3009
rect 17862 3000 17868 3052
rect 17920 3040 17926 3052
rect 18506 3040 18512 3052
rect 17920 3012 18512 3040
rect 17920 3000 17926 3012
rect 18506 3000 18512 3012
rect 18564 3040 18570 3052
rect 18693 3043 18751 3049
rect 18693 3040 18705 3043
rect 18564 3012 18705 3040
rect 18564 3000 18570 3012
rect 18693 3009 18705 3012
rect 18739 3009 18751 3043
rect 18693 3003 18751 3009
rect 21726 3000 21732 3052
rect 21784 3040 21790 3052
rect 22646 3040 22652 3052
rect 21784 3012 22652 3040
rect 21784 3000 21790 3012
rect 22646 3000 22652 3012
rect 22704 3000 22710 3052
rect 3237 2975 3295 2981
rect 3237 2941 3249 2975
rect 3283 2972 3295 2975
rect 3326 2972 3332 2984
rect 3283 2944 3332 2972
rect 3283 2941 3295 2944
rect 3237 2935 3295 2941
rect 3326 2932 3332 2944
rect 3384 2932 3390 2984
rect 3513 2975 3571 2981
rect 3513 2941 3525 2975
rect 3559 2972 3571 2975
rect 7742 2972 7748 2984
rect 3559 2944 7748 2972
rect 3559 2941 3571 2944
rect 3513 2935 3571 2941
rect 7742 2932 7748 2944
rect 7800 2932 7806 2984
rect 9030 2932 9036 2984
rect 9088 2932 9094 2984
rect 10321 2975 10379 2981
rect 10321 2941 10333 2975
rect 10367 2972 10379 2975
rect 10502 2972 10508 2984
rect 10367 2944 10508 2972
rect 10367 2941 10379 2944
rect 10321 2935 10379 2941
rect 10502 2932 10508 2944
rect 10560 2932 10566 2984
rect 13354 2932 13360 2984
rect 13412 2932 13418 2984
rect 14182 2932 14188 2984
rect 14240 2972 14246 2984
rect 14737 2975 14795 2981
rect 14737 2972 14749 2975
rect 14240 2944 14749 2972
rect 14240 2932 14246 2944
rect 14737 2941 14749 2944
rect 14783 2941 14795 2975
rect 14737 2935 14795 2941
rect 15654 2932 15660 2984
rect 15712 2972 15718 2984
rect 17313 2975 17371 2981
rect 17313 2972 17325 2975
rect 15712 2944 17325 2972
rect 15712 2932 15718 2944
rect 17313 2941 17325 2944
rect 17359 2941 17371 2975
rect 17313 2935 17371 2941
rect 19153 2975 19211 2981
rect 19153 2941 19165 2975
rect 19199 2941 19211 2975
rect 19153 2935 19211 2941
rect 2041 2907 2099 2913
rect 2041 2873 2053 2907
rect 2087 2904 2099 2907
rect 5810 2904 5816 2916
rect 2087 2876 5816 2904
rect 2087 2873 2099 2876
rect 2041 2867 2099 2873
rect 5810 2864 5816 2876
rect 5868 2864 5874 2916
rect 17126 2864 17132 2916
rect 17184 2904 17190 2916
rect 19168 2904 19196 2935
rect 20622 2932 20628 2984
rect 20680 2972 20686 2984
rect 23382 2972 23388 2984
rect 20680 2944 23388 2972
rect 20680 2932 20686 2944
rect 23382 2932 23388 2944
rect 23440 2932 23446 2984
rect 17184 2876 19196 2904
rect 17184 2864 17190 2876
rect 19702 2864 19708 2916
rect 19760 2904 19766 2916
rect 20714 2904 20720 2916
rect 19760 2876 20720 2904
rect 19760 2864 19766 2876
rect 20714 2864 20720 2876
rect 20772 2864 20778 2916
rect 1486 2796 1492 2848
rect 1544 2796 1550 2848
rect 4246 2796 4252 2848
rect 4304 2836 4310 2848
rect 4341 2839 4399 2845
rect 4341 2836 4353 2839
rect 4304 2808 4353 2836
rect 4304 2796 4310 2808
rect 4341 2805 4353 2808
rect 4387 2805 4399 2839
rect 4341 2799 4399 2805
rect 6454 2796 6460 2848
rect 6512 2796 6518 2848
rect 18598 2796 18604 2848
rect 18656 2836 18662 2848
rect 19886 2836 19892 2848
rect 18656 2808 19892 2836
rect 18656 2796 18662 2808
rect 19886 2796 19892 2808
rect 19944 2796 19950 2848
rect 20806 2796 20812 2848
rect 20864 2836 20870 2848
rect 22462 2836 22468 2848
rect 20864 2808 22468 2836
rect 20864 2796 20870 2808
rect 22462 2796 22468 2808
rect 22520 2796 22526 2848
rect 1104 2746 25852 2768
rect 1104 2694 2950 2746
rect 3002 2694 3014 2746
rect 3066 2694 3078 2746
rect 3130 2694 3142 2746
rect 3194 2694 3206 2746
rect 3258 2694 12950 2746
rect 13002 2694 13014 2746
rect 13066 2694 13078 2746
rect 13130 2694 13142 2746
rect 13194 2694 13206 2746
rect 13258 2694 22950 2746
rect 23002 2694 23014 2746
rect 23066 2694 23078 2746
rect 23130 2694 23142 2746
rect 23194 2694 23206 2746
rect 23258 2694 25852 2746
rect 1104 2672 25852 2694
rect 1854 2592 1860 2644
rect 1912 2592 1918 2644
rect 2590 2592 2596 2644
rect 2648 2592 2654 2644
rect 3329 2635 3387 2641
rect 3329 2601 3341 2635
rect 3375 2632 3387 2635
rect 4798 2632 4804 2644
rect 3375 2604 4804 2632
rect 3375 2601 3387 2604
rect 3329 2595 3387 2601
rect 4798 2592 4804 2604
rect 4856 2592 4862 2644
rect 7101 2635 7159 2641
rect 7101 2601 7113 2635
rect 7147 2632 7159 2635
rect 7650 2632 7656 2644
rect 7147 2604 7656 2632
rect 7147 2601 7159 2604
rect 7101 2595 7159 2601
rect 7650 2592 7656 2604
rect 7708 2592 7714 2644
rect 9769 2635 9827 2641
rect 9769 2601 9781 2635
rect 9815 2632 9827 2635
rect 11054 2632 11060 2644
rect 9815 2604 11060 2632
rect 9815 2601 9827 2604
rect 9769 2595 9827 2601
rect 11054 2592 11060 2604
rect 11112 2592 11118 2644
rect 11701 2635 11759 2641
rect 11701 2601 11713 2635
rect 11747 2632 11759 2635
rect 15746 2632 15752 2644
rect 11747 2604 15752 2632
rect 11747 2601 11759 2604
rect 11701 2595 11759 2601
rect 15746 2592 15752 2604
rect 15804 2592 15810 2644
rect 17402 2592 17408 2644
rect 17460 2632 17466 2644
rect 17460 2604 22048 2632
rect 17460 2592 17466 2604
rect 4157 2567 4215 2573
rect 4157 2533 4169 2567
rect 4203 2564 4215 2567
rect 7558 2564 7564 2576
rect 4203 2536 7564 2564
rect 4203 2533 4215 2536
rect 4157 2527 4215 2533
rect 7558 2524 7564 2536
rect 7616 2524 7622 2576
rect 12802 2564 12808 2576
rect 10612 2536 12808 2564
rect 4982 2456 4988 2508
rect 5040 2456 5046 2508
rect 10612 2505 10640 2536
rect 12802 2524 12808 2536
rect 12860 2524 12866 2576
rect 14826 2524 14832 2576
rect 14884 2564 14890 2576
rect 14884 2536 19472 2564
rect 14884 2524 14890 2536
rect 7929 2499 7987 2505
rect 7929 2465 7941 2499
rect 7975 2496 7987 2499
rect 10597 2499 10655 2505
rect 7975 2468 10548 2496
rect 7975 2465 7987 2468
rect 7929 2459 7987 2465
rect 1486 2388 1492 2440
rect 1544 2428 1550 2440
rect 1673 2431 1731 2437
rect 1673 2428 1685 2431
rect 1544 2400 1685 2428
rect 1544 2388 1550 2400
rect 1673 2397 1685 2400
rect 1719 2428 1731 2431
rect 2314 2428 2320 2440
rect 1719 2400 2320 2428
rect 1719 2397 1731 2400
rect 1673 2391 1731 2397
rect 2314 2388 2320 2400
rect 2372 2388 2378 2440
rect 2409 2431 2467 2437
rect 2409 2397 2421 2431
rect 2455 2428 2467 2431
rect 3510 2428 3516 2440
rect 2455 2400 3516 2428
rect 2455 2397 2467 2400
rect 2409 2391 2467 2397
rect 3510 2388 3516 2400
rect 3568 2388 3574 2440
rect 3973 2431 4031 2437
rect 3973 2397 3985 2431
rect 4019 2428 4031 2431
rect 4246 2428 4252 2440
rect 4019 2400 4252 2428
rect 4019 2397 4031 2400
rect 3973 2391 4031 2397
rect 4246 2388 4252 2400
rect 4304 2388 4310 2440
rect 4614 2388 4620 2440
rect 4672 2428 4678 2440
rect 4709 2431 4767 2437
rect 4709 2428 4721 2431
rect 4672 2400 4721 2428
rect 4672 2388 4678 2400
rect 4709 2397 4721 2400
rect 4755 2428 4767 2431
rect 5813 2431 5871 2437
rect 5813 2428 5825 2431
rect 4755 2400 5825 2428
rect 4755 2397 4767 2400
rect 4709 2391 4767 2397
rect 5813 2397 5825 2400
rect 5859 2397 5871 2431
rect 5813 2391 5871 2397
rect 6457 2431 6515 2437
rect 6457 2397 6469 2431
rect 6503 2428 6515 2431
rect 6917 2431 6975 2437
rect 6917 2428 6929 2431
rect 6503 2400 6929 2428
rect 6503 2397 6515 2400
rect 6457 2391 6515 2397
rect 6917 2397 6929 2400
rect 6963 2428 6975 2431
rect 7190 2428 7196 2440
rect 6963 2400 7196 2428
rect 6963 2397 6975 2400
rect 6917 2391 6975 2397
rect 7190 2388 7196 2400
rect 7248 2388 7254 2440
rect 7558 2388 7564 2440
rect 7616 2428 7622 2440
rect 7653 2431 7711 2437
rect 7653 2428 7665 2431
rect 7616 2400 7665 2428
rect 7616 2388 7622 2400
rect 7653 2397 7665 2400
rect 7699 2397 7711 2431
rect 7653 2391 7711 2397
rect 9125 2431 9183 2437
rect 9125 2397 9137 2431
rect 9171 2428 9183 2431
rect 9585 2431 9643 2437
rect 9585 2428 9597 2431
rect 9171 2400 9597 2428
rect 9171 2397 9183 2400
rect 9125 2391 9183 2397
rect 9585 2397 9597 2400
rect 9631 2428 9643 2431
rect 10134 2428 10140 2440
rect 9631 2400 10140 2428
rect 9631 2397 9643 2400
rect 9585 2391 9643 2397
rect 10134 2388 10140 2400
rect 10192 2388 10198 2440
rect 10321 2431 10379 2437
rect 10321 2397 10333 2431
rect 10367 2397 10379 2431
rect 10520 2428 10548 2468
rect 10597 2465 10609 2499
rect 10643 2465 10655 2499
rect 11974 2496 11980 2508
rect 10597 2459 10655 2465
rect 11900 2468 11980 2496
rect 11698 2428 11704 2440
rect 10520 2400 11704 2428
rect 10321 2391 10379 2397
rect 3237 2363 3295 2369
rect 3237 2329 3249 2363
rect 3283 2360 3295 2363
rect 3878 2360 3884 2372
rect 3283 2332 3884 2360
rect 3283 2329 3295 2332
rect 3237 2323 3295 2329
rect 3878 2320 3884 2332
rect 3936 2320 3942 2372
rect 5718 2320 5724 2372
rect 5776 2360 5782 2372
rect 6089 2363 6147 2369
rect 6089 2360 6101 2363
rect 5776 2332 6101 2360
rect 5776 2320 5782 2332
rect 6089 2329 6101 2332
rect 6135 2329 6147 2363
rect 6089 2323 6147 2329
rect 6641 2363 6699 2369
rect 6641 2329 6653 2363
rect 6687 2360 6699 2363
rect 7576 2360 7604 2388
rect 6687 2332 7604 2360
rect 9309 2363 9367 2369
rect 6687 2329 6699 2332
rect 6641 2323 6699 2329
rect 9309 2329 9321 2363
rect 9355 2360 9367 2363
rect 10336 2360 10364 2391
rect 11698 2388 11704 2400
rect 11756 2388 11762 2440
rect 11900 2437 11928 2468
rect 11974 2456 11980 2468
rect 12032 2496 12038 2508
rect 14093 2499 14151 2505
rect 14093 2496 14105 2499
rect 12032 2468 14105 2496
rect 12032 2456 12038 2468
rect 14093 2465 14105 2468
rect 14139 2465 14151 2499
rect 14093 2459 14151 2465
rect 14550 2456 14556 2508
rect 14608 2496 14614 2508
rect 15197 2499 15255 2505
rect 15197 2496 15209 2499
rect 14608 2468 15209 2496
rect 14608 2456 14614 2468
rect 15197 2465 15209 2468
rect 15243 2465 15255 2499
rect 15197 2459 15255 2465
rect 15286 2456 15292 2508
rect 15344 2496 15350 2508
rect 17313 2499 17371 2505
rect 17313 2496 17325 2499
rect 15344 2468 17325 2496
rect 15344 2456 15350 2468
rect 17313 2465 17325 2468
rect 17359 2465 17371 2499
rect 17313 2459 17371 2465
rect 18506 2456 18512 2508
rect 18564 2456 18570 2508
rect 11885 2431 11943 2437
rect 11885 2397 11897 2431
rect 11931 2397 11943 2431
rect 11885 2391 11943 2397
rect 12526 2388 12532 2440
rect 12584 2388 12590 2440
rect 14642 2388 14648 2440
rect 14700 2388 14706 2440
rect 16942 2388 16948 2440
rect 17000 2388 17006 2440
rect 19444 2437 19472 2536
rect 19889 2499 19947 2505
rect 19889 2465 19901 2499
rect 19935 2465 19947 2499
rect 19889 2459 19947 2465
rect 19429 2431 19487 2437
rect 19429 2397 19441 2431
rect 19475 2397 19487 2431
rect 19429 2391 19487 2397
rect 12342 2360 12348 2372
rect 9355 2332 12348 2360
rect 9355 2329 9367 2332
rect 9309 2323 9367 2329
rect 12342 2320 12348 2332
rect 12400 2320 12406 2372
rect 13541 2363 13599 2369
rect 13541 2329 13553 2363
rect 13587 2360 13599 2363
rect 13814 2360 13820 2372
rect 13587 2332 13820 2360
rect 13587 2329 13599 2332
rect 13541 2323 13599 2329
rect 13814 2320 13820 2332
rect 13872 2320 13878 2372
rect 16758 2320 16764 2372
rect 16816 2360 16822 2372
rect 19904 2360 19932 2459
rect 22020 2437 22048 2604
rect 22465 2499 22523 2505
rect 22465 2465 22477 2499
rect 22511 2465 22523 2499
rect 22465 2459 22523 2465
rect 22005 2431 22063 2437
rect 22005 2397 22017 2431
rect 22051 2397 22063 2431
rect 22005 2391 22063 2397
rect 16816 2332 19932 2360
rect 16816 2320 16822 2332
rect 18322 2252 18328 2304
rect 18380 2292 18386 2304
rect 22480 2292 22508 2459
rect 25314 2388 25320 2440
rect 25372 2388 25378 2440
rect 18380 2264 22508 2292
rect 18380 2252 18386 2264
rect 1104 2202 25852 2224
rect 1104 2150 7950 2202
rect 8002 2150 8014 2202
rect 8066 2150 8078 2202
rect 8130 2150 8142 2202
rect 8194 2150 8206 2202
rect 8258 2150 17950 2202
rect 18002 2150 18014 2202
rect 18066 2150 18078 2202
rect 18130 2150 18142 2202
rect 18194 2150 18206 2202
rect 18258 2150 25852 2202
rect 1104 2128 25852 2150
<< via1 >>
rect 7950 54374 8002 54426
rect 8014 54374 8066 54426
rect 8078 54374 8130 54426
rect 8142 54374 8194 54426
rect 8206 54374 8258 54426
rect 17950 54374 18002 54426
rect 18014 54374 18066 54426
rect 18078 54374 18130 54426
rect 18142 54374 18194 54426
rect 18206 54374 18258 54426
rect 9956 54272 10008 54324
rect 14740 54272 14792 54324
rect 16212 54272 16264 54324
rect 7840 54204 7892 54256
rect 11428 54204 11480 54256
rect 4344 54136 4396 54188
rect 4620 54179 4672 54188
rect 4620 54145 4629 54179
rect 4629 54145 4663 54179
rect 4663 54145 4672 54179
rect 4620 54136 4672 54145
rect 5908 54068 5960 54120
rect 9956 54179 10008 54188
rect 9956 54145 9965 54179
rect 9965 54145 9999 54179
rect 9999 54145 10008 54179
rect 9956 54136 10008 54145
rect 12900 54204 12952 54256
rect 12348 54179 12400 54188
rect 12348 54145 12357 54179
rect 12357 54145 12391 54179
rect 12391 54145 12400 54179
rect 12348 54136 12400 54145
rect 15200 54136 15252 54188
rect 24492 54315 24544 54324
rect 24492 54281 24501 54315
rect 24501 54281 24535 54315
rect 24535 54281 24544 54315
rect 24492 54272 24544 54281
rect 24676 54315 24728 54324
rect 24676 54281 24685 54315
rect 24685 54281 24719 54315
rect 24719 54281 24728 54315
rect 24676 54272 24728 54281
rect 17684 54204 17736 54256
rect 18880 54204 18932 54256
rect 16948 54136 17000 54188
rect 10232 54068 10284 54120
rect 12532 54068 12584 54120
rect 18420 54068 18472 54120
rect 19524 54136 19576 54188
rect 20720 54136 20772 54188
rect 21364 54136 21416 54188
rect 22468 54136 22520 54188
rect 25044 54179 25096 54188
rect 25044 54145 25053 54179
rect 25053 54145 25087 54179
rect 25087 54145 25096 54179
rect 25044 54136 25096 54145
rect 19708 54068 19760 54120
rect 16212 54000 16264 54052
rect 11704 53975 11756 53984
rect 11704 53941 11713 53975
rect 11713 53941 11747 53975
rect 11747 53941 11756 53975
rect 11704 53932 11756 53941
rect 15752 53975 15804 53984
rect 15752 53941 15761 53975
rect 15761 53941 15795 53975
rect 15795 53941 15804 53975
rect 15752 53932 15804 53941
rect 16120 53932 16172 53984
rect 19340 54000 19392 54052
rect 22284 54000 22336 54052
rect 17040 53975 17092 53984
rect 17040 53941 17049 53975
rect 17049 53941 17083 53975
rect 17083 53941 17092 53975
rect 17040 53932 17092 53941
rect 18420 53932 18472 53984
rect 19432 53932 19484 53984
rect 21088 53975 21140 53984
rect 21088 53941 21097 53975
rect 21097 53941 21131 53975
rect 21131 53941 21140 53975
rect 21088 53932 21140 53941
rect 22192 53975 22244 53984
rect 22192 53941 22201 53975
rect 22201 53941 22235 53975
rect 22235 53941 22244 53975
rect 22192 53932 22244 53941
rect 22376 53932 22428 53984
rect 23572 53932 23624 53984
rect 2950 53830 3002 53882
rect 3014 53830 3066 53882
rect 3078 53830 3130 53882
rect 3142 53830 3194 53882
rect 3206 53830 3258 53882
rect 12950 53830 13002 53882
rect 13014 53830 13066 53882
rect 13078 53830 13130 53882
rect 13142 53830 13194 53882
rect 13206 53830 13258 53882
rect 22950 53830 23002 53882
rect 23014 53830 23066 53882
rect 23078 53830 23130 53882
rect 23142 53830 23194 53882
rect 23206 53830 23258 53882
rect 16580 53728 16632 53780
rect 18880 53771 18932 53780
rect 18880 53737 18889 53771
rect 18889 53737 18923 53771
rect 18923 53737 18932 53771
rect 18880 53728 18932 53737
rect 5540 53660 5592 53712
rect 21916 53660 21968 53712
rect 22376 53660 22428 53712
rect 7380 53592 7432 53644
rect 8852 53592 8904 53644
rect 11060 53635 11112 53644
rect 11060 53601 11069 53635
rect 11069 53601 11103 53635
rect 11103 53601 11112 53635
rect 11060 53592 11112 53601
rect 12164 53592 12216 53644
rect 6828 53524 6880 53576
rect 9128 53524 9180 53576
rect 10324 53524 10376 53576
rect 12624 53524 12676 53576
rect 14004 53524 14056 53576
rect 15476 53524 15528 53576
rect 16580 53524 16632 53576
rect 17316 53524 17368 53576
rect 18328 53524 18380 53576
rect 19156 53524 19208 53576
rect 19892 53524 19944 53576
rect 20996 53524 21048 53576
rect 21732 53524 21784 53576
rect 22100 53524 22152 53576
rect 22836 53524 22888 53576
rect 24492 53524 24544 53576
rect 24768 53524 24820 53576
rect 7564 53456 7616 53508
rect 18512 53456 18564 53508
rect 20628 53456 20680 53508
rect 14464 53431 14516 53440
rect 14464 53397 14473 53431
rect 14473 53397 14507 53431
rect 14507 53397 14516 53431
rect 14464 53388 14516 53397
rect 15752 53431 15804 53440
rect 15752 53397 15761 53431
rect 15761 53397 15795 53431
rect 15795 53397 15804 53431
rect 15752 53388 15804 53397
rect 16856 53431 16908 53440
rect 16856 53397 16865 53431
rect 16865 53397 16899 53431
rect 16899 53397 16908 53431
rect 16856 53388 16908 53397
rect 17408 53431 17460 53440
rect 17408 53397 17417 53431
rect 17417 53397 17451 53431
rect 17451 53397 17460 53431
rect 17408 53388 17460 53397
rect 19616 53431 19668 53440
rect 19616 53397 19625 53431
rect 19625 53397 19659 53431
rect 19659 53397 19668 53431
rect 19616 53388 19668 53397
rect 20904 53388 20956 53440
rect 22468 53431 22520 53440
rect 22468 53397 22477 53431
rect 22477 53397 22511 53431
rect 22511 53397 22520 53431
rect 22468 53388 22520 53397
rect 23940 53431 23992 53440
rect 23940 53397 23949 53431
rect 23949 53397 23983 53431
rect 23983 53397 23992 53431
rect 23940 53388 23992 53397
rect 25044 53431 25096 53440
rect 25044 53397 25053 53431
rect 25053 53397 25087 53431
rect 25087 53397 25096 53431
rect 25044 53388 25096 53397
rect 7950 53286 8002 53338
rect 8014 53286 8066 53338
rect 8078 53286 8130 53338
rect 8142 53286 8194 53338
rect 8206 53286 8258 53338
rect 17950 53286 18002 53338
rect 18014 53286 18066 53338
rect 18078 53286 18130 53338
rect 18142 53286 18194 53338
rect 18206 53286 18258 53338
rect 2780 53184 2832 53236
rect 5172 53184 5224 53236
rect 5724 53184 5776 53236
rect 17316 53227 17368 53236
rect 17316 53193 17325 53227
rect 17325 53193 17359 53227
rect 17359 53193 17368 53227
rect 17316 53184 17368 53193
rect 19156 53184 19208 53236
rect 19708 53227 19760 53236
rect 19708 53193 19717 53227
rect 19717 53193 19751 53227
rect 19751 53193 19760 53227
rect 19708 53184 19760 53193
rect 20996 53227 21048 53236
rect 20996 53193 21005 53227
rect 21005 53193 21039 53227
rect 21039 53193 21048 53227
rect 20996 53184 21048 53193
rect 21732 53184 21784 53236
rect 22100 53184 22152 53236
rect 22560 53227 22612 53236
rect 22560 53193 22569 53227
rect 22569 53193 22603 53227
rect 22603 53193 22612 53227
rect 22560 53184 22612 53193
rect 23296 53184 23348 53236
rect 4436 53116 4488 53168
rect 6276 53116 6328 53168
rect 9220 53116 9272 53168
rect 6460 53048 6512 53100
rect 10968 53116 11020 53168
rect 13636 53116 13688 53168
rect 20720 53116 20772 53168
rect 9772 53091 9824 53100
rect 9772 53057 9781 53091
rect 9781 53057 9815 53091
rect 9815 53057 9824 53091
rect 9772 53048 9824 53057
rect 11888 53091 11940 53100
rect 11888 53057 11897 53091
rect 11897 53057 11931 53091
rect 11931 53057 11940 53091
rect 11888 53048 11940 53057
rect 14372 53048 14424 53100
rect 15844 53048 15896 53100
rect 18788 53048 18840 53100
rect 20260 53048 20312 53100
rect 23664 53048 23716 53100
rect 25044 53091 25096 53100
rect 25044 53057 25053 53091
rect 25053 53057 25087 53091
rect 25087 53057 25096 53091
rect 25044 53048 25096 53057
rect 5540 52980 5592 53032
rect 10416 53023 10468 53032
rect 10416 52989 10425 53023
rect 10425 52989 10459 53023
rect 10459 52989 10468 53023
rect 10416 52980 10468 52989
rect 11796 52980 11848 53032
rect 3424 52912 3476 52964
rect 9588 52912 9640 52964
rect 14004 52955 14056 52964
rect 14004 52921 14013 52955
rect 14013 52921 14047 52955
rect 14047 52921 14056 52955
rect 14004 52912 14056 52921
rect 4068 52844 4120 52896
rect 14648 52844 14700 52896
rect 15936 52887 15988 52896
rect 15936 52853 15945 52887
rect 15945 52853 15979 52887
rect 15979 52853 15988 52887
rect 15936 52844 15988 52853
rect 18604 52844 18656 52896
rect 20352 52887 20404 52896
rect 20352 52853 20361 52887
rect 20361 52853 20395 52887
rect 20395 52853 20404 52887
rect 20352 52844 20404 52853
rect 22560 52844 22612 52896
rect 23940 52887 23992 52896
rect 23940 52853 23949 52887
rect 23949 52853 23983 52887
rect 23983 52853 23992 52887
rect 23940 52844 23992 52853
rect 24860 52844 24912 52896
rect 2950 52742 3002 52794
rect 3014 52742 3066 52794
rect 3078 52742 3130 52794
rect 3142 52742 3194 52794
rect 3206 52742 3258 52794
rect 12950 52742 13002 52794
rect 13014 52742 13066 52794
rect 13078 52742 13130 52794
rect 13142 52742 13194 52794
rect 13206 52742 13258 52794
rect 22950 52742 23002 52794
rect 23014 52742 23066 52794
rect 23078 52742 23130 52794
rect 23142 52742 23194 52794
rect 23206 52742 23258 52794
rect 2228 52640 2280 52692
rect 3424 52640 3476 52692
rect 12624 52683 12676 52692
rect 12624 52649 12633 52683
rect 12633 52649 12667 52683
rect 12667 52649 12676 52683
rect 12624 52640 12676 52649
rect 13636 52640 13688 52692
rect 24768 52640 24820 52692
rect 1860 52572 1912 52624
rect 3516 52572 3568 52624
rect 25136 52572 25188 52624
rect 3700 52504 3752 52556
rect 6644 52504 6696 52556
rect 7748 52547 7800 52556
rect 7748 52513 7757 52547
rect 7757 52513 7791 52547
rect 7791 52513 7800 52547
rect 7748 52504 7800 52513
rect 10692 52504 10744 52556
rect 13636 52547 13688 52556
rect 13636 52513 13645 52547
rect 13645 52513 13679 52547
rect 13679 52513 13688 52547
rect 13636 52504 13688 52513
rect 4804 52436 4856 52488
rect 5632 52436 5684 52488
rect 7196 52479 7248 52488
rect 7196 52445 7205 52479
rect 7205 52445 7239 52479
rect 7239 52445 7248 52479
rect 7196 52436 7248 52445
rect 10784 52479 10836 52488
rect 10784 52445 10793 52479
rect 10793 52445 10827 52479
rect 10827 52445 10836 52479
rect 10784 52436 10836 52445
rect 12808 52479 12860 52488
rect 12808 52445 12817 52479
rect 12817 52445 12851 52479
rect 12851 52445 12860 52479
rect 12808 52436 12860 52445
rect 24768 52479 24820 52488
rect 24768 52445 24777 52479
rect 24777 52445 24811 52479
rect 24811 52445 24820 52479
rect 24768 52436 24820 52445
rect 13360 52368 13412 52420
rect 7950 52198 8002 52250
rect 8014 52198 8066 52250
rect 8078 52198 8130 52250
rect 8142 52198 8194 52250
rect 8206 52198 8258 52250
rect 17950 52198 18002 52250
rect 18014 52198 18066 52250
rect 18078 52198 18130 52250
rect 18142 52198 18194 52250
rect 18206 52198 18258 52250
rect 5540 52096 5592 52148
rect 11888 52096 11940 52148
rect 12348 52139 12400 52148
rect 12348 52105 12357 52139
rect 12357 52105 12391 52139
rect 12391 52105 12400 52139
rect 12348 52096 12400 52105
rect 13360 52096 13412 52148
rect 25320 52139 25372 52148
rect 25320 52105 25329 52139
rect 25329 52105 25363 52139
rect 25363 52105 25372 52139
rect 25320 52096 25372 52105
rect 9220 52028 9272 52080
rect 4528 51960 4580 52012
rect 4988 51960 5040 52012
rect 7380 51960 7432 52012
rect 9864 52003 9916 52012
rect 9864 51969 9873 52003
rect 9873 51969 9907 52003
rect 9907 51969 9916 52003
rect 9864 51960 9916 51969
rect 11888 52003 11940 52012
rect 11888 51969 11897 52003
rect 11897 51969 11931 52003
rect 11931 51969 11940 52003
rect 11888 51960 11940 51969
rect 11980 51960 12032 52012
rect 3332 51935 3384 51944
rect 3332 51901 3341 51935
rect 3341 51901 3375 51935
rect 3375 51901 3384 51935
rect 3332 51892 3384 51901
rect 4896 51892 4948 51944
rect 8484 51935 8536 51944
rect 8484 51901 8493 51935
rect 8493 51901 8527 51935
rect 8527 51901 8536 51935
rect 8484 51892 8536 51901
rect 9680 51892 9732 51944
rect 25504 51799 25556 51808
rect 25504 51765 25513 51799
rect 25513 51765 25547 51799
rect 25547 51765 25556 51799
rect 25504 51756 25556 51765
rect 2950 51654 3002 51706
rect 3014 51654 3066 51706
rect 3078 51654 3130 51706
rect 3142 51654 3194 51706
rect 3206 51654 3258 51706
rect 12950 51654 13002 51706
rect 13014 51654 13066 51706
rect 13078 51654 13130 51706
rect 13142 51654 13194 51706
rect 13206 51654 13258 51706
rect 22950 51654 23002 51706
rect 23014 51654 23066 51706
rect 23078 51654 23130 51706
rect 23142 51654 23194 51706
rect 23206 51654 23258 51706
rect 9956 51552 10008 51604
rect 2872 51459 2924 51468
rect 2872 51425 2881 51459
rect 2881 51425 2915 51459
rect 2915 51425 2924 51459
rect 2872 51416 2924 51425
rect 5724 51459 5776 51468
rect 5724 51425 5733 51459
rect 5733 51425 5767 51459
rect 5767 51425 5776 51459
rect 5724 51416 5776 51425
rect 7012 51416 7064 51468
rect 6736 51348 6788 51400
rect 7104 51391 7156 51400
rect 7104 51357 7113 51391
rect 7113 51357 7147 51391
rect 7147 51357 7156 51391
rect 7104 51348 7156 51357
rect 9312 51348 9364 51400
rect 25504 51348 25556 51400
rect 5540 51280 5592 51332
rect 24952 51212 25004 51264
rect 7950 51110 8002 51162
rect 8014 51110 8066 51162
rect 8078 51110 8130 51162
rect 8142 51110 8194 51162
rect 8206 51110 8258 51162
rect 17950 51110 18002 51162
rect 18014 51110 18066 51162
rect 18078 51110 18130 51162
rect 18142 51110 18194 51162
rect 18206 51110 18258 51162
rect 4344 51008 4396 51060
rect 5540 51008 5592 51060
rect 4160 50872 4212 50924
rect 4344 50915 4396 50924
rect 4344 50881 4353 50915
rect 4353 50881 4387 50915
rect 4387 50881 4396 50915
rect 4344 50872 4396 50881
rect 7656 50872 7708 50924
rect 10784 50940 10836 50992
rect 9404 50915 9456 50924
rect 9404 50881 9413 50915
rect 9413 50881 9447 50915
rect 9447 50881 9456 50915
rect 9404 50872 9456 50881
rect 25044 50915 25096 50924
rect 25044 50881 25053 50915
rect 25053 50881 25087 50915
rect 25087 50881 25096 50915
rect 25044 50872 25096 50881
rect 2780 50847 2832 50856
rect 2780 50813 2789 50847
rect 2789 50813 2823 50847
rect 2823 50813 2832 50847
rect 2780 50804 2832 50813
rect 4252 50804 4304 50856
rect 7472 50847 7524 50856
rect 7472 50813 7481 50847
rect 7481 50813 7515 50847
rect 7515 50813 7524 50847
rect 7472 50804 7524 50813
rect 24308 50668 24360 50720
rect 2950 50566 3002 50618
rect 3014 50566 3066 50618
rect 3078 50566 3130 50618
rect 3142 50566 3194 50618
rect 3206 50566 3258 50618
rect 12950 50566 13002 50618
rect 13014 50566 13066 50618
rect 13078 50566 13130 50618
rect 13142 50566 13194 50618
rect 13206 50566 13258 50618
rect 22950 50566 23002 50618
rect 23014 50566 23066 50618
rect 23078 50566 23130 50618
rect 23142 50566 23194 50618
rect 23206 50566 23258 50618
rect 6828 50507 6880 50516
rect 6828 50473 6837 50507
rect 6837 50473 6871 50507
rect 6871 50473 6880 50507
rect 6828 50464 6880 50473
rect 9128 50464 9180 50516
rect 21456 50396 21508 50448
rect 3424 50328 3476 50380
rect 4712 50260 4764 50312
rect 5816 50260 5868 50312
rect 8392 50260 8444 50312
rect 25320 50303 25372 50312
rect 25320 50269 25329 50303
rect 25329 50269 25363 50303
rect 25363 50269 25372 50303
rect 25320 50260 25372 50269
rect 24492 50124 24544 50176
rect 7950 50022 8002 50074
rect 8014 50022 8066 50074
rect 8078 50022 8130 50074
rect 8142 50022 8194 50074
rect 8206 50022 8258 50074
rect 17950 50022 18002 50074
rect 18014 50022 18066 50074
rect 18078 50022 18130 50074
rect 18142 50022 18194 50074
rect 18206 50022 18258 50074
rect 3516 49852 3568 49904
rect 3608 49784 3660 49836
rect 6828 49920 6880 49972
rect 8484 49852 8536 49904
rect 9772 49852 9824 49904
rect 7840 49784 7892 49836
rect 21640 49784 21692 49836
rect 8760 49716 8812 49768
rect 24492 49759 24544 49768
rect 24492 49725 24501 49759
rect 24501 49725 24535 49759
rect 24535 49725 24544 49759
rect 24492 49716 24544 49725
rect 4068 49580 4120 49632
rect 2950 49478 3002 49530
rect 3014 49478 3066 49530
rect 3078 49478 3130 49530
rect 3142 49478 3194 49530
rect 3206 49478 3258 49530
rect 12950 49478 13002 49530
rect 13014 49478 13066 49530
rect 13078 49478 13130 49530
rect 13142 49478 13194 49530
rect 13206 49478 13258 49530
rect 22950 49478 23002 49530
rect 23014 49478 23066 49530
rect 23078 49478 23130 49530
rect 23142 49478 23194 49530
rect 23206 49478 23258 49530
rect 11980 49376 12032 49428
rect 12808 49376 12860 49428
rect 1492 49240 1544 49292
rect 10692 49172 10744 49224
rect 13452 49172 13504 49224
rect 25320 49215 25372 49224
rect 25320 49181 25329 49215
rect 25329 49181 25363 49215
rect 25363 49181 25372 49215
rect 25320 49172 25372 49181
rect 10508 49036 10560 49088
rect 18788 49036 18840 49088
rect 7950 48934 8002 48986
rect 8014 48934 8066 48986
rect 8078 48934 8130 48986
rect 8142 48934 8194 48986
rect 8206 48934 8258 48986
rect 17950 48934 18002 48986
rect 18014 48934 18066 48986
rect 18078 48934 18130 48986
rect 18142 48934 18194 48986
rect 18206 48934 18258 48986
rect 24676 48628 24728 48680
rect 24768 48492 24820 48544
rect 2950 48390 3002 48442
rect 3014 48390 3066 48442
rect 3078 48390 3130 48442
rect 3142 48390 3194 48442
rect 3206 48390 3258 48442
rect 12950 48390 13002 48442
rect 13014 48390 13066 48442
rect 13078 48390 13130 48442
rect 13142 48390 13194 48442
rect 13206 48390 13258 48442
rect 22950 48390 23002 48442
rect 23014 48390 23066 48442
rect 23078 48390 23130 48442
rect 23142 48390 23194 48442
rect 23206 48390 23258 48442
rect 11704 48220 11756 48272
rect 12716 48220 12768 48272
rect 18420 48220 18472 48272
rect 18696 48084 18748 48136
rect 16028 47948 16080 48000
rect 24768 47948 24820 48000
rect 25504 47991 25556 48000
rect 25504 47957 25513 47991
rect 25513 47957 25547 47991
rect 25547 47957 25556 47991
rect 25504 47948 25556 47957
rect 7950 47846 8002 47898
rect 8014 47846 8066 47898
rect 8078 47846 8130 47898
rect 8142 47846 8194 47898
rect 8206 47846 8258 47898
rect 17950 47846 18002 47898
rect 18014 47846 18066 47898
rect 18078 47846 18130 47898
rect 18142 47846 18194 47898
rect 18206 47846 18258 47898
rect 9220 47787 9272 47796
rect 9220 47753 9229 47787
rect 9229 47753 9263 47787
rect 9263 47753 9272 47787
rect 9220 47744 9272 47753
rect 15936 47744 15988 47796
rect 17408 47744 17460 47796
rect 18512 47787 18564 47796
rect 18512 47753 18521 47787
rect 18521 47753 18555 47787
rect 18555 47753 18564 47787
rect 18512 47744 18564 47753
rect 19064 47744 19116 47796
rect 18972 47676 19024 47728
rect 11704 47608 11756 47660
rect 18420 47608 18472 47660
rect 18512 47608 18564 47660
rect 19432 47676 19484 47728
rect 25504 47608 25556 47660
rect 17408 47583 17460 47592
rect 17408 47549 17417 47583
rect 17417 47549 17451 47583
rect 17451 47549 17460 47583
rect 17408 47540 17460 47549
rect 18696 47583 18748 47592
rect 18696 47549 18705 47583
rect 18705 47549 18739 47583
rect 18739 47549 18748 47583
rect 18696 47540 18748 47549
rect 23296 47540 23348 47592
rect 11428 47404 11480 47456
rect 16580 47404 16632 47456
rect 17500 47404 17552 47456
rect 2950 47302 3002 47354
rect 3014 47302 3066 47354
rect 3078 47302 3130 47354
rect 3142 47302 3194 47354
rect 3206 47302 3258 47354
rect 12950 47302 13002 47354
rect 13014 47302 13066 47354
rect 13078 47302 13130 47354
rect 13142 47302 13194 47354
rect 13206 47302 13258 47354
rect 22950 47302 23002 47354
rect 23014 47302 23066 47354
rect 23078 47302 23130 47354
rect 23142 47302 23194 47354
rect 23206 47302 23258 47354
rect 18328 47132 18380 47184
rect 12164 47064 12216 47116
rect 16764 47064 16816 47116
rect 17592 47064 17644 47116
rect 18604 47107 18656 47116
rect 18604 47073 18613 47107
rect 18613 47073 18647 47107
rect 18647 47073 18656 47107
rect 18604 47064 18656 47073
rect 4068 46928 4120 46980
rect 9680 46928 9732 46980
rect 11428 46928 11480 46980
rect 11152 46860 11204 46912
rect 11336 46860 11388 46912
rect 18512 47039 18564 47048
rect 18512 47005 18521 47039
rect 18521 47005 18555 47039
rect 18555 47005 18564 47039
rect 18512 46996 18564 47005
rect 19984 46996 20036 47048
rect 20444 46996 20496 47048
rect 16028 46971 16080 46980
rect 16028 46937 16037 46971
rect 16037 46937 16071 46971
rect 16071 46937 16080 46971
rect 16028 46928 16080 46937
rect 18420 46928 18472 46980
rect 23756 46996 23808 47048
rect 24400 46971 24452 46980
rect 24400 46937 24409 46971
rect 24409 46937 24443 46971
rect 24443 46937 24452 46971
rect 24400 46928 24452 46937
rect 24584 46928 24636 46980
rect 12440 46860 12492 46912
rect 14188 46860 14240 46912
rect 16396 46860 16448 46912
rect 17776 46903 17828 46912
rect 17776 46869 17785 46903
rect 17785 46869 17819 46903
rect 17819 46869 17828 46903
rect 17776 46860 17828 46869
rect 21180 46903 21232 46912
rect 21180 46869 21189 46903
rect 21189 46869 21223 46903
rect 21223 46869 21232 46903
rect 21180 46860 21232 46869
rect 23848 46860 23900 46912
rect 7950 46758 8002 46810
rect 8014 46758 8066 46810
rect 8078 46758 8130 46810
rect 8142 46758 8194 46810
rect 8206 46758 8258 46810
rect 17950 46758 18002 46810
rect 18014 46758 18066 46810
rect 18078 46758 18130 46810
rect 18142 46758 18194 46810
rect 18206 46758 18258 46810
rect 7472 46656 7524 46708
rect 11152 46699 11204 46708
rect 11152 46665 11161 46699
rect 11161 46665 11195 46699
rect 11195 46665 11204 46699
rect 11152 46656 11204 46665
rect 11888 46656 11940 46708
rect 16948 46656 17000 46708
rect 17408 46656 17460 46708
rect 14188 46588 14240 46640
rect 16396 46588 16448 46640
rect 17776 46656 17828 46708
rect 18696 46656 18748 46708
rect 19616 46656 19668 46708
rect 20352 46656 20404 46708
rect 20720 46656 20772 46708
rect 22468 46699 22520 46708
rect 22468 46665 22477 46699
rect 22477 46665 22511 46699
rect 22511 46665 22520 46699
rect 22468 46656 22520 46665
rect 9496 46520 9548 46572
rect 10600 46520 10652 46572
rect 16764 46520 16816 46572
rect 10876 46452 10928 46504
rect 12164 46452 12216 46504
rect 14280 46452 14332 46504
rect 14556 46495 14608 46504
rect 14556 46461 14565 46495
rect 14565 46461 14599 46495
rect 14599 46461 14608 46495
rect 14556 46452 14608 46461
rect 16488 46452 16540 46504
rect 18880 46452 18932 46504
rect 20352 46495 20404 46504
rect 20352 46461 20361 46495
rect 20361 46461 20395 46495
rect 20395 46461 20404 46495
rect 20352 46452 20404 46461
rect 22468 46452 22520 46504
rect 24584 46452 24636 46504
rect 24768 46495 24820 46504
rect 24768 46461 24777 46495
rect 24777 46461 24811 46495
rect 24811 46461 24820 46495
rect 24768 46452 24820 46461
rect 14096 46359 14148 46368
rect 14096 46325 14105 46359
rect 14105 46325 14139 46359
rect 14139 46325 14148 46359
rect 14096 46316 14148 46325
rect 18788 46316 18840 46368
rect 19800 46316 19852 46368
rect 22744 46316 22796 46368
rect 24492 46316 24544 46368
rect 2950 46214 3002 46266
rect 3014 46214 3066 46266
rect 3078 46214 3130 46266
rect 3142 46214 3194 46266
rect 3206 46214 3258 46266
rect 12950 46214 13002 46266
rect 13014 46214 13066 46266
rect 13078 46214 13130 46266
rect 13142 46214 13194 46266
rect 13206 46214 13258 46266
rect 22950 46214 23002 46266
rect 23014 46214 23066 46266
rect 23078 46214 23130 46266
rect 23142 46214 23194 46266
rect 23206 46214 23258 46266
rect 5632 46112 5684 46164
rect 9312 46112 9364 46164
rect 10692 46155 10744 46164
rect 10692 46121 10701 46155
rect 10701 46121 10735 46155
rect 10735 46121 10744 46155
rect 10692 46112 10744 46121
rect 14188 46155 14240 46164
rect 14188 46121 14197 46155
rect 14197 46121 14231 46155
rect 14231 46121 14240 46155
rect 14188 46112 14240 46121
rect 16488 46155 16540 46164
rect 16488 46121 16497 46155
rect 16497 46121 16531 46155
rect 16531 46121 16540 46155
rect 16488 46112 16540 46121
rect 22192 46112 22244 46164
rect 7656 46044 7708 46096
rect 11336 46019 11388 46028
rect 11336 45985 11345 46019
rect 11345 45985 11379 46019
rect 11379 45985 11388 46019
rect 11336 45976 11388 45985
rect 12164 45976 12216 46028
rect 16488 45976 16540 46028
rect 16764 45976 16816 46028
rect 18420 45976 18472 46028
rect 21180 45976 21232 46028
rect 21824 45976 21876 46028
rect 7012 45908 7064 45960
rect 11520 45908 11572 45960
rect 8852 45772 8904 45824
rect 11152 45815 11204 45824
rect 11152 45781 11161 45815
rect 11161 45781 11195 45815
rect 11195 45781 11204 45815
rect 11152 45772 11204 45781
rect 12440 45840 12492 45892
rect 14188 45840 14240 45892
rect 13176 45772 13228 45824
rect 13728 45772 13780 45824
rect 19524 45951 19576 45960
rect 19524 45917 19533 45951
rect 19533 45917 19567 45951
rect 19567 45917 19576 45951
rect 19524 45908 19576 45917
rect 22192 45908 22244 45960
rect 23940 45908 23992 45960
rect 24032 45908 24084 45960
rect 18788 45840 18840 45892
rect 16764 45772 16816 45824
rect 18696 45772 18748 45824
rect 19892 45772 19944 45824
rect 21732 45772 21784 45824
rect 22836 45772 22888 45824
rect 23848 45815 23900 45824
rect 23848 45781 23857 45815
rect 23857 45781 23891 45815
rect 23891 45781 23900 45815
rect 23848 45772 23900 45781
rect 24216 45815 24268 45824
rect 24216 45781 24225 45815
rect 24225 45781 24259 45815
rect 24259 45781 24268 45815
rect 24216 45772 24268 45781
rect 25228 45815 25280 45824
rect 25228 45781 25237 45815
rect 25237 45781 25271 45815
rect 25271 45781 25280 45815
rect 25228 45772 25280 45781
rect 7950 45670 8002 45722
rect 8014 45670 8066 45722
rect 8078 45670 8130 45722
rect 8142 45670 8194 45722
rect 8206 45670 8258 45722
rect 17950 45670 18002 45722
rect 18014 45670 18066 45722
rect 18078 45670 18130 45722
rect 18142 45670 18194 45722
rect 18206 45670 18258 45722
rect 4068 45568 4120 45620
rect 8944 45568 8996 45620
rect 10232 45568 10284 45620
rect 19984 45611 20036 45620
rect 19984 45577 19993 45611
rect 19993 45577 20027 45611
rect 20027 45577 20036 45611
rect 19984 45568 20036 45577
rect 8760 45543 8812 45552
rect 8760 45509 8769 45543
rect 8769 45509 8803 45543
rect 8803 45509 8812 45543
rect 8760 45500 8812 45509
rect 9312 45500 9364 45552
rect 11428 45500 11480 45552
rect 13176 45500 13228 45552
rect 13636 45500 13688 45552
rect 6828 45432 6880 45484
rect 11796 45475 11848 45484
rect 11796 45441 11805 45475
rect 11805 45441 11839 45475
rect 11839 45441 11848 45475
rect 11796 45432 11848 45441
rect 13544 45475 13596 45484
rect 13544 45441 13553 45475
rect 13553 45441 13587 45475
rect 13587 45441 13596 45475
rect 13544 45432 13596 45441
rect 14556 45500 14608 45552
rect 16488 45500 16540 45552
rect 21732 45568 21784 45620
rect 20904 45543 20956 45552
rect 20904 45509 20913 45543
rect 20913 45509 20947 45543
rect 20947 45509 20956 45543
rect 20904 45500 20956 45509
rect 16948 45432 17000 45484
rect 22284 45500 22336 45552
rect 23848 45500 23900 45552
rect 11060 45296 11112 45348
rect 13452 45296 13504 45348
rect 10876 45271 10928 45280
rect 10876 45237 10885 45271
rect 10885 45237 10919 45271
rect 10919 45237 10928 45271
rect 10876 45228 10928 45237
rect 12072 45228 12124 45280
rect 13820 45364 13872 45416
rect 14096 45364 14148 45416
rect 14372 45407 14424 45416
rect 14372 45373 14381 45407
rect 14381 45373 14415 45407
rect 14415 45373 14424 45407
rect 14372 45364 14424 45373
rect 15292 45228 15344 45280
rect 16304 45228 16356 45280
rect 16488 45271 16540 45280
rect 16488 45237 16497 45271
rect 16497 45237 16531 45271
rect 16531 45237 16540 45271
rect 16488 45228 16540 45237
rect 18512 45407 18564 45416
rect 18512 45373 18521 45407
rect 18521 45373 18555 45407
rect 18555 45373 18564 45407
rect 18512 45364 18564 45373
rect 19248 45364 19300 45416
rect 21272 45364 21324 45416
rect 25228 45432 25280 45484
rect 23848 45364 23900 45416
rect 24492 45407 24544 45416
rect 24492 45373 24501 45407
rect 24501 45373 24535 45407
rect 24535 45373 24544 45407
rect 24492 45364 24544 45373
rect 24768 45407 24820 45416
rect 24768 45373 24777 45407
rect 24777 45373 24811 45407
rect 24811 45373 24820 45407
rect 24768 45364 24820 45373
rect 19616 45228 19668 45280
rect 20260 45228 20312 45280
rect 21732 45228 21784 45280
rect 2950 45126 3002 45178
rect 3014 45126 3066 45178
rect 3078 45126 3130 45178
rect 3142 45126 3194 45178
rect 3206 45126 3258 45178
rect 12950 45126 13002 45178
rect 13014 45126 13066 45178
rect 13078 45126 13130 45178
rect 13142 45126 13194 45178
rect 13206 45126 13258 45178
rect 22950 45126 23002 45178
rect 23014 45126 23066 45178
rect 23078 45126 23130 45178
rect 23142 45126 23194 45178
rect 23206 45126 23258 45178
rect 6460 45024 6512 45076
rect 9404 45024 9456 45076
rect 9864 45024 9916 45076
rect 18880 45067 18932 45076
rect 18880 45033 18889 45067
rect 18889 45033 18923 45067
rect 18923 45033 18932 45067
rect 18880 45024 18932 45033
rect 20352 45024 20404 45076
rect 21732 45024 21784 45076
rect 23848 45024 23900 45076
rect 10324 44956 10376 45008
rect 7288 44888 7340 44940
rect 11428 44888 11480 44940
rect 14096 44888 14148 44940
rect 14372 44888 14424 44940
rect 16856 44888 16908 44940
rect 21548 44888 21600 44940
rect 7656 44820 7708 44872
rect 13820 44820 13872 44872
rect 16488 44820 16540 44872
rect 6644 44684 6696 44736
rect 7104 44684 7156 44736
rect 14188 44752 14240 44804
rect 15384 44795 15436 44804
rect 15384 44761 15393 44795
rect 15393 44761 15427 44795
rect 15427 44761 15436 44795
rect 15384 44752 15436 44761
rect 16764 44752 16816 44804
rect 9772 44727 9824 44736
rect 9772 44693 9781 44727
rect 9781 44693 9815 44727
rect 9815 44693 9824 44727
rect 9772 44684 9824 44693
rect 11612 44727 11664 44736
rect 11612 44693 11621 44727
rect 11621 44693 11655 44727
rect 11655 44693 11664 44727
rect 11612 44684 11664 44693
rect 12808 44684 12860 44736
rect 17316 44752 17368 44804
rect 18880 44820 18932 44872
rect 18788 44684 18840 44736
rect 19340 44727 19392 44736
rect 19340 44693 19349 44727
rect 19349 44693 19383 44727
rect 19383 44693 19392 44727
rect 19340 44684 19392 44693
rect 19616 44684 19668 44736
rect 22284 44863 22336 44872
rect 22284 44829 22293 44863
rect 22293 44829 22327 44863
rect 22327 44829 22336 44863
rect 22284 44820 22336 44829
rect 24124 44820 24176 44872
rect 21732 44752 21784 44804
rect 23848 44752 23900 44804
rect 22284 44684 22336 44736
rect 23388 44684 23440 44736
rect 24032 44727 24084 44736
rect 24032 44693 24041 44727
rect 24041 44693 24075 44727
rect 24075 44693 24084 44727
rect 24032 44684 24084 44693
rect 7950 44582 8002 44634
rect 8014 44582 8066 44634
rect 8078 44582 8130 44634
rect 8142 44582 8194 44634
rect 8206 44582 8258 44634
rect 17950 44582 18002 44634
rect 18014 44582 18066 44634
rect 18078 44582 18130 44634
rect 18142 44582 18194 44634
rect 18206 44582 18258 44634
rect 5816 44523 5868 44532
rect 5816 44489 5825 44523
rect 5825 44489 5859 44523
rect 5859 44489 5868 44523
rect 5816 44480 5868 44489
rect 6736 44523 6788 44532
rect 6736 44489 6745 44523
rect 6745 44489 6779 44523
rect 6779 44489 6788 44523
rect 6736 44480 6788 44489
rect 7196 44480 7248 44532
rect 10968 44480 11020 44532
rect 11152 44480 11204 44532
rect 12440 44480 12492 44532
rect 7564 44455 7616 44464
rect 7564 44421 7573 44455
rect 7573 44421 7607 44455
rect 7607 44421 7616 44455
rect 7564 44412 7616 44421
rect 12164 44412 12216 44464
rect 13728 44480 13780 44532
rect 6552 44344 6604 44396
rect 6644 44387 6696 44396
rect 6644 44353 6653 44387
rect 6653 44353 6687 44387
rect 6687 44353 6696 44387
rect 6644 44344 6696 44353
rect 7748 44344 7800 44396
rect 9220 44344 9272 44396
rect 10232 44387 10284 44396
rect 10232 44353 10241 44387
rect 10241 44353 10275 44387
rect 10275 44353 10284 44387
rect 10232 44344 10284 44353
rect 16488 44480 16540 44532
rect 18512 44480 18564 44532
rect 7380 44208 7432 44260
rect 7748 44140 7800 44192
rect 9220 44140 9272 44192
rect 11612 44251 11664 44260
rect 11612 44217 11621 44251
rect 11621 44217 11655 44251
rect 11655 44217 11664 44251
rect 11612 44208 11664 44217
rect 10416 44140 10468 44192
rect 12072 44208 12124 44260
rect 14096 44276 14148 44328
rect 18788 44412 18840 44464
rect 23848 44412 23900 44464
rect 16856 44387 16908 44396
rect 16856 44353 16865 44387
rect 16865 44353 16899 44387
rect 16899 44353 16908 44387
rect 16856 44344 16908 44353
rect 19892 44344 19944 44396
rect 20076 44344 20128 44396
rect 24308 44344 24360 44396
rect 18512 44276 18564 44328
rect 18696 44276 18748 44328
rect 22284 44319 22336 44328
rect 22284 44285 22293 44319
rect 22293 44285 22327 44319
rect 22327 44285 22336 44319
rect 22284 44276 22336 44285
rect 22652 44276 22704 44328
rect 24584 44276 24636 44328
rect 14372 44140 14424 44192
rect 14464 44140 14516 44192
rect 14832 44183 14884 44192
rect 14832 44149 14841 44183
rect 14841 44149 14875 44183
rect 14875 44149 14884 44183
rect 14832 44140 14884 44149
rect 16212 44140 16264 44192
rect 16764 44140 16816 44192
rect 18880 44140 18932 44192
rect 19524 44140 19576 44192
rect 20812 44140 20864 44192
rect 21916 44183 21968 44192
rect 21916 44149 21925 44183
rect 21925 44149 21959 44183
rect 21959 44149 21968 44183
rect 21916 44140 21968 44149
rect 24032 44183 24084 44192
rect 24032 44149 24041 44183
rect 24041 44149 24075 44183
rect 24075 44149 24084 44183
rect 24032 44140 24084 44149
rect 2950 44038 3002 44090
rect 3014 44038 3066 44090
rect 3078 44038 3130 44090
rect 3142 44038 3194 44090
rect 3206 44038 3258 44090
rect 12950 44038 13002 44090
rect 13014 44038 13066 44090
rect 13078 44038 13130 44090
rect 13142 44038 13194 44090
rect 13206 44038 13258 44090
rect 22950 44038 23002 44090
rect 23014 44038 23066 44090
rect 23078 44038 23130 44090
rect 23142 44038 23194 44090
rect 23206 44038 23258 44090
rect 4988 43936 5040 43988
rect 8392 43979 8444 43988
rect 8392 43945 8401 43979
rect 8401 43945 8435 43979
rect 8435 43945 8444 43979
rect 8392 43936 8444 43945
rect 9956 43936 10008 43988
rect 10508 43936 10560 43988
rect 10876 43800 10928 43852
rect 9036 43732 9088 43784
rect 11428 43936 11480 43988
rect 21548 43979 21600 43988
rect 21548 43945 21557 43979
rect 21557 43945 21591 43979
rect 21591 43945 21600 43979
rect 21548 43936 21600 43945
rect 15384 43868 15436 43920
rect 17684 43868 17736 43920
rect 21640 43868 21692 43920
rect 17500 43843 17552 43852
rect 17500 43809 17509 43843
rect 17509 43809 17543 43843
rect 17543 43809 17552 43843
rect 17500 43800 17552 43809
rect 17592 43843 17644 43852
rect 17592 43809 17601 43843
rect 17601 43809 17635 43843
rect 17635 43809 17644 43843
rect 17592 43800 17644 43809
rect 25136 43868 25188 43920
rect 13820 43732 13872 43784
rect 16304 43732 16356 43784
rect 17408 43775 17460 43784
rect 17408 43741 17417 43775
rect 17417 43741 17451 43775
rect 17451 43741 17460 43775
rect 22560 43843 22612 43852
rect 22560 43809 22569 43843
rect 22569 43809 22603 43843
rect 22603 43809 22612 43843
rect 22560 43800 22612 43809
rect 24492 43800 24544 43852
rect 17408 43732 17460 43741
rect 20628 43732 20680 43784
rect 21180 43732 21232 43784
rect 21272 43732 21324 43784
rect 24216 43732 24268 43784
rect 24768 43732 24820 43784
rect 15844 43664 15896 43716
rect 21916 43664 21968 43716
rect 23848 43664 23900 43716
rect 15016 43596 15068 43648
rect 16028 43639 16080 43648
rect 16028 43605 16037 43639
rect 16037 43605 16071 43639
rect 16071 43605 16080 43639
rect 16028 43596 16080 43605
rect 17224 43596 17276 43648
rect 18788 43639 18840 43648
rect 18788 43605 18797 43639
rect 18797 43605 18831 43639
rect 18831 43605 18840 43639
rect 18788 43596 18840 43605
rect 19248 43596 19300 43648
rect 19340 43596 19392 43648
rect 20536 43639 20588 43648
rect 20536 43605 20545 43639
rect 20545 43605 20579 43639
rect 20579 43605 20588 43639
rect 20536 43596 20588 43605
rect 20904 43596 20956 43648
rect 22192 43596 22244 43648
rect 23940 43639 23992 43648
rect 23940 43605 23949 43639
rect 23949 43605 23983 43639
rect 23983 43605 23992 43639
rect 23940 43596 23992 43605
rect 24216 43596 24268 43648
rect 25228 43596 25280 43648
rect 7950 43494 8002 43546
rect 8014 43494 8066 43546
rect 8078 43494 8130 43546
rect 8142 43494 8194 43546
rect 8206 43494 8258 43546
rect 17950 43494 18002 43546
rect 18014 43494 18066 43546
rect 18078 43494 18130 43546
rect 18142 43494 18194 43546
rect 18206 43494 18258 43546
rect 7840 43392 7892 43444
rect 10416 43392 10468 43444
rect 13728 43392 13780 43444
rect 4620 43324 4672 43376
rect 9588 43324 9640 43376
rect 12808 43367 12860 43376
rect 12808 43333 12817 43367
rect 12817 43333 12851 43367
rect 12851 43333 12860 43367
rect 12808 43324 12860 43333
rect 14096 43324 14148 43376
rect 14648 43392 14700 43444
rect 17684 43392 17736 43444
rect 22376 43392 22428 43444
rect 24584 43392 24636 43444
rect 1308 43256 1360 43308
rect 7656 43256 7708 43308
rect 9312 43256 9364 43308
rect 3516 43120 3568 43172
rect 8944 43188 8996 43240
rect 10232 43256 10284 43308
rect 15936 43256 15988 43308
rect 16856 43324 16908 43376
rect 19248 43324 19300 43376
rect 22284 43324 22336 43376
rect 14648 43188 14700 43240
rect 18236 43299 18288 43308
rect 18236 43265 18245 43299
rect 18245 43265 18279 43299
rect 18279 43265 18288 43299
rect 18236 43256 18288 43265
rect 20168 43256 20220 43308
rect 20536 43299 20588 43308
rect 20536 43265 20545 43299
rect 20545 43265 20579 43299
rect 20579 43265 20588 43299
rect 20536 43256 20588 43265
rect 21916 43256 21968 43308
rect 24124 43324 24176 43376
rect 25136 43256 25188 43308
rect 25596 43256 25648 43308
rect 14096 43120 14148 43172
rect 14740 43120 14792 43172
rect 16120 43120 16172 43172
rect 7472 43095 7524 43104
rect 7472 43061 7481 43095
rect 7481 43061 7515 43095
rect 7515 43061 7524 43095
rect 7472 43052 7524 43061
rect 14924 43052 14976 43104
rect 15936 43052 15988 43104
rect 16396 43095 16448 43104
rect 16396 43061 16405 43095
rect 16405 43061 16439 43095
rect 16439 43061 16448 43095
rect 16396 43052 16448 43061
rect 16948 43095 17000 43104
rect 16948 43061 16957 43095
rect 16957 43061 16991 43095
rect 16991 43061 17000 43095
rect 16948 43052 17000 43061
rect 19524 43188 19576 43240
rect 22560 43231 22612 43240
rect 22560 43197 22569 43231
rect 22569 43197 22603 43231
rect 22603 43197 22612 43231
rect 22560 43188 22612 43197
rect 23480 43188 23532 43240
rect 23848 43231 23900 43240
rect 23848 43197 23857 43231
rect 23857 43197 23891 43231
rect 23891 43197 23900 43231
rect 23848 43188 23900 43197
rect 19524 43052 19576 43104
rect 20076 43052 20128 43104
rect 25412 43120 25464 43172
rect 25320 43095 25372 43104
rect 25320 43061 25329 43095
rect 25329 43061 25363 43095
rect 25363 43061 25372 43095
rect 25320 43052 25372 43061
rect 2950 42950 3002 43002
rect 3014 42950 3066 43002
rect 3078 42950 3130 43002
rect 3142 42950 3194 43002
rect 3206 42950 3258 43002
rect 12950 42950 13002 43002
rect 13014 42950 13066 43002
rect 13078 42950 13130 43002
rect 13142 42950 13194 43002
rect 13206 42950 13258 43002
rect 22950 42950 23002 43002
rect 23014 42950 23066 43002
rect 23078 42950 23130 43002
rect 23142 42950 23194 43002
rect 23206 42950 23258 43002
rect 8944 42891 8996 42900
rect 8944 42857 8953 42891
rect 8953 42857 8987 42891
rect 8987 42857 8996 42891
rect 8944 42848 8996 42857
rect 9588 42848 9640 42900
rect 9680 42848 9732 42900
rect 11244 42848 11296 42900
rect 16396 42848 16448 42900
rect 4528 42712 4580 42764
rect 8484 42712 8536 42764
rect 10876 42755 10928 42764
rect 10876 42721 10885 42755
rect 10885 42721 10919 42755
rect 10919 42721 10928 42755
rect 10876 42712 10928 42721
rect 12164 42712 12216 42764
rect 8300 42644 8352 42696
rect 9772 42687 9824 42696
rect 9772 42653 9781 42687
rect 9781 42653 9815 42687
rect 9815 42653 9824 42687
rect 9772 42644 9824 42653
rect 14004 42780 14056 42832
rect 16580 42780 16632 42832
rect 12348 42712 12400 42764
rect 13820 42712 13872 42764
rect 14648 42712 14700 42764
rect 16856 42712 16908 42764
rect 16120 42644 16172 42696
rect 16488 42644 16540 42696
rect 19248 42848 19300 42900
rect 23940 42848 23992 42900
rect 24124 42848 24176 42900
rect 24952 42848 25004 42900
rect 22376 42780 22428 42832
rect 17592 42712 17644 42764
rect 22008 42712 22060 42764
rect 24032 42780 24084 42832
rect 23020 42712 23072 42764
rect 18236 42644 18288 42696
rect 18788 42644 18840 42696
rect 19616 42687 19668 42696
rect 19616 42653 19625 42687
rect 19625 42653 19659 42687
rect 19659 42653 19668 42687
rect 19616 42644 19668 42653
rect 23204 42687 23256 42696
rect 23204 42653 23213 42687
rect 23213 42653 23247 42687
rect 23247 42653 23256 42687
rect 23204 42644 23256 42653
rect 25136 42644 25188 42696
rect 25320 42644 25372 42696
rect 15016 42619 15068 42628
rect 15016 42585 15025 42619
rect 15025 42585 15059 42619
rect 15059 42585 15068 42619
rect 15016 42576 15068 42585
rect 17132 42576 17184 42628
rect 20168 42576 20220 42628
rect 20904 42576 20956 42628
rect 22744 42576 22796 42628
rect 6736 42508 6788 42560
rect 7840 42508 7892 42560
rect 20628 42508 20680 42560
rect 21548 42508 21600 42560
rect 22008 42508 22060 42560
rect 23756 42508 23808 42560
rect 7950 42406 8002 42458
rect 8014 42406 8066 42458
rect 8078 42406 8130 42458
rect 8142 42406 8194 42458
rect 8206 42406 8258 42458
rect 17950 42406 18002 42458
rect 18014 42406 18066 42458
rect 18078 42406 18130 42458
rect 18142 42406 18194 42458
rect 18206 42406 18258 42458
rect 4344 42304 4396 42356
rect 9496 42304 9548 42356
rect 11060 42347 11112 42356
rect 11060 42313 11069 42347
rect 11069 42313 11103 42347
rect 11103 42313 11112 42347
rect 11060 42304 11112 42313
rect 11704 42347 11756 42356
rect 11704 42313 11713 42347
rect 11713 42313 11747 42347
rect 11747 42313 11756 42347
rect 11704 42304 11756 42313
rect 13544 42304 13596 42356
rect 15292 42347 15344 42356
rect 15292 42313 15301 42347
rect 15301 42313 15335 42347
rect 15335 42313 15344 42347
rect 15292 42304 15344 42313
rect 16948 42304 17000 42356
rect 7840 42279 7892 42288
rect 7840 42245 7849 42279
rect 7849 42245 7883 42279
rect 7883 42245 7892 42279
rect 7840 42236 7892 42245
rect 8484 42236 8536 42288
rect 12164 42236 12216 42288
rect 13452 42236 13504 42288
rect 14372 42236 14424 42288
rect 18604 42304 18656 42356
rect 22008 42304 22060 42356
rect 22192 42304 22244 42356
rect 22652 42304 22704 42356
rect 24492 42304 24544 42356
rect 5908 42168 5960 42220
rect 6828 42168 6880 42220
rect 10140 42211 10192 42220
rect 10140 42177 10149 42211
rect 10149 42177 10183 42211
rect 10183 42177 10192 42211
rect 10140 42168 10192 42177
rect 10508 42168 10560 42220
rect 17500 42211 17552 42220
rect 17500 42177 17509 42211
rect 17509 42177 17543 42211
rect 17543 42177 17552 42211
rect 17500 42168 17552 42177
rect 9772 42100 9824 42152
rect 10324 42143 10376 42152
rect 10324 42109 10333 42143
rect 10333 42109 10367 42143
rect 10367 42109 10376 42143
rect 10324 42100 10376 42109
rect 10232 42032 10284 42084
rect 12348 42143 12400 42152
rect 12348 42109 12357 42143
rect 12357 42109 12391 42143
rect 12391 42109 12400 42143
rect 12348 42100 12400 42109
rect 14832 42100 14884 42152
rect 19340 42236 19392 42288
rect 20904 42236 20956 42288
rect 23756 42279 23808 42288
rect 23756 42245 23765 42279
rect 23765 42245 23799 42279
rect 23799 42245 23808 42279
rect 23756 42236 23808 42245
rect 24216 42236 24268 42288
rect 18788 42211 18840 42220
rect 18788 42177 18797 42211
rect 18797 42177 18831 42211
rect 18831 42177 18840 42211
rect 18788 42168 18840 42177
rect 10784 42007 10836 42016
rect 10784 41973 10793 42007
rect 10793 41973 10827 42007
rect 10827 41973 10836 42007
rect 10784 41964 10836 41973
rect 15108 42032 15160 42084
rect 19432 42100 19484 42152
rect 17776 41964 17828 42016
rect 21180 42032 21232 42084
rect 22468 42168 22520 42220
rect 22652 42168 22704 42220
rect 22100 42032 22152 42084
rect 20904 42007 20956 42016
rect 20904 41973 20913 42007
rect 20913 41973 20947 42007
rect 20947 41973 20956 42007
rect 20904 41964 20956 41973
rect 22468 41964 22520 42016
rect 23296 41964 23348 42016
rect 23480 42143 23532 42152
rect 23480 42109 23489 42143
rect 23489 42109 23523 42143
rect 23523 42109 23532 42143
rect 23480 42100 23532 42109
rect 24216 41964 24268 42016
rect 2950 41862 3002 41914
rect 3014 41862 3066 41914
rect 3078 41862 3130 41914
rect 3142 41862 3194 41914
rect 3206 41862 3258 41914
rect 12950 41862 13002 41914
rect 13014 41862 13066 41914
rect 13078 41862 13130 41914
rect 13142 41862 13194 41914
rect 13206 41862 13258 41914
rect 22950 41862 23002 41914
rect 23014 41862 23066 41914
rect 23078 41862 23130 41914
rect 23142 41862 23194 41914
rect 23206 41862 23258 41914
rect 4160 41803 4212 41812
rect 4160 41769 4169 41803
rect 4169 41769 4203 41803
rect 4203 41769 4212 41803
rect 4160 41760 4212 41769
rect 4804 41760 4856 41812
rect 6460 41760 6512 41812
rect 6828 41760 6880 41812
rect 8484 41760 8536 41812
rect 8944 41760 8996 41812
rect 11520 41803 11572 41812
rect 11520 41769 11529 41803
rect 11529 41769 11563 41803
rect 11563 41769 11572 41803
rect 11520 41760 11572 41769
rect 8300 41692 8352 41744
rect 10324 41692 10376 41744
rect 7288 41624 7340 41676
rect 8944 41624 8996 41676
rect 8392 41556 8444 41608
rect 8668 41556 8720 41608
rect 9496 41556 9548 41608
rect 10784 41624 10836 41676
rect 10876 41667 10928 41676
rect 10876 41633 10885 41667
rect 10885 41633 10919 41667
rect 10919 41633 10928 41667
rect 10876 41624 10928 41633
rect 12808 41692 12860 41744
rect 12072 41667 12124 41676
rect 12072 41633 12081 41667
rect 12081 41633 12115 41667
rect 12115 41633 12124 41667
rect 12072 41624 12124 41633
rect 4068 41531 4120 41540
rect 4068 41497 4077 41531
rect 4077 41497 4111 41531
rect 4111 41497 4120 41531
rect 4068 41488 4120 41497
rect 5264 41531 5316 41540
rect 5264 41497 5273 41531
rect 5273 41497 5307 41531
rect 5307 41497 5316 41531
rect 5264 41488 5316 41497
rect 11428 41556 11480 41608
rect 12532 41556 12584 41608
rect 16304 41624 16356 41676
rect 3976 41420 4028 41472
rect 9128 41463 9180 41472
rect 9128 41429 9137 41463
rect 9137 41429 9171 41463
rect 9171 41429 9180 41463
rect 9128 41420 9180 41429
rect 11152 41488 11204 41540
rect 14464 41488 14516 41540
rect 10600 41420 10652 41472
rect 10692 41463 10744 41472
rect 10692 41429 10701 41463
rect 10701 41429 10735 41463
rect 10735 41429 10744 41463
rect 10692 41420 10744 41429
rect 11796 41420 11848 41472
rect 13360 41463 13412 41472
rect 13360 41429 13369 41463
rect 13369 41429 13403 41463
rect 13403 41429 13412 41463
rect 13360 41420 13412 41429
rect 14188 41420 14240 41472
rect 16672 41556 16724 41608
rect 16120 41488 16172 41540
rect 22468 41760 22520 41812
rect 17500 41692 17552 41744
rect 20352 41692 20404 41744
rect 18328 41624 18380 41676
rect 15292 41420 15344 41472
rect 16396 41463 16448 41472
rect 16396 41429 16405 41463
rect 16405 41429 16439 41463
rect 16439 41429 16448 41463
rect 16396 41420 16448 41429
rect 17592 41556 17644 41608
rect 18512 41556 18564 41608
rect 20168 41667 20220 41676
rect 20168 41633 20177 41667
rect 20177 41633 20211 41667
rect 20211 41633 20220 41667
rect 20168 41624 20220 41633
rect 20628 41624 20680 41676
rect 20260 41556 20312 41608
rect 22928 41692 22980 41744
rect 23204 41692 23256 41744
rect 23480 41692 23532 41744
rect 23848 41760 23900 41812
rect 25044 41692 25096 41744
rect 22376 41624 22428 41676
rect 22744 41624 22796 41676
rect 23664 41624 23716 41676
rect 18328 41488 18380 41540
rect 18420 41420 18472 41472
rect 20628 41488 20680 41540
rect 20720 41488 20772 41540
rect 18972 41420 19024 41472
rect 19156 41420 19208 41472
rect 19616 41463 19668 41472
rect 19616 41429 19625 41463
rect 19625 41429 19659 41463
rect 19659 41429 19668 41463
rect 19616 41420 19668 41429
rect 19984 41463 20036 41472
rect 19984 41429 19993 41463
rect 19993 41429 20027 41463
rect 20027 41429 20036 41463
rect 19984 41420 20036 41429
rect 21732 41463 21784 41472
rect 21732 41429 21741 41463
rect 21741 41429 21775 41463
rect 21775 41429 21784 41463
rect 21732 41420 21784 41429
rect 22744 41420 22796 41472
rect 24124 41556 24176 41608
rect 24584 41599 24636 41608
rect 24584 41565 24593 41599
rect 24593 41565 24627 41599
rect 24627 41565 24636 41599
rect 24584 41556 24636 41565
rect 7950 41318 8002 41370
rect 8014 41318 8066 41370
rect 8078 41318 8130 41370
rect 8142 41318 8194 41370
rect 8206 41318 8258 41370
rect 17950 41318 18002 41370
rect 18014 41318 18066 41370
rect 18078 41318 18130 41370
rect 18142 41318 18194 41370
rect 18206 41318 18258 41370
rect 3608 41259 3660 41268
rect 3608 41225 3617 41259
rect 3617 41225 3651 41259
rect 3651 41225 3660 41259
rect 3608 41216 3660 41225
rect 4712 41259 4764 41268
rect 4712 41225 4721 41259
rect 4721 41225 4755 41259
rect 4755 41225 4764 41259
rect 4712 41216 4764 41225
rect 1308 41080 1360 41132
rect 4528 41080 4580 41132
rect 5080 41080 5132 41132
rect 10876 41216 10928 41268
rect 11060 41259 11112 41268
rect 11060 41225 11069 41259
rect 11069 41225 11103 41259
rect 11103 41225 11112 41259
rect 11060 41216 11112 41225
rect 17132 41216 17184 41268
rect 19800 41259 19852 41268
rect 19800 41225 19809 41259
rect 19809 41225 19843 41259
rect 19843 41225 19852 41259
rect 19800 41216 19852 41225
rect 20904 41216 20956 41268
rect 16120 41191 16172 41200
rect 16120 41157 16129 41191
rect 16129 41157 16163 41191
rect 16163 41157 16172 41191
rect 16120 41148 16172 41157
rect 18972 41148 19024 41200
rect 19248 41148 19300 41200
rect 21824 41216 21876 41268
rect 10876 41080 10928 41132
rect 11060 41080 11112 41132
rect 11980 41080 12032 41132
rect 12256 41080 12308 41132
rect 15200 41080 15252 41132
rect 16488 41080 16540 41132
rect 16856 41080 16908 41132
rect 20904 41080 20956 41132
rect 22100 41080 22152 41132
rect 23204 41148 23256 41200
rect 24584 41259 24636 41268
rect 24584 41225 24593 41259
rect 24593 41225 24627 41259
rect 24627 41225 24636 41259
rect 24584 41216 24636 41225
rect 25228 41148 25280 41200
rect 24216 41080 24268 41132
rect 24400 41080 24452 41132
rect 25320 41123 25372 41132
rect 25320 41089 25329 41123
rect 25329 41089 25363 41123
rect 25363 41089 25372 41123
rect 25320 41080 25372 41089
rect 8484 41012 8536 41064
rect 13360 41012 13412 41064
rect 16028 41012 16080 41064
rect 18604 41012 18656 41064
rect 19892 41055 19944 41064
rect 19892 41021 19901 41055
rect 19901 41021 19935 41055
rect 19935 41021 19944 41055
rect 19892 41012 19944 41021
rect 20996 41012 21048 41064
rect 16488 40944 16540 40996
rect 3608 40876 3660 40928
rect 5080 40919 5132 40928
rect 5080 40885 5089 40919
rect 5089 40885 5123 40919
rect 5123 40885 5132 40919
rect 5080 40876 5132 40885
rect 8576 40919 8628 40928
rect 8576 40885 8585 40919
rect 8585 40885 8619 40919
rect 8619 40885 8628 40919
rect 8576 40876 8628 40885
rect 10876 40876 10928 40928
rect 12348 40876 12400 40928
rect 13820 40876 13872 40928
rect 16580 40876 16632 40928
rect 17868 40876 17920 40928
rect 18788 40876 18840 40928
rect 18972 40919 19024 40928
rect 18972 40885 18981 40919
rect 18981 40885 19015 40919
rect 19015 40885 19024 40919
rect 18972 40876 19024 40885
rect 19340 40919 19392 40928
rect 19340 40885 19349 40919
rect 19349 40885 19383 40919
rect 19383 40885 19392 40919
rect 19340 40876 19392 40885
rect 20444 40876 20496 40928
rect 21456 40944 21508 40996
rect 24952 41012 25004 41064
rect 21732 40876 21784 40928
rect 21916 40876 21968 40928
rect 24124 40876 24176 40928
rect 25504 40876 25556 40928
rect 2950 40774 3002 40826
rect 3014 40774 3066 40826
rect 3078 40774 3130 40826
rect 3142 40774 3194 40826
rect 3206 40774 3258 40826
rect 12950 40774 13002 40826
rect 13014 40774 13066 40826
rect 13078 40774 13130 40826
rect 13142 40774 13194 40826
rect 13206 40774 13258 40826
rect 22950 40774 23002 40826
rect 23014 40774 23066 40826
rect 23078 40774 23130 40826
rect 23142 40774 23194 40826
rect 23206 40774 23258 40826
rect 7288 40672 7340 40724
rect 8668 40715 8720 40724
rect 8668 40681 8677 40715
rect 8677 40681 8711 40715
rect 8711 40681 8720 40715
rect 8668 40672 8720 40681
rect 10232 40672 10284 40724
rect 11060 40672 11112 40724
rect 11796 40672 11848 40724
rect 15844 40672 15896 40724
rect 18604 40715 18656 40724
rect 18604 40681 18613 40715
rect 18613 40681 18647 40715
rect 18647 40681 18656 40715
rect 18604 40672 18656 40681
rect 22192 40672 22244 40724
rect 7840 40604 7892 40656
rect 10876 40647 10928 40656
rect 10876 40613 10885 40647
rect 10885 40613 10919 40647
rect 10919 40613 10928 40647
rect 10876 40604 10928 40613
rect 12624 40604 12676 40656
rect 7380 40536 7432 40588
rect 8760 40536 8812 40588
rect 6460 40511 6512 40520
rect 6460 40477 6469 40511
rect 6469 40477 6503 40511
rect 6503 40477 6512 40511
rect 6460 40468 6512 40477
rect 8484 40468 8536 40520
rect 12900 40536 12952 40588
rect 16580 40604 16632 40656
rect 17592 40604 17644 40656
rect 22008 40604 22060 40656
rect 22100 40604 22152 40656
rect 23572 40604 23624 40656
rect 23940 40604 23992 40656
rect 24032 40604 24084 40656
rect 12716 40468 12768 40520
rect 13360 40536 13412 40588
rect 17224 40579 17276 40588
rect 17224 40545 17233 40579
rect 17233 40545 17267 40579
rect 17267 40545 17276 40579
rect 17224 40536 17276 40545
rect 17316 40579 17368 40588
rect 17316 40545 17325 40579
rect 17325 40545 17359 40579
rect 17359 40545 17368 40579
rect 17316 40536 17368 40545
rect 21456 40579 21508 40588
rect 21456 40545 21465 40579
rect 21465 40545 21499 40579
rect 21499 40545 21508 40579
rect 21456 40536 21508 40545
rect 21548 40536 21600 40588
rect 23388 40536 23440 40588
rect 13728 40468 13780 40520
rect 15292 40468 15344 40520
rect 15752 40468 15804 40520
rect 17868 40468 17920 40520
rect 20628 40468 20680 40520
rect 8668 40400 8720 40452
rect 10232 40400 10284 40452
rect 8484 40375 8536 40384
rect 8484 40341 8493 40375
rect 8493 40341 8527 40375
rect 8527 40341 8536 40375
rect 8484 40332 8536 40341
rect 9404 40332 9456 40384
rect 9680 40332 9732 40384
rect 12072 40332 12124 40384
rect 13544 40400 13596 40452
rect 13820 40400 13872 40452
rect 19708 40400 19760 40452
rect 20536 40400 20588 40452
rect 22008 40468 22060 40520
rect 22652 40468 22704 40520
rect 22836 40511 22888 40520
rect 22836 40477 22845 40511
rect 22845 40477 22879 40511
rect 22879 40477 22888 40511
rect 22836 40468 22888 40477
rect 24032 40511 24084 40520
rect 24032 40477 24041 40511
rect 24041 40477 24075 40511
rect 24075 40477 24084 40511
rect 24032 40468 24084 40477
rect 24216 40468 24268 40520
rect 24492 40468 24544 40520
rect 24860 40468 24912 40520
rect 22928 40400 22980 40452
rect 23388 40400 23440 40452
rect 12900 40332 12952 40384
rect 15016 40332 15068 40384
rect 16856 40332 16908 40384
rect 21364 40332 21416 40384
rect 21824 40332 21876 40384
rect 22376 40332 22428 40384
rect 23572 40332 23624 40384
rect 24860 40332 24912 40384
rect 7950 40230 8002 40282
rect 8014 40230 8066 40282
rect 8078 40230 8130 40282
rect 8142 40230 8194 40282
rect 8206 40230 8258 40282
rect 17950 40230 18002 40282
rect 18014 40230 18066 40282
rect 18078 40230 18130 40282
rect 18142 40230 18194 40282
rect 18206 40230 18258 40282
rect 7012 40128 7064 40180
rect 8852 40128 8904 40180
rect 9680 40128 9732 40180
rect 12072 40171 12124 40180
rect 12072 40137 12081 40171
rect 12081 40137 12115 40171
rect 12115 40137 12124 40171
rect 12072 40128 12124 40137
rect 8392 40060 8444 40112
rect 8576 40060 8628 40112
rect 9496 40060 9548 40112
rect 10600 40060 10652 40112
rect 10784 40060 10836 40112
rect 14740 40171 14792 40180
rect 14740 40137 14749 40171
rect 14749 40137 14783 40171
rect 14783 40137 14792 40171
rect 14740 40128 14792 40137
rect 15108 40128 15160 40180
rect 18236 40171 18288 40180
rect 18236 40137 18245 40171
rect 18245 40137 18279 40171
rect 18279 40137 18288 40171
rect 18236 40128 18288 40137
rect 19340 40128 19392 40180
rect 19984 40128 20036 40180
rect 22100 40171 22152 40180
rect 22100 40137 22109 40171
rect 22109 40137 22143 40171
rect 22143 40137 22152 40171
rect 22100 40128 22152 40137
rect 22376 40171 22428 40180
rect 22376 40137 22385 40171
rect 22385 40137 22419 40171
rect 22419 40137 22428 40171
rect 22376 40128 22428 40137
rect 22652 40128 22704 40180
rect 11336 39992 11388 40044
rect 7748 39924 7800 39976
rect 8576 39924 8628 39976
rect 8668 39967 8720 39976
rect 8668 39933 8677 39967
rect 8677 39933 8711 39967
rect 8711 39933 8720 39967
rect 8668 39924 8720 39933
rect 12716 39992 12768 40044
rect 14372 39992 14424 40044
rect 15292 40060 15344 40112
rect 16580 40060 16632 40112
rect 15200 39992 15252 40044
rect 11520 39788 11572 39840
rect 16120 39967 16172 39976
rect 16120 39933 16129 39967
rect 16129 39933 16163 39967
rect 16163 39933 16172 39967
rect 16120 39924 16172 39933
rect 16488 39992 16540 40044
rect 16672 39924 16724 39976
rect 17776 39924 17828 39976
rect 18420 39924 18472 39976
rect 18880 39967 18932 39976
rect 18880 39933 18889 39967
rect 18889 39933 18923 39967
rect 18923 39933 18932 39967
rect 18880 39924 18932 39933
rect 22468 40060 22520 40112
rect 24400 40060 24452 40112
rect 14648 39788 14700 39840
rect 19248 39788 19300 39840
rect 22928 39992 22980 40044
rect 20076 39967 20128 39976
rect 20076 39933 20085 39967
rect 20085 39933 20119 39967
rect 20119 39933 20128 39967
rect 20076 39924 20128 39933
rect 21272 39967 21324 39976
rect 21272 39933 21281 39967
rect 21281 39933 21315 39967
rect 21315 39933 21324 39967
rect 21272 39924 21324 39933
rect 21824 39924 21876 39976
rect 22376 39924 22428 39976
rect 25228 39924 25280 39976
rect 21916 39831 21968 39840
rect 21916 39797 21925 39831
rect 21925 39797 21959 39831
rect 21959 39797 21968 39831
rect 21916 39788 21968 39797
rect 22836 39831 22888 39840
rect 22836 39797 22845 39831
rect 22845 39797 22879 39831
rect 22879 39797 22888 39831
rect 22836 39788 22888 39797
rect 25320 39856 25372 39908
rect 2950 39686 3002 39738
rect 3014 39686 3066 39738
rect 3078 39686 3130 39738
rect 3142 39686 3194 39738
rect 3206 39686 3258 39738
rect 12950 39686 13002 39738
rect 13014 39686 13066 39738
rect 13078 39686 13130 39738
rect 13142 39686 13194 39738
rect 13206 39686 13258 39738
rect 22950 39686 23002 39738
rect 23014 39686 23066 39738
rect 23078 39686 23130 39738
rect 23142 39686 23194 39738
rect 23206 39686 23258 39738
rect 5908 39584 5960 39636
rect 6460 39448 6512 39500
rect 7380 39584 7432 39636
rect 8484 39627 8536 39636
rect 8484 39593 8493 39627
rect 8493 39593 8527 39627
rect 8527 39593 8536 39627
rect 8484 39584 8536 39593
rect 8576 39584 8628 39636
rect 11888 39584 11940 39636
rect 8668 39516 8720 39568
rect 12532 39584 12584 39636
rect 13360 39584 13412 39636
rect 13820 39584 13872 39636
rect 14188 39584 14240 39636
rect 16856 39584 16908 39636
rect 22744 39584 22796 39636
rect 5172 39423 5224 39432
rect 5172 39389 5181 39423
rect 5181 39389 5215 39423
rect 5215 39389 5224 39423
rect 5172 39380 5224 39389
rect 8576 39448 8628 39500
rect 9128 39448 9180 39500
rect 13636 39516 13688 39568
rect 19156 39516 19208 39568
rect 21088 39516 21140 39568
rect 21732 39516 21784 39568
rect 8760 39380 8812 39432
rect 9312 39380 9364 39432
rect 11980 39448 12032 39500
rect 12716 39448 12768 39500
rect 13912 39448 13964 39500
rect 15384 39448 15436 39500
rect 15568 39448 15620 39500
rect 12348 39380 12400 39432
rect 13636 39380 13688 39432
rect 14372 39380 14424 39432
rect 18604 39448 18656 39500
rect 18788 39448 18840 39500
rect 21824 39491 21876 39500
rect 21824 39457 21833 39491
rect 21833 39457 21867 39491
rect 21867 39457 21876 39491
rect 21824 39448 21876 39457
rect 23664 39448 23716 39500
rect 25044 39491 25096 39500
rect 25044 39457 25053 39491
rect 25053 39457 25087 39491
rect 25087 39457 25096 39491
rect 25044 39448 25096 39457
rect 25136 39491 25188 39500
rect 25136 39457 25145 39491
rect 25145 39457 25179 39491
rect 25179 39457 25188 39491
rect 25136 39448 25188 39457
rect 20444 39380 20496 39432
rect 20628 39380 20680 39432
rect 5448 39355 5500 39364
rect 5448 39321 5457 39355
rect 5457 39321 5491 39355
rect 5491 39321 5500 39355
rect 5448 39312 5500 39321
rect 8668 39355 8720 39364
rect 6460 39244 6512 39296
rect 8668 39321 8677 39355
rect 8677 39321 8711 39355
rect 8711 39321 8720 39355
rect 8668 39312 8720 39321
rect 9404 39312 9456 39364
rect 10048 39244 10100 39296
rect 12992 39244 13044 39296
rect 13084 39287 13136 39296
rect 13084 39253 13093 39287
rect 13093 39253 13127 39287
rect 13127 39253 13136 39287
rect 13084 39244 13136 39253
rect 13820 39244 13872 39296
rect 14004 39244 14056 39296
rect 14832 39287 14884 39296
rect 14832 39253 14841 39287
rect 14841 39253 14875 39287
rect 14875 39253 14884 39287
rect 14832 39244 14884 39253
rect 15200 39244 15252 39296
rect 17224 39244 17276 39296
rect 19984 39312 20036 39364
rect 21364 39312 21416 39364
rect 20076 39244 20128 39296
rect 24768 39244 24820 39296
rect 7950 39142 8002 39194
rect 8014 39142 8066 39194
rect 8078 39142 8130 39194
rect 8142 39142 8194 39194
rect 8206 39142 8258 39194
rect 17950 39142 18002 39194
rect 18014 39142 18066 39194
rect 18078 39142 18130 39194
rect 18142 39142 18194 39194
rect 18206 39142 18258 39194
rect 5448 39040 5500 39092
rect 6552 39083 6604 39092
rect 6552 39049 6561 39083
rect 6561 39049 6595 39083
rect 6595 39049 6604 39083
rect 6552 39040 6604 39049
rect 8392 39040 8444 39092
rect 10692 39040 10744 39092
rect 12164 39040 12216 39092
rect 12624 39040 12676 39092
rect 5816 38972 5868 39024
rect 5448 38904 5500 38956
rect 8944 38972 8996 39024
rect 9588 38972 9640 39024
rect 10968 38972 11020 39024
rect 16120 39040 16172 39092
rect 18604 39083 18656 39092
rect 18604 39049 18613 39083
rect 18613 39049 18647 39083
rect 18647 39049 18656 39083
rect 18604 39040 18656 39049
rect 19432 39083 19484 39092
rect 19432 39049 19441 39083
rect 19441 39049 19475 39083
rect 19475 39049 19484 39083
rect 19432 39040 19484 39049
rect 20996 39083 21048 39092
rect 20996 39049 21005 39083
rect 21005 39049 21039 39083
rect 21039 39049 21048 39083
rect 20996 39040 21048 39049
rect 21088 39083 21140 39092
rect 21088 39049 21097 39083
rect 21097 39049 21131 39083
rect 21131 39049 21140 39083
rect 21088 39040 21140 39049
rect 22836 39040 22888 39092
rect 14648 38972 14700 39024
rect 15476 38972 15528 39024
rect 7748 38947 7800 38956
rect 7748 38913 7757 38947
rect 7757 38913 7791 38947
rect 7791 38913 7800 38947
rect 7748 38904 7800 38913
rect 7840 38904 7892 38956
rect 9588 38879 9640 38888
rect 9588 38845 9597 38879
rect 9597 38845 9631 38879
rect 9631 38845 9640 38879
rect 9588 38836 9640 38845
rect 11704 38904 11756 38956
rect 12716 38904 12768 38956
rect 13084 38904 13136 38956
rect 14740 38904 14792 38956
rect 16672 38904 16724 38956
rect 17224 38972 17276 39024
rect 18972 38972 19024 39024
rect 19892 38972 19944 39024
rect 25228 39083 25280 39092
rect 25228 39049 25237 39083
rect 25237 39049 25271 39083
rect 25271 39049 25280 39083
rect 25228 39040 25280 39049
rect 24400 38972 24452 39024
rect 19524 38904 19576 38956
rect 8944 38768 8996 38820
rect 10140 38768 10192 38820
rect 10876 38879 10928 38888
rect 10876 38845 10885 38879
rect 10885 38845 10919 38879
rect 10919 38845 10928 38879
rect 10876 38836 10928 38845
rect 12532 38836 12584 38888
rect 12992 38836 13044 38888
rect 15108 38836 15160 38888
rect 15384 38879 15436 38888
rect 15384 38845 15393 38879
rect 15393 38845 15427 38879
rect 15427 38845 15436 38879
rect 15384 38836 15436 38845
rect 15752 38836 15804 38888
rect 24492 38904 24544 38956
rect 13820 38768 13872 38820
rect 15660 38768 15712 38820
rect 21272 38879 21324 38888
rect 21272 38845 21281 38879
rect 21281 38845 21315 38879
rect 21315 38845 21324 38879
rect 21272 38836 21324 38845
rect 22376 38879 22428 38888
rect 22376 38845 22385 38879
rect 22385 38845 22419 38879
rect 22419 38845 22428 38879
rect 22376 38836 22428 38845
rect 24860 38836 24912 38888
rect 20536 38768 20588 38820
rect 22008 38768 22060 38820
rect 6828 38700 6880 38752
rect 9588 38700 9640 38752
rect 12164 38700 12216 38752
rect 14004 38700 14056 38752
rect 14096 38743 14148 38752
rect 14096 38709 14105 38743
rect 14105 38709 14139 38743
rect 14139 38709 14148 38743
rect 14096 38700 14148 38709
rect 14188 38700 14240 38752
rect 15384 38700 15436 38752
rect 15936 38743 15988 38752
rect 15936 38709 15945 38743
rect 15945 38709 15979 38743
rect 15979 38709 15988 38743
rect 15936 38700 15988 38709
rect 21364 38700 21416 38752
rect 24032 38700 24084 38752
rect 24860 38700 24912 38752
rect 2950 38598 3002 38650
rect 3014 38598 3066 38650
rect 3078 38598 3130 38650
rect 3142 38598 3194 38650
rect 3206 38598 3258 38650
rect 12950 38598 13002 38650
rect 13014 38598 13066 38650
rect 13078 38598 13130 38650
rect 13142 38598 13194 38650
rect 13206 38598 13258 38650
rect 22950 38598 23002 38650
rect 23014 38598 23066 38650
rect 23078 38598 23130 38650
rect 23142 38598 23194 38650
rect 23206 38598 23258 38650
rect 6092 38496 6144 38548
rect 5172 38360 5224 38412
rect 7564 38496 7616 38548
rect 10508 38496 10560 38548
rect 14096 38496 14148 38548
rect 15108 38496 15160 38548
rect 9220 38428 9272 38480
rect 1308 38292 1360 38344
rect 9680 38403 9732 38412
rect 9680 38369 9689 38403
rect 9689 38369 9723 38403
rect 9723 38369 9732 38403
rect 9680 38360 9732 38369
rect 9864 38360 9916 38412
rect 10968 38403 11020 38412
rect 10968 38369 10977 38403
rect 10977 38369 11011 38403
rect 11011 38369 11020 38403
rect 10968 38360 11020 38369
rect 11980 38403 12032 38412
rect 11980 38369 11989 38403
rect 11989 38369 12023 38403
rect 12023 38369 12032 38403
rect 11980 38360 12032 38369
rect 13360 38428 13412 38480
rect 12624 38360 12676 38412
rect 16580 38496 16632 38548
rect 18696 38496 18748 38548
rect 21548 38496 21600 38548
rect 24676 38496 24728 38548
rect 14832 38360 14884 38412
rect 18512 38428 18564 38480
rect 22100 38428 22152 38480
rect 24584 38471 24636 38480
rect 24584 38437 24593 38471
rect 24593 38437 24627 38471
rect 24627 38437 24636 38471
rect 24584 38428 24636 38437
rect 17500 38360 17552 38412
rect 18420 38403 18472 38412
rect 18420 38369 18429 38403
rect 18429 38369 18463 38403
rect 18463 38369 18472 38403
rect 18420 38360 18472 38369
rect 21548 38360 21600 38412
rect 22284 38360 22336 38412
rect 6000 38224 6052 38276
rect 6460 38224 6512 38276
rect 7012 38224 7064 38276
rect 10048 38292 10100 38344
rect 15844 38292 15896 38344
rect 17132 38292 17184 38344
rect 24032 38360 24084 38412
rect 24400 38360 24452 38412
rect 23480 38292 23532 38344
rect 25412 38292 25464 38344
rect 11244 38224 11296 38276
rect 13636 38224 13688 38276
rect 3884 38156 3936 38208
rect 7748 38156 7800 38208
rect 7840 38156 7892 38208
rect 9864 38156 9916 38208
rect 10692 38156 10744 38208
rect 10968 38156 11020 38208
rect 17500 38224 17552 38276
rect 18788 38224 18840 38276
rect 20168 38267 20220 38276
rect 20168 38233 20177 38267
rect 20177 38233 20211 38267
rect 20211 38233 20220 38267
rect 20168 38224 20220 38233
rect 22008 38224 22060 38276
rect 22376 38224 22428 38276
rect 22836 38224 22888 38276
rect 23204 38224 23256 38276
rect 24676 38224 24728 38276
rect 15384 38199 15436 38208
rect 15384 38165 15393 38199
rect 15393 38165 15427 38199
rect 15427 38165 15436 38199
rect 15384 38156 15436 38165
rect 16580 38199 16632 38208
rect 16580 38165 16589 38199
rect 16589 38165 16623 38199
rect 16623 38165 16632 38199
rect 16580 38156 16632 38165
rect 18420 38156 18472 38208
rect 18880 38156 18932 38208
rect 19064 38156 19116 38208
rect 22744 38199 22796 38208
rect 22744 38165 22753 38199
rect 22753 38165 22787 38199
rect 22787 38165 22796 38199
rect 22744 38156 22796 38165
rect 22928 38156 22980 38208
rect 25596 38156 25648 38208
rect 7950 38054 8002 38106
rect 8014 38054 8066 38106
rect 8078 38054 8130 38106
rect 8142 38054 8194 38106
rect 8206 38054 8258 38106
rect 17950 38054 18002 38106
rect 18014 38054 18066 38106
rect 18078 38054 18130 38106
rect 18142 38054 18194 38106
rect 18206 38054 18258 38106
rect 6000 37995 6052 38004
rect 6000 37961 6009 37995
rect 6009 37961 6043 37995
rect 6043 37961 6052 37995
rect 6000 37952 6052 37961
rect 6644 37952 6696 38004
rect 6828 37927 6880 37936
rect 6828 37893 6837 37927
rect 6837 37893 6871 37927
rect 6871 37893 6880 37927
rect 6828 37884 6880 37893
rect 8208 37884 8260 37936
rect 8668 37884 8720 37936
rect 9036 37952 9088 38004
rect 9496 37952 9548 38004
rect 10600 37952 10652 38004
rect 10968 37952 11020 38004
rect 11428 37952 11480 38004
rect 11704 37995 11756 38004
rect 11704 37961 11713 37995
rect 11713 37961 11747 37995
rect 11747 37961 11756 37995
rect 11704 37952 11756 37961
rect 13636 37952 13688 38004
rect 14004 37952 14056 38004
rect 15384 37995 15436 38004
rect 15384 37961 15393 37995
rect 15393 37961 15427 37995
rect 15427 37961 15436 37995
rect 15384 37952 15436 37961
rect 16580 37952 16632 38004
rect 17500 37995 17552 38004
rect 17500 37961 17509 37995
rect 17509 37961 17543 37995
rect 17543 37961 17552 37995
rect 17500 37952 17552 37961
rect 18696 37952 18748 38004
rect 19616 37952 19668 38004
rect 22008 37995 22060 38004
rect 22008 37961 22017 37995
rect 22017 37961 22051 37995
rect 22051 37961 22060 37995
rect 22008 37952 22060 37961
rect 22100 37952 22152 38004
rect 22652 37952 22704 38004
rect 10508 37884 10560 37936
rect 10692 37927 10744 37936
rect 10692 37893 10701 37927
rect 10701 37893 10735 37927
rect 10735 37893 10744 37927
rect 10692 37884 10744 37893
rect 11520 37884 11572 37936
rect 9404 37816 9456 37868
rect 11336 37816 11388 37868
rect 15108 37816 15160 37868
rect 6552 37791 6604 37800
rect 6552 37757 6561 37791
rect 6561 37757 6595 37791
rect 6595 37757 6604 37791
rect 6552 37748 6604 37757
rect 7196 37748 7248 37800
rect 8576 37612 8628 37664
rect 9588 37680 9640 37732
rect 11428 37748 11480 37800
rect 13636 37748 13688 37800
rect 15292 37748 15344 37800
rect 11520 37680 11572 37732
rect 11704 37680 11756 37732
rect 12256 37655 12308 37664
rect 12256 37621 12265 37655
rect 12265 37621 12299 37655
rect 12299 37621 12308 37655
rect 12256 37612 12308 37621
rect 12532 37655 12584 37664
rect 12532 37621 12541 37655
rect 12541 37621 12575 37655
rect 12575 37621 12584 37655
rect 12532 37612 12584 37621
rect 12716 37612 12768 37664
rect 14280 37612 14332 37664
rect 15384 37612 15436 37664
rect 16212 37816 16264 37868
rect 21916 37884 21968 37936
rect 22928 37884 22980 37936
rect 23388 37884 23440 37936
rect 18880 37816 18932 37868
rect 19340 37816 19392 37868
rect 20444 37816 20496 37868
rect 15752 37748 15804 37800
rect 21456 37816 21508 37868
rect 24216 37952 24268 38004
rect 24860 37884 24912 37936
rect 16028 37680 16080 37732
rect 18420 37680 18472 37732
rect 21180 37791 21232 37800
rect 21180 37757 21189 37791
rect 21189 37757 21223 37791
rect 21223 37757 21232 37791
rect 21180 37748 21232 37757
rect 22836 37748 22888 37800
rect 23848 37791 23900 37800
rect 23848 37757 23857 37791
rect 23857 37757 23891 37791
rect 23891 37757 23900 37791
rect 23848 37748 23900 37757
rect 20720 37680 20772 37732
rect 22192 37680 22244 37732
rect 23204 37680 23256 37732
rect 17868 37612 17920 37664
rect 18696 37612 18748 37664
rect 19064 37612 19116 37664
rect 20260 37612 20312 37664
rect 21916 37612 21968 37664
rect 22376 37612 22428 37664
rect 23388 37612 23440 37664
rect 23940 37612 23992 37664
rect 24492 37612 24544 37664
rect 2950 37510 3002 37562
rect 3014 37510 3066 37562
rect 3078 37510 3130 37562
rect 3142 37510 3194 37562
rect 3206 37510 3258 37562
rect 12950 37510 13002 37562
rect 13014 37510 13066 37562
rect 13078 37510 13130 37562
rect 13142 37510 13194 37562
rect 13206 37510 13258 37562
rect 22950 37510 23002 37562
rect 23014 37510 23066 37562
rect 23078 37510 23130 37562
rect 23142 37510 23194 37562
rect 23206 37510 23258 37562
rect 6460 37408 6512 37460
rect 6920 37408 6972 37460
rect 6644 37340 6696 37392
rect 8576 37451 8628 37460
rect 8576 37417 8585 37451
rect 8585 37417 8619 37451
rect 8619 37417 8628 37451
rect 8576 37408 8628 37417
rect 9312 37408 9364 37460
rect 9864 37340 9916 37392
rect 5632 37272 5684 37324
rect 6552 37272 6604 37324
rect 8576 37272 8628 37324
rect 8208 37204 8260 37256
rect 10416 37408 10468 37460
rect 10968 37408 11020 37460
rect 12256 37408 12308 37460
rect 13084 37408 13136 37460
rect 13820 37408 13872 37460
rect 16304 37408 16356 37460
rect 18696 37408 18748 37460
rect 19248 37408 19300 37460
rect 19340 37451 19392 37460
rect 19340 37417 19349 37451
rect 19349 37417 19383 37451
rect 19383 37417 19392 37451
rect 19340 37408 19392 37417
rect 20904 37408 20956 37460
rect 21640 37408 21692 37460
rect 22100 37408 22152 37460
rect 23848 37408 23900 37460
rect 16488 37340 16540 37392
rect 10324 37272 10376 37324
rect 10600 37315 10652 37324
rect 10600 37281 10609 37315
rect 10609 37281 10643 37315
rect 10643 37281 10652 37315
rect 10600 37272 10652 37281
rect 10968 37272 11020 37324
rect 13084 37272 13136 37324
rect 13360 37272 13412 37324
rect 16396 37272 16448 37324
rect 17868 37315 17920 37324
rect 17868 37281 17877 37315
rect 17877 37281 17911 37315
rect 17911 37281 17920 37315
rect 17868 37272 17920 37281
rect 11152 37204 11204 37256
rect 11704 37247 11756 37256
rect 11704 37213 11713 37247
rect 11713 37213 11747 37247
rect 11747 37213 11756 37247
rect 11704 37204 11756 37213
rect 14188 37204 14240 37256
rect 15384 37204 15436 37256
rect 18788 37204 18840 37256
rect 6460 37136 6512 37188
rect 10508 37136 10560 37188
rect 10692 37136 10744 37188
rect 5632 37068 5684 37120
rect 5816 37111 5868 37120
rect 5816 37077 5825 37111
rect 5825 37077 5859 37111
rect 5859 37077 5868 37111
rect 5816 37068 5868 37077
rect 11152 37068 11204 37120
rect 12808 37136 12860 37188
rect 12716 37068 12768 37120
rect 13084 37136 13136 37188
rect 17776 37136 17828 37188
rect 23664 37340 23716 37392
rect 19156 37272 19208 37324
rect 19294 37204 19346 37256
rect 18972 37179 19024 37188
rect 14280 37111 14332 37120
rect 14280 37077 14289 37111
rect 14289 37077 14323 37111
rect 14323 37077 14332 37111
rect 14280 37068 14332 37077
rect 14464 37068 14516 37120
rect 15936 37068 15988 37120
rect 16120 37111 16172 37120
rect 16120 37077 16129 37111
rect 16129 37077 16163 37111
rect 16163 37077 16172 37111
rect 16120 37068 16172 37077
rect 17316 37111 17368 37120
rect 17316 37077 17325 37111
rect 17325 37077 17359 37111
rect 17359 37077 17368 37111
rect 17316 37068 17368 37077
rect 18512 37111 18564 37120
rect 18512 37077 18521 37111
rect 18521 37077 18555 37111
rect 18555 37077 18564 37111
rect 18512 37068 18564 37077
rect 18972 37145 18981 37179
rect 18981 37145 19015 37179
rect 19015 37145 19024 37179
rect 18972 37136 19024 37145
rect 20536 37247 20588 37256
rect 20536 37213 20545 37247
rect 20545 37213 20579 37247
rect 20579 37213 20588 37247
rect 20536 37204 20588 37213
rect 20904 37204 20956 37256
rect 21916 37247 21968 37256
rect 21916 37213 21925 37247
rect 21925 37213 21959 37247
rect 21959 37213 21968 37247
rect 21916 37204 21968 37213
rect 22560 37272 22612 37324
rect 23112 37272 23164 37324
rect 22100 37204 22152 37256
rect 21824 37068 21876 37120
rect 22652 37068 22704 37120
rect 23296 37204 23348 37256
rect 24400 37204 24452 37256
rect 24952 37204 25004 37256
rect 25044 37204 25096 37256
rect 24676 37136 24728 37188
rect 23480 37068 23532 37120
rect 23848 37068 23900 37120
rect 24584 37068 24636 37120
rect 7950 36966 8002 37018
rect 8014 36966 8066 37018
rect 8078 36966 8130 37018
rect 8142 36966 8194 37018
rect 8206 36966 8258 37018
rect 17950 36966 18002 37018
rect 18014 36966 18066 37018
rect 18078 36966 18130 37018
rect 18142 36966 18194 37018
rect 18206 36966 18258 37018
rect 6460 36864 6512 36916
rect 7288 36907 7340 36916
rect 7288 36873 7297 36907
rect 7297 36873 7331 36907
rect 7331 36873 7340 36907
rect 7288 36864 7340 36873
rect 11060 36864 11112 36916
rect 13084 36864 13136 36916
rect 14280 36864 14332 36916
rect 14924 36907 14976 36916
rect 14924 36873 14933 36907
rect 14933 36873 14967 36907
rect 14967 36873 14976 36907
rect 14924 36864 14976 36873
rect 17132 36864 17184 36916
rect 18512 36864 18564 36916
rect 18696 36864 18748 36916
rect 10784 36796 10836 36848
rect 9680 36660 9732 36712
rect 12440 36728 12492 36780
rect 13360 36728 13412 36780
rect 12808 36660 12860 36712
rect 13268 36660 13320 36712
rect 14096 36728 14148 36780
rect 14832 36771 14884 36780
rect 14832 36737 14841 36771
rect 14841 36737 14875 36771
rect 14875 36737 14884 36771
rect 14832 36728 14884 36737
rect 13820 36660 13872 36712
rect 17224 36796 17276 36848
rect 19156 36796 19208 36848
rect 20628 36864 20680 36916
rect 21640 36864 21692 36916
rect 22560 36864 22612 36916
rect 23204 36864 23256 36916
rect 24400 36864 24452 36916
rect 16672 36771 16724 36780
rect 16672 36737 16681 36771
rect 16681 36737 16715 36771
rect 16715 36737 16724 36771
rect 16672 36728 16724 36737
rect 18604 36728 18656 36780
rect 18788 36728 18840 36780
rect 19248 36728 19300 36780
rect 19616 36728 19668 36780
rect 20444 36771 20496 36780
rect 20444 36737 20453 36771
rect 20453 36737 20487 36771
rect 20487 36737 20496 36771
rect 20444 36728 20496 36737
rect 21088 36728 21140 36780
rect 23388 36796 23440 36848
rect 24860 36864 24912 36916
rect 24400 36728 24452 36780
rect 24860 36728 24912 36780
rect 19800 36660 19852 36712
rect 21732 36660 21784 36712
rect 22652 36660 22704 36712
rect 22836 36703 22888 36712
rect 22836 36669 22845 36703
rect 22845 36669 22879 36703
rect 22879 36669 22888 36703
rect 22836 36660 22888 36669
rect 23112 36703 23164 36712
rect 23112 36669 23121 36703
rect 23121 36669 23155 36703
rect 23155 36669 23164 36703
rect 23112 36660 23164 36669
rect 23480 36660 23532 36712
rect 11244 36592 11296 36644
rect 17316 36592 17368 36644
rect 7196 36567 7248 36576
rect 7196 36533 7205 36567
rect 7205 36533 7239 36567
rect 7239 36533 7248 36567
rect 7196 36524 7248 36533
rect 8576 36524 8628 36576
rect 9496 36524 9548 36576
rect 12440 36524 12492 36576
rect 14372 36524 14424 36576
rect 14464 36567 14516 36576
rect 14464 36533 14473 36567
rect 14473 36533 14507 36567
rect 14507 36533 14516 36567
rect 14464 36524 14516 36533
rect 14832 36524 14884 36576
rect 19984 36592 20036 36644
rect 18328 36524 18380 36576
rect 19616 36567 19668 36576
rect 19616 36533 19625 36567
rect 19625 36533 19659 36567
rect 19659 36533 19668 36567
rect 19616 36524 19668 36533
rect 20444 36524 20496 36576
rect 21088 36567 21140 36576
rect 21088 36533 21097 36567
rect 21097 36533 21131 36567
rect 21131 36533 21140 36567
rect 21088 36524 21140 36533
rect 2950 36422 3002 36474
rect 3014 36422 3066 36474
rect 3078 36422 3130 36474
rect 3142 36422 3194 36474
rect 3206 36422 3258 36474
rect 12950 36422 13002 36474
rect 13014 36422 13066 36474
rect 13078 36422 13130 36474
rect 13142 36422 13194 36474
rect 13206 36422 13258 36474
rect 22950 36422 23002 36474
rect 23014 36422 23066 36474
rect 23078 36422 23130 36474
rect 23142 36422 23194 36474
rect 23206 36422 23258 36474
rect 7012 36363 7064 36372
rect 7012 36329 7021 36363
rect 7021 36329 7055 36363
rect 7055 36329 7064 36363
rect 7012 36320 7064 36329
rect 7288 36363 7340 36372
rect 7288 36329 7297 36363
rect 7297 36329 7331 36363
rect 7331 36329 7340 36363
rect 7288 36320 7340 36329
rect 7656 36320 7708 36372
rect 8944 36320 8996 36372
rect 9956 36320 10008 36372
rect 10324 36320 10376 36372
rect 11060 36363 11112 36372
rect 11060 36329 11069 36363
rect 11069 36329 11103 36363
rect 11103 36329 11112 36363
rect 11060 36320 11112 36329
rect 11244 36363 11296 36372
rect 11244 36329 11253 36363
rect 11253 36329 11287 36363
rect 11287 36329 11296 36363
rect 11244 36320 11296 36329
rect 5632 36184 5684 36236
rect 7656 36184 7708 36236
rect 8760 36184 8812 36236
rect 1768 36159 1820 36168
rect 1768 36125 1777 36159
rect 1777 36125 1811 36159
rect 1811 36125 1820 36159
rect 1768 36116 1820 36125
rect 12532 36184 12584 36236
rect 11060 36116 11112 36168
rect 1584 36023 1636 36032
rect 1584 35989 1593 36023
rect 1593 35989 1627 36023
rect 1627 35989 1636 36023
rect 1584 35980 1636 35989
rect 6828 36048 6880 36100
rect 7288 36048 7340 36100
rect 7196 35980 7248 36032
rect 7564 35980 7616 36032
rect 10232 35980 10284 36032
rect 11704 36048 11756 36100
rect 12624 35980 12676 36032
rect 13452 36320 13504 36372
rect 15200 36320 15252 36372
rect 16212 36363 16264 36372
rect 16212 36329 16221 36363
rect 16221 36329 16255 36363
rect 16255 36329 16264 36363
rect 16212 36320 16264 36329
rect 17040 36320 17092 36372
rect 17592 36320 17644 36372
rect 22652 36320 22704 36372
rect 25044 36320 25096 36372
rect 15016 36252 15068 36304
rect 13360 36184 13412 36236
rect 15568 36184 15620 36236
rect 16948 36184 17000 36236
rect 15660 36116 15712 36168
rect 21364 36227 21416 36236
rect 21364 36193 21373 36227
rect 21373 36193 21407 36227
rect 21407 36193 21416 36227
rect 21364 36184 21416 36193
rect 21272 36116 21324 36168
rect 24492 36252 24544 36304
rect 23940 36227 23992 36236
rect 23940 36193 23949 36227
rect 23949 36193 23983 36227
rect 23983 36193 23992 36227
rect 23940 36184 23992 36193
rect 23848 36116 23900 36168
rect 21180 36048 21232 36100
rect 22100 36048 22152 36100
rect 25504 36184 25556 36236
rect 24676 36116 24728 36168
rect 13820 35980 13872 36032
rect 14372 35980 14424 36032
rect 16672 36023 16724 36032
rect 16672 35989 16681 36023
rect 16681 35989 16715 36023
rect 16715 35989 16724 36023
rect 16672 35980 16724 35989
rect 19984 35980 20036 36032
rect 20996 35980 21048 36032
rect 22652 36023 22704 36032
rect 22652 35989 22661 36023
rect 22661 35989 22695 36023
rect 22695 35989 22704 36023
rect 22652 35980 22704 35989
rect 23664 36023 23716 36032
rect 23664 35989 23673 36023
rect 23673 35989 23707 36023
rect 23707 35989 23716 36023
rect 23664 35980 23716 35989
rect 24400 36023 24452 36032
rect 24400 35989 24409 36023
rect 24409 35989 24443 36023
rect 24443 35989 24452 36023
rect 24400 35980 24452 35989
rect 24676 36023 24728 36032
rect 24676 35989 24685 36023
rect 24685 35989 24719 36023
rect 24719 35989 24728 36023
rect 24676 35980 24728 35989
rect 24860 36023 24912 36032
rect 24860 35989 24869 36023
rect 24869 35989 24903 36023
rect 24903 35989 24912 36023
rect 24860 35980 24912 35989
rect 25136 36023 25188 36032
rect 25136 35989 25145 36023
rect 25145 35989 25179 36023
rect 25179 35989 25188 36023
rect 25136 35980 25188 35989
rect 7950 35878 8002 35930
rect 8014 35878 8066 35930
rect 8078 35878 8130 35930
rect 8142 35878 8194 35930
rect 8206 35878 8258 35930
rect 17950 35878 18002 35930
rect 18014 35878 18066 35930
rect 18078 35878 18130 35930
rect 18142 35878 18194 35930
rect 18206 35878 18258 35930
rect 6092 35776 6144 35828
rect 6828 35776 6880 35828
rect 13360 35776 13412 35828
rect 13636 35776 13688 35828
rect 13912 35776 13964 35828
rect 15936 35776 15988 35828
rect 7288 35708 7340 35760
rect 8116 35708 8168 35760
rect 13452 35708 13504 35760
rect 14004 35708 14056 35760
rect 11704 35683 11756 35692
rect 11704 35649 11713 35683
rect 11713 35649 11747 35683
rect 11747 35649 11756 35683
rect 11704 35640 11756 35649
rect 7012 35504 7064 35556
rect 5632 35436 5684 35488
rect 6552 35436 6604 35488
rect 9772 35572 9824 35624
rect 14740 35572 14792 35624
rect 8392 35436 8444 35488
rect 9864 35436 9916 35488
rect 12348 35436 12400 35488
rect 12532 35436 12584 35488
rect 13636 35504 13688 35556
rect 15476 35640 15528 35692
rect 16488 35640 16540 35692
rect 18052 35708 18104 35760
rect 18696 35708 18748 35760
rect 20352 35819 20404 35828
rect 20352 35785 20361 35819
rect 20361 35785 20395 35819
rect 20395 35785 20404 35819
rect 20352 35776 20404 35785
rect 22652 35776 22704 35828
rect 22928 35776 22980 35828
rect 23480 35776 23532 35828
rect 21916 35708 21968 35760
rect 22836 35708 22888 35760
rect 23388 35708 23440 35760
rect 25412 35708 25464 35760
rect 15016 35615 15068 35624
rect 15016 35581 15025 35615
rect 15025 35581 15059 35615
rect 15059 35581 15068 35615
rect 15016 35572 15068 35581
rect 18328 35572 18380 35624
rect 18604 35572 18656 35624
rect 17316 35504 17368 35556
rect 14188 35436 14240 35488
rect 15660 35436 15712 35488
rect 16672 35436 16724 35488
rect 19524 35436 19576 35488
rect 22468 35615 22520 35624
rect 22468 35581 22477 35615
rect 22477 35581 22511 35615
rect 22511 35581 22520 35615
rect 22468 35572 22520 35581
rect 23112 35572 23164 35624
rect 25228 35572 25280 35624
rect 20720 35436 20772 35488
rect 20996 35479 21048 35488
rect 20996 35445 21005 35479
rect 21005 35445 21039 35479
rect 21039 35445 21048 35479
rect 20996 35436 21048 35445
rect 23664 35436 23716 35488
rect 25412 35479 25464 35488
rect 25412 35445 25421 35479
rect 25421 35445 25455 35479
rect 25455 35445 25464 35479
rect 25412 35436 25464 35445
rect 2950 35334 3002 35386
rect 3014 35334 3066 35386
rect 3078 35334 3130 35386
rect 3142 35334 3194 35386
rect 3206 35334 3258 35386
rect 12950 35334 13002 35386
rect 13014 35334 13066 35386
rect 13078 35334 13130 35386
rect 13142 35334 13194 35386
rect 13206 35334 13258 35386
rect 22950 35334 23002 35386
rect 23014 35334 23066 35386
rect 23078 35334 23130 35386
rect 23142 35334 23194 35386
rect 23206 35334 23258 35386
rect 6644 35232 6696 35284
rect 8760 35232 8812 35284
rect 8852 35232 8904 35284
rect 11060 35232 11112 35284
rect 11336 35232 11388 35284
rect 8116 35164 8168 35216
rect 8392 35164 8444 35216
rect 9496 35164 9548 35216
rect 6092 35096 6144 35148
rect 6552 35139 6604 35148
rect 6552 35105 6561 35139
rect 6561 35105 6595 35139
rect 6595 35105 6604 35139
rect 6552 35096 6604 35105
rect 7748 35096 7800 35148
rect 5632 35028 5684 35080
rect 9312 35096 9364 35148
rect 11704 35164 11756 35216
rect 12716 35164 12768 35216
rect 14188 35164 14240 35216
rect 14740 35232 14792 35284
rect 15752 35232 15804 35284
rect 17316 35232 17368 35284
rect 8484 35028 8536 35080
rect 9864 35028 9916 35080
rect 11980 35028 12032 35080
rect 15476 35139 15528 35148
rect 15476 35105 15485 35139
rect 15485 35105 15519 35139
rect 15519 35105 15528 35139
rect 15476 35096 15528 35105
rect 19248 35164 19300 35216
rect 20996 35232 21048 35284
rect 22008 35164 22060 35216
rect 18052 35096 18104 35148
rect 18328 35096 18380 35148
rect 20168 35096 20220 35148
rect 23296 35096 23348 35148
rect 25228 35275 25280 35284
rect 25228 35241 25237 35275
rect 25237 35241 25271 35275
rect 25271 35241 25280 35275
rect 25228 35232 25280 35241
rect 14280 35071 14332 35080
rect 14280 35037 14289 35071
rect 14289 35037 14323 35071
rect 14323 35037 14332 35071
rect 14280 35028 14332 35037
rect 5816 34935 5868 34944
rect 5816 34901 5825 34935
rect 5825 34901 5859 34935
rect 5859 34901 5868 34935
rect 5816 34892 5868 34901
rect 7288 34892 7340 34944
rect 12348 34960 12400 35012
rect 13452 34960 13504 35012
rect 15752 35003 15804 35012
rect 15752 34969 15761 35003
rect 15761 34969 15795 35003
rect 15795 34969 15804 35003
rect 15752 34960 15804 34969
rect 11244 34892 11296 34944
rect 12072 34935 12124 34944
rect 12072 34901 12081 34935
rect 12081 34901 12115 34935
rect 12115 34901 12124 34935
rect 12072 34892 12124 34901
rect 14924 34892 14976 34944
rect 16580 34892 16632 34944
rect 24400 35096 24452 35148
rect 20996 34960 21048 35012
rect 22192 34960 22244 35012
rect 18512 34892 18564 34944
rect 21088 34892 21140 34944
rect 21272 34892 21324 34944
rect 22376 34892 22428 34944
rect 24032 34935 24084 34944
rect 24032 34901 24041 34935
rect 24041 34901 24075 34935
rect 24075 34901 24084 34935
rect 24032 34892 24084 34901
rect 7950 34790 8002 34842
rect 8014 34790 8066 34842
rect 8078 34790 8130 34842
rect 8142 34790 8194 34842
rect 8206 34790 8258 34842
rect 17950 34790 18002 34842
rect 18014 34790 18066 34842
rect 18078 34790 18130 34842
rect 18142 34790 18194 34842
rect 18206 34790 18258 34842
rect 7748 34688 7800 34740
rect 8392 34688 8444 34740
rect 9588 34688 9640 34740
rect 9864 34731 9916 34740
rect 9864 34697 9873 34731
rect 9873 34697 9907 34731
rect 9907 34697 9916 34731
rect 9864 34688 9916 34697
rect 11060 34688 11112 34740
rect 12716 34688 12768 34740
rect 13544 34731 13596 34740
rect 13544 34697 13553 34731
rect 13553 34697 13587 34731
rect 13587 34697 13596 34731
rect 13544 34688 13596 34697
rect 15200 34688 15252 34740
rect 15752 34688 15804 34740
rect 18788 34731 18840 34740
rect 18788 34697 18797 34731
rect 18797 34697 18831 34731
rect 18831 34697 18840 34731
rect 18788 34688 18840 34697
rect 18972 34688 19024 34740
rect 22560 34688 22612 34740
rect 8484 34620 8536 34672
rect 7380 34484 7432 34536
rect 15660 34620 15712 34672
rect 19524 34620 19576 34672
rect 21548 34620 21600 34672
rect 24400 34620 24452 34672
rect 25412 34620 25464 34672
rect 12532 34552 12584 34604
rect 13544 34552 13596 34604
rect 16856 34552 16908 34604
rect 20076 34552 20128 34604
rect 6000 34416 6052 34468
rect 6828 34416 6880 34468
rect 11060 34416 11112 34468
rect 12072 34416 12124 34468
rect 16028 34527 16080 34536
rect 16028 34493 16037 34527
rect 16037 34493 16071 34527
rect 16071 34493 16080 34527
rect 16028 34484 16080 34493
rect 15752 34416 15804 34468
rect 17868 34416 17920 34468
rect 20904 34484 20956 34536
rect 8392 34348 8444 34400
rect 15292 34348 15344 34400
rect 16396 34348 16448 34400
rect 18420 34391 18472 34400
rect 18420 34357 18429 34391
rect 18429 34357 18463 34391
rect 18463 34357 18472 34391
rect 18420 34348 18472 34357
rect 20628 34391 20680 34400
rect 20628 34357 20637 34391
rect 20637 34357 20671 34391
rect 20671 34357 20680 34391
rect 20628 34348 20680 34357
rect 21088 34348 21140 34400
rect 21640 34484 21692 34536
rect 22100 34484 22152 34536
rect 23572 34552 23624 34604
rect 25320 34595 25372 34604
rect 25320 34561 25329 34595
rect 25329 34561 25363 34595
rect 25363 34561 25372 34595
rect 25320 34552 25372 34561
rect 24676 34484 24728 34536
rect 22008 34391 22060 34400
rect 22008 34357 22017 34391
rect 22017 34357 22051 34391
rect 22051 34357 22060 34391
rect 22008 34348 22060 34357
rect 22560 34348 22612 34400
rect 23572 34348 23624 34400
rect 2950 34246 3002 34298
rect 3014 34246 3066 34298
rect 3078 34246 3130 34298
rect 3142 34246 3194 34298
rect 3206 34246 3258 34298
rect 12950 34246 13002 34298
rect 13014 34246 13066 34298
rect 13078 34246 13130 34298
rect 13142 34246 13194 34298
rect 13206 34246 13258 34298
rect 22950 34246 23002 34298
rect 23014 34246 23066 34298
rect 23078 34246 23130 34298
rect 23142 34246 23194 34298
rect 23206 34246 23258 34298
rect 7840 34187 7892 34196
rect 7840 34153 7849 34187
rect 7849 34153 7883 34187
rect 7883 34153 7892 34187
rect 7840 34144 7892 34153
rect 9772 34187 9824 34196
rect 9772 34153 9781 34187
rect 9781 34153 9815 34187
rect 9815 34153 9824 34187
rect 9772 34144 9824 34153
rect 10232 34187 10284 34196
rect 10232 34153 10241 34187
rect 10241 34153 10275 34187
rect 10275 34153 10284 34187
rect 10232 34144 10284 34153
rect 8300 34076 8352 34128
rect 5816 34051 5868 34060
rect 5816 34017 5825 34051
rect 5825 34017 5859 34051
rect 5859 34017 5868 34051
rect 5816 34008 5868 34017
rect 7104 34008 7156 34060
rect 10692 34051 10744 34060
rect 10692 34017 10701 34051
rect 10701 34017 10735 34051
rect 10735 34017 10744 34051
rect 10692 34008 10744 34017
rect 5540 33983 5592 33992
rect 5540 33949 5549 33983
rect 5549 33949 5583 33983
rect 5583 33949 5592 33983
rect 5540 33940 5592 33949
rect 6920 33940 6972 33992
rect 7748 33940 7800 33992
rect 9588 33940 9640 33992
rect 16304 34144 16356 34196
rect 16396 34144 16448 34196
rect 14280 34076 14332 34128
rect 14832 34076 14884 34128
rect 18512 34144 18564 34196
rect 20996 34076 21048 34128
rect 21548 34144 21600 34196
rect 21916 34144 21968 34196
rect 23848 34144 23900 34196
rect 25320 34187 25372 34196
rect 25320 34153 25329 34187
rect 25329 34153 25363 34187
rect 25363 34153 25372 34187
rect 25320 34144 25372 34153
rect 25412 34187 25464 34196
rect 25412 34153 25421 34187
rect 25421 34153 25455 34187
rect 25455 34153 25464 34187
rect 25412 34144 25464 34153
rect 22652 34076 22704 34128
rect 11704 34008 11756 34060
rect 16580 34008 16632 34060
rect 18696 34008 18748 34060
rect 13452 33983 13504 33992
rect 13452 33949 13461 33983
rect 13461 33949 13495 33983
rect 13495 33949 13504 33983
rect 13452 33940 13504 33949
rect 13728 33940 13780 33992
rect 21272 34008 21324 34060
rect 22928 34008 22980 34060
rect 24032 34008 24084 34060
rect 20720 33940 20772 33992
rect 8576 33872 8628 33924
rect 7472 33804 7524 33856
rect 10508 33804 10560 33856
rect 15936 33915 15988 33924
rect 15936 33881 15945 33915
rect 15945 33881 15979 33915
rect 15979 33881 15988 33915
rect 15936 33872 15988 33881
rect 16580 33872 16632 33924
rect 20536 33872 20588 33924
rect 24768 33983 24820 33992
rect 24768 33949 24777 33983
rect 24777 33949 24811 33983
rect 24811 33949 24820 33983
rect 24768 33940 24820 33949
rect 12440 33804 12492 33856
rect 14280 33804 14332 33856
rect 20168 33804 20220 33856
rect 20444 33847 20496 33856
rect 20444 33813 20453 33847
rect 20453 33813 20487 33847
rect 20487 33813 20496 33847
rect 20444 33804 20496 33813
rect 22100 33804 22152 33856
rect 23940 33804 23992 33856
rect 24584 33847 24636 33856
rect 24584 33813 24593 33847
rect 24593 33813 24627 33847
rect 24627 33813 24636 33847
rect 24584 33804 24636 33813
rect 7950 33702 8002 33754
rect 8014 33702 8066 33754
rect 8078 33702 8130 33754
rect 8142 33702 8194 33754
rect 8206 33702 8258 33754
rect 17950 33702 18002 33754
rect 18014 33702 18066 33754
rect 18078 33702 18130 33754
rect 18142 33702 18194 33754
rect 18206 33702 18258 33754
rect 7748 33600 7800 33652
rect 8852 33600 8904 33652
rect 10968 33600 11020 33652
rect 12624 33600 12676 33652
rect 13452 33532 13504 33584
rect 1308 33464 1360 33516
rect 7656 33464 7708 33516
rect 12532 33464 12584 33516
rect 13728 33464 13780 33516
rect 5540 33396 5592 33448
rect 9772 33439 9824 33448
rect 9772 33405 9781 33439
rect 9781 33405 9815 33439
rect 9815 33405 9824 33439
rect 9772 33396 9824 33405
rect 13360 33439 13412 33448
rect 13360 33405 13369 33439
rect 13369 33405 13403 33439
rect 13403 33405 13412 33439
rect 13360 33396 13412 33405
rect 13452 33396 13504 33448
rect 13636 33396 13688 33448
rect 16120 33396 16172 33448
rect 20444 33600 20496 33652
rect 20536 33643 20588 33652
rect 20536 33609 20545 33643
rect 20545 33609 20579 33643
rect 20579 33609 20588 33643
rect 20536 33600 20588 33609
rect 20904 33643 20956 33652
rect 20904 33609 20913 33643
rect 20913 33609 20947 33643
rect 20947 33609 20956 33643
rect 20904 33600 20956 33609
rect 22376 33643 22428 33652
rect 22376 33609 22385 33643
rect 22385 33609 22419 33643
rect 22419 33609 22428 33643
rect 22376 33600 22428 33609
rect 25044 33600 25096 33652
rect 18696 33532 18748 33584
rect 20168 33532 20220 33584
rect 21456 33532 21508 33584
rect 23480 33532 23532 33584
rect 18328 33507 18380 33516
rect 18328 33473 18337 33507
rect 18337 33473 18371 33507
rect 18371 33473 18380 33507
rect 18328 33464 18380 33473
rect 21272 33464 21324 33516
rect 19800 33396 19852 33448
rect 20076 33439 20128 33448
rect 20076 33405 20085 33439
rect 20085 33405 20119 33439
rect 20119 33405 20128 33439
rect 20076 33396 20128 33405
rect 22192 33396 22244 33448
rect 20168 33328 20220 33380
rect 20996 33328 21048 33380
rect 24860 33464 24912 33516
rect 23388 33396 23440 33448
rect 23756 33439 23808 33448
rect 23756 33405 23765 33439
rect 23765 33405 23799 33439
rect 23799 33405 23808 33439
rect 23756 33396 23808 33405
rect 3424 33260 3476 33312
rect 7840 33260 7892 33312
rect 12532 33303 12584 33312
rect 12532 33269 12541 33303
rect 12541 33269 12575 33303
rect 12575 33269 12584 33303
rect 12532 33260 12584 33269
rect 13636 33260 13688 33312
rect 15752 33303 15804 33312
rect 15752 33269 15761 33303
rect 15761 33269 15795 33303
rect 15795 33269 15804 33303
rect 15752 33260 15804 33269
rect 16028 33303 16080 33312
rect 16028 33269 16037 33303
rect 16037 33269 16071 33303
rect 16071 33269 16080 33303
rect 16028 33260 16080 33269
rect 16580 33260 16632 33312
rect 21640 33260 21692 33312
rect 2950 33158 3002 33210
rect 3014 33158 3066 33210
rect 3078 33158 3130 33210
rect 3142 33158 3194 33210
rect 3206 33158 3258 33210
rect 12950 33158 13002 33210
rect 13014 33158 13066 33210
rect 13078 33158 13130 33210
rect 13142 33158 13194 33210
rect 13206 33158 13258 33210
rect 22950 33158 23002 33210
rect 23014 33158 23066 33210
rect 23078 33158 23130 33210
rect 23142 33158 23194 33210
rect 23206 33158 23258 33210
rect 7564 33099 7616 33108
rect 7564 33065 7573 33099
rect 7573 33065 7607 33099
rect 7607 33065 7616 33099
rect 7564 33056 7616 33065
rect 9404 33099 9456 33108
rect 9404 33065 9413 33099
rect 9413 33065 9447 33099
rect 9447 33065 9456 33099
rect 9404 33056 9456 33065
rect 10876 33099 10928 33108
rect 10876 33065 10885 33099
rect 10885 33065 10919 33099
rect 10919 33065 10928 33099
rect 10876 33056 10928 33065
rect 11888 33099 11940 33108
rect 11888 33065 11897 33099
rect 11897 33065 11931 33099
rect 11931 33065 11940 33099
rect 11888 33056 11940 33065
rect 15936 33056 15988 33108
rect 16580 33099 16632 33108
rect 16580 33065 16589 33099
rect 16589 33065 16623 33099
rect 16623 33065 16632 33099
rect 16580 33056 16632 33065
rect 17040 33056 17092 33108
rect 17684 33099 17736 33108
rect 17684 33065 17693 33099
rect 17693 33065 17727 33099
rect 17727 33065 17736 33099
rect 17684 33056 17736 33065
rect 22468 33056 22520 33108
rect 22652 33056 22704 33108
rect 7656 32988 7708 33040
rect 8484 32988 8536 33040
rect 9956 32988 10008 33040
rect 5632 32920 5684 32972
rect 6276 32920 6328 32972
rect 6920 32920 6972 32972
rect 8300 32920 8352 32972
rect 8392 32920 8444 32972
rect 11336 32963 11388 32972
rect 9772 32895 9824 32904
rect 9772 32861 9781 32895
rect 9781 32861 9815 32895
rect 9815 32861 9824 32895
rect 9772 32852 9824 32861
rect 11336 32929 11345 32963
rect 11345 32929 11379 32963
rect 11379 32929 11388 32963
rect 11336 32920 11388 32929
rect 18696 32988 18748 33040
rect 14464 32920 14516 32972
rect 14832 32963 14884 32972
rect 14832 32929 14841 32963
rect 14841 32929 14875 32963
rect 14875 32929 14884 32963
rect 14832 32920 14884 32929
rect 17040 32963 17092 32972
rect 17040 32929 17049 32963
rect 17049 32929 17083 32963
rect 17083 32929 17092 32963
rect 17040 32920 17092 32929
rect 17224 32963 17276 32972
rect 17224 32929 17233 32963
rect 17233 32929 17267 32963
rect 17267 32929 17276 32963
rect 17224 32920 17276 32929
rect 17408 32920 17460 32972
rect 22836 32988 22888 33040
rect 23020 33031 23072 33040
rect 23020 32997 23029 33031
rect 23029 32997 23063 33031
rect 23063 32997 23072 33031
rect 23020 32988 23072 32997
rect 23664 33031 23716 33040
rect 23664 32997 23673 33031
rect 23673 32997 23707 33031
rect 23707 32997 23716 33031
rect 23664 32988 23716 32997
rect 20720 32920 20772 32972
rect 22652 32920 22704 32972
rect 11980 32852 12032 32904
rect 14372 32852 14424 32904
rect 16304 32852 16356 32904
rect 7748 32784 7800 32836
rect 8576 32784 8628 32836
rect 12256 32784 12308 32836
rect 16672 32784 16724 32836
rect 21456 32852 21508 32904
rect 21732 32852 21784 32904
rect 21916 32852 21968 32904
rect 25320 32895 25372 32904
rect 25320 32861 25329 32895
rect 25329 32861 25363 32895
rect 25363 32861 25372 32895
rect 25320 32852 25372 32861
rect 7656 32716 7708 32768
rect 9772 32716 9824 32768
rect 10968 32716 11020 32768
rect 11336 32716 11388 32768
rect 14280 32716 14332 32768
rect 14648 32759 14700 32768
rect 14648 32725 14657 32759
rect 14657 32725 14691 32759
rect 14691 32725 14700 32759
rect 14648 32716 14700 32725
rect 14740 32716 14792 32768
rect 16948 32759 17000 32768
rect 16948 32725 16957 32759
rect 16957 32725 16991 32759
rect 16991 32725 17000 32759
rect 16948 32716 17000 32725
rect 20904 32716 20956 32768
rect 21364 32784 21416 32836
rect 21916 32716 21968 32768
rect 22284 32716 22336 32768
rect 22468 32759 22520 32768
rect 22468 32725 22477 32759
rect 22477 32725 22511 32759
rect 22511 32725 22520 32759
rect 22468 32716 22520 32725
rect 22652 32716 22704 32768
rect 23204 32759 23256 32768
rect 23204 32725 23213 32759
rect 23213 32725 23247 32759
rect 23247 32725 23256 32759
rect 23204 32716 23256 32725
rect 7950 32614 8002 32666
rect 8014 32614 8066 32666
rect 8078 32614 8130 32666
rect 8142 32614 8194 32666
rect 8206 32614 8258 32666
rect 17950 32614 18002 32666
rect 18014 32614 18066 32666
rect 18078 32614 18130 32666
rect 18142 32614 18194 32666
rect 18206 32614 18258 32666
rect 4528 32512 4580 32564
rect 5448 32512 5500 32564
rect 5540 32555 5592 32564
rect 5540 32521 5549 32555
rect 5549 32521 5583 32555
rect 5583 32521 5592 32555
rect 5540 32512 5592 32521
rect 7656 32512 7708 32564
rect 9680 32512 9732 32564
rect 11244 32512 11296 32564
rect 5540 32376 5592 32428
rect 6276 32376 6328 32428
rect 7840 32444 7892 32496
rect 8024 32444 8076 32496
rect 9588 32444 9640 32496
rect 9404 32376 9456 32428
rect 10232 32419 10284 32428
rect 10232 32385 10241 32419
rect 10241 32385 10275 32419
rect 10275 32385 10284 32419
rect 10232 32376 10284 32385
rect 10692 32376 10744 32428
rect 6644 32308 6696 32360
rect 6920 32308 6972 32360
rect 8024 32308 8076 32360
rect 8300 32308 8352 32360
rect 12440 32308 12492 32360
rect 10232 32240 10284 32292
rect 14188 32376 14240 32428
rect 15936 32376 15988 32428
rect 16120 32555 16172 32564
rect 16120 32521 16129 32555
rect 16129 32521 16163 32555
rect 16163 32521 16172 32555
rect 16120 32512 16172 32521
rect 17776 32555 17828 32564
rect 17776 32521 17785 32555
rect 17785 32521 17819 32555
rect 17819 32521 17828 32555
rect 17776 32512 17828 32521
rect 19432 32512 19484 32564
rect 19708 32512 19760 32564
rect 20260 32512 20312 32564
rect 16672 32444 16724 32496
rect 17040 32444 17092 32496
rect 17500 32444 17552 32496
rect 18788 32376 18840 32428
rect 19800 32444 19852 32496
rect 20352 32444 20404 32496
rect 21364 32444 21416 32496
rect 21824 32444 21876 32496
rect 23204 32444 23256 32496
rect 16580 32308 16632 32360
rect 22192 32419 22244 32428
rect 22192 32385 22201 32419
rect 22201 32385 22235 32419
rect 22235 32385 22244 32419
rect 22192 32376 22244 32385
rect 22376 32376 22428 32428
rect 25412 32376 25464 32428
rect 15016 32240 15068 32292
rect 8668 32172 8720 32224
rect 9588 32172 9640 32224
rect 9864 32172 9916 32224
rect 13268 32215 13320 32224
rect 13268 32181 13277 32215
rect 13277 32181 13311 32215
rect 13311 32181 13320 32215
rect 13268 32172 13320 32181
rect 14004 32172 14056 32224
rect 14188 32172 14240 32224
rect 14740 32172 14792 32224
rect 14832 32172 14884 32224
rect 16948 32240 17000 32292
rect 17776 32240 17828 32292
rect 16856 32172 16908 32224
rect 17684 32172 17736 32224
rect 19248 32351 19300 32360
rect 19248 32317 19257 32351
rect 19257 32317 19291 32351
rect 19291 32317 19300 32351
rect 19248 32308 19300 32317
rect 19340 32308 19392 32360
rect 20444 32351 20496 32360
rect 20444 32317 20453 32351
rect 20453 32317 20487 32351
rect 20487 32317 20496 32351
rect 20444 32308 20496 32317
rect 18512 32172 18564 32224
rect 19524 32172 19576 32224
rect 20720 32240 20772 32292
rect 20996 32215 21048 32224
rect 20996 32181 21005 32215
rect 21005 32181 21039 32215
rect 21039 32181 21048 32215
rect 20996 32172 21048 32181
rect 21824 32172 21876 32224
rect 22468 32172 22520 32224
rect 22836 32172 22888 32224
rect 2950 32070 3002 32122
rect 3014 32070 3066 32122
rect 3078 32070 3130 32122
rect 3142 32070 3194 32122
rect 3206 32070 3258 32122
rect 12950 32070 13002 32122
rect 13014 32070 13066 32122
rect 13078 32070 13130 32122
rect 13142 32070 13194 32122
rect 13206 32070 13258 32122
rect 22950 32070 23002 32122
rect 23014 32070 23066 32122
rect 23078 32070 23130 32122
rect 23142 32070 23194 32122
rect 23206 32070 23258 32122
rect 8392 31968 8444 32020
rect 8576 32011 8628 32020
rect 8576 31977 8585 32011
rect 8585 31977 8619 32011
rect 8619 31977 8628 32011
rect 8576 31968 8628 31977
rect 9956 31968 10008 32020
rect 7840 31900 7892 31952
rect 11980 31968 12032 32020
rect 14648 31968 14700 32020
rect 15936 31968 15988 32020
rect 18604 31968 18656 32020
rect 19248 31968 19300 32020
rect 20720 31968 20772 32020
rect 21272 31968 21324 32020
rect 23756 31968 23808 32020
rect 6276 31875 6328 31884
rect 6276 31841 6285 31875
rect 6285 31841 6319 31875
rect 6319 31841 6328 31875
rect 6276 31832 6328 31841
rect 8024 31832 8076 31884
rect 9404 31832 9456 31884
rect 9496 31875 9548 31884
rect 9496 31841 9505 31875
rect 9505 31841 9539 31875
rect 9539 31841 9548 31875
rect 9496 31832 9548 31841
rect 9864 31832 9916 31884
rect 11612 31671 11664 31680
rect 11612 31637 11621 31671
rect 11621 31637 11655 31671
rect 11655 31637 11664 31671
rect 11612 31628 11664 31637
rect 14096 31900 14148 31952
rect 16948 31900 17000 31952
rect 12808 31832 12860 31884
rect 13452 31832 13504 31884
rect 17684 31832 17736 31884
rect 12440 31807 12492 31816
rect 12440 31773 12449 31807
rect 12449 31773 12483 31807
rect 12483 31773 12492 31807
rect 12440 31764 12492 31773
rect 15292 31807 15344 31816
rect 15292 31773 15301 31807
rect 15301 31773 15335 31807
rect 15335 31773 15344 31807
rect 15292 31764 15344 31773
rect 15568 31739 15620 31748
rect 15568 31705 15577 31739
rect 15577 31705 15611 31739
rect 15611 31705 15620 31739
rect 15568 31696 15620 31705
rect 15660 31696 15712 31748
rect 16028 31696 16080 31748
rect 15292 31628 15344 31680
rect 16488 31628 16540 31680
rect 16580 31628 16632 31680
rect 19616 31900 19668 31952
rect 18052 31875 18104 31884
rect 18052 31841 18061 31875
rect 18061 31841 18095 31875
rect 18095 31841 18104 31875
rect 18052 31832 18104 31841
rect 18604 31832 18656 31884
rect 19432 31832 19484 31884
rect 21548 31900 21600 31952
rect 23296 31900 23348 31952
rect 23480 31900 23532 31952
rect 20352 31875 20404 31884
rect 20352 31841 20361 31875
rect 20361 31841 20395 31875
rect 20395 31841 20404 31875
rect 20352 31832 20404 31841
rect 20904 31832 20956 31884
rect 23664 31832 23716 31884
rect 20168 31807 20220 31816
rect 20168 31773 20177 31807
rect 20177 31773 20211 31807
rect 20211 31773 20220 31807
rect 20168 31764 20220 31773
rect 22652 31764 22704 31816
rect 25320 31807 25372 31816
rect 25320 31773 25329 31807
rect 25329 31773 25363 31807
rect 25363 31773 25372 31807
rect 25320 31764 25372 31773
rect 20996 31696 21048 31748
rect 21272 31696 21324 31748
rect 22284 31696 22336 31748
rect 18328 31628 18380 31680
rect 20260 31628 20312 31680
rect 20444 31628 20496 31680
rect 7950 31526 8002 31578
rect 8014 31526 8066 31578
rect 8078 31526 8130 31578
rect 8142 31526 8194 31578
rect 8206 31526 8258 31578
rect 17950 31526 18002 31578
rect 18014 31526 18066 31578
rect 18078 31526 18130 31578
rect 18142 31526 18194 31578
rect 18206 31526 18258 31578
rect 7472 31424 7524 31476
rect 11060 31356 11112 31408
rect 11612 31356 11664 31408
rect 12808 31356 12860 31408
rect 13636 31424 13688 31476
rect 15568 31424 15620 31476
rect 16396 31424 16448 31476
rect 19800 31424 19852 31476
rect 19984 31467 20036 31476
rect 19984 31433 19993 31467
rect 19993 31433 20027 31467
rect 20027 31433 20036 31467
rect 19984 31424 20036 31433
rect 20168 31424 20220 31476
rect 22192 31424 22244 31476
rect 22560 31424 22612 31476
rect 23848 31424 23900 31476
rect 19708 31356 19760 31408
rect 21640 31356 21692 31408
rect 22100 31356 22152 31408
rect 3608 31331 3660 31340
rect 3608 31297 3617 31331
rect 3617 31297 3651 31331
rect 3651 31297 3660 31331
rect 3608 31288 3660 31297
rect 9404 31331 9456 31340
rect 9404 31297 9413 31331
rect 9413 31297 9447 31331
rect 9447 31297 9456 31331
rect 9404 31288 9456 31297
rect 3792 31263 3844 31272
rect 3792 31229 3801 31263
rect 3801 31229 3835 31263
rect 3835 31229 3844 31263
rect 3792 31220 3844 31229
rect 4988 31263 5040 31272
rect 4988 31229 4997 31263
rect 4997 31229 5031 31263
rect 5031 31229 5040 31263
rect 4988 31220 5040 31229
rect 6736 31220 6788 31272
rect 7564 31220 7616 31272
rect 7932 31263 7984 31272
rect 7932 31229 7941 31263
rect 7941 31229 7975 31263
rect 7975 31229 7984 31263
rect 7932 31220 7984 31229
rect 10968 31220 11020 31272
rect 12624 31263 12676 31272
rect 12624 31229 12633 31263
rect 12633 31229 12667 31263
rect 12667 31229 12676 31263
rect 12624 31220 12676 31229
rect 7196 31152 7248 31204
rect 12440 31152 12492 31204
rect 11612 31127 11664 31136
rect 11612 31093 11621 31127
rect 11621 31093 11655 31127
rect 11655 31093 11664 31127
rect 17132 31288 17184 31340
rect 20444 31288 20496 31340
rect 23848 31288 23900 31340
rect 24492 31331 24544 31340
rect 24492 31297 24501 31331
rect 24501 31297 24535 31331
rect 24535 31297 24544 31331
rect 24492 31288 24544 31297
rect 25320 31331 25372 31340
rect 25320 31297 25329 31331
rect 25329 31297 25363 31331
rect 25363 31297 25372 31331
rect 25320 31288 25372 31297
rect 15568 31220 15620 31272
rect 16304 31220 16356 31272
rect 17040 31220 17092 31272
rect 14924 31152 14976 31204
rect 11612 31084 11664 31093
rect 14096 31084 14148 31136
rect 14372 31127 14424 31136
rect 14372 31093 14381 31127
rect 14381 31093 14415 31127
rect 14415 31093 14424 31127
rect 14372 31084 14424 31093
rect 15016 31084 15068 31136
rect 20076 31263 20128 31272
rect 20076 31229 20085 31263
rect 20085 31229 20119 31263
rect 20119 31229 20128 31263
rect 20076 31220 20128 31229
rect 19524 31127 19576 31136
rect 19524 31093 19533 31127
rect 19533 31093 19567 31127
rect 19567 31093 19576 31127
rect 19524 31084 19576 31093
rect 23388 31084 23440 31136
rect 23664 31084 23716 31136
rect 24308 31127 24360 31136
rect 24308 31093 24317 31127
rect 24317 31093 24351 31127
rect 24351 31093 24360 31127
rect 24308 31084 24360 31093
rect 24952 31084 25004 31136
rect 2950 30982 3002 31034
rect 3014 30982 3066 31034
rect 3078 30982 3130 31034
rect 3142 30982 3194 31034
rect 3206 30982 3258 31034
rect 12950 30982 13002 31034
rect 13014 30982 13066 31034
rect 13078 30982 13130 31034
rect 13142 30982 13194 31034
rect 13206 30982 13258 31034
rect 22950 30982 23002 31034
rect 23014 30982 23066 31034
rect 23078 30982 23130 31034
rect 23142 30982 23194 31034
rect 23206 30982 23258 31034
rect 7288 30880 7340 30932
rect 8668 30880 8720 30932
rect 10508 30880 10560 30932
rect 10876 30812 10928 30864
rect 11980 30787 12032 30796
rect 11980 30753 11989 30787
rect 11989 30753 12023 30787
rect 12023 30753 12032 30787
rect 11980 30744 12032 30753
rect 7932 30676 7984 30728
rect 8300 30608 8352 30660
rect 12440 30676 12492 30728
rect 12992 30676 13044 30728
rect 14004 30676 14056 30728
rect 14280 30676 14332 30728
rect 15752 30880 15804 30932
rect 15936 30880 15988 30932
rect 19800 30880 19852 30932
rect 22744 30880 22796 30932
rect 25320 30880 25372 30932
rect 16488 30744 16540 30796
rect 20720 30812 20772 30864
rect 22192 30812 22244 30864
rect 17776 30744 17828 30796
rect 20168 30744 20220 30796
rect 22744 30744 22796 30796
rect 19708 30676 19760 30728
rect 25136 30744 25188 30796
rect 23940 30719 23992 30728
rect 23940 30685 23949 30719
rect 23949 30685 23983 30719
rect 23983 30685 23992 30719
rect 23940 30676 23992 30685
rect 25504 30676 25556 30728
rect 5264 30540 5316 30592
rect 7472 30583 7524 30592
rect 7472 30549 7481 30583
rect 7481 30549 7515 30583
rect 7515 30549 7524 30583
rect 7472 30540 7524 30549
rect 9956 30540 10008 30592
rect 11980 30540 12032 30592
rect 16212 30608 16264 30660
rect 17408 30651 17460 30660
rect 17408 30617 17417 30651
rect 17417 30617 17451 30651
rect 17451 30617 17460 30651
rect 17408 30608 17460 30617
rect 14004 30540 14056 30592
rect 15384 30583 15436 30592
rect 15384 30549 15393 30583
rect 15393 30549 15427 30583
rect 15427 30549 15436 30583
rect 15384 30540 15436 30549
rect 15568 30540 15620 30592
rect 18328 30540 18380 30592
rect 18788 30608 18840 30660
rect 20168 30608 20220 30660
rect 19892 30583 19944 30592
rect 19892 30549 19901 30583
rect 19901 30549 19935 30583
rect 19935 30549 19944 30583
rect 19892 30540 19944 30549
rect 24492 30540 24544 30592
rect 25136 30583 25188 30592
rect 25136 30549 25145 30583
rect 25145 30549 25179 30583
rect 25179 30549 25188 30583
rect 25136 30540 25188 30549
rect 7950 30438 8002 30490
rect 8014 30438 8066 30490
rect 8078 30438 8130 30490
rect 8142 30438 8194 30490
rect 8206 30438 8258 30490
rect 17950 30438 18002 30490
rect 18014 30438 18066 30490
rect 18078 30438 18130 30490
rect 18142 30438 18194 30490
rect 18206 30438 18258 30490
rect 15660 30336 15712 30388
rect 10876 30268 10928 30320
rect 12624 30268 12676 30320
rect 13728 30268 13780 30320
rect 18328 30336 18380 30388
rect 18696 30336 18748 30388
rect 19432 30336 19484 30388
rect 19892 30336 19944 30388
rect 21364 30336 21416 30388
rect 18788 30268 18840 30320
rect 23664 30311 23716 30320
rect 23664 30277 23673 30311
rect 23673 30277 23707 30311
rect 23707 30277 23716 30311
rect 23664 30268 23716 30277
rect 23940 30268 23992 30320
rect 24952 30336 25004 30388
rect 10324 30132 10376 30184
rect 10968 30175 11020 30184
rect 10968 30141 10977 30175
rect 10977 30141 11011 30175
rect 11011 30141 11020 30175
rect 10968 30132 11020 30141
rect 12716 30132 12768 30184
rect 13084 30175 13136 30184
rect 13084 30141 13093 30175
rect 13093 30141 13127 30175
rect 13127 30141 13136 30175
rect 13084 30132 13136 30141
rect 15568 30132 15620 30184
rect 8300 29996 8352 30048
rect 12716 29996 12768 30048
rect 14556 29996 14608 30048
rect 19800 30243 19852 30252
rect 19800 30209 19809 30243
rect 19809 30209 19843 30243
rect 19843 30209 19852 30243
rect 19800 30200 19852 30209
rect 23388 30243 23440 30252
rect 23388 30209 23397 30243
rect 23397 30209 23431 30243
rect 23431 30209 23440 30243
rect 23388 30200 23440 30209
rect 20904 30132 20956 30184
rect 16304 30039 16356 30048
rect 16304 30005 16313 30039
rect 16313 30005 16347 30039
rect 16347 30005 16356 30039
rect 16304 29996 16356 30005
rect 18328 29996 18380 30048
rect 19800 30064 19852 30116
rect 20168 30064 20220 30116
rect 18696 29996 18748 30048
rect 25412 30132 25464 30184
rect 22652 29996 22704 30048
rect 23388 29996 23440 30048
rect 2950 29894 3002 29946
rect 3014 29894 3066 29946
rect 3078 29894 3130 29946
rect 3142 29894 3194 29946
rect 3206 29894 3258 29946
rect 12950 29894 13002 29946
rect 13014 29894 13066 29946
rect 13078 29894 13130 29946
rect 13142 29894 13194 29946
rect 13206 29894 13258 29946
rect 22950 29894 23002 29946
rect 23014 29894 23066 29946
rect 23078 29894 23130 29946
rect 23142 29894 23194 29946
rect 23206 29894 23258 29946
rect 15844 29792 15896 29844
rect 16212 29792 16264 29844
rect 23940 29792 23992 29844
rect 15568 29724 15620 29776
rect 3884 29656 3936 29708
rect 9680 29699 9732 29708
rect 9680 29665 9689 29699
rect 9689 29665 9723 29699
rect 9723 29665 9732 29699
rect 9680 29656 9732 29665
rect 9956 29699 10008 29708
rect 9956 29665 9965 29699
rect 9965 29665 9999 29699
rect 9999 29665 10008 29699
rect 9956 29656 10008 29665
rect 10508 29656 10560 29708
rect 15660 29656 15712 29708
rect 16396 29724 16448 29776
rect 19892 29724 19944 29776
rect 20076 29724 20128 29776
rect 17776 29656 17828 29708
rect 18328 29656 18380 29708
rect 20904 29656 20956 29708
rect 23296 29699 23348 29708
rect 23296 29665 23305 29699
rect 23305 29665 23339 29699
rect 23339 29665 23348 29699
rect 23296 29656 23348 29665
rect 23388 29699 23440 29708
rect 23388 29665 23397 29699
rect 23397 29665 23431 29699
rect 23431 29665 23440 29699
rect 23388 29656 23440 29665
rect 11060 29588 11112 29640
rect 3884 29520 3936 29572
rect 6184 29520 6236 29572
rect 16672 29588 16724 29640
rect 17316 29588 17368 29640
rect 17500 29588 17552 29640
rect 20628 29588 20680 29640
rect 22560 29588 22612 29640
rect 25320 29631 25372 29640
rect 25320 29597 25329 29631
rect 25329 29597 25363 29631
rect 25363 29597 25372 29631
rect 25320 29588 25372 29597
rect 20260 29520 20312 29572
rect 7288 29452 7340 29504
rect 11428 29495 11480 29504
rect 11428 29461 11437 29495
rect 11437 29461 11471 29495
rect 11471 29461 11480 29495
rect 11428 29452 11480 29461
rect 12256 29452 12308 29504
rect 15292 29452 15344 29504
rect 16764 29495 16816 29504
rect 16764 29461 16773 29495
rect 16773 29461 16807 29495
rect 16807 29461 16816 29495
rect 16764 29452 16816 29461
rect 17040 29495 17092 29504
rect 17040 29461 17049 29495
rect 17049 29461 17083 29495
rect 17083 29461 17092 29495
rect 17040 29452 17092 29461
rect 17500 29495 17552 29504
rect 17500 29461 17509 29495
rect 17509 29461 17543 29495
rect 17543 29461 17552 29495
rect 17500 29452 17552 29461
rect 19800 29452 19852 29504
rect 24768 29520 24820 29572
rect 7950 29350 8002 29402
rect 8014 29350 8066 29402
rect 8078 29350 8130 29402
rect 8142 29350 8194 29402
rect 8206 29350 8258 29402
rect 17950 29350 18002 29402
rect 18014 29350 18066 29402
rect 18078 29350 18130 29402
rect 18142 29350 18194 29402
rect 18206 29350 18258 29402
rect 3792 29248 3844 29300
rect 5080 29248 5132 29300
rect 8944 29248 8996 29300
rect 9220 29291 9272 29300
rect 9220 29257 9229 29291
rect 9229 29257 9263 29291
rect 9263 29257 9272 29291
rect 9220 29248 9272 29257
rect 9772 29291 9824 29300
rect 9772 29257 9781 29291
rect 9781 29257 9815 29291
rect 9815 29257 9824 29291
rect 9772 29248 9824 29257
rect 11060 29291 11112 29300
rect 11060 29257 11069 29291
rect 11069 29257 11103 29291
rect 11103 29257 11112 29291
rect 11060 29248 11112 29257
rect 15200 29248 15252 29300
rect 16948 29248 17000 29300
rect 17316 29248 17368 29300
rect 17500 29248 17552 29300
rect 18420 29248 18472 29300
rect 20076 29248 20128 29300
rect 8576 29180 8628 29232
rect 2228 29112 2280 29164
rect 8668 29112 8720 29164
rect 9220 29112 9272 29164
rect 6460 29044 6512 29096
rect 8760 29019 8812 29028
rect 8760 28985 8769 29019
rect 8769 28985 8803 29019
rect 8803 28985 8812 29019
rect 8760 28976 8812 28985
rect 9680 28976 9732 29028
rect 10140 28976 10192 29028
rect 10692 29044 10744 29096
rect 11336 29180 11388 29232
rect 12256 29180 12308 29232
rect 15660 29180 15712 29232
rect 21824 29248 21876 29300
rect 22008 29248 22060 29300
rect 23940 29291 23992 29300
rect 23940 29257 23949 29291
rect 23949 29257 23983 29291
rect 23983 29257 23992 29291
rect 23940 29248 23992 29257
rect 25320 29291 25372 29300
rect 25320 29257 25329 29291
rect 25329 29257 25363 29291
rect 25363 29257 25372 29291
rect 25320 29248 25372 29257
rect 25504 29291 25556 29300
rect 25504 29257 25513 29291
rect 25513 29257 25547 29291
rect 25547 29257 25556 29291
rect 25504 29248 25556 29257
rect 13360 29112 13412 29164
rect 17684 29112 17736 29164
rect 17960 29112 18012 29164
rect 14096 29087 14148 29096
rect 14096 29053 14105 29087
rect 14105 29053 14139 29087
rect 14139 29053 14148 29087
rect 14096 29044 14148 29053
rect 14740 29044 14792 29096
rect 17408 29087 17460 29096
rect 17408 29053 17417 29087
rect 17417 29053 17451 29087
rect 17451 29053 17460 29087
rect 17408 29044 17460 29053
rect 17592 29044 17644 29096
rect 20720 29180 20772 29232
rect 24584 29180 24636 29232
rect 19800 29112 19852 29164
rect 20812 29155 20864 29164
rect 20812 29121 20821 29155
rect 20821 29121 20855 29155
rect 20855 29121 20864 29155
rect 20812 29112 20864 29121
rect 20260 29087 20312 29096
rect 20260 29053 20269 29087
rect 20269 29053 20303 29087
rect 20303 29053 20312 29087
rect 20260 29044 20312 29053
rect 20536 29044 20588 29096
rect 22744 29112 22796 29164
rect 24124 29155 24176 29164
rect 24124 29121 24133 29155
rect 24133 29121 24167 29155
rect 24167 29121 24176 29155
rect 24124 29112 24176 29121
rect 21272 29087 21324 29096
rect 21272 29053 21281 29087
rect 21281 29053 21315 29087
rect 21315 29053 21324 29087
rect 21272 29044 21324 29053
rect 10784 28976 10836 29028
rect 12624 28976 12676 29028
rect 15476 29019 15528 29028
rect 15476 28985 15485 29019
rect 15485 28985 15519 29019
rect 15519 28985 15528 29019
rect 15476 28976 15528 28985
rect 18420 28976 18472 29028
rect 22468 29044 22520 29096
rect 23296 29044 23348 29096
rect 21916 28976 21968 29028
rect 25044 28976 25096 29028
rect 8300 28908 8352 28960
rect 8668 28908 8720 28960
rect 10968 28908 11020 28960
rect 11612 28908 11664 28960
rect 15016 28908 15068 28960
rect 17960 28908 18012 28960
rect 2950 28806 3002 28858
rect 3014 28806 3066 28858
rect 3078 28806 3130 28858
rect 3142 28806 3194 28858
rect 3206 28806 3258 28858
rect 12950 28806 13002 28858
rect 13014 28806 13066 28858
rect 13078 28806 13130 28858
rect 13142 28806 13194 28858
rect 13206 28806 13258 28858
rect 22950 28806 23002 28858
rect 23014 28806 23066 28858
rect 23078 28806 23130 28858
rect 23142 28806 23194 28858
rect 23206 28806 23258 28858
rect 4068 28704 4120 28756
rect 7656 28704 7708 28756
rect 7748 28704 7800 28756
rect 10876 28747 10928 28756
rect 10876 28713 10885 28747
rect 10885 28713 10919 28747
rect 10919 28713 10928 28747
rect 10876 28704 10928 28713
rect 13360 28704 13412 28756
rect 17960 28747 18012 28756
rect 17960 28713 17969 28747
rect 17969 28713 18003 28747
rect 18003 28713 18012 28747
rect 17960 28704 18012 28713
rect 1584 28568 1636 28620
rect 7748 28568 7800 28620
rect 7840 28568 7892 28620
rect 13452 28636 13504 28688
rect 8760 28500 8812 28552
rect 9128 28543 9180 28552
rect 9128 28509 9137 28543
rect 9137 28509 9171 28543
rect 9171 28509 9180 28543
rect 9128 28500 9180 28509
rect 12808 28500 12860 28552
rect 17592 28636 17644 28688
rect 19156 28704 19208 28756
rect 22560 28704 22612 28756
rect 18880 28636 18932 28688
rect 13820 28568 13872 28620
rect 16304 28568 16356 28620
rect 23664 28568 23716 28620
rect 15292 28500 15344 28552
rect 16120 28500 16172 28552
rect 17040 28500 17092 28552
rect 21272 28500 21324 28552
rect 3516 28432 3568 28484
rect 5724 28432 5776 28484
rect 7288 28432 7340 28484
rect 9404 28475 9456 28484
rect 9404 28441 9413 28475
rect 9413 28441 9447 28475
rect 9447 28441 9456 28475
rect 9404 28432 9456 28441
rect 10968 28432 11020 28484
rect 12348 28432 12400 28484
rect 16488 28432 16540 28484
rect 16856 28432 16908 28484
rect 24768 28543 24820 28552
rect 24768 28509 24777 28543
rect 24777 28509 24811 28543
rect 24811 28509 24820 28543
rect 24768 28500 24820 28509
rect 25228 28432 25280 28484
rect 6828 28364 6880 28416
rect 7656 28364 7708 28416
rect 9588 28364 9640 28416
rect 11060 28364 11112 28416
rect 13728 28364 13780 28416
rect 13912 28364 13964 28416
rect 14464 28364 14516 28416
rect 16212 28407 16264 28416
rect 16212 28373 16221 28407
rect 16221 28373 16255 28407
rect 16255 28373 16264 28407
rect 16212 28364 16264 28373
rect 17316 28407 17368 28416
rect 17316 28373 17325 28407
rect 17325 28373 17359 28407
rect 17359 28373 17368 28407
rect 17316 28364 17368 28373
rect 17684 28407 17736 28416
rect 17684 28373 17693 28407
rect 17693 28373 17727 28407
rect 17727 28373 17736 28407
rect 17684 28364 17736 28373
rect 20720 28407 20772 28416
rect 20720 28373 20729 28407
rect 20729 28373 20763 28407
rect 20763 28373 20772 28407
rect 20720 28364 20772 28373
rect 21824 28364 21876 28416
rect 23756 28364 23808 28416
rect 24768 28364 24820 28416
rect 7950 28262 8002 28314
rect 8014 28262 8066 28314
rect 8078 28262 8130 28314
rect 8142 28262 8194 28314
rect 8206 28262 8258 28314
rect 17950 28262 18002 28314
rect 18014 28262 18066 28314
rect 18078 28262 18130 28314
rect 18142 28262 18194 28314
rect 18206 28262 18258 28314
rect 8576 28160 8628 28212
rect 8668 28203 8720 28212
rect 8668 28169 8677 28203
rect 8677 28169 8711 28203
rect 8711 28169 8720 28203
rect 8668 28160 8720 28169
rect 9404 28160 9456 28212
rect 13636 28160 13688 28212
rect 14740 28203 14792 28212
rect 14740 28169 14749 28203
rect 14749 28169 14783 28203
rect 14783 28169 14792 28203
rect 14740 28160 14792 28169
rect 15660 28160 15712 28212
rect 17684 28160 17736 28212
rect 6828 28135 6880 28144
rect 6828 28101 6837 28135
rect 6837 28101 6871 28135
rect 6871 28101 6880 28135
rect 6828 28092 6880 28101
rect 10968 28092 11020 28144
rect 11428 28092 11480 28144
rect 11704 28067 11756 28076
rect 11704 28033 11713 28067
rect 11713 28033 11747 28067
rect 11747 28033 11756 28067
rect 11704 28024 11756 28033
rect 2228 27999 2280 28008
rect 2228 27965 2237 27999
rect 2237 27965 2271 27999
rect 2271 27965 2280 27999
rect 2228 27956 2280 27965
rect 2780 27999 2832 28008
rect 2780 27965 2789 27999
rect 2789 27965 2823 27999
rect 2823 27965 2832 27999
rect 2780 27956 2832 27965
rect 6460 27956 6512 28008
rect 9220 27999 9272 28008
rect 9220 27965 9229 27999
rect 9229 27965 9263 27999
rect 9263 27965 9272 27999
rect 9220 27956 9272 27965
rect 10508 27956 10560 28008
rect 12808 27956 12860 28008
rect 13360 27956 13412 28008
rect 4068 27888 4120 27940
rect 5724 27820 5776 27872
rect 11612 27888 11664 27940
rect 11060 27820 11112 27872
rect 15384 28067 15436 28076
rect 15384 28033 15393 28067
rect 15393 28033 15427 28067
rect 15427 28033 15436 28067
rect 15384 28024 15436 28033
rect 21456 28160 21508 28212
rect 21640 28092 21692 28144
rect 16120 27956 16172 28008
rect 14464 27888 14516 27940
rect 17776 27888 17828 27940
rect 17960 27888 18012 27940
rect 19156 27999 19208 28008
rect 19156 27965 19165 27999
rect 19165 27965 19199 27999
rect 19199 27965 19208 27999
rect 19156 27956 19208 27965
rect 19800 27956 19852 28008
rect 20996 28024 21048 28076
rect 20904 27999 20956 28008
rect 20904 27965 20913 27999
rect 20913 27965 20947 27999
rect 20947 27965 20956 27999
rect 20904 27956 20956 27965
rect 18788 27888 18840 27940
rect 15936 27820 15988 27872
rect 16028 27863 16080 27872
rect 16028 27829 16037 27863
rect 16037 27829 16071 27863
rect 16071 27829 16080 27863
rect 16028 27820 16080 27829
rect 18328 27820 18380 27872
rect 19248 27820 19300 27872
rect 22192 28092 22244 28144
rect 22560 28092 22612 28144
rect 23756 28203 23808 28212
rect 23756 28169 23765 28203
rect 23765 28169 23799 28203
rect 23799 28169 23808 28203
rect 23756 28160 23808 28169
rect 25228 28203 25280 28212
rect 25228 28169 25237 28203
rect 25237 28169 25271 28203
rect 25271 28169 25280 28203
rect 25228 28160 25280 28169
rect 24676 28135 24728 28144
rect 24676 28101 24685 28135
rect 24685 28101 24719 28135
rect 24719 28101 24728 28135
rect 24676 28092 24728 28101
rect 22008 27999 22060 28008
rect 22008 27965 22017 27999
rect 22017 27965 22051 27999
rect 22051 27965 22060 27999
rect 22008 27956 22060 27965
rect 25136 27956 25188 28008
rect 25228 27888 25280 27940
rect 22836 27820 22888 27872
rect 23848 27820 23900 27872
rect 2950 27718 3002 27770
rect 3014 27718 3066 27770
rect 3078 27718 3130 27770
rect 3142 27718 3194 27770
rect 3206 27718 3258 27770
rect 12950 27718 13002 27770
rect 13014 27718 13066 27770
rect 13078 27718 13130 27770
rect 13142 27718 13194 27770
rect 13206 27718 13258 27770
rect 22950 27718 23002 27770
rect 23014 27718 23066 27770
rect 23078 27718 23130 27770
rect 23142 27718 23194 27770
rect 23206 27718 23258 27770
rect 7840 27616 7892 27668
rect 10968 27616 11020 27668
rect 16028 27616 16080 27668
rect 14556 27548 14608 27600
rect 8760 27480 8812 27532
rect 12072 27480 12124 27532
rect 3792 27412 3844 27464
rect 8300 27412 8352 27464
rect 14096 27480 14148 27532
rect 16396 27480 16448 27532
rect 19156 27616 19208 27668
rect 22100 27616 22152 27668
rect 17960 27548 18012 27600
rect 13820 27412 13872 27464
rect 14740 27412 14792 27464
rect 17868 27412 17920 27464
rect 18420 27412 18472 27464
rect 22192 27548 22244 27600
rect 19984 27480 20036 27532
rect 20352 27480 20404 27532
rect 21088 27523 21140 27532
rect 21088 27489 21097 27523
rect 21097 27489 21131 27523
rect 21131 27489 21140 27523
rect 21088 27480 21140 27489
rect 22652 27480 22704 27532
rect 23296 27480 23348 27532
rect 22008 27412 22060 27464
rect 3884 27344 3936 27396
rect 9128 27344 9180 27396
rect 6736 27276 6788 27328
rect 9496 27276 9548 27328
rect 12256 27276 12308 27328
rect 12440 27276 12492 27328
rect 14464 27344 14516 27396
rect 15936 27344 15988 27396
rect 13268 27276 13320 27328
rect 13544 27276 13596 27328
rect 17316 27276 17368 27328
rect 17684 27319 17736 27328
rect 17684 27285 17693 27319
rect 17693 27285 17727 27319
rect 17727 27285 17736 27319
rect 17684 27276 17736 27285
rect 19340 27344 19392 27396
rect 22652 27344 22704 27396
rect 22836 27344 22888 27396
rect 19708 27276 19760 27328
rect 20444 27276 20496 27328
rect 20628 27276 20680 27328
rect 22376 27276 22428 27328
rect 25320 27344 25372 27396
rect 7950 27174 8002 27226
rect 8014 27174 8066 27226
rect 8078 27174 8130 27226
rect 8142 27174 8194 27226
rect 8206 27174 8258 27226
rect 17950 27174 18002 27226
rect 18014 27174 18066 27226
rect 18078 27174 18130 27226
rect 18142 27174 18194 27226
rect 18206 27174 18258 27226
rect 7840 27072 7892 27124
rect 8576 27072 8628 27124
rect 8668 27115 8720 27124
rect 8668 27081 8677 27115
rect 8677 27081 8711 27115
rect 8711 27081 8720 27115
rect 8668 27072 8720 27081
rect 9128 27115 9180 27124
rect 9128 27081 9137 27115
rect 9137 27081 9171 27115
rect 9171 27081 9180 27115
rect 9128 27072 9180 27081
rect 9496 27115 9548 27124
rect 9496 27081 9505 27115
rect 9505 27081 9539 27115
rect 9539 27081 9548 27115
rect 9496 27072 9548 27081
rect 15108 27072 15160 27124
rect 15384 27072 15436 27124
rect 16304 27072 16356 27124
rect 17776 27072 17828 27124
rect 18880 27072 18932 27124
rect 20444 27115 20496 27124
rect 20444 27081 20453 27115
rect 20453 27081 20487 27115
rect 20487 27081 20496 27115
rect 20444 27072 20496 27081
rect 22652 27072 22704 27124
rect 11152 27004 11204 27056
rect 13544 27047 13596 27056
rect 13544 27013 13553 27047
rect 13553 27013 13587 27047
rect 13587 27013 13596 27047
rect 13544 27004 13596 27013
rect 17316 27004 17368 27056
rect 3424 26979 3476 26988
rect 3424 26945 3433 26979
rect 3433 26945 3467 26979
rect 3467 26945 3476 26979
rect 3424 26936 3476 26945
rect 10968 26936 11020 26988
rect 12072 26936 12124 26988
rect 12808 26936 12860 26988
rect 3608 26911 3660 26920
rect 3608 26877 3617 26911
rect 3617 26877 3651 26911
rect 3651 26877 3660 26911
rect 3608 26868 3660 26877
rect 5172 26911 5224 26920
rect 5172 26877 5181 26911
rect 5181 26877 5215 26911
rect 5215 26877 5224 26911
rect 5172 26868 5224 26877
rect 6460 26868 6512 26920
rect 8576 26868 8628 26920
rect 8852 26868 8904 26920
rect 10876 26868 10928 26920
rect 8300 26843 8352 26852
rect 8300 26809 8309 26843
rect 8309 26809 8343 26843
rect 8343 26809 8352 26843
rect 8300 26800 8352 26809
rect 10692 26800 10744 26852
rect 10048 26732 10100 26784
rect 11244 26732 11296 26784
rect 13268 26732 13320 26784
rect 14096 26732 14148 26784
rect 17224 26979 17276 26988
rect 17224 26945 17233 26979
rect 17233 26945 17267 26979
rect 17267 26945 17276 26979
rect 17224 26936 17276 26945
rect 17960 26936 18012 26988
rect 16120 26868 16172 26920
rect 17316 26911 17368 26920
rect 17316 26877 17325 26911
rect 17325 26877 17359 26911
rect 17359 26877 17368 26911
rect 17316 26868 17368 26877
rect 19800 27004 19852 27056
rect 22836 27004 22888 27056
rect 24308 27004 24360 27056
rect 19432 26979 19484 26988
rect 19432 26945 19441 26979
rect 19441 26945 19475 26979
rect 19475 26945 19484 26979
rect 19432 26936 19484 26945
rect 20904 26936 20956 26988
rect 14648 26800 14700 26852
rect 19800 26868 19852 26920
rect 22008 26911 22060 26920
rect 22008 26877 22017 26911
rect 22017 26877 22051 26911
rect 22051 26877 22060 26911
rect 22008 26868 22060 26877
rect 22284 26911 22336 26920
rect 22284 26877 22293 26911
rect 22293 26877 22327 26911
rect 22327 26877 22336 26911
rect 22284 26868 22336 26877
rect 22836 26868 22888 26920
rect 21272 26800 21324 26852
rect 15936 26732 15988 26784
rect 16120 26732 16172 26784
rect 16856 26775 16908 26784
rect 16856 26741 16865 26775
rect 16865 26741 16899 26775
rect 16899 26741 16908 26775
rect 16856 26732 16908 26741
rect 18052 26775 18104 26784
rect 18052 26741 18061 26775
rect 18061 26741 18095 26775
rect 18095 26741 18104 26775
rect 18052 26732 18104 26741
rect 20720 26732 20772 26784
rect 24952 26800 25004 26852
rect 22836 26732 22888 26784
rect 2950 26630 3002 26682
rect 3014 26630 3066 26682
rect 3078 26630 3130 26682
rect 3142 26630 3194 26682
rect 3206 26630 3258 26682
rect 12950 26630 13002 26682
rect 13014 26630 13066 26682
rect 13078 26630 13130 26682
rect 13142 26630 13194 26682
rect 13206 26630 13258 26682
rect 22950 26630 23002 26682
rect 23014 26630 23066 26682
rect 23078 26630 23130 26682
rect 23142 26630 23194 26682
rect 23206 26630 23258 26682
rect 3700 26528 3752 26580
rect 4804 26528 4856 26580
rect 6184 26528 6236 26580
rect 6828 26528 6880 26580
rect 7748 26528 7800 26580
rect 8668 26528 8720 26580
rect 10232 26528 10284 26580
rect 2228 26392 2280 26444
rect 6736 26435 6788 26444
rect 6736 26401 6745 26435
rect 6745 26401 6779 26435
rect 6779 26401 6788 26435
rect 6736 26392 6788 26401
rect 6828 26392 6880 26444
rect 14832 26528 14884 26580
rect 17224 26528 17276 26580
rect 11796 26460 11848 26512
rect 3700 26324 3752 26376
rect 6460 26367 6512 26376
rect 6460 26333 6469 26367
rect 6469 26333 6503 26367
rect 6503 26333 6512 26367
rect 6460 26324 6512 26333
rect 8668 26324 8720 26376
rect 9312 26324 9364 26376
rect 11428 26435 11480 26444
rect 11428 26401 11437 26435
rect 11437 26401 11471 26435
rect 11471 26401 11480 26435
rect 11428 26392 11480 26401
rect 12348 26435 12400 26444
rect 12348 26401 12357 26435
rect 12357 26401 12391 26435
rect 12391 26401 12400 26435
rect 12348 26392 12400 26401
rect 17960 26571 18012 26580
rect 17960 26537 17969 26571
rect 17969 26537 18003 26571
rect 18003 26537 18012 26571
rect 17960 26528 18012 26537
rect 18604 26528 18656 26580
rect 18696 26528 18748 26580
rect 20628 26528 20680 26580
rect 20812 26571 20864 26580
rect 20812 26537 20821 26571
rect 20821 26537 20855 26571
rect 20855 26537 20864 26571
rect 20812 26528 20864 26537
rect 22100 26528 22152 26580
rect 25136 26528 25188 26580
rect 13820 26392 13872 26444
rect 14096 26392 14148 26444
rect 5172 26256 5224 26308
rect 11060 26256 11112 26308
rect 12072 26256 12124 26308
rect 13360 26324 13412 26376
rect 13544 26324 13596 26376
rect 16304 26392 16356 26444
rect 16120 26367 16172 26376
rect 16120 26333 16129 26367
rect 16129 26333 16163 26367
rect 16163 26333 16172 26367
rect 16120 26324 16172 26333
rect 16672 26392 16724 26444
rect 18052 26392 18104 26444
rect 20904 26392 20956 26444
rect 21548 26460 21600 26512
rect 19156 26324 19208 26376
rect 19800 26367 19852 26376
rect 19800 26333 19809 26367
rect 19809 26333 19843 26367
rect 19843 26333 19852 26367
rect 19800 26324 19852 26333
rect 20444 26324 20496 26376
rect 20812 26324 20864 26376
rect 9772 26188 9824 26240
rect 11152 26231 11204 26240
rect 11152 26197 11161 26231
rect 11161 26197 11195 26231
rect 11195 26197 11204 26231
rect 11152 26188 11204 26197
rect 13360 26231 13412 26240
rect 13360 26197 13369 26231
rect 13369 26197 13403 26231
rect 13403 26197 13412 26231
rect 13360 26188 13412 26197
rect 15568 26256 15620 26308
rect 16672 26256 16724 26308
rect 18696 26256 18748 26308
rect 21824 26435 21876 26444
rect 21824 26401 21833 26435
rect 21833 26401 21867 26435
rect 21867 26401 21876 26435
rect 21824 26392 21876 26401
rect 22468 26392 22520 26444
rect 24032 26392 24084 26444
rect 22744 26324 22796 26376
rect 24584 26367 24636 26376
rect 24584 26333 24593 26367
rect 24593 26333 24627 26367
rect 24627 26333 24636 26367
rect 24584 26324 24636 26333
rect 22376 26256 22428 26308
rect 22560 26256 22612 26308
rect 16764 26231 16816 26240
rect 16764 26197 16773 26231
rect 16773 26197 16807 26231
rect 16807 26197 16816 26231
rect 16764 26188 16816 26197
rect 19432 26231 19484 26240
rect 19432 26197 19441 26231
rect 19441 26197 19475 26231
rect 19475 26197 19484 26231
rect 19432 26188 19484 26197
rect 19800 26188 19852 26240
rect 22468 26231 22520 26240
rect 22468 26197 22477 26231
rect 22477 26197 22511 26231
rect 22511 26197 22520 26231
rect 22468 26188 22520 26197
rect 7950 26086 8002 26138
rect 8014 26086 8066 26138
rect 8078 26086 8130 26138
rect 8142 26086 8194 26138
rect 8206 26086 8258 26138
rect 17950 26086 18002 26138
rect 18014 26086 18066 26138
rect 18078 26086 18130 26138
rect 18142 26086 18194 26138
rect 18206 26086 18258 26138
rect 3516 25984 3568 26036
rect 8484 25984 8536 26036
rect 8668 25984 8720 26036
rect 7748 25959 7800 25968
rect 7748 25925 7757 25959
rect 7757 25925 7791 25959
rect 7791 25925 7800 25959
rect 7748 25916 7800 25925
rect 10784 25984 10836 26036
rect 11152 25984 11204 26036
rect 11796 25984 11848 26036
rect 13912 25984 13964 26036
rect 12072 25916 12124 25968
rect 16764 25984 16816 26036
rect 18328 26027 18380 26036
rect 18328 25993 18337 26027
rect 18337 25993 18371 26027
rect 18371 25993 18380 26027
rect 18328 25984 18380 25993
rect 19616 26027 19668 26036
rect 19616 25993 19625 26027
rect 19625 25993 19659 26027
rect 19659 25993 19668 26027
rect 19616 25984 19668 25993
rect 19708 26027 19760 26036
rect 19708 25993 19717 26027
rect 19717 25993 19751 26027
rect 19751 25993 19760 26027
rect 19708 25984 19760 25993
rect 22192 25984 22244 26036
rect 16304 25959 16356 25968
rect 16304 25925 16313 25959
rect 16313 25925 16347 25959
rect 16347 25925 16356 25959
rect 16304 25916 16356 25925
rect 18420 25916 18472 25968
rect 2688 25848 2740 25900
rect 3700 25848 3752 25900
rect 6552 25848 6604 25900
rect 10508 25891 10560 25900
rect 10508 25857 10517 25891
rect 10517 25857 10551 25891
rect 10551 25857 10560 25891
rect 10508 25848 10560 25857
rect 11152 25848 11204 25900
rect 11704 25848 11756 25900
rect 6828 25823 6880 25832
rect 6828 25789 6837 25823
rect 6837 25789 6871 25823
rect 6871 25789 6880 25823
rect 6828 25780 6880 25789
rect 10692 25823 10744 25832
rect 10692 25789 10701 25823
rect 10701 25789 10735 25823
rect 10735 25789 10744 25823
rect 10692 25780 10744 25789
rect 15936 25848 15988 25900
rect 16580 25848 16632 25900
rect 19156 25848 19208 25900
rect 19616 25848 19668 25900
rect 23388 25916 23440 25968
rect 24124 25891 24176 25900
rect 24124 25857 24133 25891
rect 24133 25857 24167 25891
rect 24167 25857 24176 25891
rect 24124 25848 24176 25857
rect 3792 25712 3844 25764
rect 4344 25644 4396 25696
rect 9312 25644 9364 25696
rect 10692 25644 10744 25696
rect 11152 25644 11204 25696
rect 12348 25644 12400 25696
rect 14096 25644 14148 25696
rect 18880 25780 18932 25832
rect 20628 25780 20680 25832
rect 23204 25780 23256 25832
rect 25136 25823 25188 25832
rect 25136 25789 25145 25823
rect 25145 25789 25179 25823
rect 25179 25789 25188 25823
rect 25136 25780 25188 25789
rect 17132 25712 17184 25764
rect 16396 25644 16448 25696
rect 16580 25644 16632 25696
rect 17776 25644 17828 25696
rect 19248 25687 19300 25696
rect 19248 25653 19257 25687
rect 19257 25653 19291 25687
rect 19291 25653 19300 25687
rect 19248 25644 19300 25653
rect 22376 25644 22428 25696
rect 2950 25542 3002 25594
rect 3014 25542 3066 25594
rect 3078 25542 3130 25594
rect 3142 25542 3194 25594
rect 3206 25542 3258 25594
rect 12950 25542 13002 25594
rect 13014 25542 13066 25594
rect 13078 25542 13130 25594
rect 13142 25542 13194 25594
rect 13206 25542 13258 25594
rect 22950 25542 23002 25594
rect 23014 25542 23066 25594
rect 23078 25542 23130 25594
rect 23142 25542 23194 25594
rect 23206 25542 23258 25594
rect 4068 25483 4120 25492
rect 4068 25449 4077 25483
rect 4077 25449 4111 25483
rect 4111 25449 4120 25483
rect 4068 25440 4120 25449
rect 10508 25440 10560 25492
rect 10600 25440 10652 25492
rect 10968 25483 11020 25492
rect 10968 25449 10977 25483
rect 10977 25449 11011 25483
rect 11011 25449 11020 25483
rect 10968 25440 11020 25449
rect 13360 25440 13412 25492
rect 14096 25440 14148 25492
rect 18420 25440 18472 25492
rect 22284 25440 22336 25492
rect 7840 25372 7892 25424
rect 4896 25304 4948 25356
rect 7472 25304 7524 25356
rect 9220 25347 9272 25356
rect 9220 25313 9229 25347
rect 9229 25313 9263 25347
rect 9263 25313 9272 25347
rect 9220 25304 9272 25313
rect 9864 25304 9916 25356
rect 4804 25279 4856 25288
rect 4804 25245 4813 25279
rect 4813 25245 4847 25279
rect 4847 25245 4856 25279
rect 4804 25236 4856 25245
rect 4988 25236 5040 25288
rect 6460 25168 6512 25220
rect 4252 25100 4304 25152
rect 6828 25236 6880 25288
rect 11152 25372 11204 25424
rect 12440 25372 12492 25424
rect 13268 25372 13320 25424
rect 21732 25372 21784 25424
rect 23572 25372 23624 25424
rect 12532 25304 12584 25356
rect 13544 25304 13596 25356
rect 15108 25347 15160 25356
rect 15108 25313 15117 25347
rect 15117 25313 15151 25347
rect 15151 25313 15160 25347
rect 15108 25304 15160 25313
rect 17132 25304 17184 25356
rect 17500 25304 17552 25356
rect 20720 25304 20772 25356
rect 21364 25304 21416 25356
rect 9772 25168 9824 25220
rect 13912 25236 13964 25288
rect 13544 25168 13596 25220
rect 13728 25168 13780 25220
rect 14832 25236 14884 25288
rect 15476 25236 15528 25288
rect 19708 25236 19760 25288
rect 18604 25168 18656 25220
rect 21640 25168 21692 25220
rect 24492 25236 24544 25288
rect 12072 25100 12124 25152
rect 12440 25100 12492 25152
rect 14924 25100 14976 25152
rect 16764 25143 16816 25152
rect 16764 25109 16773 25143
rect 16773 25109 16807 25143
rect 16807 25109 16816 25143
rect 16764 25100 16816 25109
rect 17408 25100 17460 25152
rect 17592 25100 17644 25152
rect 22100 25143 22152 25152
rect 22100 25109 22109 25143
rect 22109 25109 22143 25143
rect 22143 25109 22152 25143
rect 22100 25100 22152 25109
rect 23940 25143 23992 25152
rect 23940 25109 23949 25143
rect 23949 25109 23983 25143
rect 23983 25109 23992 25143
rect 23940 25100 23992 25109
rect 24676 25143 24728 25152
rect 24676 25109 24685 25143
rect 24685 25109 24719 25143
rect 24719 25109 24728 25143
rect 24676 25100 24728 25109
rect 7950 24998 8002 25050
rect 8014 24998 8066 25050
rect 8078 24998 8130 25050
rect 8142 24998 8194 25050
rect 8206 24998 8258 25050
rect 17950 24998 18002 25050
rect 18014 24998 18066 25050
rect 18078 24998 18130 25050
rect 18142 24998 18194 25050
rect 18206 24998 18258 25050
rect 7748 24896 7800 24948
rect 9956 24939 10008 24948
rect 9956 24905 9965 24939
rect 9965 24905 9999 24939
rect 9999 24905 10008 24939
rect 9956 24896 10008 24905
rect 11428 24896 11480 24948
rect 12072 24896 12124 24948
rect 12716 24896 12768 24948
rect 18328 24896 18380 24948
rect 19432 24896 19484 24948
rect 21640 24896 21692 24948
rect 23664 24896 23716 24948
rect 25136 24896 25188 24948
rect 4252 24871 4304 24880
rect 4252 24837 4261 24871
rect 4261 24837 4295 24871
rect 4295 24837 4304 24871
rect 4252 24828 4304 24837
rect 1952 24692 2004 24744
rect 2872 24735 2924 24744
rect 2872 24701 2881 24735
rect 2881 24701 2915 24735
rect 2915 24701 2924 24735
rect 2872 24692 2924 24701
rect 3976 24735 4028 24744
rect 3976 24701 3985 24735
rect 3985 24701 4019 24735
rect 4019 24701 4028 24735
rect 3976 24692 4028 24701
rect 4344 24692 4396 24744
rect 3884 24624 3936 24676
rect 7748 24760 7800 24812
rect 8668 24803 8720 24812
rect 8668 24769 8677 24803
rect 8677 24769 8711 24803
rect 8711 24769 8720 24803
rect 8668 24760 8720 24769
rect 9312 24828 9364 24880
rect 7564 24692 7616 24744
rect 8760 24735 8812 24744
rect 8760 24701 8769 24735
rect 8769 24701 8803 24735
rect 8803 24701 8812 24735
rect 8760 24692 8812 24701
rect 12440 24828 12492 24880
rect 17500 24828 17552 24880
rect 18052 24828 18104 24880
rect 23296 24871 23348 24880
rect 23296 24837 23305 24871
rect 23305 24837 23339 24871
rect 23339 24837 23348 24871
rect 23296 24828 23348 24837
rect 9404 24692 9456 24744
rect 10324 24692 10376 24744
rect 7656 24624 7708 24676
rect 1952 24556 2004 24608
rect 3792 24556 3844 24608
rect 6092 24599 6144 24608
rect 6092 24565 6101 24599
rect 6101 24565 6135 24599
rect 6135 24565 6144 24599
rect 6092 24556 6144 24565
rect 6828 24556 6880 24608
rect 13452 24735 13504 24744
rect 13452 24701 13461 24735
rect 13461 24701 13495 24735
rect 13495 24701 13504 24735
rect 13452 24692 13504 24701
rect 15384 24760 15436 24812
rect 15752 24692 15804 24744
rect 16396 24760 16448 24812
rect 17132 24760 17184 24812
rect 19892 24760 19944 24812
rect 22560 24803 22612 24812
rect 22560 24769 22569 24803
rect 22569 24769 22603 24803
rect 22603 24769 22612 24803
rect 22560 24760 22612 24769
rect 16764 24692 16816 24744
rect 17960 24692 18012 24744
rect 22100 24692 22152 24744
rect 22836 24692 22888 24744
rect 10784 24556 10836 24608
rect 15200 24556 15252 24608
rect 17224 24556 17276 24608
rect 18696 24624 18748 24676
rect 20352 24624 20404 24676
rect 17960 24556 18012 24608
rect 23756 24556 23808 24608
rect 24584 24556 24636 24608
rect 2950 24454 3002 24506
rect 3014 24454 3066 24506
rect 3078 24454 3130 24506
rect 3142 24454 3194 24506
rect 3206 24454 3258 24506
rect 12950 24454 13002 24506
rect 13014 24454 13066 24506
rect 13078 24454 13130 24506
rect 13142 24454 13194 24506
rect 13206 24454 13258 24506
rect 22950 24454 23002 24506
rect 23014 24454 23066 24506
rect 23078 24454 23130 24506
rect 23142 24454 23194 24506
rect 23206 24454 23258 24506
rect 4804 24352 4856 24404
rect 6460 24395 6512 24404
rect 6460 24361 6469 24395
rect 6469 24361 6503 24395
rect 6503 24361 6512 24395
rect 6460 24352 6512 24361
rect 7472 24352 7524 24404
rect 8576 24352 8628 24404
rect 9956 24352 10008 24404
rect 11336 24352 11388 24404
rect 12440 24352 12492 24404
rect 12992 24352 13044 24404
rect 16120 24352 16172 24404
rect 25136 24395 25188 24404
rect 25136 24361 25145 24395
rect 25145 24361 25179 24395
rect 25179 24361 25188 24395
rect 25136 24352 25188 24361
rect 6092 24327 6144 24336
rect 6092 24293 6101 24327
rect 6101 24293 6135 24327
rect 6135 24293 6144 24327
rect 6092 24284 6144 24293
rect 8484 24284 8536 24336
rect 9588 24284 9640 24336
rect 14096 24284 14148 24336
rect 23480 24284 23532 24336
rect 2228 24191 2280 24200
rect 2228 24157 2237 24191
rect 2237 24157 2271 24191
rect 2271 24157 2280 24191
rect 2228 24148 2280 24157
rect 3976 24191 4028 24200
rect 3976 24157 3985 24191
rect 3985 24157 4019 24191
rect 4019 24157 4028 24191
rect 3976 24148 4028 24157
rect 7104 24259 7156 24268
rect 7104 24225 7113 24259
rect 7113 24225 7147 24259
rect 7147 24225 7156 24259
rect 7104 24216 7156 24225
rect 8668 24216 8720 24268
rect 9956 24216 10008 24268
rect 11244 24259 11296 24268
rect 11244 24225 11253 24259
rect 11253 24225 11287 24259
rect 11287 24225 11296 24259
rect 11244 24216 11296 24225
rect 12440 24216 12492 24268
rect 16396 24216 16448 24268
rect 20352 24216 20404 24268
rect 20536 24259 20588 24268
rect 20536 24225 20545 24259
rect 20545 24225 20579 24259
rect 20579 24225 20588 24259
rect 20536 24216 20588 24225
rect 21916 24259 21968 24268
rect 21916 24225 21925 24259
rect 21925 24225 21959 24259
rect 21959 24225 21968 24259
rect 21916 24216 21968 24225
rect 23756 24216 23808 24268
rect 24860 24216 24912 24268
rect 12348 24148 12400 24200
rect 14096 24148 14148 24200
rect 14832 24148 14884 24200
rect 17868 24191 17920 24200
rect 17868 24157 17877 24191
rect 17877 24157 17911 24191
rect 17911 24157 17920 24191
rect 17868 24148 17920 24157
rect 19156 24148 19208 24200
rect 4252 24123 4304 24132
rect 4252 24089 4261 24123
rect 4261 24089 4295 24123
rect 4295 24089 4304 24123
rect 4252 24080 4304 24089
rect 9680 24080 9732 24132
rect 1860 24012 1912 24064
rect 6736 24012 6788 24064
rect 9128 24012 9180 24064
rect 12992 24123 13044 24132
rect 12992 24089 13001 24123
rect 13001 24089 13035 24123
rect 13035 24089 13044 24123
rect 12992 24080 13044 24089
rect 13360 24012 13412 24064
rect 13452 24055 13504 24064
rect 13452 24021 13461 24055
rect 13461 24021 13495 24055
rect 13495 24021 13504 24055
rect 13452 24012 13504 24021
rect 13728 24012 13780 24064
rect 16580 24080 16632 24132
rect 17868 24012 17920 24064
rect 18052 24012 18104 24064
rect 22376 24148 22428 24200
rect 19892 24080 19944 24132
rect 23572 24148 23624 24200
rect 21732 24012 21784 24064
rect 25044 24080 25096 24132
rect 22652 24012 22704 24064
rect 24400 24012 24452 24064
rect 7950 23910 8002 23962
rect 8014 23910 8066 23962
rect 8078 23910 8130 23962
rect 8142 23910 8194 23962
rect 8206 23910 8258 23962
rect 17950 23910 18002 23962
rect 18014 23910 18066 23962
rect 18078 23910 18130 23962
rect 18142 23910 18194 23962
rect 18206 23910 18258 23962
rect 3608 23808 3660 23860
rect 4252 23808 4304 23860
rect 7104 23808 7156 23860
rect 8484 23808 8536 23860
rect 9588 23808 9640 23860
rect 9680 23851 9732 23860
rect 9680 23817 9689 23851
rect 9689 23817 9723 23851
rect 9723 23817 9732 23851
rect 9680 23808 9732 23817
rect 6828 23783 6880 23792
rect 6828 23749 6837 23783
rect 6837 23749 6871 23783
rect 6871 23749 6880 23783
rect 6828 23740 6880 23749
rect 9312 23740 9364 23792
rect 13452 23808 13504 23860
rect 14004 23808 14056 23860
rect 14464 23808 14516 23860
rect 2320 23672 2372 23724
rect 5908 23672 5960 23724
rect 9588 23715 9640 23724
rect 9588 23681 9597 23715
rect 9597 23681 9631 23715
rect 9631 23681 9640 23715
rect 9588 23672 9640 23681
rect 11704 23672 11756 23724
rect 3976 23604 4028 23656
rect 6552 23647 6604 23656
rect 6552 23613 6561 23647
rect 6561 23613 6595 23647
rect 6595 23613 6604 23647
rect 6552 23604 6604 23613
rect 7196 23604 7248 23656
rect 9864 23647 9916 23656
rect 9864 23613 9873 23647
rect 9873 23613 9907 23647
rect 9907 23613 9916 23647
rect 9864 23604 9916 23613
rect 10600 23604 10652 23656
rect 11060 23604 11112 23656
rect 11980 23536 12032 23588
rect 7840 23468 7892 23520
rect 9036 23468 9088 23520
rect 9772 23468 9824 23520
rect 12164 23604 12216 23656
rect 14740 23808 14792 23860
rect 15016 23851 15068 23860
rect 15016 23817 15025 23851
rect 15025 23817 15059 23851
rect 15059 23817 15068 23851
rect 15016 23808 15068 23817
rect 15384 23851 15436 23860
rect 15384 23817 15393 23851
rect 15393 23817 15427 23851
rect 15427 23817 15436 23851
rect 15384 23808 15436 23817
rect 15752 23851 15804 23860
rect 15752 23817 15761 23851
rect 15761 23817 15795 23851
rect 15795 23817 15804 23851
rect 15752 23808 15804 23817
rect 17224 23851 17276 23860
rect 17224 23817 17233 23851
rect 17233 23817 17267 23851
rect 17267 23817 17276 23851
rect 17224 23808 17276 23817
rect 17684 23808 17736 23860
rect 19892 23808 19944 23860
rect 20260 23808 20312 23860
rect 20628 23808 20680 23860
rect 21640 23808 21692 23860
rect 24032 23808 24084 23860
rect 24584 23851 24636 23860
rect 24584 23817 24593 23851
rect 24593 23817 24627 23851
rect 24627 23817 24636 23851
rect 24584 23808 24636 23817
rect 19156 23740 19208 23792
rect 19984 23783 20036 23792
rect 19984 23749 19993 23783
rect 19993 23749 20027 23783
rect 20027 23749 20036 23783
rect 19984 23740 20036 23749
rect 22744 23740 22796 23792
rect 23664 23740 23716 23792
rect 25412 23740 25464 23792
rect 12992 23672 13044 23724
rect 17316 23672 17368 23724
rect 18328 23672 18380 23724
rect 18604 23672 18656 23724
rect 18788 23672 18840 23724
rect 22100 23672 22152 23724
rect 22836 23715 22888 23724
rect 22836 23681 22845 23715
rect 22845 23681 22879 23715
rect 22879 23681 22888 23715
rect 22836 23672 22888 23681
rect 13728 23536 13780 23588
rect 16120 23604 16172 23656
rect 17868 23604 17920 23656
rect 17500 23536 17552 23588
rect 12164 23511 12216 23520
rect 12164 23477 12173 23511
rect 12173 23477 12207 23511
rect 12207 23477 12216 23511
rect 12164 23468 12216 23477
rect 16856 23511 16908 23520
rect 16856 23477 16865 23511
rect 16865 23477 16899 23511
rect 16899 23477 16908 23511
rect 16856 23468 16908 23477
rect 19708 23647 19760 23656
rect 19708 23613 19717 23647
rect 19717 23613 19751 23647
rect 19751 23613 19760 23647
rect 19708 23604 19760 23613
rect 20536 23604 20588 23656
rect 22744 23604 22796 23656
rect 23664 23604 23716 23656
rect 19156 23468 19208 23520
rect 20720 23468 20772 23520
rect 2950 23366 3002 23418
rect 3014 23366 3066 23418
rect 3078 23366 3130 23418
rect 3142 23366 3194 23418
rect 3206 23366 3258 23418
rect 12950 23366 13002 23418
rect 13014 23366 13066 23418
rect 13078 23366 13130 23418
rect 13142 23366 13194 23418
rect 13206 23366 13258 23418
rect 22950 23366 23002 23418
rect 23014 23366 23066 23418
rect 23078 23366 23130 23418
rect 23142 23366 23194 23418
rect 23206 23366 23258 23418
rect 2780 23264 2832 23316
rect 2780 23128 2832 23180
rect 7748 23264 7800 23316
rect 8484 23264 8536 23316
rect 11520 23264 11572 23316
rect 15844 23264 15896 23316
rect 18880 23307 18932 23316
rect 18880 23273 18889 23307
rect 18889 23273 18923 23307
rect 18923 23273 18932 23307
rect 18880 23264 18932 23273
rect 20076 23264 20128 23316
rect 11796 23196 11848 23248
rect 17040 23196 17092 23248
rect 9956 23128 10008 23180
rect 12808 23128 12860 23180
rect 14556 23128 14608 23180
rect 14832 23171 14884 23180
rect 14832 23137 14841 23171
rect 14841 23137 14875 23171
rect 14875 23137 14884 23171
rect 14832 23128 14884 23137
rect 17132 23171 17184 23180
rect 17132 23137 17141 23171
rect 17141 23137 17175 23171
rect 17175 23137 17184 23171
rect 17132 23128 17184 23137
rect 19340 23128 19392 23180
rect 19708 23128 19760 23180
rect 21088 23128 21140 23180
rect 4344 23060 4396 23112
rect 9588 23103 9640 23112
rect 9588 23069 9597 23103
rect 9597 23069 9631 23103
rect 9631 23069 9640 23103
rect 9588 23060 9640 23069
rect 2044 22992 2096 23044
rect 4436 22924 4488 22976
rect 8484 22992 8536 23044
rect 8852 22992 8904 23044
rect 10232 23035 10284 23044
rect 10232 23001 10241 23035
rect 10241 23001 10275 23035
rect 10275 23001 10284 23035
rect 10232 22992 10284 23001
rect 12348 22992 12400 23044
rect 7564 22924 7616 22976
rect 11520 22924 11572 22976
rect 11980 22924 12032 22976
rect 20812 23060 20864 23112
rect 21640 23264 21692 23316
rect 24584 23264 24636 23316
rect 23480 23196 23532 23248
rect 13820 22924 13872 22976
rect 14556 22924 14608 22976
rect 16580 22992 16632 23044
rect 17868 22992 17920 23044
rect 23848 23103 23900 23112
rect 23848 23069 23857 23103
rect 23857 23069 23891 23103
rect 23891 23069 23900 23103
rect 23848 23060 23900 23069
rect 15568 22924 15620 22976
rect 24676 22992 24728 23044
rect 20720 22924 20772 22976
rect 23572 22924 23624 22976
rect 7950 22822 8002 22874
rect 8014 22822 8066 22874
rect 8078 22822 8130 22874
rect 8142 22822 8194 22874
rect 8206 22822 8258 22874
rect 17950 22822 18002 22874
rect 18014 22822 18066 22874
rect 18078 22822 18130 22874
rect 18142 22822 18194 22874
rect 18206 22822 18258 22874
rect 2044 22720 2096 22772
rect 2688 22720 2740 22772
rect 7748 22720 7800 22772
rect 8116 22720 8168 22772
rect 9772 22720 9824 22772
rect 11796 22720 11848 22772
rect 12532 22763 12584 22772
rect 12532 22729 12541 22763
rect 12541 22729 12575 22763
rect 12575 22729 12584 22763
rect 12532 22720 12584 22729
rect 13912 22763 13964 22772
rect 13912 22729 13921 22763
rect 13921 22729 13955 22763
rect 13955 22729 13964 22763
rect 13912 22720 13964 22729
rect 15844 22720 15896 22772
rect 3700 22652 3752 22704
rect 10232 22652 10284 22704
rect 10416 22652 10468 22704
rect 11704 22695 11756 22704
rect 11704 22661 11713 22695
rect 11713 22661 11747 22695
rect 11747 22661 11756 22695
rect 11704 22652 11756 22661
rect 12256 22652 12308 22704
rect 6368 22584 6420 22636
rect 7104 22627 7156 22636
rect 7104 22593 7113 22627
rect 7113 22593 7147 22627
rect 7147 22593 7156 22627
rect 7104 22584 7156 22593
rect 7840 22584 7892 22636
rect 10692 22584 10744 22636
rect 12072 22584 12124 22636
rect 12624 22584 12676 22636
rect 14648 22627 14700 22636
rect 14648 22593 14657 22627
rect 14657 22593 14691 22627
rect 14691 22593 14700 22627
rect 14648 22584 14700 22593
rect 24124 22720 24176 22772
rect 25136 22763 25188 22772
rect 25136 22729 25145 22763
rect 25145 22729 25179 22763
rect 25179 22729 25188 22763
rect 25136 22720 25188 22729
rect 17132 22652 17184 22704
rect 18328 22652 18380 22704
rect 10968 22559 11020 22568
rect 10968 22525 10977 22559
rect 10977 22525 11011 22559
rect 11011 22525 11020 22559
rect 10968 22516 11020 22525
rect 14096 22559 14148 22568
rect 14096 22525 14105 22559
rect 14105 22525 14139 22559
rect 14139 22525 14148 22559
rect 14096 22516 14148 22525
rect 17500 22516 17552 22568
rect 18880 22584 18932 22636
rect 20536 22627 20588 22636
rect 20536 22593 20547 22627
rect 20547 22593 20581 22627
rect 20581 22593 20588 22627
rect 20536 22584 20588 22593
rect 24768 22627 24820 22636
rect 24768 22593 24777 22627
rect 24777 22593 24811 22627
rect 24811 22593 24820 22627
rect 24768 22584 24820 22593
rect 9220 22448 9272 22500
rect 11980 22448 12032 22500
rect 17592 22448 17644 22500
rect 21088 22516 21140 22568
rect 22100 22559 22152 22568
rect 22100 22525 22109 22559
rect 22109 22525 22143 22559
rect 22143 22525 22152 22559
rect 22100 22516 22152 22525
rect 24032 22516 24084 22568
rect 5816 22380 5868 22432
rect 7748 22423 7800 22432
rect 7748 22389 7757 22423
rect 7757 22389 7791 22423
rect 7791 22389 7800 22423
rect 7748 22380 7800 22389
rect 10416 22423 10468 22432
rect 10416 22389 10425 22423
rect 10425 22389 10459 22423
rect 10459 22389 10468 22423
rect 10416 22380 10468 22389
rect 12624 22380 12676 22432
rect 14556 22380 14608 22432
rect 16120 22423 16172 22432
rect 16120 22389 16129 22423
rect 16129 22389 16163 22423
rect 16163 22389 16172 22423
rect 16120 22380 16172 22389
rect 20076 22423 20128 22432
rect 20076 22389 20085 22423
rect 20085 22389 20119 22423
rect 20119 22389 20128 22423
rect 20076 22380 20128 22389
rect 2950 22278 3002 22330
rect 3014 22278 3066 22330
rect 3078 22278 3130 22330
rect 3142 22278 3194 22330
rect 3206 22278 3258 22330
rect 12950 22278 13002 22330
rect 13014 22278 13066 22330
rect 13078 22278 13130 22330
rect 13142 22278 13194 22330
rect 13206 22278 13258 22330
rect 22950 22278 23002 22330
rect 23014 22278 23066 22330
rect 23078 22278 23130 22330
rect 23142 22278 23194 22330
rect 23206 22278 23258 22330
rect 5632 22176 5684 22228
rect 3976 22040 4028 22092
rect 4160 22083 4212 22092
rect 4160 22049 4169 22083
rect 4169 22049 4203 22083
rect 4203 22049 4212 22083
rect 4160 22040 4212 22049
rect 5908 22083 5960 22092
rect 5908 22049 5917 22083
rect 5917 22049 5951 22083
rect 5951 22049 5960 22083
rect 5908 22040 5960 22049
rect 8852 22108 8904 22160
rect 14648 22176 14700 22228
rect 1952 21972 2004 22024
rect 3332 22015 3384 22024
rect 3332 21981 3341 22015
rect 3341 21981 3375 22015
rect 3375 21981 3384 22015
rect 3332 21972 3384 21981
rect 8116 22083 8168 22092
rect 8116 22049 8125 22083
rect 8125 22049 8159 22083
rect 8159 22049 8168 22083
rect 8116 22040 8168 22049
rect 9404 22040 9456 22092
rect 10692 22040 10744 22092
rect 11704 22083 11756 22092
rect 11704 22049 11713 22083
rect 11713 22049 11747 22083
rect 11747 22049 11756 22083
rect 11704 22040 11756 22049
rect 12532 22040 12584 22092
rect 13820 22108 13872 22160
rect 20812 22219 20864 22228
rect 20812 22185 20821 22219
rect 20821 22185 20855 22219
rect 20855 22185 20864 22219
rect 20812 22176 20864 22185
rect 22100 22176 22152 22228
rect 23204 22176 23256 22228
rect 25136 22219 25188 22228
rect 25136 22185 25145 22219
rect 25145 22185 25179 22219
rect 25179 22185 25188 22219
rect 25136 22176 25188 22185
rect 7656 21972 7708 22024
rect 8392 21972 8444 22024
rect 8760 21972 8812 22024
rect 12256 21972 12308 22024
rect 13912 22040 13964 22092
rect 14188 22083 14240 22092
rect 14188 22049 14197 22083
rect 14197 22049 14231 22083
rect 14231 22049 14240 22083
rect 14188 22040 14240 22049
rect 15108 22040 15160 22092
rect 16488 22083 16540 22092
rect 16488 22049 16497 22083
rect 16497 22049 16531 22083
rect 16531 22049 16540 22083
rect 16488 22040 16540 22049
rect 17776 22040 17828 22092
rect 19984 22108 20036 22160
rect 18604 22040 18656 22092
rect 19340 22040 19392 22092
rect 22744 22040 22796 22092
rect 24032 22083 24084 22092
rect 24032 22049 24041 22083
rect 24041 22049 24075 22083
rect 24075 22049 24084 22083
rect 24032 22040 24084 22049
rect 15016 21972 15068 22024
rect 1768 21836 1820 21888
rect 2136 21836 2188 21888
rect 6092 21836 6144 21888
rect 6736 21836 6788 21888
rect 8392 21836 8444 21888
rect 9588 21879 9640 21888
rect 9588 21845 9597 21879
rect 9597 21845 9631 21879
rect 9631 21845 9640 21879
rect 9588 21836 9640 21845
rect 11152 21879 11204 21888
rect 11152 21845 11161 21879
rect 11161 21845 11195 21879
rect 11195 21845 11204 21879
rect 11152 21836 11204 21845
rect 11612 21836 11664 21888
rect 16580 21972 16632 22024
rect 16764 21972 16816 22024
rect 12808 21879 12860 21888
rect 12808 21845 12817 21879
rect 12817 21845 12851 21879
rect 12851 21845 12860 21879
rect 12808 21836 12860 21845
rect 14096 21836 14148 21888
rect 15016 21836 15068 21888
rect 15660 21836 15712 21888
rect 15936 21879 15988 21888
rect 15936 21845 15945 21879
rect 15945 21845 15979 21879
rect 15979 21845 15988 21879
rect 15936 21836 15988 21845
rect 16580 21836 16632 21888
rect 16764 21836 16816 21888
rect 17500 21836 17552 21888
rect 17868 21836 17920 21888
rect 20812 21972 20864 22024
rect 21088 22015 21140 22024
rect 21088 21981 21097 22015
rect 21097 21981 21131 22015
rect 21131 21981 21140 22015
rect 21088 21972 21140 21981
rect 23388 22015 23440 22024
rect 23388 21981 23397 22015
rect 23397 21981 23431 22015
rect 23431 21981 23440 22015
rect 23388 21972 23440 21981
rect 20536 21947 20588 21956
rect 20536 21913 20545 21947
rect 20545 21913 20579 21947
rect 20579 21913 20588 21947
rect 20536 21904 20588 21913
rect 21364 21947 21416 21956
rect 21364 21913 21373 21947
rect 21373 21913 21407 21947
rect 21407 21913 21416 21947
rect 21364 21904 21416 21913
rect 21640 21904 21692 21956
rect 20904 21836 20956 21888
rect 21272 21836 21324 21888
rect 24124 21836 24176 21888
rect 7950 21734 8002 21786
rect 8014 21734 8066 21786
rect 8078 21734 8130 21786
rect 8142 21734 8194 21786
rect 8206 21734 8258 21786
rect 17950 21734 18002 21786
rect 18014 21734 18066 21786
rect 18078 21734 18130 21786
rect 18142 21734 18194 21786
rect 18206 21734 18258 21786
rect 3332 21632 3384 21684
rect 7196 21632 7248 21684
rect 2136 21564 2188 21616
rect 6276 21564 6328 21616
rect 10692 21632 10744 21684
rect 10784 21675 10836 21684
rect 10784 21641 10793 21675
rect 10793 21641 10827 21675
rect 10827 21641 10836 21675
rect 10784 21632 10836 21641
rect 7748 21564 7800 21616
rect 8852 21564 8904 21616
rect 11704 21632 11756 21684
rect 12808 21632 12860 21684
rect 10968 21564 11020 21616
rect 6920 21496 6972 21548
rect 7840 21539 7892 21548
rect 7840 21505 7849 21539
rect 7849 21505 7883 21539
rect 7883 21505 7892 21539
rect 7840 21496 7892 21505
rect 12348 21496 12400 21548
rect 12716 21564 12768 21616
rect 17500 21632 17552 21684
rect 17592 21675 17644 21684
rect 17592 21641 17601 21675
rect 17601 21641 17635 21675
rect 17635 21641 17644 21675
rect 17592 21632 17644 21641
rect 19984 21632 20036 21684
rect 17868 21564 17920 21616
rect 19156 21564 19208 21616
rect 14096 21496 14148 21548
rect 2320 21428 2372 21480
rect 2872 21471 2924 21480
rect 2872 21437 2881 21471
rect 2881 21437 2915 21471
rect 2915 21437 2924 21471
rect 2872 21428 2924 21437
rect 5908 21428 5960 21480
rect 7104 21471 7156 21480
rect 7104 21437 7113 21471
rect 7113 21437 7147 21471
rect 7147 21437 7156 21471
rect 7104 21428 7156 21437
rect 7012 21360 7064 21412
rect 9956 21428 10008 21480
rect 11612 21428 11664 21480
rect 13636 21428 13688 21480
rect 13912 21428 13964 21480
rect 14280 21428 14332 21480
rect 20720 21632 20772 21684
rect 22468 21675 22520 21684
rect 22468 21641 22477 21675
rect 22477 21641 22511 21675
rect 22511 21641 22520 21675
rect 22468 21632 22520 21641
rect 18052 21428 18104 21480
rect 18328 21471 18380 21480
rect 18328 21437 18337 21471
rect 18337 21437 18371 21471
rect 18371 21437 18380 21471
rect 18328 21428 18380 21437
rect 20076 21428 20128 21480
rect 9496 21360 9548 21412
rect 12256 21403 12308 21412
rect 12256 21369 12265 21403
rect 12265 21369 12299 21403
rect 12299 21369 12308 21403
rect 12256 21360 12308 21369
rect 13820 21360 13872 21412
rect 8484 21292 8536 21344
rect 13912 21335 13964 21344
rect 13912 21301 13921 21335
rect 13921 21301 13955 21335
rect 13955 21301 13964 21335
rect 13912 21292 13964 21301
rect 14188 21292 14240 21344
rect 15108 21292 15160 21344
rect 15660 21335 15712 21344
rect 15660 21301 15669 21335
rect 15669 21301 15703 21335
rect 15703 21301 15712 21335
rect 15660 21292 15712 21301
rect 16580 21292 16632 21344
rect 16672 21292 16724 21344
rect 17776 21292 17828 21344
rect 17868 21292 17920 21344
rect 19892 21292 19944 21344
rect 21824 21292 21876 21344
rect 23388 21632 23440 21684
rect 25136 21564 25188 21616
rect 23204 21539 23256 21548
rect 23204 21505 23213 21539
rect 23213 21505 23247 21539
rect 23247 21505 23256 21539
rect 23204 21496 23256 21505
rect 24492 21428 24544 21480
rect 23572 21292 23624 21344
rect 2950 21190 3002 21242
rect 3014 21190 3066 21242
rect 3078 21190 3130 21242
rect 3142 21190 3194 21242
rect 3206 21190 3258 21242
rect 12950 21190 13002 21242
rect 13014 21190 13066 21242
rect 13078 21190 13130 21242
rect 13142 21190 13194 21242
rect 13206 21190 13258 21242
rect 22950 21190 23002 21242
rect 23014 21190 23066 21242
rect 23078 21190 23130 21242
rect 23142 21190 23194 21242
rect 23206 21190 23258 21242
rect 5632 21088 5684 21140
rect 7564 21088 7616 21140
rect 9128 21131 9180 21140
rect 9128 21097 9137 21131
rect 9137 21097 9171 21131
rect 9171 21097 9180 21131
rect 9128 21088 9180 21097
rect 13636 21088 13688 21140
rect 15844 21088 15896 21140
rect 16028 21131 16080 21140
rect 16028 21097 16037 21131
rect 16037 21097 16071 21131
rect 16071 21097 16080 21131
rect 16028 21088 16080 21097
rect 16488 21088 16540 21140
rect 16580 21088 16632 21140
rect 19800 21088 19852 21140
rect 21640 21088 21692 21140
rect 22560 21088 22612 21140
rect 9404 21020 9456 21072
rect 19156 21020 19208 21072
rect 1308 20952 1360 21004
rect 4160 20995 4212 21004
rect 4160 20961 4169 20995
rect 4169 20961 4203 20995
rect 4203 20961 4212 20995
rect 4160 20952 4212 20961
rect 4436 20995 4488 21004
rect 4436 20961 4445 20995
rect 4445 20961 4479 20995
rect 4479 20961 4488 20995
rect 4436 20952 4488 20961
rect 8208 20952 8260 21004
rect 11796 20995 11848 21004
rect 11796 20961 11805 20995
rect 11805 20961 11839 20995
rect 11839 20961 11848 20995
rect 11796 20952 11848 20961
rect 14556 20995 14608 21004
rect 14556 20961 14565 20995
rect 14565 20961 14599 20995
rect 14599 20961 14608 20995
rect 14556 20952 14608 20961
rect 15016 20952 15068 21004
rect 15568 20952 15620 21004
rect 17776 20995 17828 21004
rect 17776 20961 17785 20995
rect 17785 20961 17819 20995
rect 17819 20961 17828 20995
rect 17776 20952 17828 20961
rect 1860 20884 1912 20936
rect 7012 20884 7064 20936
rect 9404 20884 9456 20936
rect 11244 20884 11296 20936
rect 12164 20884 12216 20936
rect 13820 20884 13872 20936
rect 16212 20884 16264 20936
rect 17684 20927 17736 20936
rect 17684 20893 17693 20927
rect 17693 20893 17727 20927
rect 17727 20893 17736 20927
rect 17684 20884 17736 20893
rect 6092 20816 6144 20868
rect 5908 20791 5960 20800
rect 5908 20757 5917 20791
rect 5917 20757 5951 20791
rect 5951 20757 5960 20791
rect 5908 20748 5960 20757
rect 10232 20791 10284 20800
rect 10232 20757 10241 20791
rect 10241 20757 10275 20791
rect 10275 20757 10284 20791
rect 10232 20748 10284 20757
rect 14004 20816 14056 20868
rect 15016 20816 15068 20868
rect 18052 20952 18104 21004
rect 18880 20952 18932 21004
rect 20812 20952 20864 21004
rect 24860 20952 24912 21004
rect 18420 20884 18472 20936
rect 21640 20884 21692 20936
rect 25228 20884 25280 20936
rect 20260 20816 20312 20868
rect 14280 20748 14332 20800
rect 15844 20748 15896 20800
rect 20444 20748 20496 20800
rect 21640 20791 21692 20800
rect 21640 20757 21649 20791
rect 21649 20757 21683 20791
rect 21683 20757 21692 20791
rect 21640 20748 21692 20757
rect 7950 20646 8002 20698
rect 8014 20646 8066 20698
rect 8078 20646 8130 20698
rect 8142 20646 8194 20698
rect 8206 20646 8258 20698
rect 17950 20646 18002 20698
rect 18014 20646 18066 20698
rect 18078 20646 18130 20698
rect 18142 20646 18194 20698
rect 18206 20646 18258 20698
rect 2780 20544 2832 20596
rect 3884 20544 3936 20596
rect 7104 20544 7156 20596
rect 8944 20544 8996 20596
rect 9312 20587 9364 20596
rect 9312 20553 9321 20587
rect 9321 20553 9355 20587
rect 9355 20553 9364 20587
rect 9312 20544 9364 20553
rect 9496 20544 9548 20596
rect 13544 20544 13596 20596
rect 13728 20544 13780 20596
rect 9404 20519 9456 20528
rect 9404 20485 9413 20519
rect 9413 20485 9447 20519
rect 9447 20485 9456 20519
rect 9404 20476 9456 20485
rect 4252 20408 4304 20460
rect 6460 20408 6512 20460
rect 9220 20408 9272 20460
rect 13820 20476 13872 20528
rect 14004 20476 14056 20528
rect 19064 20544 19116 20596
rect 19248 20544 19300 20596
rect 21364 20544 21416 20596
rect 23388 20476 23440 20528
rect 16028 20408 16080 20460
rect 9864 20340 9916 20392
rect 12256 20383 12308 20392
rect 12256 20349 12265 20383
rect 12265 20349 12299 20383
rect 12299 20349 12308 20383
rect 12256 20340 12308 20349
rect 19156 20408 19208 20460
rect 21640 20408 21692 20460
rect 22284 20451 22336 20460
rect 22284 20417 22293 20451
rect 22293 20417 22327 20451
rect 22327 20417 22336 20451
rect 22284 20408 22336 20417
rect 24952 20408 25004 20460
rect 9312 20272 9364 20324
rect 23296 20340 23348 20392
rect 6092 20247 6144 20256
rect 6092 20213 6101 20247
rect 6101 20213 6135 20247
rect 6135 20213 6144 20247
rect 6092 20204 6144 20213
rect 6736 20204 6788 20256
rect 7748 20247 7800 20256
rect 7748 20213 7757 20247
rect 7757 20213 7791 20247
rect 7791 20213 7800 20247
rect 7748 20204 7800 20213
rect 12072 20204 12124 20256
rect 22836 20272 22888 20324
rect 17868 20204 17920 20256
rect 18052 20204 18104 20256
rect 2950 20102 3002 20154
rect 3014 20102 3066 20154
rect 3078 20102 3130 20154
rect 3142 20102 3194 20154
rect 3206 20102 3258 20154
rect 12950 20102 13002 20154
rect 13014 20102 13066 20154
rect 13078 20102 13130 20154
rect 13142 20102 13194 20154
rect 13206 20102 13258 20154
rect 22950 20102 23002 20154
rect 23014 20102 23066 20154
rect 23078 20102 23130 20154
rect 23142 20102 23194 20154
rect 23206 20102 23258 20154
rect 6920 20000 6972 20052
rect 10140 20000 10192 20052
rect 10876 20000 10928 20052
rect 11244 20043 11296 20052
rect 11244 20009 11253 20043
rect 11253 20009 11287 20043
rect 11287 20009 11296 20043
rect 11244 20000 11296 20009
rect 16580 20000 16632 20052
rect 18052 20000 18104 20052
rect 18972 20043 19024 20052
rect 18972 20009 18981 20043
rect 18981 20009 19015 20043
rect 19015 20009 19024 20043
rect 18972 20000 19024 20009
rect 6736 19932 6788 19984
rect 7564 19932 7616 19984
rect 10232 19932 10284 19984
rect 14004 19932 14056 19984
rect 19064 19932 19116 19984
rect 4160 19864 4212 19916
rect 7748 19864 7800 19916
rect 6736 19796 6788 19848
rect 7012 19660 7064 19712
rect 9404 19864 9456 19916
rect 11060 19864 11112 19916
rect 11796 19907 11848 19916
rect 11796 19873 11805 19907
rect 11805 19873 11839 19907
rect 11839 19873 11848 19907
rect 11796 19864 11848 19873
rect 15200 19864 15252 19916
rect 8484 19796 8536 19848
rect 9496 19839 9548 19848
rect 9496 19805 9505 19839
rect 9505 19805 9539 19839
rect 9539 19805 9548 19839
rect 9496 19796 9548 19805
rect 10416 19796 10468 19848
rect 13728 19796 13780 19848
rect 16856 19796 16908 19848
rect 18972 19864 19024 19916
rect 24952 19864 25004 19916
rect 19524 19796 19576 19848
rect 20444 19839 20496 19848
rect 20444 19805 20453 19839
rect 20453 19805 20487 19839
rect 20487 19805 20496 19839
rect 20444 19796 20496 19805
rect 21456 19796 21508 19848
rect 25320 19796 25372 19848
rect 12808 19728 12860 19780
rect 16028 19771 16080 19780
rect 16028 19737 16037 19771
rect 16037 19737 16071 19771
rect 16071 19737 16080 19771
rect 16028 19728 16080 19737
rect 10140 19660 10192 19712
rect 10324 19660 10376 19712
rect 12164 19660 12216 19712
rect 13636 19703 13688 19712
rect 13636 19669 13645 19703
rect 13645 19669 13679 19703
rect 13679 19669 13688 19703
rect 13636 19660 13688 19669
rect 20260 19728 20312 19780
rect 22744 19728 22796 19780
rect 18512 19660 18564 19712
rect 22192 19703 22244 19712
rect 22192 19669 22201 19703
rect 22201 19669 22235 19703
rect 22235 19669 22244 19703
rect 22192 19660 22244 19669
rect 22652 19660 22704 19712
rect 24308 19660 24360 19712
rect 7950 19558 8002 19610
rect 8014 19558 8066 19610
rect 8078 19558 8130 19610
rect 8142 19558 8194 19610
rect 8206 19558 8258 19610
rect 17950 19558 18002 19610
rect 18014 19558 18066 19610
rect 18078 19558 18130 19610
rect 18142 19558 18194 19610
rect 18206 19558 18258 19610
rect 9680 19456 9732 19508
rect 10508 19456 10560 19508
rect 10876 19499 10928 19508
rect 10876 19465 10885 19499
rect 10885 19465 10919 19499
rect 10919 19465 10928 19499
rect 10876 19456 10928 19465
rect 12716 19456 12768 19508
rect 2044 19388 2096 19440
rect 8668 19388 8720 19440
rect 8852 19388 8904 19440
rect 10140 19320 10192 19372
rect 10876 19320 10928 19372
rect 12072 19363 12124 19372
rect 12072 19329 12081 19363
rect 12081 19329 12115 19363
rect 12115 19329 12124 19363
rect 12072 19320 12124 19329
rect 12348 19388 12400 19440
rect 14004 19388 14056 19440
rect 21732 19456 21784 19508
rect 22008 19456 22060 19508
rect 12624 19320 12676 19372
rect 11612 19252 11664 19304
rect 10232 19184 10284 19236
rect 13728 19295 13780 19304
rect 13728 19261 13737 19295
rect 13737 19261 13771 19295
rect 13771 19261 13780 19295
rect 13728 19252 13780 19261
rect 17132 19320 17184 19372
rect 18696 19320 18748 19372
rect 21180 19388 21232 19440
rect 22560 19388 22612 19440
rect 13452 19184 13504 19236
rect 15936 19252 15988 19304
rect 16028 19252 16080 19304
rect 16948 19252 17000 19304
rect 20628 19252 20680 19304
rect 20720 19252 20772 19304
rect 21180 19295 21232 19304
rect 21180 19261 21189 19295
rect 21189 19261 21223 19295
rect 21223 19261 21232 19295
rect 21180 19252 21232 19261
rect 21732 19252 21784 19304
rect 2228 19159 2280 19168
rect 2228 19125 2237 19159
rect 2237 19125 2271 19159
rect 2271 19125 2280 19159
rect 2228 19116 2280 19125
rect 6368 19116 6420 19168
rect 6828 19159 6880 19168
rect 6828 19125 6837 19159
rect 6837 19125 6871 19159
rect 6871 19125 6880 19159
rect 6828 19116 6880 19125
rect 8576 19116 8628 19168
rect 9864 19159 9916 19168
rect 9864 19125 9873 19159
rect 9873 19125 9907 19159
rect 9907 19125 9916 19159
rect 9864 19116 9916 19125
rect 11704 19159 11756 19168
rect 11704 19125 11713 19159
rect 11713 19125 11747 19159
rect 11747 19125 11756 19159
rect 11704 19116 11756 19125
rect 11980 19116 12032 19168
rect 13728 19116 13780 19168
rect 14004 19116 14056 19168
rect 15016 19184 15068 19236
rect 15108 19184 15160 19236
rect 14740 19159 14792 19168
rect 14740 19125 14749 19159
rect 14749 19125 14783 19159
rect 14783 19125 14792 19159
rect 14740 19116 14792 19125
rect 17500 19159 17552 19168
rect 17500 19125 17509 19159
rect 17509 19125 17543 19159
rect 17543 19125 17552 19159
rect 17500 19116 17552 19125
rect 21916 19184 21968 19236
rect 22652 19252 22704 19304
rect 23572 19252 23624 19304
rect 19248 19116 19300 19168
rect 20904 19116 20956 19168
rect 2950 19014 3002 19066
rect 3014 19014 3066 19066
rect 3078 19014 3130 19066
rect 3142 19014 3194 19066
rect 3206 19014 3258 19066
rect 12950 19014 13002 19066
rect 13014 19014 13066 19066
rect 13078 19014 13130 19066
rect 13142 19014 13194 19066
rect 13206 19014 13258 19066
rect 22950 19014 23002 19066
rect 23014 19014 23066 19066
rect 23078 19014 23130 19066
rect 23142 19014 23194 19066
rect 23206 19014 23258 19066
rect 8576 18912 8628 18964
rect 11060 18912 11112 18964
rect 12808 18912 12860 18964
rect 13544 18912 13596 18964
rect 14280 18955 14332 18964
rect 14280 18921 14289 18955
rect 14289 18921 14323 18955
rect 14323 18921 14332 18955
rect 14280 18912 14332 18921
rect 15936 18912 15988 18964
rect 2320 18844 2372 18896
rect 10692 18844 10744 18896
rect 14372 18844 14424 18896
rect 1308 18776 1360 18828
rect 5908 18776 5960 18828
rect 1768 18751 1820 18760
rect 1768 18717 1777 18751
rect 1777 18717 1811 18751
rect 1811 18717 1820 18751
rect 1768 18708 1820 18717
rect 6092 18708 6144 18760
rect 6828 18708 6880 18760
rect 8668 18776 8720 18828
rect 10968 18776 11020 18828
rect 11888 18776 11940 18828
rect 12256 18776 12308 18828
rect 13544 18776 13596 18828
rect 6736 18640 6788 18692
rect 6828 18572 6880 18624
rect 10876 18708 10928 18760
rect 11980 18708 12032 18760
rect 13728 18776 13780 18828
rect 15108 18708 15160 18760
rect 20352 18912 20404 18964
rect 21364 18912 21416 18964
rect 21916 18912 21968 18964
rect 22284 18844 22336 18896
rect 16856 18776 16908 18828
rect 21548 18819 21600 18828
rect 21548 18785 21557 18819
rect 21557 18785 21591 18819
rect 21591 18785 21600 18819
rect 21548 18776 21600 18785
rect 22008 18776 22060 18828
rect 18604 18708 18656 18760
rect 20996 18708 21048 18760
rect 21732 18708 21784 18760
rect 24584 18751 24636 18760
rect 24584 18717 24593 18751
rect 24593 18717 24627 18751
rect 24627 18717 24636 18751
rect 24584 18708 24636 18717
rect 9680 18572 9732 18624
rect 14004 18640 14056 18692
rect 10140 18572 10192 18624
rect 11244 18615 11296 18624
rect 11244 18581 11253 18615
rect 11253 18581 11287 18615
rect 11287 18581 11296 18615
rect 11244 18572 11296 18581
rect 12532 18572 12584 18624
rect 13176 18572 13228 18624
rect 16028 18640 16080 18692
rect 17408 18640 17460 18692
rect 18972 18640 19024 18692
rect 19156 18640 19208 18692
rect 23572 18640 23624 18692
rect 14740 18615 14792 18624
rect 14740 18581 14749 18615
rect 14749 18581 14783 18615
rect 14783 18581 14792 18615
rect 14740 18572 14792 18581
rect 15016 18572 15068 18624
rect 17592 18572 17644 18624
rect 19524 18572 19576 18624
rect 19984 18572 20036 18624
rect 7950 18470 8002 18522
rect 8014 18470 8066 18522
rect 8078 18470 8130 18522
rect 8142 18470 8194 18522
rect 8206 18470 8258 18522
rect 17950 18470 18002 18522
rect 18014 18470 18066 18522
rect 18078 18470 18130 18522
rect 18142 18470 18194 18522
rect 18206 18470 18258 18522
rect 4252 18368 4304 18420
rect 7104 18368 7156 18420
rect 10048 18411 10100 18420
rect 10048 18377 10057 18411
rect 10057 18377 10091 18411
rect 10091 18377 10100 18411
rect 10048 18368 10100 18377
rect 10324 18368 10376 18420
rect 13176 18411 13228 18420
rect 13176 18377 13185 18411
rect 13185 18377 13219 18411
rect 13219 18377 13228 18411
rect 13176 18368 13228 18377
rect 6828 18343 6880 18352
rect 6828 18309 6837 18343
rect 6837 18309 6871 18343
rect 6871 18309 6880 18343
rect 6828 18300 6880 18309
rect 6920 18300 6972 18352
rect 10232 18300 10284 18352
rect 12348 18343 12400 18352
rect 12348 18309 12357 18343
rect 12357 18309 12391 18343
rect 12391 18309 12400 18343
rect 12348 18300 12400 18309
rect 13544 18368 13596 18420
rect 14004 18411 14056 18420
rect 14004 18377 14013 18411
rect 14013 18377 14047 18411
rect 14047 18377 14056 18411
rect 14004 18368 14056 18377
rect 18328 18368 18380 18420
rect 20720 18368 20772 18420
rect 20536 18300 20588 18352
rect 9404 18275 9456 18284
rect 9404 18241 9413 18275
rect 9413 18241 9447 18275
rect 9447 18241 9456 18275
rect 9404 18232 9456 18241
rect 11980 18232 12032 18284
rect 23664 18232 23716 18284
rect 24400 18232 24452 18284
rect 6092 18164 6144 18216
rect 6552 18207 6604 18216
rect 6552 18173 6561 18207
rect 6561 18173 6595 18207
rect 6595 18173 6604 18207
rect 6552 18164 6604 18173
rect 7380 18164 7432 18216
rect 9036 18164 9088 18216
rect 9496 18164 9548 18216
rect 9864 18164 9916 18216
rect 13452 18207 13504 18216
rect 13452 18173 13461 18207
rect 13461 18173 13495 18207
rect 13495 18173 13504 18207
rect 13452 18164 13504 18173
rect 13820 18164 13872 18216
rect 14648 18207 14700 18216
rect 14648 18173 14657 18207
rect 14657 18173 14691 18207
rect 14691 18173 14700 18207
rect 14648 18164 14700 18173
rect 15108 18164 15160 18216
rect 11612 18096 11664 18148
rect 7472 18028 7524 18080
rect 9036 18071 9088 18080
rect 9036 18037 9045 18071
rect 9045 18037 9079 18071
rect 9079 18037 9088 18071
rect 9036 18028 9088 18037
rect 18144 18207 18196 18216
rect 18144 18173 18153 18207
rect 18153 18173 18187 18207
rect 18187 18173 18196 18207
rect 18144 18164 18196 18173
rect 21732 18164 21784 18216
rect 23388 18164 23440 18216
rect 24768 18207 24820 18216
rect 24768 18173 24777 18207
rect 24777 18173 24811 18207
rect 24811 18173 24820 18207
rect 24768 18164 24820 18173
rect 20996 18096 21048 18148
rect 18696 18028 18748 18080
rect 2950 17926 3002 17978
rect 3014 17926 3066 17978
rect 3078 17926 3130 17978
rect 3142 17926 3194 17978
rect 3206 17926 3258 17978
rect 12950 17926 13002 17978
rect 13014 17926 13066 17978
rect 13078 17926 13130 17978
rect 13142 17926 13194 17978
rect 13206 17926 13258 17978
rect 22950 17926 23002 17978
rect 23014 17926 23066 17978
rect 23078 17926 23130 17978
rect 23142 17926 23194 17978
rect 23206 17926 23258 17978
rect 5540 17824 5592 17876
rect 5816 17824 5868 17876
rect 6092 17824 6144 17876
rect 7104 17867 7156 17876
rect 7104 17833 7113 17867
rect 7113 17833 7147 17867
rect 7147 17833 7156 17867
rect 7104 17824 7156 17833
rect 7564 17731 7616 17740
rect 7564 17697 7573 17731
rect 7573 17697 7607 17731
rect 7607 17697 7616 17731
rect 7564 17688 7616 17697
rect 7748 17731 7800 17740
rect 7748 17697 7757 17731
rect 7757 17697 7791 17731
rect 7791 17697 7800 17731
rect 7748 17688 7800 17697
rect 9404 17688 9456 17740
rect 4804 17663 4856 17672
rect 4804 17629 4813 17663
rect 4813 17629 4847 17663
rect 4847 17629 4856 17663
rect 4804 17620 4856 17629
rect 9036 17620 9088 17672
rect 11520 17824 11572 17876
rect 18144 17824 18196 17876
rect 11060 17731 11112 17740
rect 11060 17697 11069 17731
rect 11069 17697 11103 17731
rect 11103 17697 11112 17731
rect 11060 17688 11112 17697
rect 13636 17688 13688 17740
rect 14924 17620 14976 17672
rect 16764 17620 16816 17672
rect 16856 17663 16908 17672
rect 16856 17629 16865 17663
rect 16865 17629 16899 17663
rect 16899 17629 16908 17663
rect 16856 17620 16908 17629
rect 20536 17824 20588 17876
rect 21456 17867 21508 17876
rect 21456 17833 21465 17867
rect 21465 17833 21499 17867
rect 21499 17833 21508 17867
rect 21456 17824 21508 17833
rect 23664 17867 23716 17876
rect 23664 17833 23673 17867
rect 23673 17833 23707 17867
rect 23707 17833 23716 17867
rect 23664 17824 23716 17833
rect 24584 17824 24636 17876
rect 19708 17731 19760 17740
rect 19708 17697 19717 17731
rect 19717 17697 19751 17731
rect 19751 17697 19760 17731
rect 19708 17688 19760 17697
rect 22192 17731 22244 17740
rect 22192 17697 22201 17731
rect 22201 17697 22235 17731
rect 22235 17697 22244 17731
rect 22192 17688 22244 17697
rect 21732 17620 21784 17672
rect 23572 17756 23624 17808
rect 5080 17595 5132 17604
rect 5080 17561 5089 17595
rect 5089 17561 5123 17595
rect 5123 17561 5132 17595
rect 5080 17552 5132 17561
rect 6920 17552 6972 17604
rect 9864 17595 9916 17604
rect 9864 17561 9873 17595
rect 9873 17561 9907 17595
rect 9907 17561 9916 17595
rect 9864 17552 9916 17561
rect 9312 17484 9364 17536
rect 10508 17527 10560 17536
rect 10508 17493 10517 17527
rect 10517 17493 10551 17527
rect 10551 17493 10560 17527
rect 10508 17484 10560 17493
rect 18696 17595 18748 17604
rect 18696 17561 18705 17595
rect 18705 17561 18739 17595
rect 18739 17561 18748 17595
rect 18696 17552 18748 17561
rect 19984 17595 20036 17604
rect 19984 17561 19993 17595
rect 19993 17561 20027 17595
rect 20027 17561 20036 17595
rect 19984 17552 20036 17561
rect 20720 17552 20772 17604
rect 13636 17484 13688 17536
rect 13820 17527 13872 17536
rect 13820 17493 13829 17527
rect 13829 17493 13863 17527
rect 13863 17493 13872 17527
rect 13820 17484 13872 17493
rect 15476 17484 15528 17536
rect 15568 17484 15620 17536
rect 7950 17382 8002 17434
rect 8014 17382 8066 17434
rect 8078 17382 8130 17434
rect 8142 17382 8194 17434
rect 8206 17382 8258 17434
rect 17950 17382 18002 17434
rect 18014 17382 18066 17434
rect 18078 17382 18130 17434
rect 18142 17382 18194 17434
rect 18206 17382 18258 17434
rect 5080 17280 5132 17332
rect 6920 17280 6972 17332
rect 7472 17323 7524 17332
rect 7472 17289 7481 17323
rect 7481 17289 7515 17323
rect 7515 17289 7524 17323
rect 7472 17280 7524 17289
rect 2320 17212 2372 17264
rect 7748 17212 7800 17264
rect 9220 17280 9272 17332
rect 10140 17280 10192 17332
rect 10508 17280 10560 17332
rect 11704 17280 11756 17332
rect 12072 17280 12124 17332
rect 15384 17280 15436 17332
rect 15660 17280 15712 17332
rect 16304 17280 16356 17332
rect 11060 17212 11112 17264
rect 11796 17212 11848 17264
rect 15752 17212 15804 17264
rect 19708 17280 19760 17332
rect 20628 17280 20680 17332
rect 5816 17008 5868 17060
rect 1768 16940 1820 16992
rect 5908 16940 5960 16992
rect 6552 16940 6604 16992
rect 7840 17008 7892 17060
rect 9128 17187 9180 17196
rect 9128 17153 9137 17187
rect 9137 17153 9171 17187
rect 9171 17153 9180 17187
rect 9128 17144 9180 17153
rect 9312 17119 9364 17128
rect 9312 17085 9321 17119
rect 9321 17085 9355 17119
rect 9355 17085 9364 17119
rect 9312 17076 9364 17085
rect 10324 17076 10376 17128
rect 10508 17008 10560 17060
rect 11520 17144 11572 17196
rect 10784 17076 10836 17128
rect 12808 17076 12860 17128
rect 14096 17144 14148 17196
rect 19616 17212 19668 17264
rect 20720 17212 20772 17264
rect 22192 17212 22244 17264
rect 22836 17212 22888 17264
rect 8484 16940 8536 16992
rect 14280 17008 14332 17060
rect 14464 17008 14516 17060
rect 13820 16940 13872 16992
rect 18236 17144 18288 17196
rect 19432 17187 19484 17196
rect 19432 17153 19441 17187
rect 19441 17153 19475 17187
rect 19475 17153 19484 17187
rect 19432 17144 19484 17153
rect 20628 17187 20680 17196
rect 20628 17153 20637 17187
rect 20637 17153 20671 17187
rect 20671 17153 20680 17187
rect 20628 17144 20680 17153
rect 22008 17187 22060 17196
rect 22008 17153 22017 17187
rect 22017 17153 22051 17187
rect 22051 17153 22060 17187
rect 22008 17144 22060 17153
rect 23940 17187 23992 17196
rect 23940 17153 23949 17187
rect 23949 17153 23983 17187
rect 23983 17153 23992 17187
rect 23940 17144 23992 17153
rect 15660 17076 15712 17128
rect 18604 17076 18656 17128
rect 21456 17076 21508 17128
rect 24676 17119 24728 17128
rect 24676 17085 24685 17119
rect 24685 17085 24719 17119
rect 24719 17085 24728 17119
rect 24676 17076 24728 17085
rect 23388 17051 23440 17060
rect 23388 17017 23397 17051
rect 23397 17017 23431 17051
rect 23431 17017 23440 17051
rect 23388 17008 23440 17017
rect 16488 16940 16540 16992
rect 16856 16940 16908 16992
rect 20444 16940 20496 16992
rect 22008 16940 22060 16992
rect 2950 16838 3002 16890
rect 3014 16838 3066 16890
rect 3078 16838 3130 16890
rect 3142 16838 3194 16890
rect 3206 16838 3258 16890
rect 12950 16838 13002 16890
rect 13014 16838 13066 16890
rect 13078 16838 13130 16890
rect 13142 16838 13194 16890
rect 13206 16838 13258 16890
rect 22950 16838 23002 16890
rect 23014 16838 23066 16890
rect 23078 16838 23130 16890
rect 23142 16838 23194 16890
rect 23206 16838 23258 16890
rect 7932 16736 7984 16788
rect 8484 16779 8536 16788
rect 8484 16745 8493 16779
rect 8493 16745 8527 16779
rect 8527 16745 8536 16779
rect 8484 16736 8536 16745
rect 11520 16736 11572 16788
rect 12808 16736 12860 16788
rect 16304 16736 16356 16788
rect 19432 16736 19484 16788
rect 23848 16736 23900 16788
rect 4804 16600 4856 16652
rect 5908 16600 5960 16652
rect 6644 16600 6696 16652
rect 9864 16668 9916 16720
rect 7748 16643 7800 16652
rect 7748 16609 7757 16643
rect 7757 16609 7791 16643
rect 7791 16609 7800 16643
rect 7748 16600 7800 16609
rect 8944 16600 8996 16652
rect 9588 16600 9640 16652
rect 9956 16600 10008 16652
rect 15200 16668 15252 16720
rect 2228 16532 2280 16584
rect 9220 16532 9272 16584
rect 10692 16575 10744 16584
rect 10692 16541 10701 16575
rect 10701 16541 10735 16575
rect 10735 16541 10744 16575
rect 10692 16532 10744 16541
rect 11520 16575 11572 16584
rect 11520 16541 11529 16575
rect 11529 16541 11563 16575
rect 11563 16541 11572 16575
rect 11520 16532 11572 16541
rect 12072 16532 12124 16584
rect 14924 16600 14976 16652
rect 18788 16668 18840 16720
rect 15200 16532 15252 16584
rect 15752 16600 15804 16652
rect 17592 16600 17644 16652
rect 16028 16532 16080 16584
rect 17776 16532 17828 16584
rect 18236 16600 18288 16652
rect 20812 16600 20864 16652
rect 20904 16600 20956 16652
rect 21732 16643 21784 16652
rect 21732 16609 21741 16643
rect 21741 16609 21775 16643
rect 21775 16609 21784 16643
rect 21732 16600 21784 16609
rect 22008 16643 22060 16652
rect 22008 16609 22017 16643
rect 22017 16609 22051 16643
rect 22051 16609 22060 16643
rect 22008 16600 22060 16609
rect 22468 16600 22520 16652
rect 18328 16532 18380 16584
rect 18604 16575 18656 16584
rect 18604 16541 18613 16575
rect 18613 16541 18647 16575
rect 18647 16541 18656 16575
rect 18604 16532 18656 16541
rect 20260 16532 20312 16584
rect 1308 16464 1360 16516
rect 6920 16396 6972 16448
rect 7932 16464 7984 16516
rect 14556 16464 14608 16516
rect 19892 16464 19944 16516
rect 21088 16507 21140 16516
rect 21088 16473 21097 16507
rect 21097 16473 21131 16507
rect 21131 16473 21140 16507
rect 21088 16464 21140 16473
rect 22652 16464 22704 16516
rect 8484 16396 8536 16448
rect 9128 16439 9180 16448
rect 9128 16405 9137 16439
rect 9137 16405 9171 16439
rect 9171 16405 9180 16439
rect 9128 16396 9180 16405
rect 9588 16439 9640 16448
rect 9588 16405 9597 16439
rect 9597 16405 9631 16439
rect 9631 16405 9640 16439
rect 9588 16396 9640 16405
rect 10324 16439 10376 16448
rect 10324 16405 10333 16439
rect 10333 16405 10367 16439
rect 10367 16405 10376 16439
rect 10324 16396 10376 16405
rect 11060 16396 11112 16448
rect 11244 16396 11296 16448
rect 13636 16396 13688 16448
rect 15108 16439 15160 16448
rect 15108 16405 15117 16439
rect 15117 16405 15151 16439
rect 15151 16405 15160 16439
rect 15108 16396 15160 16405
rect 16120 16396 16172 16448
rect 18420 16396 18472 16448
rect 19524 16396 19576 16448
rect 20536 16396 20588 16448
rect 24584 16396 24636 16448
rect 7950 16294 8002 16346
rect 8014 16294 8066 16346
rect 8078 16294 8130 16346
rect 8142 16294 8194 16346
rect 8206 16294 8258 16346
rect 17950 16294 18002 16346
rect 18014 16294 18066 16346
rect 18078 16294 18130 16346
rect 18142 16294 18194 16346
rect 18206 16294 18258 16346
rect 6368 16192 6420 16244
rect 9128 16192 9180 16244
rect 9588 16235 9640 16244
rect 9588 16201 9597 16235
rect 9597 16201 9631 16235
rect 9631 16201 9640 16235
rect 9588 16192 9640 16201
rect 11152 16192 11204 16244
rect 10324 16124 10376 16176
rect 8208 16099 8260 16108
rect 8208 16065 8217 16099
rect 8217 16065 8251 16099
rect 8251 16065 8260 16099
rect 8208 16056 8260 16065
rect 7748 15920 7800 15972
rect 11888 16192 11940 16244
rect 13544 16192 13596 16244
rect 16212 16235 16264 16244
rect 16212 16201 16221 16235
rect 16221 16201 16255 16235
rect 16255 16201 16264 16235
rect 16212 16192 16264 16201
rect 16672 16192 16724 16244
rect 18788 16235 18840 16244
rect 18788 16201 18797 16235
rect 18797 16201 18831 16235
rect 18831 16201 18840 16235
rect 18788 16192 18840 16201
rect 19156 16235 19208 16244
rect 19156 16201 19165 16235
rect 19165 16201 19199 16235
rect 19199 16201 19208 16235
rect 19156 16192 19208 16201
rect 19524 16235 19576 16244
rect 19524 16201 19533 16235
rect 19533 16201 19567 16235
rect 19567 16201 19576 16235
rect 19524 16192 19576 16201
rect 20352 16192 20404 16244
rect 22192 16192 22244 16244
rect 22468 16192 22520 16244
rect 22652 16192 22704 16244
rect 12072 16167 12124 16176
rect 12072 16133 12081 16167
rect 12081 16133 12115 16167
rect 12115 16133 12124 16167
rect 12072 16124 12124 16133
rect 13636 16056 13688 16108
rect 10876 15988 10928 16040
rect 11796 16031 11848 16040
rect 11796 15997 11805 16031
rect 11805 15997 11839 16031
rect 11839 15997 11848 16031
rect 11796 15988 11848 15997
rect 11704 15920 11756 15972
rect 8392 15852 8444 15904
rect 13544 15895 13596 15904
rect 13544 15861 13553 15895
rect 13553 15861 13587 15895
rect 13587 15861 13596 15895
rect 13544 15852 13596 15861
rect 21364 16124 21416 16176
rect 21272 16056 21324 16108
rect 24124 16099 24176 16108
rect 24124 16065 24133 16099
rect 24133 16065 24167 16099
rect 24167 16065 24176 16099
rect 24124 16056 24176 16065
rect 20996 16031 21048 16040
rect 20996 15997 21005 16031
rect 21005 15997 21039 16031
rect 21039 15997 21048 16031
rect 20996 15988 21048 15997
rect 16304 15920 16356 15972
rect 17408 15920 17460 15972
rect 20444 15920 20496 15972
rect 23664 15988 23716 16040
rect 24768 16031 24820 16040
rect 24768 15997 24777 16031
rect 24777 15997 24811 16031
rect 24811 15997 24820 16031
rect 24768 15988 24820 15997
rect 17040 15852 17092 15904
rect 17776 15852 17828 15904
rect 18236 15852 18288 15904
rect 21548 15852 21600 15904
rect 23480 15852 23532 15904
rect 2950 15750 3002 15802
rect 3014 15750 3066 15802
rect 3078 15750 3130 15802
rect 3142 15750 3194 15802
rect 3206 15750 3258 15802
rect 12950 15750 13002 15802
rect 13014 15750 13066 15802
rect 13078 15750 13130 15802
rect 13142 15750 13194 15802
rect 13206 15750 13258 15802
rect 22950 15750 23002 15802
rect 23014 15750 23066 15802
rect 23078 15750 23130 15802
rect 23142 15750 23194 15802
rect 23206 15750 23258 15802
rect 8208 15648 8260 15700
rect 10140 15648 10192 15700
rect 12164 15648 12216 15700
rect 15016 15691 15068 15700
rect 15016 15657 15025 15691
rect 15025 15657 15059 15691
rect 15059 15657 15068 15691
rect 15016 15648 15068 15657
rect 15292 15648 15344 15700
rect 14096 15623 14148 15632
rect 14096 15589 14105 15623
rect 14105 15589 14139 15623
rect 14139 15589 14148 15623
rect 14096 15580 14148 15589
rect 18328 15648 18380 15700
rect 18420 15648 18472 15700
rect 20996 15648 21048 15700
rect 8576 15512 8628 15564
rect 10876 15512 10928 15564
rect 13728 15512 13780 15564
rect 6736 15487 6788 15496
rect 6736 15453 6745 15487
rect 6745 15453 6779 15487
rect 6779 15453 6788 15487
rect 6736 15444 6788 15453
rect 9036 15444 9088 15496
rect 13636 15444 13688 15496
rect 18236 15512 18288 15564
rect 21180 15580 21232 15632
rect 18880 15512 18932 15564
rect 19892 15555 19944 15564
rect 19892 15521 19901 15555
rect 19901 15521 19935 15555
rect 19935 15521 19944 15555
rect 19892 15512 19944 15521
rect 20536 15512 20588 15564
rect 21272 15555 21324 15564
rect 21272 15521 21281 15555
rect 21281 15521 21315 15555
rect 21315 15521 21324 15555
rect 21272 15512 21324 15521
rect 15016 15444 15068 15496
rect 15200 15444 15252 15496
rect 17040 15444 17092 15496
rect 17408 15444 17460 15496
rect 20720 15444 20772 15496
rect 21640 15444 21692 15496
rect 22744 15487 22796 15496
rect 22744 15453 22753 15487
rect 22753 15453 22787 15487
rect 22787 15453 22796 15487
rect 22744 15444 22796 15453
rect 24584 15487 24636 15496
rect 24584 15453 24593 15487
rect 24593 15453 24627 15487
rect 24627 15453 24636 15487
rect 24584 15444 24636 15453
rect 7656 15308 7708 15360
rect 8484 15376 8536 15428
rect 8760 15376 8812 15428
rect 10140 15376 10192 15428
rect 10784 15376 10836 15428
rect 11244 15376 11296 15428
rect 13268 15376 13320 15428
rect 15568 15376 15620 15428
rect 15844 15376 15896 15428
rect 15936 15419 15988 15428
rect 15936 15385 15945 15419
rect 15945 15385 15979 15419
rect 15979 15385 15988 15419
rect 15936 15376 15988 15385
rect 9128 15308 9180 15360
rect 11520 15308 11572 15360
rect 12348 15308 12400 15360
rect 14648 15351 14700 15360
rect 14648 15317 14657 15351
rect 14657 15317 14691 15351
rect 14691 15317 14700 15351
rect 14648 15308 14700 15317
rect 20536 15376 20588 15428
rect 24952 15376 25004 15428
rect 18236 15308 18288 15360
rect 21088 15308 21140 15360
rect 21364 15308 21416 15360
rect 22284 15308 22336 15360
rect 7950 15206 8002 15258
rect 8014 15206 8066 15258
rect 8078 15206 8130 15258
rect 8142 15206 8194 15258
rect 8206 15206 8258 15258
rect 17950 15206 18002 15258
rect 18014 15206 18066 15258
rect 18078 15206 18130 15258
rect 18142 15206 18194 15258
rect 18206 15206 18258 15258
rect 7840 15104 7892 15156
rect 11980 15104 12032 15156
rect 13268 15104 13320 15156
rect 13728 15104 13780 15156
rect 14004 15104 14056 15156
rect 14096 15104 14148 15156
rect 15292 15147 15344 15156
rect 15292 15113 15301 15147
rect 15301 15113 15335 15147
rect 15335 15113 15344 15147
rect 15292 15104 15344 15113
rect 15936 15104 15988 15156
rect 16488 15104 16540 15156
rect 20628 15104 20680 15156
rect 21456 15147 21508 15156
rect 7656 15036 7708 15088
rect 8392 15079 8444 15088
rect 8392 15045 8401 15079
rect 8401 15045 8435 15079
rect 8435 15045 8444 15079
rect 8392 15036 8444 15045
rect 10784 15036 10836 15088
rect 13452 15036 13504 15088
rect 8484 14900 8536 14952
rect 11244 14968 11296 15020
rect 12808 14968 12860 15020
rect 8392 14764 8444 14816
rect 12348 14943 12400 14952
rect 12348 14909 12357 14943
rect 12357 14909 12391 14943
rect 12391 14909 12400 14943
rect 12348 14900 12400 14909
rect 16672 15036 16724 15088
rect 21456 15113 21465 15147
rect 21465 15113 21499 15147
rect 21499 15113 21508 15147
rect 21456 15104 21508 15113
rect 21088 15036 21140 15088
rect 13636 14832 13688 14884
rect 14740 14943 14792 14952
rect 14740 14909 14749 14943
rect 14749 14909 14783 14943
rect 14783 14909 14792 14943
rect 14740 14900 14792 14909
rect 15660 15011 15712 15020
rect 15660 14977 15669 15011
rect 15669 14977 15703 15011
rect 15703 14977 15712 15011
rect 15660 14968 15712 14977
rect 17960 15011 18012 15020
rect 17960 14977 17969 15011
rect 17969 14977 18003 15011
rect 18003 14977 18012 15011
rect 17960 14968 18012 14977
rect 21824 14968 21876 15020
rect 21916 14968 21968 15020
rect 24308 14968 24360 15020
rect 16120 14900 16172 14952
rect 18236 14943 18288 14952
rect 18236 14909 18245 14943
rect 18245 14909 18279 14943
rect 18279 14909 18288 14943
rect 18236 14900 18288 14909
rect 18328 14900 18380 14952
rect 18696 14900 18748 14952
rect 19156 14900 19208 14952
rect 19800 14900 19852 14952
rect 16212 14832 16264 14884
rect 22192 14900 22244 14952
rect 24676 14943 24728 14952
rect 24676 14909 24685 14943
rect 24685 14909 24719 14943
rect 24719 14909 24728 14943
rect 24676 14900 24728 14909
rect 22744 14875 22796 14884
rect 22744 14841 22753 14875
rect 22753 14841 22787 14875
rect 22787 14841 22796 14875
rect 22744 14832 22796 14841
rect 23940 14832 23992 14884
rect 16764 14764 16816 14816
rect 19432 14764 19484 14816
rect 19524 14764 19576 14816
rect 21456 14764 21508 14816
rect 22652 14764 22704 14816
rect 2950 14662 3002 14714
rect 3014 14662 3066 14714
rect 3078 14662 3130 14714
rect 3142 14662 3194 14714
rect 3206 14662 3258 14714
rect 12950 14662 13002 14714
rect 13014 14662 13066 14714
rect 13078 14662 13130 14714
rect 13142 14662 13194 14714
rect 13206 14662 13258 14714
rect 22950 14662 23002 14714
rect 23014 14662 23066 14714
rect 23078 14662 23130 14714
rect 23142 14662 23194 14714
rect 23206 14662 23258 14714
rect 8576 14603 8628 14612
rect 8576 14569 8585 14603
rect 8585 14569 8619 14603
rect 8619 14569 8628 14603
rect 8576 14560 8628 14569
rect 11060 14560 11112 14612
rect 14832 14603 14884 14612
rect 14832 14569 14841 14603
rect 14841 14569 14875 14603
rect 14875 14569 14884 14603
rect 14832 14560 14884 14569
rect 15660 14560 15712 14612
rect 17500 14560 17552 14612
rect 21916 14560 21968 14612
rect 11796 14492 11848 14544
rect 13820 14492 13872 14544
rect 19892 14492 19944 14544
rect 10876 14424 10928 14476
rect 11336 14424 11388 14476
rect 9956 14356 10008 14408
rect 13544 14467 13596 14476
rect 13544 14433 13553 14467
rect 13553 14433 13587 14467
rect 13587 14433 13596 14467
rect 13544 14424 13596 14433
rect 17960 14424 18012 14476
rect 22284 14424 22336 14476
rect 15108 14356 15160 14408
rect 15200 14356 15252 14408
rect 17316 14356 17368 14408
rect 18420 14399 18472 14408
rect 18420 14365 18429 14399
rect 18429 14365 18463 14399
rect 18463 14365 18472 14399
rect 18420 14356 18472 14365
rect 20904 14356 20956 14408
rect 9680 14288 9732 14340
rect 12716 14331 12768 14340
rect 12716 14297 12725 14331
rect 12725 14297 12759 14331
rect 12759 14297 12768 14331
rect 12716 14288 12768 14297
rect 13636 14288 13688 14340
rect 14832 14288 14884 14340
rect 15568 14331 15620 14340
rect 15568 14297 15577 14331
rect 15577 14297 15611 14331
rect 15611 14297 15620 14331
rect 15568 14288 15620 14297
rect 17040 14288 17092 14340
rect 17500 14288 17552 14340
rect 18788 14288 18840 14340
rect 22652 14288 22704 14340
rect 8668 14220 8720 14272
rect 11612 14220 11664 14272
rect 13452 14263 13504 14272
rect 13452 14229 13461 14263
rect 13461 14229 13495 14263
rect 13495 14229 13504 14263
rect 13452 14220 13504 14229
rect 13820 14220 13872 14272
rect 17684 14263 17736 14272
rect 17684 14229 17693 14263
rect 17693 14229 17727 14263
rect 17727 14229 17736 14263
rect 17684 14220 17736 14229
rect 22100 14220 22152 14272
rect 7950 14118 8002 14170
rect 8014 14118 8066 14170
rect 8078 14118 8130 14170
rect 8142 14118 8194 14170
rect 8206 14118 8258 14170
rect 17950 14118 18002 14170
rect 18014 14118 18066 14170
rect 18078 14118 18130 14170
rect 18142 14118 18194 14170
rect 18206 14118 18258 14170
rect 9956 14016 10008 14068
rect 11336 14016 11388 14068
rect 11704 14016 11756 14068
rect 1768 13923 1820 13932
rect 1768 13889 1777 13923
rect 1777 13889 1811 13923
rect 1811 13889 1820 13923
rect 1768 13880 1820 13889
rect 12532 14016 12584 14068
rect 12900 14059 12952 14068
rect 12900 14025 12909 14059
rect 12909 14025 12943 14059
rect 12943 14025 12952 14059
rect 12900 14016 12952 14025
rect 13360 14016 13412 14068
rect 14924 14059 14976 14068
rect 14924 14025 14933 14059
rect 14933 14025 14967 14059
rect 14967 14025 14976 14059
rect 14924 14016 14976 14025
rect 15568 14016 15620 14068
rect 19156 14059 19208 14068
rect 19156 14025 19165 14059
rect 19165 14025 19199 14059
rect 19199 14025 19208 14059
rect 19156 14016 19208 14025
rect 21916 14016 21968 14068
rect 22836 14016 22888 14068
rect 15660 13948 15712 14000
rect 17316 13948 17368 14000
rect 20536 13991 20588 14000
rect 20536 13957 20545 13991
rect 20545 13957 20579 13991
rect 20579 13957 20588 13991
rect 20536 13948 20588 13957
rect 25136 13991 25188 14000
rect 25136 13957 25145 13991
rect 25145 13957 25179 13991
rect 25179 13957 25188 13991
rect 25136 13948 25188 13957
rect 12900 13880 12952 13932
rect 1308 13812 1360 13864
rect 5264 13812 5316 13864
rect 6736 13812 6788 13864
rect 8484 13812 8536 13864
rect 14924 13880 14976 13932
rect 11704 13744 11756 13796
rect 14648 13812 14700 13864
rect 15568 13812 15620 13864
rect 16580 13880 16632 13932
rect 17040 13880 17092 13932
rect 18880 13880 18932 13932
rect 22560 13880 22612 13932
rect 23848 13880 23900 13932
rect 18144 13812 18196 13864
rect 19064 13812 19116 13864
rect 19248 13812 19300 13864
rect 19432 13812 19484 13864
rect 20260 13812 20312 13864
rect 20628 13855 20680 13864
rect 20628 13821 20637 13855
rect 20637 13821 20671 13855
rect 20671 13821 20680 13855
rect 20628 13812 20680 13821
rect 8392 13676 8444 13728
rect 8852 13676 8904 13728
rect 17500 13676 17552 13728
rect 2950 13574 3002 13626
rect 3014 13574 3066 13626
rect 3078 13574 3130 13626
rect 3142 13574 3194 13626
rect 3206 13574 3258 13626
rect 12950 13574 13002 13626
rect 13014 13574 13066 13626
rect 13078 13574 13130 13626
rect 13142 13574 13194 13626
rect 13206 13574 13258 13626
rect 22950 13574 23002 13626
rect 23014 13574 23066 13626
rect 23078 13574 23130 13626
rect 23142 13574 23194 13626
rect 23206 13574 23258 13626
rect 8484 13472 8536 13524
rect 19616 13472 19668 13524
rect 17776 13404 17828 13456
rect 20812 13404 20864 13456
rect 10508 13336 10560 13388
rect 10968 13379 11020 13388
rect 10968 13345 10977 13379
rect 10977 13345 11011 13379
rect 11011 13345 11020 13379
rect 10968 13336 11020 13345
rect 13544 13336 13596 13388
rect 14004 13336 14056 13388
rect 14280 13311 14332 13320
rect 14280 13277 14289 13311
rect 14289 13277 14323 13311
rect 14323 13277 14332 13311
rect 14280 13268 14332 13277
rect 15384 13268 15436 13320
rect 16212 13336 16264 13388
rect 17040 13379 17092 13388
rect 17040 13345 17049 13379
rect 17049 13345 17083 13379
rect 17083 13345 17092 13379
rect 17040 13336 17092 13345
rect 18144 13379 18196 13388
rect 18144 13345 18153 13379
rect 18153 13345 18187 13379
rect 18187 13345 18196 13379
rect 18144 13336 18196 13345
rect 18696 13336 18748 13388
rect 19708 13336 19760 13388
rect 19984 13336 20036 13388
rect 19340 13268 19392 13320
rect 19892 13268 19944 13320
rect 22100 13268 22152 13320
rect 7104 13200 7156 13252
rect 13360 13200 13412 13252
rect 16304 13200 16356 13252
rect 18420 13200 18472 13252
rect 19984 13200 20036 13252
rect 20536 13200 20588 13252
rect 24952 13200 25004 13252
rect 12348 13132 12400 13184
rect 13636 13175 13688 13184
rect 13636 13141 13645 13175
rect 13645 13141 13679 13175
rect 13679 13141 13688 13175
rect 13636 13132 13688 13141
rect 14924 13175 14976 13184
rect 14924 13141 14933 13175
rect 14933 13141 14967 13175
rect 14967 13141 14976 13175
rect 14924 13132 14976 13141
rect 16856 13175 16908 13184
rect 16856 13141 16865 13175
rect 16865 13141 16899 13175
rect 16899 13141 16908 13175
rect 16856 13132 16908 13141
rect 20812 13132 20864 13184
rect 7950 13030 8002 13082
rect 8014 13030 8066 13082
rect 8078 13030 8130 13082
rect 8142 13030 8194 13082
rect 8206 13030 8258 13082
rect 17950 13030 18002 13082
rect 18014 13030 18066 13082
rect 18078 13030 18130 13082
rect 18142 13030 18194 13082
rect 18206 13030 18258 13082
rect 10968 12928 11020 12980
rect 12808 12928 12860 12980
rect 9128 12903 9180 12912
rect 9128 12869 9137 12903
rect 9137 12869 9171 12903
rect 9171 12869 9180 12903
rect 9128 12860 9180 12869
rect 4988 12792 5040 12844
rect 8760 12792 8812 12844
rect 11704 12835 11756 12844
rect 11704 12801 11713 12835
rect 11713 12801 11747 12835
rect 11747 12801 11756 12835
rect 11704 12792 11756 12801
rect 8852 12767 8904 12776
rect 8852 12733 8861 12767
rect 8861 12733 8895 12767
rect 8895 12733 8904 12767
rect 8852 12724 8904 12733
rect 9588 12724 9640 12776
rect 10324 12724 10376 12776
rect 11888 12656 11940 12708
rect 14004 12928 14056 12980
rect 15200 12928 15252 12980
rect 15292 12860 15344 12912
rect 16856 12860 16908 12912
rect 18328 12928 18380 12980
rect 18880 12928 18932 12980
rect 19892 12971 19944 12980
rect 19892 12937 19901 12971
rect 19901 12937 19935 12971
rect 19935 12937 19944 12971
rect 19892 12928 19944 12937
rect 21180 12971 21232 12980
rect 21180 12937 21189 12971
rect 21189 12937 21223 12971
rect 21223 12937 21232 12971
rect 21180 12928 21232 12937
rect 20352 12860 20404 12912
rect 14188 12724 14240 12776
rect 13728 12656 13780 12708
rect 12072 12588 12124 12640
rect 22192 12792 22244 12844
rect 23388 12792 23440 12844
rect 15476 12724 15528 12776
rect 17040 12724 17092 12776
rect 20628 12724 20680 12776
rect 22008 12724 22060 12776
rect 24768 12767 24820 12776
rect 24768 12733 24777 12767
rect 24777 12733 24811 12767
rect 24811 12733 24820 12767
rect 24768 12724 24820 12733
rect 15200 12588 15252 12640
rect 15384 12588 15436 12640
rect 16120 12588 16172 12640
rect 17500 12631 17552 12640
rect 17500 12597 17509 12631
rect 17509 12597 17543 12631
rect 17543 12597 17552 12631
rect 17500 12588 17552 12597
rect 20352 12588 20404 12640
rect 20720 12631 20772 12640
rect 20720 12597 20729 12631
rect 20729 12597 20763 12631
rect 20763 12597 20772 12631
rect 20720 12588 20772 12597
rect 22100 12588 22152 12640
rect 2950 12486 3002 12538
rect 3014 12486 3066 12538
rect 3078 12486 3130 12538
rect 3142 12486 3194 12538
rect 3206 12486 3258 12538
rect 12950 12486 13002 12538
rect 13014 12486 13066 12538
rect 13078 12486 13130 12538
rect 13142 12486 13194 12538
rect 13206 12486 13258 12538
rect 22950 12486 23002 12538
rect 23014 12486 23066 12538
rect 23078 12486 23130 12538
rect 23142 12486 23194 12538
rect 23206 12486 23258 12538
rect 1860 12384 1912 12436
rect 9496 12384 9548 12436
rect 11704 12384 11756 12436
rect 13452 12384 13504 12436
rect 16212 12384 16264 12436
rect 14188 12316 14240 12368
rect 9588 12291 9640 12300
rect 9588 12257 9597 12291
rect 9597 12257 9631 12291
rect 9631 12257 9640 12291
rect 9588 12248 9640 12257
rect 10876 12248 10928 12300
rect 12072 12291 12124 12300
rect 12072 12257 12081 12291
rect 12081 12257 12115 12291
rect 12115 12257 12124 12291
rect 12072 12248 12124 12257
rect 14280 12248 14332 12300
rect 15016 12248 15068 12300
rect 11796 12223 11848 12232
rect 11796 12189 11805 12223
rect 11805 12189 11839 12223
rect 11839 12189 11848 12223
rect 11796 12180 11848 12189
rect 14372 12223 14424 12232
rect 14372 12189 14381 12223
rect 14381 12189 14415 12223
rect 14415 12189 14424 12223
rect 14372 12180 14424 12189
rect 15752 12316 15804 12368
rect 18420 12316 18472 12368
rect 16028 12248 16080 12300
rect 18696 12180 18748 12232
rect 24860 12316 24912 12368
rect 20904 12248 20956 12300
rect 21548 12248 21600 12300
rect 21824 12180 21876 12232
rect 23480 12223 23532 12232
rect 23480 12189 23489 12223
rect 23489 12189 23523 12223
rect 23523 12189 23532 12223
rect 23480 12180 23532 12189
rect 9864 12155 9916 12164
rect 9864 12121 9873 12155
rect 9873 12121 9907 12155
rect 9907 12121 9916 12155
rect 9864 12112 9916 12121
rect 2780 12044 2832 12096
rect 5172 12044 5224 12096
rect 10324 12112 10376 12164
rect 13728 12044 13780 12096
rect 15292 12112 15344 12164
rect 16212 12112 16264 12164
rect 19524 12112 19576 12164
rect 19800 12112 19852 12164
rect 14280 12044 14332 12096
rect 15568 12087 15620 12096
rect 15568 12053 15577 12087
rect 15577 12053 15611 12087
rect 15611 12053 15620 12087
rect 15568 12044 15620 12053
rect 15752 12044 15804 12096
rect 16856 12087 16908 12096
rect 16856 12053 16865 12087
rect 16865 12053 16899 12087
rect 16899 12053 16908 12087
rect 16856 12044 16908 12053
rect 17408 12044 17460 12096
rect 17592 12087 17644 12096
rect 17592 12053 17601 12087
rect 17601 12053 17635 12087
rect 17635 12053 17644 12087
rect 17592 12044 17644 12053
rect 18880 12087 18932 12096
rect 18880 12053 18889 12087
rect 18889 12053 18923 12087
rect 18923 12053 18932 12087
rect 18880 12044 18932 12053
rect 21180 12112 21232 12164
rect 20812 12044 20864 12096
rect 22008 12044 22060 12096
rect 22652 12044 22704 12096
rect 23296 12087 23348 12096
rect 23296 12053 23305 12087
rect 23305 12053 23339 12087
rect 23339 12053 23348 12087
rect 23296 12044 23348 12053
rect 7950 11942 8002 11994
rect 8014 11942 8066 11994
rect 8078 11942 8130 11994
rect 8142 11942 8194 11994
rect 8206 11942 8258 11994
rect 17950 11942 18002 11994
rect 18014 11942 18066 11994
rect 18078 11942 18130 11994
rect 18142 11942 18194 11994
rect 18206 11942 18258 11994
rect 9864 11840 9916 11892
rect 14740 11883 14792 11892
rect 14740 11849 14749 11883
rect 14749 11849 14783 11883
rect 14783 11849 14792 11883
rect 14740 11840 14792 11849
rect 17592 11840 17644 11892
rect 20628 11840 20680 11892
rect 21180 11883 21232 11892
rect 21180 11849 21189 11883
rect 21189 11849 21223 11883
rect 21223 11849 21232 11883
rect 21180 11840 21232 11849
rect 5908 11772 5960 11824
rect 10416 11772 10468 11824
rect 13728 11772 13780 11824
rect 15660 11815 15712 11824
rect 15660 11781 15669 11815
rect 15669 11781 15703 11815
rect 15703 11781 15712 11815
rect 15660 11772 15712 11781
rect 16212 11815 16264 11824
rect 16212 11781 16221 11815
rect 16221 11781 16255 11815
rect 16255 11781 16264 11815
rect 16212 11772 16264 11781
rect 10968 11704 11020 11756
rect 11796 11704 11848 11756
rect 15016 11704 15068 11756
rect 18328 11772 18380 11824
rect 20260 11772 20312 11824
rect 21824 11772 21876 11824
rect 25136 11815 25188 11824
rect 25136 11781 25145 11815
rect 25145 11781 25179 11815
rect 25179 11781 25188 11815
rect 25136 11772 25188 11781
rect 10324 11636 10376 11688
rect 14924 11636 14976 11688
rect 18880 11636 18932 11688
rect 19708 11704 19760 11756
rect 20352 11704 20404 11756
rect 21180 11704 21232 11756
rect 22744 11704 22796 11756
rect 11612 11568 11664 11620
rect 11796 11568 11848 11620
rect 11980 11500 12032 11552
rect 16856 11500 16908 11552
rect 18328 11500 18380 11552
rect 19708 11543 19760 11552
rect 19708 11509 19717 11543
rect 19717 11509 19751 11543
rect 19751 11509 19760 11543
rect 19708 11500 19760 11509
rect 2950 11398 3002 11450
rect 3014 11398 3066 11450
rect 3078 11398 3130 11450
rect 3142 11398 3194 11450
rect 3206 11398 3258 11450
rect 12950 11398 13002 11450
rect 13014 11398 13066 11450
rect 13078 11398 13130 11450
rect 13142 11398 13194 11450
rect 13206 11398 13258 11450
rect 22950 11398 23002 11450
rect 23014 11398 23066 11450
rect 23078 11398 23130 11450
rect 23142 11398 23194 11450
rect 23206 11398 23258 11450
rect 15476 11339 15528 11348
rect 15476 11305 15485 11339
rect 15485 11305 15519 11339
rect 15519 11305 15528 11339
rect 15476 11296 15528 11305
rect 21732 11296 21784 11348
rect 16028 11228 16080 11280
rect 17776 11228 17828 11280
rect 12348 11160 12400 11212
rect 14740 11092 14792 11144
rect 16028 11135 16080 11144
rect 16028 11101 16037 11135
rect 16037 11101 16071 11135
rect 16071 11101 16080 11135
rect 16028 11092 16080 11101
rect 18604 11160 18656 11212
rect 22192 11228 22244 11280
rect 23388 11228 23440 11280
rect 21732 11135 21784 11144
rect 21732 11101 21741 11135
rect 21741 11101 21775 11135
rect 21775 11101 21784 11135
rect 21732 11092 21784 11101
rect 16764 11024 16816 11076
rect 18696 11024 18748 11076
rect 21088 11024 21140 11076
rect 23848 11024 23900 11076
rect 19524 10999 19576 11008
rect 19524 10965 19533 10999
rect 19533 10965 19567 10999
rect 19567 10965 19576 10999
rect 19524 10956 19576 10965
rect 7950 10854 8002 10906
rect 8014 10854 8066 10906
rect 8078 10854 8130 10906
rect 8142 10854 8194 10906
rect 8206 10854 8258 10906
rect 17950 10854 18002 10906
rect 18014 10854 18066 10906
rect 18078 10854 18130 10906
rect 18142 10854 18194 10906
rect 18206 10854 18258 10906
rect 19524 10795 19576 10804
rect 19524 10761 19533 10795
rect 19533 10761 19567 10795
rect 19567 10761 19576 10795
rect 19524 10752 19576 10761
rect 19616 10795 19668 10804
rect 19616 10761 19625 10795
rect 19625 10761 19659 10795
rect 19659 10761 19668 10795
rect 19616 10752 19668 10761
rect 21088 10752 21140 10804
rect 10048 10684 10100 10736
rect 18328 10616 18380 10668
rect 20720 10616 20772 10668
rect 23940 10659 23992 10668
rect 23940 10625 23949 10659
rect 23949 10625 23983 10659
rect 23983 10625 23992 10659
rect 23940 10616 23992 10625
rect 18788 10548 18840 10600
rect 19156 10548 19208 10600
rect 19708 10591 19760 10600
rect 19708 10557 19717 10591
rect 19717 10557 19751 10591
rect 19751 10557 19760 10591
rect 19708 10548 19760 10557
rect 24768 10591 24820 10600
rect 24768 10557 24777 10591
rect 24777 10557 24811 10591
rect 24811 10557 24820 10591
rect 24768 10548 24820 10557
rect 12532 10480 12584 10532
rect 20628 10480 20680 10532
rect 21180 10412 21232 10464
rect 22560 10412 22612 10464
rect 2950 10310 3002 10362
rect 3014 10310 3066 10362
rect 3078 10310 3130 10362
rect 3142 10310 3194 10362
rect 3206 10310 3258 10362
rect 12950 10310 13002 10362
rect 13014 10310 13066 10362
rect 13078 10310 13130 10362
rect 13142 10310 13194 10362
rect 13206 10310 13258 10362
rect 22950 10310 23002 10362
rect 23014 10310 23066 10362
rect 23078 10310 23130 10362
rect 23142 10310 23194 10362
rect 23206 10310 23258 10362
rect 12624 10004 12676 10056
rect 18512 10004 18564 10056
rect 21916 10004 21968 10056
rect 22652 10047 22704 10056
rect 22652 10013 22661 10047
rect 22661 10013 22695 10047
rect 22695 10013 22704 10047
rect 22652 10004 22704 10013
rect 22836 10004 22888 10056
rect 14832 9936 14884 9988
rect 24952 9936 25004 9988
rect 16948 9911 17000 9920
rect 16948 9877 16957 9911
rect 16957 9877 16991 9911
rect 16991 9877 17000 9911
rect 16948 9868 17000 9877
rect 21824 9868 21876 9920
rect 23572 9868 23624 9920
rect 7950 9766 8002 9818
rect 8014 9766 8066 9818
rect 8078 9766 8130 9818
rect 8142 9766 8194 9818
rect 8206 9766 8258 9818
rect 17950 9766 18002 9818
rect 18014 9766 18066 9818
rect 18078 9766 18130 9818
rect 18142 9766 18194 9818
rect 18206 9766 18258 9818
rect 22652 9664 22704 9716
rect 10048 9596 10100 9648
rect 14096 9596 14148 9648
rect 17500 9596 17552 9648
rect 19064 9596 19116 9648
rect 22008 9596 22060 9648
rect 7656 9528 7708 9580
rect 12440 9528 12492 9580
rect 20628 9528 20680 9580
rect 23848 9528 23900 9580
rect 2872 9460 2924 9512
rect 5724 9460 5776 9512
rect 7472 9460 7524 9512
rect 24676 9503 24728 9512
rect 24676 9469 24685 9503
rect 24685 9469 24719 9503
rect 24719 9469 24728 9503
rect 24676 9460 24728 9469
rect 17408 9392 17460 9444
rect 22836 9392 22888 9444
rect 23480 9324 23532 9376
rect 2950 9222 3002 9274
rect 3014 9222 3066 9274
rect 3078 9222 3130 9274
rect 3142 9222 3194 9274
rect 3206 9222 3258 9274
rect 12950 9222 13002 9274
rect 13014 9222 13066 9274
rect 13078 9222 13130 9274
rect 13142 9222 13194 9274
rect 13206 9222 13258 9274
rect 22950 9222 23002 9274
rect 23014 9222 23066 9274
rect 23078 9222 23130 9274
rect 23142 9222 23194 9274
rect 23206 9222 23258 9274
rect 7104 9163 7156 9172
rect 7104 9129 7113 9163
rect 7113 9129 7147 9163
rect 7147 9129 7156 9163
rect 7104 9120 7156 9129
rect 9036 8984 9088 9036
rect 7472 8959 7524 8968
rect 7472 8925 7481 8959
rect 7481 8925 7515 8959
rect 7515 8925 7524 8959
rect 7472 8916 7524 8925
rect 23296 8916 23348 8968
rect 24860 8959 24912 8968
rect 24860 8925 24869 8959
rect 24869 8925 24903 8959
rect 24903 8925 24912 8959
rect 24860 8916 24912 8925
rect 5632 8780 5684 8832
rect 9496 8848 9548 8900
rect 13912 8848 13964 8900
rect 23296 8780 23348 8832
rect 23940 8823 23992 8832
rect 23940 8789 23949 8823
rect 23949 8789 23983 8823
rect 23983 8789 23992 8823
rect 23940 8780 23992 8789
rect 7950 8678 8002 8730
rect 8014 8678 8066 8730
rect 8078 8678 8130 8730
rect 8142 8678 8194 8730
rect 8206 8678 8258 8730
rect 17950 8678 18002 8730
rect 18014 8678 18066 8730
rect 18078 8678 18130 8730
rect 18142 8678 18194 8730
rect 18206 8678 18258 8730
rect 5264 8576 5316 8628
rect 10324 8508 10376 8560
rect 17040 8508 17092 8560
rect 21364 8508 21416 8560
rect 25136 8551 25188 8560
rect 25136 8517 25145 8551
rect 25145 8517 25179 8551
rect 25179 8517 25188 8551
rect 25136 8508 25188 8517
rect 6828 8440 6880 8492
rect 22376 8440 22428 8492
rect 23388 8440 23440 8492
rect 2780 8372 2832 8424
rect 22744 8415 22796 8424
rect 22744 8381 22753 8415
rect 22753 8381 22787 8415
rect 22787 8381 22796 8415
rect 22744 8372 22796 8381
rect 20444 8304 20496 8356
rect 21272 8304 21324 8356
rect 2950 8134 3002 8186
rect 3014 8134 3066 8186
rect 3078 8134 3130 8186
rect 3142 8134 3194 8186
rect 3206 8134 3258 8186
rect 12950 8134 13002 8186
rect 13014 8134 13066 8186
rect 13078 8134 13130 8186
rect 13142 8134 13194 8186
rect 13206 8134 13258 8186
rect 22950 8134 23002 8186
rect 23014 8134 23066 8186
rect 23078 8134 23130 8186
rect 23142 8134 23194 8186
rect 23206 8134 23258 8186
rect 23296 7939 23348 7948
rect 23296 7905 23305 7939
rect 23305 7905 23339 7939
rect 23339 7905 23348 7939
rect 23296 7896 23348 7905
rect 19800 7828 19852 7880
rect 21180 7828 21232 7880
rect 23572 7828 23624 7880
rect 20260 7692 20312 7744
rect 24676 7692 24728 7744
rect 7950 7590 8002 7642
rect 8014 7590 8066 7642
rect 8078 7590 8130 7642
rect 8142 7590 8194 7642
rect 8206 7590 8258 7642
rect 17950 7590 18002 7642
rect 18014 7590 18066 7642
rect 18078 7590 18130 7642
rect 18142 7590 18194 7642
rect 18206 7590 18258 7642
rect 15200 7420 15252 7472
rect 15844 7352 15896 7404
rect 20444 7420 20496 7472
rect 20720 7352 20772 7404
rect 25136 7463 25188 7472
rect 25136 7429 25145 7463
rect 25145 7429 25179 7463
rect 25179 7429 25188 7463
rect 25136 7420 25188 7429
rect 16212 7284 16264 7336
rect 17684 7216 17736 7268
rect 21640 7284 21692 7336
rect 22284 7284 22336 7336
rect 20628 7148 20680 7200
rect 2950 7046 3002 7098
rect 3014 7046 3066 7098
rect 3078 7046 3130 7098
rect 3142 7046 3194 7098
rect 3206 7046 3258 7098
rect 12950 7046 13002 7098
rect 13014 7046 13066 7098
rect 13078 7046 13130 7098
rect 13142 7046 13194 7098
rect 13206 7046 13258 7098
rect 22950 7046 23002 7098
rect 23014 7046 23066 7098
rect 23078 7046 23130 7098
rect 23142 7046 23194 7098
rect 23206 7046 23258 7098
rect 15568 6740 15620 6792
rect 3056 6672 3108 6724
rect 6092 6672 6144 6724
rect 23388 6740 23440 6792
rect 22008 6715 22060 6724
rect 22008 6681 22017 6715
rect 22017 6681 22051 6715
rect 22051 6681 22060 6715
rect 22008 6672 22060 6681
rect 25780 6672 25832 6724
rect 7950 6502 8002 6554
rect 8014 6502 8066 6554
rect 8078 6502 8130 6554
rect 8142 6502 8194 6554
rect 8206 6502 8258 6554
rect 17950 6502 18002 6554
rect 18014 6502 18066 6554
rect 18078 6502 18130 6554
rect 18142 6502 18194 6554
rect 18206 6502 18258 6554
rect 11796 6400 11848 6452
rect 5540 6264 5592 6316
rect 9772 6264 9824 6316
rect 20260 6307 20312 6316
rect 20260 6273 20269 6307
rect 20269 6273 20303 6307
rect 20303 6273 20312 6307
rect 20260 6264 20312 6273
rect 22192 6307 22244 6316
rect 22192 6273 22201 6307
rect 22201 6273 22235 6307
rect 22235 6273 22244 6307
rect 22192 6264 22244 6273
rect 23480 6264 23532 6316
rect 21732 6196 21784 6248
rect 21916 6196 21968 6248
rect 24768 6239 24820 6248
rect 24768 6205 24777 6239
rect 24777 6205 24811 6239
rect 24811 6205 24820 6239
rect 24768 6196 24820 6205
rect 22192 6128 22244 6180
rect 2950 5958 3002 6010
rect 3014 5958 3066 6010
rect 3078 5958 3130 6010
rect 3142 5958 3194 6010
rect 3206 5958 3258 6010
rect 12950 5958 13002 6010
rect 13014 5958 13066 6010
rect 13078 5958 13130 6010
rect 13142 5958 13194 6010
rect 13206 5958 13258 6010
rect 22950 5958 23002 6010
rect 23014 5958 23066 6010
rect 23078 5958 23130 6010
rect 23142 5958 23194 6010
rect 23206 5958 23258 6010
rect 20720 5856 20772 5908
rect 10600 5788 10652 5840
rect 11888 5788 11940 5840
rect 20444 5720 20496 5772
rect 21548 5720 21600 5772
rect 9312 5652 9364 5704
rect 13452 5652 13504 5704
rect 20536 5695 20588 5704
rect 20536 5661 20545 5695
rect 20545 5661 20579 5695
rect 20579 5661 20588 5695
rect 20536 5652 20588 5661
rect 20628 5652 20680 5704
rect 2688 5584 2740 5636
rect 9404 5584 9456 5636
rect 21824 5584 21876 5636
rect 5172 5516 5224 5568
rect 6276 5516 6328 5568
rect 12624 5516 12676 5568
rect 14556 5516 14608 5568
rect 7950 5414 8002 5466
rect 8014 5414 8066 5466
rect 8078 5414 8130 5466
rect 8142 5414 8194 5466
rect 8206 5414 8258 5466
rect 17950 5414 18002 5466
rect 18014 5414 18066 5466
rect 18078 5414 18130 5466
rect 18142 5414 18194 5466
rect 18206 5414 18258 5466
rect 19524 5244 19576 5296
rect 17776 5219 17828 5228
rect 17776 5185 17785 5219
rect 17785 5185 17819 5219
rect 17819 5185 17828 5219
rect 17776 5176 17828 5185
rect 19064 5176 19116 5228
rect 22100 5219 22152 5228
rect 22100 5185 22109 5219
rect 22109 5185 22143 5219
rect 22143 5185 22152 5219
rect 22100 5176 22152 5185
rect 23940 5219 23992 5228
rect 23940 5185 23949 5219
rect 23949 5185 23983 5219
rect 23983 5185 23992 5219
rect 23940 5176 23992 5185
rect 19340 5108 19392 5160
rect 22468 5151 22520 5160
rect 22468 5117 22477 5151
rect 22477 5117 22511 5151
rect 22511 5117 22520 5151
rect 22468 5108 22520 5117
rect 24768 5151 24820 5160
rect 24768 5117 24777 5151
rect 24777 5117 24811 5151
rect 24811 5117 24820 5151
rect 24768 5108 24820 5117
rect 2950 4870 3002 4922
rect 3014 4870 3066 4922
rect 3078 4870 3130 4922
rect 3142 4870 3194 4922
rect 3206 4870 3258 4922
rect 12950 4870 13002 4922
rect 13014 4870 13066 4922
rect 13078 4870 13130 4922
rect 13142 4870 13194 4922
rect 13206 4870 13258 4922
rect 22950 4870 23002 4922
rect 23014 4870 23066 4922
rect 23078 4870 23130 4922
rect 23142 4870 23194 4922
rect 23206 4870 23258 4922
rect 22376 4768 22428 4820
rect 17776 4700 17828 4752
rect 19892 4675 19944 4684
rect 19892 4641 19901 4675
rect 19901 4641 19935 4675
rect 19935 4641 19944 4675
rect 19892 4632 19944 4641
rect 20720 4632 20772 4684
rect 22560 4632 22612 4684
rect 17684 4607 17736 4616
rect 17684 4573 17693 4607
rect 17693 4573 17727 4607
rect 17727 4573 17736 4607
rect 17684 4564 17736 4573
rect 18696 4564 18748 4616
rect 21272 4607 21324 4616
rect 21272 4573 21281 4607
rect 21281 4573 21315 4607
rect 21315 4573 21324 4607
rect 21272 4564 21324 4573
rect 24676 4607 24728 4616
rect 24676 4573 24685 4607
rect 24685 4573 24719 4607
rect 24719 4573 24728 4607
rect 24676 4564 24728 4573
rect 20628 4496 20680 4548
rect 7950 4326 8002 4378
rect 8014 4326 8066 4378
rect 8078 4326 8130 4378
rect 8142 4326 8194 4378
rect 8206 4326 8258 4378
rect 17950 4326 18002 4378
rect 18014 4326 18066 4378
rect 18078 4326 18130 4378
rect 18142 4326 18194 4378
rect 18206 4326 18258 4378
rect 2596 4224 2648 4276
rect 8300 4224 8352 4276
rect 15108 4156 15160 4208
rect 16488 4156 16540 4208
rect 11980 4131 12032 4140
rect 11980 4097 11989 4131
rect 11989 4097 12023 4131
rect 12023 4097 12032 4131
rect 11980 4088 12032 4097
rect 13544 4131 13596 4140
rect 13544 4097 13553 4131
rect 13553 4097 13587 4131
rect 13587 4097 13596 4131
rect 13544 4088 13596 4097
rect 16120 4131 16172 4140
rect 16120 4097 16129 4131
rect 16129 4097 16163 4131
rect 16163 4097 16172 4131
rect 16120 4088 16172 4097
rect 16212 4088 16264 4140
rect 16672 4088 16724 4140
rect 19248 4088 19300 4140
rect 19984 4088 20036 4140
rect 22836 4088 22888 4140
rect 2872 4020 2924 4072
rect 5080 4020 5132 4072
rect 11612 4020 11664 4072
rect 13452 4020 13504 4072
rect 16396 4020 16448 4072
rect 17500 4020 17552 4072
rect 20076 4020 20128 4072
rect 2780 3952 2832 4004
rect 9036 3952 9088 4004
rect 21180 3952 21232 4004
rect 2872 3884 2924 3936
rect 6092 3884 6144 3936
rect 9404 3884 9456 3936
rect 9772 3927 9824 3936
rect 9772 3893 9781 3927
rect 9781 3893 9815 3927
rect 9815 3893 9824 3927
rect 9772 3884 9824 3893
rect 10508 3884 10560 3936
rect 19524 3884 19576 3936
rect 22100 3884 22152 3936
rect 2950 3782 3002 3834
rect 3014 3782 3066 3834
rect 3078 3782 3130 3834
rect 3142 3782 3194 3834
rect 3206 3782 3258 3834
rect 12950 3782 13002 3834
rect 13014 3782 13066 3834
rect 13078 3782 13130 3834
rect 13142 3782 13194 3834
rect 13206 3782 13258 3834
rect 22950 3782 23002 3834
rect 23014 3782 23066 3834
rect 23078 3782 23130 3834
rect 23142 3782 23194 3834
rect 23206 3782 23258 3834
rect 5540 3680 5592 3732
rect 6000 3680 6052 3732
rect 7380 3680 7432 3732
rect 9496 3680 9548 3732
rect 10048 3723 10100 3732
rect 10048 3689 10057 3723
rect 10057 3689 10091 3723
rect 10091 3689 10100 3723
rect 10048 3680 10100 3689
rect 5632 3612 5684 3664
rect 16120 3612 16172 3664
rect 19156 3612 19208 3664
rect 8300 3544 8352 3596
rect 12716 3544 12768 3596
rect 14924 3544 14976 3596
rect 16028 3544 16080 3596
rect 17776 3544 17828 3596
rect 1676 3476 1728 3528
rect 3332 3408 3384 3460
rect 6092 3519 6144 3528
rect 6092 3485 6101 3519
rect 6101 3485 6135 3519
rect 6135 3485 6144 3519
rect 6092 3476 6144 3485
rect 6460 3476 6512 3528
rect 9404 3476 9456 3528
rect 9772 3476 9824 3528
rect 10876 3476 10928 3528
rect 13636 3476 13688 3528
rect 15108 3519 15160 3528
rect 15108 3485 15117 3519
rect 15117 3485 15151 3519
rect 15151 3485 15160 3519
rect 15108 3476 15160 3485
rect 16304 3476 16356 3528
rect 17592 3476 17644 3528
rect 14740 3408 14792 3460
rect 18972 3408 19024 3460
rect 22192 3408 22244 3460
rect 24952 3408 25004 3460
rect 2044 3340 2096 3392
rect 2780 3340 2832 3392
rect 3516 3340 3568 3392
rect 3884 3340 3936 3392
rect 4896 3340 4948 3392
rect 6828 3340 6880 3392
rect 7840 3340 7892 3392
rect 8668 3383 8720 3392
rect 8668 3349 8677 3383
rect 8677 3349 8711 3383
rect 8711 3349 8720 3383
rect 8668 3340 8720 3349
rect 11244 3340 11296 3392
rect 22008 3340 22060 3392
rect 22836 3340 22888 3392
rect 23572 3340 23624 3392
rect 24124 3340 24176 3392
rect 7950 3238 8002 3290
rect 8014 3238 8066 3290
rect 8078 3238 8130 3290
rect 8142 3238 8194 3290
rect 8206 3238 8258 3290
rect 17950 3238 18002 3290
rect 18014 3238 18066 3290
rect 18078 3238 18130 3290
rect 18142 3238 18194 3290
rect 18206 3238 18258 3290
rect 2688 3179 2740 3188
rect 2688 3145 2697 3179
rect 2697 3145 2731 3179
rect 2731 3145 2740 3179
rect 2688 3136 2740 3145
rect 5172 3179 5224 3188
rect 5172 3145 5181 3179
rect 5181 3145 5215 3179
rect 5215 3145 5224 3179
rect 5172 3136 5224 3145
rect 5908 3179 5960 3188
rect 5908 3145 5917 3179
rect 5917 3145 5951 3179
rect 5951 3145 5960 3179
rect 5908 3136 5960 3145
rect 7012 3179 7064 3188
rect 7012 3145 7021 3179
rect 7021 3145 7055 3179
rect 7055 3145 7064 3179
rect 7012 3136 7064 3145
rect 7288 3136 7340 3188
rect 8484 3179 8536 3188
rect 8484 3145 8493 3179
rect 8493 3145 8527 3179
rect 8527 3145 8536 3179
rect 8484 3136 8536 3145
rect 11888 3179 11940 3188
rect 11888 3145 11897 3179
rect 11897 3145 11931 3179
rect 11931 3145 11940 3179
rect 11888 3136 11940 3145
rect 22652 3136 22704 3188
rect 23572 3111 23624 3120
rect 23572 3077 23581 3111
rect 23581 3077 23615 3111
rect 23615 3077 23624 3111
rect 23572 3068 23624 3077
rect 2044 3000 2096 3052
rect 2780 3000 2832 3052
rect 5356 3000 5408 3052
rect 5724 3043 5776 3052
rect 5724 3009 5733 3043
rect 5733 3009 5767 3043
rect 5767 3009 5776 3043
rect 5724 3000 5776 3009
rect 6828 3043 6880 3052
rect 6828 3009 6837 3043
rect 6837 3009 6871 3043
rect 6871 3009 6880 3043
rect 6828 3000 6880 3009
rect 8208 3000 8260 3052
rect 8668 3000 8720 3052
rect 9312 3043 9364 3052
rect 9312 3009 9321 3043
rect 9321 3009 9355 3043
rect 9355 3009 9364 3043
rect 9312 3000 9364 3009
rect 10600 3043 10652 3052
rect 10600 3009 10609 3043
rect 10609 3009 10643 3043
rect 10643 3009 10652 3043
rect 10600 3000 10652 3009
rect 11244 3000 11296 3052
rect 12624 3043 12676 3052
rect 12624 3009 12633 3043
rect 12633 3009 12667 3043
rect 12667 3009 12676 3043
rect 12624 3000 12676 3009
rect 14280 3043 14332 3052
rect 14280 3009 14289 3043
rect 14289 3009 14323 3043
rect 14323 3009 14332 3043
rect 14280 3000 14332 3009
rect 16764 3000 16816 3052
rect 17868 3000 17920 3052
rect 18512 3000 18564 3052
rect 21732 3000 21784 3052
rect 22652 3000 22704 3052
rect 3332 2932 3384 2984
rect 7748 2932 7800 2984
rect 9036 2975 9088 2984
rect 9036 2941 9045 2975
rect 9045 2941 9079 2975
rect 9079 2941 9088 2975
rect 9036 2932 9088 2941
rect 10508 2932 10560 2984
rect 13360 2975 13412 2984
rect 13360 2941 13369 2975
rect 13369 2941 13403 2975
rect 13403 2941 13412 2975
rect 13360 2932 13412 2941
rect 14188 2932 14240 2984
rect 15660 2932 15712 2984
rect 5816 2864 5868 2916
rect 17132 2864 17184 2916
rect 20628 2932 20680 2984
rect 23388 2932 23440 2984
rect 19708 2864 19760 2916
rect 20720 2864 20772 2916
rect 1492 2839 1544 2848
rect 1492 2805 1501 2839
rect 1501 2805 1535 2839
rect 1535 2805 1544 2839
rect 1492 2796 1544 2805
rect 4252 2796 4304 2848
rect 6460 2839 6512 2848
rect 6460 2805 6469 2839
rect 6469 2805 6503 2839
rect 6503 2805 6512 2839
rect 6460 2796 6512 2805
rect 18604 2796 18656 2848
rect 19892 2796 19944 2848
rect 20812 2796 20864 2848
rect 22468 2796 22520 2848
rect 2950 2694 3002 2746
rect 3014 2694 3066 2746
rect 3078 2694 3130 2746
rect 3142 2694 3194 2746
rect 3206 2694 3258 2746
rect 12950 2694 13002 2746
rect 13014 2694 13066 2746
rect 13078 2694 13130 2746
rect 13142 2694 13194 2746
rect 13206 2694 13258 2746
rect 22950 2694 23002 2746
rect 23014 2694 23066 2746
rect 23078 2694 23130 2746
rect 23142 2694 23194 2746
rect 23206 2694 23258 2746
rect 1860 2635 1912 2644
rect 1860 2601 1869 2635
rect 1869 2601 1903 2635
rect 1903 2601 1912 2635
rect 1860 2592 1912 2601
rect 2596 2635 2648 2644
rect 2596 2601 2605 2635
rect 2605 2601 2639 2635
rect 2639 2601 2648 2635
rect 2596 2592 2648 2601
rect 4804 2592 4856 2644
rect 7656 2592 7708 2644
rect 11060 2592 11112 2644
rect 15752 2592 15804 2644
rect 17408 2592 17460 2644
rect 7564 2524 7616 2576
rect 4988 2499 5040 2508
rect 4988 2465 4997 2499
rect 4997 2465 5031 2499
rect 5031 2465 5040 2499
rect 4988 2456 5040 2465
rect 12808 2524 12860 2576
rect 14832 2524 14884 2576
rect 1492 2388 1544 2440
rect 2320 2388 2372 2440
rect 3516 2388 3568 2440
rect 4252 2388 4304 2440
rect 4620 2388 4672 2440
rect 7196 2388 7248 2440
rect 7564 2388 7616 2440
rect 10140 2388 10192 2440
rect 3884 2320 3936 2372
rect 5724 2320 5776 2372
rect 11704 2388 11756 2440
rect 11980 2456 12032 2508
rect 14556 2456 14608 2508
rect 15292 2456 15344 2508
rect 18512 2499 18564 2508
rect 18512 2465 18521 2499
rect 18521 2465 18555 2499
rect 18555 2465 18564 2499
rect 18512 2456 18564 2465
rect 12532 2431 12584 2440
rect 12532 2397 12541 2431
rect 12541 2397 12575 2431
rect 12575 2397 12584 2431
rect 12532 2388 12584 2397
rect 14648 2431 14700 2440
rect 14648 2397 14657 2431
rect 14657 2397 14691 2431
rect 14691 2397 14700 2431
rect 14648 2388 14700 2397
rect 16948 2431 17000 2440
rect 16948 2397 16957 2431
rect 16957 2397 16991 2431
rect 16991 2397 17000 2431
rect 16948 2388 17000 2397
rect 12348 2320 12400 2372
rect 13820 2320 13872 2372
rect 16764 2320 16816 2372
rect 18328 2252 18380 2304
rect 25320 2431 25372 2440
rect 25320 2397 25329 2431
rect 25329 2397 25363 2431
rect 25363 2397 25372 2431
rect 25320 2388 25372 2397
rect 7950 2150 8002 2202
rect 8014 2150 8066 2202
rect 8078 2150 8130 2202
rect 8142 2150 8194 2202
rect 8206 2150 8258 2202
rect 17950 2150 18002 2202
rect 18014 2150 18066 2202
rect 18078 2150 18130 2202
rect 18142 2150 18194 2202
rect 18206 2150 18258 2202
<< metal2 >>
rect 1490 56200 1546 57000
rect 1858 56200 1914 57000
rect 2226 56200 2282 57000
rect 2594 56200 2650 57000
rect 2962 56200 3018 57000
rect 3330 56200 3386 57000
rect 3698 56200 3754 57000
rect 4066 56200 4122 57000
rect 4434 56200 4490 57000
rect 4802 56200 4858 57000
rect 5170 56200 5226 57000
rect 5538 56200 5594 57000
rect 5906 56200 5962 57000
rect 6274 56200 6330 57000
rect 6642 56200 6698 57000
rect 7010 56200 7066 57000
rect 7378 56200 7434 57000
rect 7746 56200 7802 57000
rect 7852 56222 8064 56250
rect 1504 49298 1532 56200
rect 1872 52630 1900 56200
rect 2240 52698 2268 56200
rect 2608 52986 2636 56200
rect 2778 55448 2834 55457
rect 2778 55383 2834 55392
rect 2792 53242 2820 55383
rect 2976 55214 3004 56200
rect 2884 55186 3004 55214
rect 2780 53236 2832 53242
rect 2780 53178 2832 53184
rect 2608 52958 2820 52986
rect 2228 52692 2280 52698
rect 2228 52634 2280 52640
rect 1860 52624 1912 52630
rect 1860 52566 1912 52572
rect 2792 50862 2820 52958
rect 2884 51474 2912 55186
rect 2950 53884 3258 53893
rect 2950 53882 2956 53884
rect 3012 53882 3036 53884
rect 3092 53882 3116 53884
rect 3172 53882 3196 53884
rect 3252 53882 3258 53884
rect 3012 53830 3014 53882
rect 3194 53830 3196 53882
rect 2950 53828 2956 53830
rect 3012 53828 3036 53830
rect 3092 53828 3116 53830
rect 3172 53828 3196 53830
rect 3252 53828 3258 53830
rect 2950 53819 3258 53828
rect 2950 52796 3258 52805
rect 2950 52794 2956 52796
rect 3012 52794 3036 52796
rect 3092 52794 3116 52796
rect 3172 52794 3196 52796
rect 3252 52794 3258 52796
rect 3012 52742 3014 52794
rect 3194 52742 3196 52794
rect 2950 52740 2956 52742
rect 3012 52740 3036 52742
rect 3092 52740 3116 52742
rect 3172 52740 3196 52742
rect 3252 52740 3258 52742
rect 2950 52731 3258 52740
rect 3344 51950 3372 56200
rect 3422 53000 3478 53009
rect 3422 52935 3424 52944
rect 3476 52935 3478 52944
rect 3424 52906 3476 52912
rect 3424 52692 3476 52698
rect 3424 52634 3476 52640
rect 3332 51944 3384 51950
rect 3332 51886 3384 51892
rect 2950 51708 3258 51717
rect 2950 51706 2956 51708
rect 3012 51706 3036 51708
rect 3092 51706 3116 51708
rect 3172 51706 3196 51708
rect 3252 51706 3258 51708
rect 3012 51654 3014 51706
rect 3194 51654 3196 51706
rect 2950 51652 2956 51654
rect 3012 51652 3036 51654
rect 3092 51652 3116 51654
rect 3172 51652 3196 51654
rect 3252 51652 3258 51654
rect 2950 51643 3258 51652
rect 2872 51468 2924 51474
rect 2872 51410 2924 51416
rect 2780 50856 2832 50862
rect 2780 50798 2832 50804
rect 2950 50620 3258 50629
rect 2950 50618 2956 50620
rect 3012 50618 3036 50620
rect 3092 50618 3116 50620
rect 3172 50618 3196 50620
rect 3252 50618 3258 50620
rect 3012 50566 3014 50618
rect 3194 50566 3196 50618
rect 2950 50564 2956 50566
rect 3012 50564 3036 50566
rect 3092 50564 3116 50566
rect 3172 50564 3196 50566
rect 3252 50564 3258 50566
rect 2950 50555 3258 50564
rect 3436 50386 3464 52634
rect 3516 52624 3568 52630
rect 3516 52566 3568 52572
rect 3424 50380 3476 50386
rect 3424 50322 3476 50328
rect 3528 49910 3556 52566
rect 3712 52562 3740 56200
rect 4080 52986 4108 56200
rect 4344 54188 4396 54194
rect 4344 54130 4396 54136
rect 4080 52958 4292 52986
rect 4068 52896 4120 52902
rect 4068 52838 4120 52844
rect 3700 52556 3752 52562
rect 3700 52498 3752 52504
rect 3974 50416 4030 50425
rect 3974 50351 4030 50360
rect 3516 49904 3568 49910
rect 3516 49846 3568 49852
rect 3608 49836 3660 49842
rect 3608 49778 3660 49784
rect 2950 49532 3258 49541
rect 2950 49530 2956 49532
rect 3012 49530 3036 49532
rect 3092 49530 3116 49532
rect 3172 49530 3196 49532
rect 3252 49530 3258 49532
rect 3012 49478 3014 49530
rect 3194 49478 3196 49530
rect 2950 49476 2956 49478
rect 3012 49476 3036 49478
rect 3092 49476 3116 49478
rect 3172 49476 3196 49478
rect 3252 49476 3258 49478
rect 2950 49467 3258 49476
rect 1492 49292 1544 49298
rect 1492 49234 1544 49240
rect 2950 48444 3258 48453
rect 2950 48442 2956 48444
rect 3012 48442 3036 48444
rect 3092 48442 3116 48444
rect 3172 48442 3196 48444
rect 3252 48442 3258 48444
rect 3012 48390 3014 48442
rect 3194 48390 3196 48442
rect 2950 48388 2956 48390
rect 3012 48388 3036 48390
rect 3092 48388 3116 48390
rect 3172 48388 3196 48390
rect 3252 48388 3258 48390
rect 2950 48379 3258 48388
rect 2950 47356 3258 47365
rect 2950 47354 2956 47356
rect 3012 47354 3036 47356
rect 3092 47354 3116 47356
rect 3172 47354 3196 47356
rect 3252 47354 3258 47356
rect 3012 47302 3014 47354
rect 3194 47302 3196 47354
rect 2950 47300 2956 47302
rect 3012 47300 3036 47302
rect 3092 47300 3116 47302
rect 3172 47300 3196 47302
rect 3252 47300 3258 47302
rect 2950 47291 3258 47300
rect 2950 46268 3258 46277
rect 2950 46266 2956 46268
rect 3012 46266 3036 46268
rect 3092 46266 3116 46268
rect 3172 46266 3196 46268
rect 3252 46266 3258 46268
rect 3012 46214 3014 46266
rect 3194 46214 3196 46266
rect 2950 46212 2956 46214
rect 3012 46212 3036 46214
rect 3092 46212 3116 46214
rect 3172 46212 3196 46214
rect 3252 46212 3258 46214
rect 2950 46203 3258 46212
rect 2950 45180 3258 45189
rect 2950 45178 2956 45180
rect 3012 45178 3036 45180
rect 3092 45178 3116 45180
rect 3172 45178 3196 45180
rect 3252 45178 3258 45180
rect 3012 45126 3014 45178
rect 3194 45126 3196 45178
rect 2950 45124 2956 45126
rect 3012 45124 3036 45126
rect 3092 45124 3116 45126
rect 3172 45124 3196 45126
rect 3252 45124 3258 45126
rect 2950 45115 3258 45124
rect 2950 44092 3258 44101
rect 2950 44090 2956 44092
rect 3012 44090 3036 44092
rect 3092 44090 3116 44092
rect 3172 44090 3196 44092
rect 3252 44090 3258 44092
rect 3012 44038 3014 44090
rect 3194 44038 3196 44090
rect 2950 44036 2956 44038
rect 3012 44036 3036 44038
rect 3092 44036 3116 44038
rect 3172 44036 3196 44038
rect 3252 44036 3258 44038
rect 2950 44027 3258 44036
rect 1308 43308 1360 43314
rect 1308 43250 1360 43256
rect 1320 43217 1348 43250
rect 1306 43208 1362 43217
rect 1306 43143 1362 43152
rect 3516 43172 3568 43178
rect 3516 43114 3568 43120
rect 2950 43004 3258 43013
rect 2950 43002 2956 43004
rect 3012 43002 3036 43004
rect 3092 43002 3116 43004
rect 3172 43002 3196 43004
rect 3252 43002 3258 43004
rect 3012 42950 3014 43002
rect 3194 42950 3196 43002
rect 2950 42948 2956 42950
rect 3012 42948 3036 42950
rect 3092 42948 3116 42950
rect 3172 42948 3196 42950
rect 3252 42948 3258 42950
rect 2950 42939 3258 42948
rect 2950 41916 3258 41925
rect 2950 41914 2956 41916
rect 3012 41914 3036 41916
rect 3092 41914 3116 41916
rect 3172 41914 3196 41916
rect 3252 41914 3258 41916
rect 3012 41862 3014 41914
rect 3194 41862 3196 41914
rect 2950 41860 2956 41862
rect 3012 41860 3036 41862
rect 3092 41860 3116 41862
rect 3172 41860 3196 41862
rect 3252 41860 3258 41862
rect 2950 41851 3258 41860
rect 1308 41132 1360 41138
rect 1308 41074 1360 41080
rect 1320 40769 1348 41074
rect 2950 40828 3258 40837
rect 2950 40826 2956 40828
rect 3012 40826 3036 40828
rect 3092 40826 3116 40828
rect 3172 40826 3196 40828
rect 3252 40826 3258 40828
rect 3012 40774 3014 40826
rect 3194 40774 3196 40826
rect 2950 40772 2956 40774
rect 3012 40772 3036 40774
rect 3092 40772 3116 40774
rect 3172 40772 3196 40774
rect 3252 40772 3258 40774
rect 1306 40760 1362 40769
rect 2950 40763 3258 40772
rect 1306 40695 1362 40704
rect 2950 39740 3258 39749
rect 2950 39738 2956 39740
rect 3012 39738 3036 39740
rect 3092 39738 3116 39740
rect 3172 39738 3196 39740
rect 3252 39738 3258 39740
rect 3012 39686 3014 39738
rect 3194 39686 3196 39738
rect 2950 39684 2956 39686
rect 3012 39684 3036 39686
rect 3092 39684 3116 39686
rect 3172 39684 3196 39686
rect 3252 39684 3258 39686
rect 2950 39675 3258 39684
rect 2950 38652 3258 38661
rect 2950 38650 2956 38652
rect 3012 38650 3036 38652
rect 3092 38650 3116 38652
rect 3172 38650 3196 38652
rect 3252 38650 3258 38652
rect 3012 38598 3014 38650
rect 3194 38598 3196 38650
rect 2950 38596 2956 38598
rect 3012 38596 3036 38598
rect 3092 38596 3116 38598
rect 3172 38596 3196 38598
rect 3252 38596 3258 38598
rect 2950 38587 3258 38596
rect 1308 38344 1360 38350
rect 1306 38312 1308 38321
rect 1360 38312 1362 38321
rect 1306 38247 1362 38256
rect 2950 37564 3258 37573
rect 2950 37562 2956 37564
rect 3012 37562 3036 37564
rect 3092 37562 3116 37564
rect 3172 37562 3196 37564
rect 3252 37562 3258 37564
rect 3012 37510 3014 37562
rect 3194 37510 3196 37562
rect 2950 37508 2956 37510
rect 3012 37508 3036 37510
rect 3092 37508 3116 37510
rect 3172 37508 3196 37510
rect 3252 37508 3258 37510
rect 2950 37499 3258 37508
rect 2950 36476 3258 36485
rect 2950 36474 2956 36476
rect 3012 36474 3036 36476
rect 3092 36474 3116 36476
rect 3172 36474 3196 36476
rect 3252 36474 3258 36476
rect 3012 36422 3014 36474
rect 3194 36422 3196 36474
rect 2950 36420 2956 36422
rect 3012 36420 3036 36422
rect 3092 36420 3116 36422
rect 3172 36420 3196 36422
rect 3252 36420 3258 36422
rect 2950 36411 3258 36420
rect 1768 36168 1820 36174
rect 1768 36110 1820 36116
rect 1584 36032 1636 36038
rect 1584 35974 1636 35980
rect 1308 33516 1360 33522
rect 1308 33458 1360 33464
rect 1320 33425 1348 33458
rect 1306 33416 1362 33425
rect 1306 33351 1362 33360
rect 1596 28626 1624 35974
rect 1780 35873 1808 36110
rect 1766 35864 1822 35873
rect 1766 35799 1822 35808
rect 2950 35388 3258 35397
rect 2950 35386 2956 35388
rect 3012 35386 3036 35388
rect 3092 35386 3116 35388
rect 3172 35386 3196 35388
rect 3252 35386 3258 35388
rect 3012 35334 3014 35386
rect 3194 35334 3196 35386
rect 2950 35332 2956 35334
rect 3012 35332 3036 35334
rect 3092 35332 3116 35334
rect 3172 35332 3196 35334
rect 3252 35332 3258 35334
rect 2950 35323 3258 35332
rect 2950 34300 3258 34309
rect 2950 34298 2956 34300
rect 3012 34298 3036 34300
rect 3092 34298 3116 34300
rect 3172 34298 3196 34300
rect 3252 34298 3258 34300
rect 3012 34246 3014 34298
rect 3194 34246 3196 34298
rect 2950 34244 2956 34246
rect 3012 34244 3036 34246
rect 3092 34244 3116 34246
rect 3172 34244 3196 34246
rect 3252 34244 3258 34246
rect 2950 34235 3258 34244
rect 3424 33312 3476 33318
rect 3424 33254 3476 33260
rect 2950 33212 3258 33221
rect 2950 33210 2956 33212
rect 3012 33210 3036 33212
rect 3092 33210 3116 33212
rect 3172 33210 3196 33212
rect 3252 33210 3258 33212
rect 3012 33158 3014 33210
rect 3194 33158 3196 33210
rect 2950 33156 2956 33158
rect 3012 33156 3036 33158
rect 3092 33156 3116 33158
rect 3172 33156 3196 33158
rect 3252 33156 3258 33158
rect 2950 33147 3258 33156
rect 2950 32124 3258 32133
rect 2950 32122 2956 32124
rect 3012 32122 3036 32124
rect 3092 32122 3116 32124
rect 3172 32122 3196 32124
rect 3252 32122 3258 32124
rect 3012 32070 3014 32122
rect 3194 32070 3196 32122
rect 2950 32068 2956 32070
rect 3012 32068 3036 32070
rect 3092 32068 3116 32070
rect 3172 32068 3196 32070
rect 3252 32068 3258 32070
rect 2950 32059 3258 32068
rect 2950 31036 3258 31045
rect 2950 31034 2956 31036
rect 3012 31034 3036 31036
rect 3092 31034 3116 31036
rect 3172 31034 3196 31036
rect 3252 31034 3258 31036
rect 3012 30982 3014 31034
rect 3194 30982 3196 31034
rect 2950 30980 2956 30982
rect 3012 30980 3036 30982
rect 3092 30980 3116 30982
rect 3172 30980 3196 30982
rect 3252 30980 3258 30982
rect 2778 30968 2834 30977
rect 2950 30971 3258 30980
rect 2778 30903 2834 30912
rect 2228 29164 2280 29170
rect 2228 29106 2280 29112
rect 1584 28620 1636 28626
rect 1584 28562 1636 28568
rect 2240 28014 2268 29106
rect 2792 28014 2820 30903
rect 2950 29948 3258 29957
rect 2950 29946 2956 29948
rect 3012 29946 3036 29948
rect 3092 29946 3116 29948
rect 3172 29946 3196 29948
rect 3252 29946 3258 29948
rect 3012 29894 3014 29946
rect 3194 29894 3196 29946
rect 2950 29892 2956 29894
rect 3012 29892 3036 29894
rect 3092 29892 3116 29894
rect 3172 29892 3196 29894
rect 3252 29892 3258 29894
rect 2950 29883 3258 29892
rect 2950 28860 3258 28869
rect 2950 28858 2956 28860
rect 3012 28858 3036 28860
rect 3092 28858 3116 28860
rect 3172 28858 3196 28860
rect 3252 28858 3258 28860
rect 3012 28806 3014 28858
rect 3194 28806 3196 28858
rect 2950 28804 2956 28806
rect 3012 28804 3036 28806
rect 3092 28804 3116 28806
rect 3172 28804 3196 28806
rect 3252 28804 3258 28806
rect 2950 28795 3258 28804
rect 2870 28520 2926 28529
rect 2870 28455 2926 28464
rect 2228 28008 2280 28014
rect 2228 27950 2280 27956
rect 2780 28008 2832 28014
rect 2780 27950 2832 27956
rect 2240 26450 2268 27950
rect 2228 26444 2280 26450
rect 2228 26386 2280 26392
rect 1952 24744 2004 24750
rect 1952 24686 2004 24692
rect 1964 24614 1992 24686
rect 1952 24608 2004 24614
rect 1952 24550 2004 24556
rect 1860 24064 1912 24070
rect 1860 24006 1912 24012
rect 1768 21888 1820 21894
rect 1768 21830 1820 21836
rect 1306 21176 1362 21185
rect 1306 21111 1362 21120
rect 1320 21010 1348 21111
rect 1308 21004 1360 21010
rect 1308 20946 1360 20952
rect 1308 18828 1360 18834
rect 1308 18770 1360 18776
rect 1320 18737 1348 18770
rect 1780 18766 1808 21830
rect 1872 20942 1900 24006
rect 1964 22030 1992 24550
rect 2240 24206 2268 26386
rect 2778 26072 2834 26081
rect 2778 26007 2834 26016
rect 2688 25900 2740 25906
rect 2688 25842 2740 25848
rect 2228 24200 2280 24206
rect 2228 24142 2280 24148
rect 2320 23724 2372 23730
rect 2320 23666 2372 23672
rect 2044 23044 2096 23050
rect 2044 22986 2096 22992
rect 2056 22778 2084 22986
rect 2044 22772 2096 22778
rect 2044 22714 2096 22720
rect 1952 22024 2004 22030
rect 1952 21966 2004 21972
rect 1860 20936 1912 20942
rect 1860 20878 1912 20884
rect 2056 19446 2084 22714
rect 2136 21888 2188 21894
rect 2136 21830 2188 21836
rect 2148 21622 2176 21830
rect 2136 21616 2188 21622
rect 2136 21558 2188 21564
rect 2332 21486 2360 23666
rect 2700 22778 2728 25842
rect 2792 23322 2820 26007
rect 2884 24750 2912 28455
rect 2950 27772 3258 27781
rect 2950 27770 2956 27772
rect 3012 27770 3036 27772
rect 3092 27770 3116 27772
rect 3172 27770 3196 27772
rect 3252 27770 3258 27772
rect 3012 27718 3014 27770
rect 3194 27718 3196 27770
rect 2950 27716 2956 27718
rect 3012 27716 3036 27718
rect 3092 27716 3116 27718
rect 3172 27716 3196 27718
rect 3252 27716 3258 27718
rect 2950 27707 3258 27716
rect 3436 26994 3464 33254
rect 3528 28642 3556 43114
rect 3620 41274 3648 49778
rect 3988 41478 4016 50351
rect 4080 49638 4108 52838
rect 4160 50924 4212 50930
rect 4160 50866 4212 50872
rect 4068 49632 4120 49638
rect 4068 49574 4120 49580
rect 4066 48104 4122 48113
rect 4066 48039 4122 48048
rect 4080 46986 4108 48039
rect 4068 46980 4120 46986
rect 4068 46922 4120 46928
rect 4066 45656 4122 45665
rect 4066 45591 4068 45600
rect 4120 45591 4122 45600
rect 4068 45562 4120 45568
rect 4172 41818 4200 50866
rect 4264 50862 4292 52958
rect 4356 51066 4384 54130
rect 4448 53174 4476 56200
rect 4816 55214 4844 56200
rect 4816 55186 4936 55214
rect 4620 54188 4672 54194
rect 4620 54130 4672 54136
rect 4436 53168 4488 53174
rect 4436 53110 4488 53116
rect 4528 52012 4580 52018
rect 4528 51954 4580 51960
rect 4344 51060 4396 51066
rect 4344 51002 4396 51008
rect 4344 50924 4396 50930
rect 4344 50866 4396 50872
rect 4252 50856 4304 50862
rect 4252 50798 4304 50804
rect 4356 42362 4384 50866
rect 4540 42770 4568 51954
rect 4632 43382 4660 54130
rect 4804 52488 4856 52494
rect 4804 52430 4856 52436
rect 4712 50312 4764 50318
rect 4712 50254 4764 50260
rect 4620 43376 4672 43382
rect 4620 43318 4672 43324
rect 4528 42764 4580 42770
rect 4528 42706 4580 42712
rect 4344 42356 4396 42362
rect 4344 42298 4396 42304
rect 4160 41812 4212 41818
rect 4160 41754 4212 41760
rect 4068 41540 4120 41546
rect 4068 41482 4120 41488
rect 3976 41472 4028 41478
rect 3976 41414 4028 41420
rect 3608 41268 3660 41274
rect 3608 41210 3660 41216
rect 3608 40928 3660 40934
rect 3608 40870 3660 40876
rect 3620 31346 3648 40870
rect 3884 38208 3936 38214
rect 3884 38150 3936 38156
rect 3608 31340 3660 31346
rect 3608 31282 3660 31288
rect 3792 31272 3844 31278
rect 3792 31214 3844 31220
rect 3804 29306 3832 31214
rect 3896 29714 3924 38150
rect 3884 29708 3936 29714
rect 3884 29650 3936 29656
rect 3884 29572 3936 29578
rect 3884 29514 3936 29520
rect 3792 29300 3844 29306
rect 3792 29242 3844 29248
rect 3528 28614 3740 28642
rect 3516 28484 3568 28490
rect 3516 28426 3568 28432
rect 3424 26988 3476 26994
rect 3424 26930 3476 26936
rect 2950 26684 3258 26693
rect 2950 26682 2956 26684
rect 3012 26682 3036 26684
rect 3092 26682 3116 26684
rect 3172 26682 3196 26684
rect 3252 26682 3258 26684
rect 3012 26630 3014 26682
rect 3194 26630 3196 26682
rect 2950 26628 2956 26630
rect 3012 26628 3036 26630
rect 3092 26628 3116 26630
rect 3172 26628 3196 26630
rect 3252 26628 3258 26630
rect 2950 26619 3258 26628
rect 3528 26042 3556 28426
rect 3608 26920 3660 26926
rect 3608 26862 3660 26868
rect 3516 26036 3568 26042
rect 3516 25978 3568 25984
rect 2950 25596 3258 25605
rect 2950 25594 2956 25596
rect 3012 25594 3036 25596
rect 3092 25594 3116 25596
rect 3172 25594 3196 25596
rect 3252 25594 3258 25596
rect 3012 25542 3014 25594
rect 3194 25542 3196 25594
rect 2950 25540 2956 25542
rect 3012 25540 3036 25542
rect 3092 25540 3116 25542
rect 3172 25540 3196 25542
rect 3252 25540 3258 25542
rect 2950 25531 3258 25540
rect 2872 24744 2924 24750
rect 2872 24686 2924 24692
rect 2950 24508 3258 24517
rect 2950 24506 2956 24508
rect 3012 24506 3036 24508
rect 3092 24506 3116 24508
rect 3172 24506 3196 24508
rect 3252 24506 3258 24508
rect 3012 24454 3014 24506
rect 3194 24454 3196 24506
rect 2950 24452 2956 24454
rect 3012 24452 3036 24454
rect 3092 24452 3116 24454
rect 3172 24452 3196 24454
rect 3252 24452 3258 24454
rect 2950 24443 3258 24452
rect 3620 23866 3648 26862
rect 3712 26586 3740 28614
rect 3792 27464 3844 27470
rect 3792 27406 3844 27412
rect 3700 26580 3752 26586
rect 3700 26522 3752 26528
rect 3712 26382 3740 26522
rect 3700 26376 3752 26382
rect 3700 26318 3752 26324
rect 3712 25906 3740 26318
rect 3700 25900 3752 25906
rect 3700 25842 3752 25848
rect 3608 23860 3660 23866
rect 3608 23802 3660 23808
rect 2870 23624 2926 23633
rect 2870 23559 2926 23568
rect 2780 23316 2832 23322
rect 2780 23258 2832 23264
rect 2780 23180 2832 23186
rect 2780 23122 2832 23128
rect 2688 22772 2740 22778
rect 2688 22714 2740 22720
rect 2320 21480 2372 21486
rect 2320 21422 2372 21428
rect 2044 19440 2096 19446
rect 2044 19382 2096 19388
rect 2228 19168 2280 19174
rect 2228 19110 2280 19116
rect 1768 18760 1820 18766
rect 1306 18728 1362 18737
rect 1768 18702 1820 18708
rect 1306 18663 1362 18672
rect 1768 16992 1820 16998
rect 1768 16934 1820 16940
rect 1308 16516 1360 16522
rect 1308 16458 1360 16464
rect 1320 16289 1348 16458
rect 1306 16280 1362 16289
rect 1306 16215 1362 16224
rect 1780 13938 1808 16934
rect 2240 16590 2268 19110
rect 2332 18902 2360 21422
rect 2792 20602 2820 23122
rect 2884 21486 2912 23559
rect 2950 23420 3258 23429
rect 2950 23418 2956 23420
rect 3012 23418 3036 23420
rect 3092 23418 3116 23420
rect 3172 23418 3196 23420
rect 3252 23418 3258 23420
rect 3012 23366 3014 23418
rect 3194 23366 3196 23418
rect 2950 23364 2956 23366
rect 3012 23364 3036 23366
rect 3092 23364 3116 23366
rect 3172 23364 3196 23366
rect 3252 23364 3258 23366
rect 2950 23355 3258 23364
rect 3712 22710 3740 25842
rect 3804 25770 3832 27406
rect 3896 27402 3924 29514
rect 4080 28762 4108 41482
rect 4724 41274 4752 50254
rect 4816 41818 4844 52430
rect 4908 51950 4936 55186
rect 5184 53242 5212 56200
rect 5552 53718 5580 56200
rect 5920 54126 5948 56200
rect 5908 54120 5960 54126
rect 5908 54062 5960 54068
rect 5540 53712 5592 53718
rect 5540 53654 5592 53660
rect 5172 53236 5224 53242
rect 5172 53178 5224 53184
rect 5724 53236 5776 53242
rect 5724 53178 5776 53184
rect 5540 53032 5592 53038
rect 5540 52974 5592 52980
rect 5552 52154 5580 52974
rect 5632 52488 5684 52494
rect 5632 52430 5684 52436
rect 5540 52148 5592 52154
rect 5540 52090 5592 52096
rect 4988 52012 5040 52018
rect 4988 51954 5040 51960
rect 4896 51944 4948 51950
rect 4896 51886 4948 51892
rect 5000 43994 5028 51954
rect 5540 51332 5592 51338
rect 5540 51274 5592 51280
rect 5552 51066 5580 51274
rect 5540 51060 5592 51066
rect 5540 51002 5592 51008
rect 5644 46170 5672 52430
rect 5736 51474 5764 53178
rect 6288 53174 6316 56200
rect 6276 53168 6328 53174
rect 6276 53110 6328 53116
rect 6460 53100 6512 53106
rect 6460 53042 6512 53048
rect 5724 51468 5776 51474
rect 5724 51410 5776 51416
rect 5816 50312 5868 50318
rect 5816 50254 5868 50260
rect 5632 46164 5684 46170
rect 5632 46106 5684 46112
rect 5828 44538 5856 50254
rect 6472 45082 6500 53042
rect 6656 52562 6684 56200
rect 6828 53576 6880 53582
rect 6828 53518 6880 53524
rect 6644 52556 6696 52562
rect 6644 52498 6696 52504
rect 6736 51400 6788 51406
rect 6736 51342 6788 51348
rect 6460 45076 6512 45082
rect 6460 45018 6512 45024
rect 6644 44736 6696 44742
rect 6644 44678 6696 44684
rect 5816 44532 5868 44538
rect 5816 44474 5868 44480
rect 6656 44402 6684 44678
rect 6748 44538 6776 51342
rect 6840 50522 6868 53518
rect 7024 51474 7052 56200
rect 7392 53650 7420 56200
rect 7380 53644 7432 53650
rect 7380 53586 7432 53592
rect 7564 53508 7616 53514
rect 7564 53450 7616 53456
rect 7196 52488 7248 52494
rect 7196 52430 7248 52436
rect 7012 51468 7064 51474
rect 7012 51410 7064 51416
rect 7104 51400 7156 51406
rect 7104 51342 7156 51348
rect 6828 50516 6880 50522
rect 6828 50458 6880 50464
rect 6828 49972 6880 49978
rect 6828 49914 6880 49920
rect 6840 45490 6868 49914
rect 7116 47682 7144 51342
rect 7208 51074 7236 52430
rect 7380 52012 7432 52018
rect 7380 51954 7432 51960
rect 7208 51046 7328 51074
rect 7116 47654 7236 47682
rect 7012 45960 7064 45966
rect 7012 45902 7064 45908
rect 6828 45484 6880 45490
rect 6828 45426 6880 45432
rect 6736 44532 6788 44538
rect 6736 44474 6788 44480
rect 6552 44396 6604 44402
rect 6552 44338 6604 44344
rect 6644 44396 6696 44402
rect 6644 44338 6696 44344
rect 4988 43988 5040 43994
rect 4988 43930 5040 43936
rect 5908 42220 5960 42226
rect 5908 42162 5960 42168
rect 4804 41812 4856 41818
rect 4804 41754 4856 41760
rect 5264 41540 5316 41546
rect 5264 41482 5316 41488
rect 4712 41268 4764 41274
rect 4712 41210 4764 41216
rect 4528 41132 4580 41138
rect 4528 41074 4580 41080
rect 5080 41132 5132 41138
rect 5080 41074 5132 41080
rect 4540 32570 4568 41074
rect 5092 40934 5120 41074
rect 5080 40928 5132 40934
rect 5080 40870 5132 40876
rect 4528 32564 4580 32570
rect 4528 32506 4580 32512
rect 4988 31272 5040 31278
rect 4988 31214 5040 31220
rect 4068 28756 4120 28762
rect 4068 28698 4120 28704
rect 4068 27940 4120 27946
rect 4068 27882 4120 27888
rect 3884 27396 3936 27402
rect 3884 27338 3936 27344
rect 3792 25764 3844 25770
rect 3792 25706 3844 25712
rect 3804 24614 3832 25706
rect 4080 25498 4108 27882
rect 4804 26580 4856 26586
rect 4804 26522 4856 26528
rect 4344 25696 4396 25702
rect 4344 25638 4396 25644
rect 4068 25492 4120 25498
rect 4068 25434 4120 25440
rect 4252 25152 4304 25158
rect 4252 25094 4304 25100
rect 4264 24886 4292 25094
rect 4252 24880 4304 24886
rect 4252 24822 4304 24828
rect 4356 24750 4384 25638
rect 4816 25294 4844 26522
rect 4896 25356 4948 25362
rect 4896 25298 4948 25304
rect 4804 25288 4856 25294
rect 4804 25230 4856 25236
rect 3976 24744 4028 24750
rect 3976 24686 4028 24692
rect 4344 24744 4396 24750
rect 4344 24686 4396 24692
rect 3884 24676 3936 24682
rect 3884 24618 3936 24624
rect 3792 24608 3844 24614
rect 3792 24550 3844 24556
rect 3700 22704 3752 22710
rect 3700 22646 3752 22652
rect 2950 22332 3258 22341
rect 2950 22330 2956 22332
rect 3012 22330 3036 22332
rect 3092 22330 3116 22332
rect 3172 22330 3196 22332
rect 3252 22330 3258 22332
rect 3012 22278 3014 22330
rect 3194 22278 3196 22330
rect 2950 22276 2956 22278
rect 3012 22276 3036 22278
rect 3092 22276 3116 22278
rect 3172 22276 3196 22278
rect 3252 22276 3258 22278
rect 2950 22267 3258 22276
rect 3332 22024 3384 22030
rect 3332 21966 3384 21972
rect 3344 21690 3372 21966
rect 3332 21684 3384 21690
rect 3332 21626 3384 21632
rect 2872 21480 2924 21486
rect 2872 21422 2924 21428
rect 2950 21244 3258 21253
rect 2950 21242 2956 21244
rect 3012 21242 3036 21244
rect 3092 21242 3116 21244
rect 3172 21242 3196 21244
rect 3252 21242 3258 21244
rect 3012 21190 3014 21242
rect 3194 21190 3196 21242
rect 2950 21188 2956 21190
rect 3012 21188 3036 21190
rect 3092 21188 3116 21190
rect 3172 21188 3196 21190
rect 3252 21188 3258 21190
rect 2950 21179 3258 21188
rect 3896 20602 3924 24618
rect 3988 24206 4016 24686
rect 3976 24200 4028 24206
rect 3976 24142 4028 24148
rect 3988 23662 4016 24142
rect 4252 24132 4304 24138
rect 4252 24074 4304 24080
rect 4264 23866 4292 24074
rect 4252 23860 4304 23866
rect 4252 23802 4304 23808
rect 3976 23656 4028 23662
rect 3976 23598 4028 23604
rect 3988 22098 4016 23598
rect 4356 23118 4384 24686
rect 4816 24410 4844 25230
rect 4804 24404 4856 24410
rect 4804 24346 4856 24352
rect 4344 23112 4396 23118
rect 4344 23054 4396 23060
rect 4436 22976 4488 22982
rect 4436 22918 4488 22924
rect 3976 22092 4028 22098
rect 3976 22034 4028 22040
rect 4160 22092 4212 22098
rect 4160 22034 4212 22040
rect 4172 21010 4200 22034
rect 4448 21010 4476 22918
rect 4160 21004 4212 21010
rect 4160 20946 4212 20952
rect 4436 21004 4488 21010
rect 4436 20946 4488 20952
rect 2780 20596 2832 20602
rect 2780 20538 2832 20544
rect 3884 20596 3936 20602
rect 3884 20538 3936 20544
rect 2950 20156 3258 20165
rect 2950 20154 2956 20156
rect 3012 20154 3036 20156
rect 3092 20154 3116 20156
rect 3172 20154 3196 20156
rect 3252 20154 3258 20156
rect 3012 20102 3014 20154
rect 3194 20102 3196 20154
rect 2950 20100 2956 20102
rect 3012 20100 3036 20102
rect 3092 20100 3116 20102
rect 3172 20100 3196 20102
rect 3252 20100 3258 20102
rect 2950 20091 3258 20100
rect 4172 19922 4200 20946
rect 4252 20460 4304 20466
rect 4252 20402 4304 20408
rect 4160 19916 4212 19922
rect 4160 19858 4212 19864
rect 2950 19068 3258 19077
rect 2950 19066 2956 19068
rect 3012 19066 3036 19068
rect 3092 19066 3116 19068
rect 3172 19066 3196 19068
rect 3252 19066 3258 19068
rect 3012 19014 3014 19066
rect 3194 19014 3196 19066
rect 2950 19012 2956 19014
rect 3012 19012 3036 19014
rect 3092 19012 3116 19014
rect 3172 19012 3196 19014
rect 3252 19012 3258 19014
rect 2950 19003 3258 19012
rect 2320 18896 2372 18902
rect 2320 18838 2372 18844
rect 2332 17270 2360 18838
rect 4264 18426 4292 20402
rect 4252 18420 4304 18426
rect 4252 18362 4304 18368
rect 2950 17980 3258 17989
rect 2950 17978 2956 17980
rect 3012 17978 3036 17980
rect 3092 17978 3116 17980
rect 3172 17978 3196 17980
rect 3252 17978 3258 17980
rect 3012 17926 3014 17978
rect 3194 17926 3196 17978
rect 2950 17924 2956 17926
rect 3012 17924 3036 17926
rect 3092 17924 3116 17926
rect 3172 17924 3196 17926
rect 3252 17924 3258 17926
rect 2950 17915 3258 17924
rect 4804 17672 4856 17678
rect 4804 17614 4856 17620
rect 2320 17264 2372 17270
rect 2320 17206 2372 17212
rect 2950 16892 3258 16901
rect 2950 16890 2956 16892
rect 3012 16890 3036 16892
rect 3092 16890 3116 16892
rect 3172 16890 3196 16892
rect 3252 16890 3258 16892
rect 3012 16838 3014 16890
rect 3194 16838 3196 16890
rect 2950 16836 2956 16838
rect 3012 16836 3036 16838
rect 3092 16836 3116 16838
rect 3172 16836 3196 16838
rect 3252 16836 3258 16838
rect 2950 16827 3258 16836
rect 4816 16658 4844 17614
rect 4804 16652 4856 16658
rect 4804 16594 4856 16600
rect 2228 16584 2280 16590
rect 2228 16526 2280 16532
rect 2950 15804 3258 15813
rect 2950 15802 2956 15804
rect 3012 15802 3036 15804
rect 3092 15802 3116 15804
rect 3172 15802 3196 15804
rect 3252 15802 3258 15804
rect 3012 15750 3014 15802
rect 3194 15750 3196 15802
rect 2950 15748 2956 15750
rect 3012 15748 3036 15750
rect 3092 15748 3116 15750
rect 3172 15748 3196 15750
rect 3252 15748 3258 15750
rect 2950 15739 3258 15748
rect 2950 14716 3258 14725
rect 2950 14714 2956 14716
rect 3012 14714 3036 14716
rect 3092 14714 3116 14716
rect 3172 14714 3196 14716
rect 3252 14714 3258 14716
rect 3012 14662 3014 14714
rect 3194 14662 3196 14714
rect 2950 14660 2956 14662
rect 3012 14660 3036 14662
rect 3092 14660 3116 14662
rect 3172 14660 3196 14662
rect 3252 14660 3258 14662
rect 2950 14651 3258 14660
rect 1768 13932 1820 13938
rect 1768 13874 1820 13880
rect 1308 13864 1360 13870
rect 1306 13832 1308 13841
rect 1360 13832 1362 13841
rect 1306 13767 1362 13776
rect 2950 13628 3258 13637
rect 2950 13626 2956 13628
rect 3012 13626 3036 13628
rect 3092 13626 3116 13628
rect 3172 13626 3196 13628
rect 3252 13626 3258 13628
rect 3012 13574 3014 13626
rect 3194 13574 3196 13626
rect 2950 13572 2956 13574
rect 3012 13572 3036 13574
rect 3092 13572 3116 13574
rect 3172 13572 3196 13574
rect 3252 13572 3258 13574
rect 2950 13563 3258 13572
rect 2950 12540 3258 12549
rect 2950 12538 2956 12540
rect 3012 12538 3036 12540
rect 3092 12538 3116 12540
rect 3172 12538 3196 12540
rect 3252 12538 3258 12540
rect 3012 12486 3014 12538
rect 3194 12486 3196 12538
rect 2950 12484 2956 12486
rect 3012 12484 3036 12486
rect 3092 12484 3116 12486
rect 3172 12484 3196 12486
rect 3252 12484 3258 12486
rect 2950 12475 3258 12484
rect 1860 12436 1912 12442
rect 1860 12378 1912 12384
rect 1676 3528 1728 3534
rect 1676 3470 1728 3476
rect 1492 2848 1544 2854
rect 1492 2790 1544 2796
rect 1504 2446 1532 2790
rect 1492 2440 1544 2446
rect 1492 2382 1544 2388
rect 1688 800 1716 3470
rect 1872 2650 1900 12378
rect 2780 12096 2832 12102
rect 2780 12038 2832 12044
rect 2792 11393 2820 12038
rect 2950 11452 3258 11461
rect 2950 11450 2956 11452
rect 3012 11450 3036 11452
rect 3092 11450 3116 11452
rect 3172 11450 3196 11452
rect 3252 11450 3258 11452
rect 3012 11398 3014 11450
rect 3194 11398 3196 11450
rect 2950 11396 2956 11398
rect 3012 11396 3036 11398
rect 3092 11396 3116 11398
rect 3172 11396 3196 11398
rect 3252 11396 3258 11398
rect 2778 11384 2834 11393
rect 2950 11387 3258 11396
rect 2778 11319 2834 11328
rect 2950 10364 3258 10373
rect 2950 10362 2956 10364
rect 3012 10362 3036 10364
rect 3092 10362 3116 10364
rect 3172 10362 3196 10364
rect 3252 10362 3258 10364
rect 3012 10310 3014 10362
rect 3194 10310 3196 10362
rect 2950 10308 2956 10310
rect 3012 10308 3036 10310
rect 3092 10308 3116 10310
rect 3172 10308 3196 10310
rect 3252 10308 3258 10310
rect 2950 10299 3258 10308
rect 2872 9512 2924 9518
rect 2872 9454 2924 9460
rect 2884 8945 2912 9454
rect 2950 9276 3258 9285
rect 2950 9274 2956 9276
rect 3012 9274 3036 9276
rect 3092 9274 3116 9276
rect 3172 9274 3196 9276
rect 3252 9274 3258 9276
rect 3012 9222 3014 9274
rect 3194 9222 3196 9274
rect 2950 9220 2956 9222
rect 3012 9220 3036 9222
rect 3092 9220 3116 9222
rect 3172 9220 3196 9222
rect 3252 9220 3258 9222
rect 2950 9211 3258 9220
rect 2870 8936 2926 8945
rect 2870 8871 2926 8880
rect 2780 8424 2832 8430
rect 2780 8366 2832 8372
rect 2688 5636 2740 5642
rect 2688 5578 2740 5584
rect 2596 4276 2648 4282
rect 2596 4218 2648 4224
rect 2044 3392 2096 3398
rect 2044 3334 2096 3340
rect 2056 3058 2084 3334
rect 2044 3052 2096 3058
rect 2044 2994 2096 3000
rect 1860 2644 1912 2650
rect 1860 2586 1912 2592
rect 2056 800 2084 2994
rect 2608 2650 2636 4218
rect 2700 3194 2728 5578
rect 2792 4010 2820 8366
rect 2950 8188 3258 8197
rect 2950 8186 2956 8188
rect 3012 8186 3036 8188
rect 3092 8186 3116 8188
rect 3172 8186 3196 8188
rect 3252 8186 3258 8188
rect 3012 8134 3014 8186
rect 3194 8134 3196 8186
rect 2950 8132 2956 8134
rect 3012 8132 3036 8134
rect 3092 8132 3116 8134
rect 3172 8132 3196 8134
rect 3252 8132 3258 8134
rect 2950 8123 3258 8132
rect 2950 7100 3258 7109
rect 2950 7098 2956 7100
rect 3012 7098 3036 7100
rect 3092 7098 3116 7100
rect 3172 7098 3196 7100
rect 3252 7098 3258 7100
rect 3012 7046 3014 7098
rect 3194 7046 3196 7098
rect 2950 7044 2956 7046
rect 3012 7044 3036 7046
rect 3092 7044 3116 7046
rect 3172 7044 3196 7046
rect 3252 7044 3258 7046
rect 2950 7035 3258 7044
rect 4908 6914 4936 25298
rect 5000 25294 5028 31214
rect 5092 29306 5120 40870
rect 5172 39432 5224 39438
rect 5172 39374 5224 39380
rect 5184 38418 5212 39374
rect 5172 38412 5224 38418
rect 5172 38354 5224 38360
rect 5276 30598 5304 41482
rect 5920 39642 5948 42162
rect 6460 41812 6512 41818
rect 6460 41754 6512 41760
rect 6472 40526 6500 41754
rect 6460 40520 6512 40526
rect 6460 40462 6512 40468
rect 5908 39636 5960 39642
rect 5908 39578 5960 39584
rect 6472 39506 6500 40462
rect 6460 39500 6512 39506
rect 6460 39442 6512 39448
rect 5448 39364 5500 39370
rect 5448 39306 5500 39312
rect 5460 39098 5488 39306
rect 6460 39296 6512 39302
rect 6460 39238 6512 39244
rect 5448 39092 5500 39098
rect 5448 39034 5500 39040
rect 5816 39024 5868 39030
rect 5816 38966 5868 38972
rect 5448 38956 5500 38962
rect 5448 38898 5500 38904
rect 5460 32570 5488 38898
rect 5632 37324 5684 37330
rect 5632 37266 5684 37272
rect 5644 37126 5672 37266
rect 5828 37126 5856 38966
rect 6092 38548 6144 38554
rect 6092 38490 6144 38496
rect 6000 38276 6052 38282
rect 6000 38218 6052 38224
rect 6012 38010 6040 38218
rect 6000 38004 6052 38010
rect 6000 37946 6052 37952
rect 5632 37120 5684 37126
rect 5632 37062 5684 37068
rect 5816 37120 5868 37126
rect 5816 37062 5868 37068
rect 5644 36242 5672 37062
rect 5632 36236 5684 36242
rect 5632 36178 5684 36184
rect 5644 35494 5672 36178
rect 6104 35834 6132 38490
rect 6472 38282 6500 39238
rect 6564 39098 6592 44338
rect 6552 39092 6604 39098
rect 6552 39034 6604 39040
rect 6460 38276 6512 38282
rect 6460 38218 6512 38224
rect 6472 37466 6500 38218
rect 6656 38010 6684 44338
rect 6736 42560 6788 42566
rect 6736 42502 6788 42508
rect 6748 41698 6776 42502
rect 6840 42226 6868 45426
rect 6828 42220 6880 42226
rect 6828 42162 6880 42168
rect 6840 41818 6868 42162
rect 6828 41812 6880 41818
rect 6828 41754 6880 41760
rect 6748 41670 6868 41698
rect 6840 41414 6868 41670
rect 6748 41386 6868 41414
rect 6644 38004 6696 38010
rect 6644 37946 6696 37952
rect 6552 37800 6604 37806
rect 6552 37742 6604 37748
rect 6460 37460 6512 37466
rect 6460 37402 6512 37408
rect 6472 37194 6500 37402
rect 6564 37330 6592 37742
rect 6644 37392 6696 37398
rect 6644 37334 6696 37340
rect 6552 37324 6604 37330
rect 6552 37266 6604 37272
rect 6460 37188 6512 37194
rect 6460 37130 6512 37136
rect 6472 36922 6500 37130
rect 6460 36916 6512 36922
rect 6460 36858 6512 36864
rect 6092 35828 6144 35834
rect 6092 35770 6144 35776
rect 5632 35488 5684 35494
rect 5632 35430 5684 35436
rect 5644 35086 5672 35430
rect 6104 35154 6132 35770
rect 6552 35488 6604 35494
rect 6552 35430 6604 35436
rect 6564 35154 6592 35430
rect 6656 35290 6684 37334
rect 6644 35284 6696 35290
rect 6644 35226 6696 35232
rect 6092 35148 6144 35154
rect 6092 35090 6144 35096
rect 6552 35148 6604 35154
rect 6552 35090 6604 35096
rect 5632 35080 5684 35086
rect 5632 35022 5684 35028
rect 5540 33992 5592 33998
rect 5644 33946 5672 35022
rect 5816 34944 5868 34950
rect 5816 34886 5868 34892
rect 5828 34066 5856 34886
rect 6000 34468 6052 34474
rect 6000 34410 6052 34416
rect 5816 34060 5868 34066
rect 5816 34002 5868 34008
rect 5592 33940 5672 33946
rect 5540 33934 5672 33940
rect 5552 33918 5672 33934
rect 5540 33448 5592 33454
rect 5540 33390 5592 33396
rect 5552 32570 5580 33390
rect 5644 32978 5672 33918
rect 5632 32972 5684 32978
rect 5632 32914 5684 32920
rect 5448 32564 5500 32570
rect 5448 32506 5500 32512
rect 5540 32564 5592 32570
rect 5540 32506 5592 32512
rect 5540 32428 5592 32434
rect 5540 32370 5592 32376
rect 5264 30592 5316 30598
rect 5264 30534 5316 30540
rect 5080 29300 5132 29306
rect 5080 29242 5132 29248
rect 5172 26920 5224 26926
rect 5172 26862 5224 26868
rect 5184 26314 5212 26862
rect 5172 26308 5224 26314
rect 5172 26250 5224 26256
rect 4988 25288 5040 25294
rect 4988 25230 5040 25236
rect 5000 16574 5028 25230
rect 5080 17604 5132 17610
rect 5080 17546 5132 17552
rect 5092 17338 5120 17546
rect 5080 17332 5132 17338
rect 5080 17274 5132 17280
rect 5000 16546 5120 16574
rect 4988 12844 5040 12850
rect 4988 12786 5040 12792
rect 4816 6886 4936 6914
rect 3056 6724 3108 6730
rect 3056 6666 3108 6672
rect 3068 6497 3096 6666
rect 3054 6488 3110 6497
rect 3054 6423 3110 6432
rect 2950 6012 3258 6021
rect 2950 6010 2956 6012
rect 3012 6010 3036 6012
rect 3092 6010 3116 6012
rect 3172 6010 3196 6012
rect 3252 6010 3258 6012
rect 3012 5958 3014 6010
rect 3194 5958 3196 6010
rect 2950 5956 2956 5958
rect 3012 5956 3036 5958
rect 3092 5956 3116 5958
rect 3172 5956 3196 5958
rect 3252 5956 3258 5958
rect 2950 5947 3258 5956
rect 2950 4924 3258 4933
rect 2950 4922 2956 4924
rect 3012 4922 3036 4924
rect 3092 4922 3116 4924
rect 3172 4922 3196 4924
rect 3252 4922 3258 4924
rect 3012 4870 3014 4922
rect 3194 4870 3196 4922
rect 2950 4868 2956 4870
rect 3012 4868 3036 4870
rect 3092 4868 3116 4870
rect 3172 4868 3196 4870
rect 3252 4868 3258 4870
rect 2950 4859 3258 4868
rect 2872 4072 2924 4078
rect 2870 4040 2872 4049
rect 2924 4040 2926 4049
rect 2780 4004 2832 4010
rect 2870 3975 2926 3984
rect 2780 3946 2832 3952
rect 2872 3936 2924 3942
rect 2872 3878 2924 3884
rect 2780 3392 2832 3398
rect 2780 3334 2832 3340
rect 2688 3188 2740 3194
rect 2688 3130 2740 3136
rect 2792 3058 2820 3334
rect 2780 3052 2832 3058
rect 2780 2994 2832 3000
rect 2596 2644 2648 2650
rect 2596 2586 2648 2592
rect 2320 2440 2372 2446
rect 2372 2400 2452 2428
rect 2320 2382 2372 2388
rect 2424 800 2452 2400
rect 2792 800 2820 2994
rect 2884 1601 2912 3878
rect 2950 3836 3258 3845
rect 2950 3834 2956 3836
rect 3012 3834 3036 3836
rect 3092 3834 3116 3836
rect 3172 3834 3196 3836
rect 3252 3834 3258 3836
rect 3012 3782 3014 3834
rect 3194 3782 3196 3834
rect 2950 3780 2956 3782
rect 3012 3780 3036 3782
rect 3092 3780 3116 3782
rect 3172 3780 3196 3782
rect 3252 3780 3258 3782
rect 2950 3771 3258 3780
rect 3332 3460 3384 3466
rect 3332 3402 3384 3408
rect 3344 2990 3372 3402
rect 3516 3392 3568 3398
rect 3516 3334 3568 3340
rect 3884 3392 3936 3398
rect 3884 3334 3936 3340
rect 3332 2984 3384 2990
rect 3332 2926 3384 2932
rect 2950 2748 3258 2757
rect 2950 2746 2956 2748
rect 3012 2746 3036 2748
rect 3092 2746 3116 2748
rect 3172 2746 3196 2748
rect 3252 2746 3258 2748
rect 3012 2694 3014 2746
rect 3194 2694 3196 2746
rect 2950 2692 2956 2694
rect 3012 2692 3036 2694
rect 3092 2692 3116 2694
rect 3172 2692 3196 2694
rect 3252 2692 3258 2694
rect 2950 2683 3258 2692
rect 3344 2122 3372 2926
rect 3528 2446 3556 3334
rect 3516 2440 3568 2446
rect 3516 2382 3568 2388
rect 3160 2094 3372 2122
rect 2870 1592 2926 1601
rect 2870 1527 2926 1536
rect 3160 800 3188 2094
rect 3528 800 3556 2382
rect 3896 2378 3924 3334
rect 4252 2848 4304 2854
rect 4252 2790 4304 2796
rect 4264 2446 4292 2790
rect 4816 2650 4844 6886
rect 4896 3392 4948 3398
rect 4896 3334 4948 3340
rect 4804 2644 4856 2650
rect 4804 2586 4856 2592
rect 4252 2440 4304 2446
rect 4252 2382 4304 2388
rect 4620 2440 4672 2446
rect 4620 2382 4672 2388
rect 4908 2394 4936 3334
rect 5000 2514 5028 12786
rect 5092 4078 5120 16546
rect 5184 12102 5212 26250
rect 5552 17882 5580 32370
rect 5724 28484 5776 28490
rect 5724 28426 5776 28432
rect 5736 27878 5764 28426
rect 5724 27872 5776 27878
rect 5724 27814 5776 27820
rect 5632 22228 5684 22234
rect 5632 22170 5684 22176
rect 5644 21146 5672 22170
rect 5632 21140 5684 21146
rect 5632 21082 5684 21088
rect 5540 17876 5592 17882
rect 5540 17818 5592 17824
rect 5264 13864 5316 13870
rect 5264 13806 5316 13812
rect 5172 12096 5224 12102
rect 5172 12038 5224 12044
rect 5276 8634 5304 13806
rect 5736 9518 5764 27814
rect 5908 23724 5960 23730
rect 5908 23666 5960 23672
rect 5816 22432 5868 22438
rect 5816 22374 5868 22380
rect 5828 21298 5856 22374
rect 5920 22098 5948 23666
rect 5908 22092 5960 22098
rect 5908 22034 5960 22040
rect 5920 21486 5948 22034
rect 5908 21480 5960 21486
rect 5908 21422 5960 21428
rect 5828 21270 5948 21298
rect 5920 20806 5948 21270
rect 5908 20800 5960 20806
rect 5908 20742 5960 20748
rect 5920 18834 5948 20742
rect 5908 18828 5960 18834
rect 5908 18770 5960 18776
rect 5816 17876 5868 17882
rect 5816 17818 5868 17824
rect 5828 17066 5856 17818
rect 5816 17060 5868 17066
rect 5816 17002 5868 17008
rect 5724 9512 5776 9518
rect 5724 9454 5776 9460
rect 5632 8832 5684 8838
rect 5632 8774 5684 8780
rect 5264 8628 5316 8634
rect 5264 8570 5316 8576
rect 5540 6316 5592 6322
rect 5540 6258 5592 6264
rect 5172 5568 5224 5574
rect 5172 5510 5224 5516
rect 5080 4072 5132 4078
rect 5080 4014 5132 4020
rect 5184 3194 5212 5510
rect 5552 3738 5580 6258
rect 5540 3732 5592 3738
rect 5540 3674 5592 3680
rect 5644 3670 5672 8774
rect 5632 3664 5684 3670
rect 5632 3606 5684 3612
rect 5172 3188 5224 3194
rect 5172 3130 5224 3136
rect 5356 3052 5408 3058
rect 5356 2994 5408 3000
rect 5724 3052 5776 3058
rect 5724 2994 5776 3000
rect 4988 2508 5040 2514
rect 4988 2450 5040 2456
rect 3884 2372 3936 2378
rect 3884 2314 3936 2320
rect 3896 800 3924 2314
rect 4264 800 4292 2382
rect 4632 800 4660 2382
rect 4908 2366 5028 2394
rect 5000 800 5028 2366
rect 5368 800 5396 2994
rect 5736 2378 5764 2994
rect 5828 2922 5856 17002
rect 5908 16992 5960 16998
rect 5908 16934 5960 16940
rect 5920 16658 5948 16934
rect 5908 16652 5960 16658
rect 5908 16594 5960 16600
rect 5908 11824 5960 11830
rect 5908 11766 5960 11772
rect 5920 3194 5948 11766
rect 6012 3738 6040 34410
rect 6276 32972 6328 32978
rect 6276 32914 6328 32920
rect 6288 32434 6316 32914
rect 6276 32428 6328 32434
rect 6276 32370 6328 32376
rect 6288 31890 6316 32370
rect 6656 32366 6684 35226
rect 6644 32360 6696 32366
rect 6644 32302 6696 32308
rect 6276 31884 6328 31890
rect 6276 31826 6328 31832
rect 6748 31278 6776 41386
rect 7024 40186 7052 45902
rect 7104 44736 7156 44742
rect 7104 44678 7156 44684
rect 7012 40180 7064 40186
rect 7012 40122 7064 40128
rect 7116 40066 7144 44678
rect 7208 44538 7236 47654
rect 7300 44946 7328 51046
rect 7288 44940 7340 44946
rect 7288 44882 7340 44888
rect 7196 44532 7248 44538
rect 7196 44474 7248 44480
rect 7392 44266 7420 51954
rect 7472 50856 7524 50862
rect 7472 50798 7524 50804
rect 7484 46714 7512 50798
rect 7472 46708 7524 46714
rect 7472 46650 7524 46656
rect 7576 44470 7604 53450
rect 7760 52562 7788 56200
rect 7852 54262 7880 56222
rect 8036 56114 8064 56222
rect 8114 56200 8170 57000
rect 8482 56200 8538 57000
rect 8850 56200 8906 57000
rect 9218 56200 9274 57000
rect 9586 56200 9642 57000
rect 9954 56200 10010 57000
rect 10322 56200 10378 57000
rect 10690 56200 10746 57000
rect 11058 56200 11114 57000
rect 11426 56200 11482 57000
rect 11794 56200 11850 57000
rect 12162 56200 12218 57000
rect 12530 56200 12586 57000
rect 12898 56200 12954 57000
rect 13266 56200 13322 57000
rect 13634 56200 13690 57000
rect 14002 56200 14058 57000
rect 14370 56200 14426 57000
rect 14738 56200 14794 57000
rect 15106 56200 15162 57000
rect 15474 56200 15530 57000
rect 15842 56200 15898 57000
rect 16210 56200 16266 57000
rect 16578 56200 16634 57000
rect 16946 56200 17002 57000
rect 17314 56200 17370 57000
rect 17682 56200 17738 57000
rect 18050 56200 18106 57000
rect 18156 56222 18368 56250
rect 8128 56114 8156 56200
rect 8036 56086 8156 56114
rect 7950 54428 8258 54437
rect 7950 54426 7956 54428
rect 8012 54426 8036 54428
rect 8092 54426 8116 54428
rect 8172 54426 8196 54428
rect 8252 54426 8258 54428
rect 8012 54374 8014 54426
rect 8194 54374 8196 54426
rect 7950 54372 7956 54374
rect 8012 54372 8036 54374
rect 8092 54372 8116 54374
rect 8172 54372 8196 54374
rect 8252 54372 8258 54374
rect 7950 54363 8258 54372
rect 7840 54256 7892 54262
rect 7840 54198 7892 54204
rect 7950 53340 8258 53349
rect 7950 53338 7956 53340
rect 8012 53338 8036 53340
rect 8092 53338 8116 53340
rect 8172 53338 8196 53340
rect 8252 53338 8258 53340
rect 8012 53286 8014 53338
rect 8194 53286 8196 53338
rect 7950 53284 7956 53286
rect 8012 53284 8036 53286
rect 8092 53284 8116 53286
rect 8172 53284 8196 53286
rect 8252 53284 8258 53286
rect 7950 53275 8258 53284
rect 7748 52556 7800 52562
rect 7748 52498 7800 52504
rect 7950 52252 8258 52261
rect 7950 52250 7956 52252
rect 8012 52250 8036 52252
rect 8092 52250 8116 52252
rect 8172 52250 8196 52252
rect 8252 52250 8258 52252
rect 8012 52198 8014 52250
rect 8194 52198 8196 52250
rect 7950 52196 7956 52198
rect 8012 52196 8036 52198
rect 8092 52196 8116 52198
rect 8172 52196 8196 52198
rect 8252 52196 8258 52198
rect 7950 52187 8258 52196
rect 8496 51950 8524 56200
rect 8864 53650 8892 56200
rect 8852 53644 8904 53650
rect 8852 53586 8904 53592
rect 9128 53576 9180 53582
rect 9128 53518 9180 53524
rect 8484 51944 8536 51950
rect 8484 51886 8536 51892
rect 7950 51164 8258 51173
rect 7950 51162 7956 51164
rect 8012 51162 8036 51164
rect 8092 51162 8116 51164
rect 8172 51162 8196 51164
rect 8252 51162 8258 51164
rect 8012 51110 8014 51162
rect 8194 51110 8196 51162
rect 7950 51108 7956 51110
rect 8012 51108 8036 51110
rect 8092 51108 8116 51110
rect 8172 51108 8196 51110
rect 8252 51108 8258 51110
rect 7950 51099 8258 51108
rect 7656 50924 7708 50930
rect 7656 50866 7708 50872
rect 7668 46102 7696 50866
rect 9140 50522 9168 53518
rect 9232 53174 9260 56200
rect 9600 53564 9628 56200
rect 9968 54330 9996 56200
rect 10336 55214 10364 56200
rect 10336 55186 10456 55214
rect 9956 54324 10008 54330
rect 9956 54266 10008 54272
rect 9956 54188 10008 54194
rect 9956 54130 10008 54136
rect 9600 53536 9720 53564
rect 9220 53168 9272 53174
rect 9220 53110 9272 53116
rect 9588 52964 9640 52970
rect 9588 52906 9640 52912
rect 9220 52080 9272 52086
rect 9220 52022 9272 52028
rect 9128 50516 9180 50522
rect 9128 50458 9180 50464
rect 8392 50312 8444 50318
rect 8392 50254 8444 50260
rect 7950 50076 8258 50085
rect 7950 50074 7956 50076
rect 8012 50074 8036 50076
rect 8092 50074 8116 50076
rect 8172 50074 8196 50076
rect 8252 50074 8258 50076
rect 8012 50022 8014 50074
rect 8194 50022 8196 50074
rect 7950 50020 7956 50022
rect 8012 50020 8036 50022
rect 8092 50020 8116 50022
rect 8172 50020 8196 50022
rect 8252 50020 8258 50022
rect 7950 50011 8258 50020
rect 7840 49836 7892 49842
rect 7840 49778 7892 49784
rect 7656 46096 7708 46102
rect 7656 46038 7708 46044
rect 7656 44872 7708 44878
rect 7656 44814 7708 44820
rect 7564 44464 7616 44470
rect 7564 44406 7616 44412
rect 7380 44260 7432 44266
rect 7380 44202 7432 44208
rect 7668 43466 7696 44814
rect 7748 44396 7800 44402
rect 7748 44338 7800 44344
rect 7760 44198 7788 44338
rect 7748 44192 7800 44198
rect 7748 44134 7800 44140
rect 7576 43438 7696 43466
rect 7472 43104 7524 43110
rect 7472 43046 7524 43052
rect 7288 41676 7340 41682
rect 7288 41618 7340 41624
rect 7300 40730 7328 41618
rect 7288 40724 7340 40730
rect 7288 40666 7340 40672
rect 7380 40588 7432 40594
rect 7380 40530 7432 40536
rect 6932 40038 7144 40066
rect 6828 38752 6880 38758
rect 6828 38694 6880 38700
rect 6840 37942 6868 38694
rect 6828 37936 6880 37942
rect 6828 37878 6880 37884
rect 6932 37466 6960 40038
rect 7392 39642 7420 40530
rect 7380 39636 7432 39642
rect 7380 39578 7432 39584
rect 7012 38276 7064 38282
rect 7012 38218 7064 38224
rect 6920 37460 6972 37466
rect 6920 37402 6972 37408
rect 6828 36100 6880 36106
rect 6828 36042 6880 36048
rect 6840 35834 6868 36042
rect 6828 35828 6880 35834
rect 6828 35770 6880 35776
rect 6932 34490 6960 37402
rect 7024 36378 7052 38218
rect 7196 37800 7248 37806
rect 7196 37742 7248 37748
rect 7208 36582 7236 37742
rect 7288 36916 7340 36922
rect 7288 36858 7340 36864
rect 7196 36576 7248 36582
rect 7196 36518 7248 36524
rect 7012 36372 7064 36378
rect 7012 36314 7064 36320
rect 7024 35562 7052 36314
rect 7208 36038 7236 36518
rect 7300 36378 7328 36858
rect 7288 36372 7340 36378
rect 7288 36314 7340 36320
rect 7300 36106 7328 36314
rect 7288 36100 7340 36106
rect 7288 36042 7340 36048
rect 7196 36032 7248 36038
rect 7196 35974 7248 35980
rect 7012 35556 7064 35562
rect 7012 35498 7064 35504
rect 7024 35170 7052 35498
rect 7024 35142 7144 35170
rect 6840 34474 6960 34490
rect 6828 34468 6960 34474
rect 6880 34462 6960 34468
rect 6828 34410 6880 34416
rect 7116 34066 7144 35142
rect 7104 34060 7156 34066
rect 7104 34002 7156 34008
rect 6920 33992 6972 33998
rect 6920 33934 6972 33940
rect 6932 32978 6960 33934
rect 6920 32972 6972 32978
rect 6920 32914 6972 32920
rect 6932 32366 6960 32914
rect 6920 32360 6972 32366
rect 6920 32302 6972 32308
rect 6736 31272 6788 31278
rect 6736 31214 6788 31220
rect 7208 31210 7236 35974
rect 7300 35766 7328 36042
rect 7484 35986 7512 43046
rect 7576 38554 7604 43438
rect 7656 43308 7708 43314
rect 7656 43250 7708 43256
rect 7564 38548 7616 38554
rect 7564 38490 7616 38496
rect 7668 36378 7696 43250
rect 7760 41414 7788 44134
rect 7852 43450 7880 49778
rect 7950 48988 8258 48997
rect 7950 48986 7956 48988
rect 8012 48986 8036 48988
rect 8092 48986 8116 48988
rect 8172 48986 8196 48988
rect 8252 48986 8258 48988
rect 8012 48934 8014 48986
rect 8194 48934 8196 48986
rect 7950 48932 7956 48934
rect 8012 48932 8036 48934
rect 8092 48932 8116 48934
rect 8172 48932 8196 48934
rect 8252 48932 8258 48934
rect 7950 48923 8258 48932
rect 7950 47900 8258 47909
rect 7950 47898 7956 47900
rect 8012 47898 8036 47900
rect 8092 47898 8116 47900
rect 8172 47898 8196 47900
rect 8252 47898 8258 47900
rect 8012 47846 8014 47898
rect 8194 47846 8196 47898
rect 7950 47844 7956 47846
rect 8012 47844 8036 47846
rect 8092 47844 8116 47846
rect 8172 47844 8196 47846
rect 8252 47844 8258 47846
rect 7950 47835 8258 47844
rect 7950 46812 8258 46821
rect 7950 46810 7956 46812
rect 8012 46810 8036 46812
rect 8092 46810 8116 46812
rect 8172 46810 8196 46812
rect 8252 46810 8258 46812
rect 8012 46758 8014 46810
rect 8194 46758 8196 46810
rect 7950 46756 7956 46758
rect 8012 46756 8036 46758
rect 8092 46756 8116 46758
rect 8172 46756 8196 46758
rect 8252 46756 8258 46758
rect 7950 46747 8258 46756
rect 7950 45724 8258 45733
rect 7950 45722 7956 45724
rect 8012 45722 8036 45724
rect 8092 45722 8116 45724
rect 8172 45722 8196 45724
rect 8252 45722 8258 45724
rect 8012 45670 8014 45722
rect 8194 45670 8196 45722
rect 7950 45668 7956 45670
rect 8012 45668 8036 45670
rect 8092 45668 8116 45670
rect 8172 45668 8196 45670
rect 8252 45668 8258 45670
rect 7950 45659 8258 45668
rect 7950 44636 8258 44645
rect 7950 44634 7956 44636
rect 8012 44634 8036 44636
rect 8092 44634 8116 44636
rect 8172 44634 8196 44636
rect 8252 44634 8258 44636
rect 8012 44582 8014 44634
rect 8194 44582 8196 44634
rect 7950 44580 7956 44582
rect 8012 44580 8036 44582
rect 8092 44580 8116 44582
rect 8172 44580 8196 44582
rect 8252 44580 8258 44582
rect 7950 44571 8258 44580
rect 8404 43994 8432 50254
rect 8484 49904 8536 49910
rect 8484 49846 8536 49852
rect 8392 43988 8444 43994
rect 8392 43930 8444 43936
rect 7950 43548 8258 43557
rect 7950 43546 7956 43548
rect 8012 43546 8036 43548
rect 8092 43546 8116 43548
rect 8172 43546 8196 43548
rect 8252 43546 8258 43548
rect 8012 43494 8014 43546
rect 8194 43494 8196 43546
rect 7950 43492 7956 43494
rect 8012 43492 8036 43494
rect 8092 43492 8116 43494
rect 8172 43492 8196 43494
rect 8252 43492 8258 43494
rect 7950 43483 8258 43492
rect 7840 43444 7892 43450
rect 7840 43386 7892 43392
rect 8496 42770 8524 49846
rect 8760 49768 8812 49774
rect 8760 49710 8812 49716
rect 8772 45558 8800 49710
rect 9232 47802 9260 52022
rect 9312 51400 9364 51406
rect 9312 51342 9364 51348
rect 9220 47796 9272 47802
rect 9220 47738 9272 47744
rect 9324 46170 9352 51342
rect 9404 50924 9456 50930
rect 9404 50866 9456 50872
rect 9312 46164 9364 46170
rect 9312 46106 9364 46112
rect 8852 45824 8904 45830
rect 8852 45766 8904 45772
rect 8760 45552 8812 45558
rect 8760 45494 8812 45500
rect 8484 42764 8536 42770
rect 8484 42706 8536 42712
rect 8300 42696 8352 42702
rect 8300 42638 8352 42644
rect 7840 42560 7892 42566
rect 7840 42502 7892 42508
rect 7852 42294 7880 42502
rect 7950 42460 8258 42469
rect 7950 42458 7956 42460
rect 8012 42458 8036 42460
rect 8092 42458 8116 42460
rect 8172 42458 8196 42460
rect 8252 42458 8258 42460
rect 8012 42406 8014 42458
rect 8194 42406 8196 42458
rect 7950 42404 7956 42406
rect 8012 42404 8036 42406
rect 8092 42404 8116 42406
rect 8172 42404 8196 42406
rect 8252 42404 8258 42406
rect 7950 42395 8258 42404
rect 7840 42288 7892 42294
rect 7840 42230 7892 42236
rect 8312 41750 8340 42638
rect 8496 42294 8524 42706
rect 8484 42288 8536 42294
rect 8484 42230 8536 42236
rect 8496 41970 8524 42230
rect 8404 41942 8524 41970
rect 8300 41744 8352 41750
rect 8300 41686 8352 41692
rect 8404 41614 8432 41942
rect 8484 41812 8536 41818
rect 8484 41754 8536 41760
rect 8392 41608 8444 41614
rect 8392 41550 8444 41556
rect 7760 41386 7880 41414
rect 7852 40746 7880 41386
rect 7950 41372 8258 41381
rect 7950 41370 7956 41372
rect 8012 41370 8036 41372
rect 8092 41370 8116 41372
rect 8172 41370 8196 41372
rect 8252 41370 8258 41372
rect 8012 41318 8014 41370
rect 8194 41318 8196 41370
rect 7950 41316 7956 41318
rect 8012 41316 8036 41318
rect 8092 41316 8116 41318
rect 8172 41316 8196 41318
rect 8252 41316 8258 41318
rect 7950 41307 8258 41316
rect 8496 41070 8524 41754
rect 8668 41608 8720 41614
rect 8668 41550 8720 41556
rect 8484 41064 8536 41070
rect 8484 41006 8536 41012
rect 7852 40718 8248 40746
rect 7840 40656 7892 40662
rect 7840 40598 7892 40604
rect 7748 39976 7800 39982
rect 7748 39918 7800 39924
rect 7760 38962 7788 39918
rect 7852 38962 7880 40598
rect 8220 40474 8248 40718
rect 8496 40526 8524 41006
rect 8576 40928 8628 40934
rect 8576 40870 8628 40876
rect 8484 40520 8536 40526
rect 8220 40446 8340 40474
rect 8484 40462 8536 40468
rect 7950 40284 8258 40293
rect 7950 40282 7956 40284
rect 8012 40282 8036 40284
rect 8092 40282 8116 40284
rect 8172 40282 8196 40284
rect 8252 40282 8258 40284
rect 8012 40230 8014 40282
rect 8194 40230 8196 40282
rect 7950 40228 7956 40230
rect 8012 40228 8036 40230
rect 8092 40228 8116 40230
rect 8172 40228 8196 40230
rect 8252 40228 8258 40230
rect 7950 40219 8258 40228
rect 7950 39196 8258 39205
rect 7950 39194 7956 39196
rect 8012 39194 8036 39196
rect 8092 39194 8116 39196
rect 8172 39194 8196 39196
rect 8252 39194 8258 39196
rect 8012 39142 8014 39194
rect 8194 39142 8196 39194
rect 7950 39140 7956 39142
rect 8012 39140 8036 39142
rect 8092 39140 8116 39142
rect 8172 39140 8196 39142
rect 8252 39140 8258 39142
rect 7950 39131 8258 39140
rect 7748 38956 7800 38962
rect 7748 38898 7800 38904
rect 7840 38956 7892 38962
rect 7840 38898 7892 38904
rect 7760 38214 7788 38898
rect 7748 38208 7800 38214
rect 7748 38150 7800 38156
rect 7840 38208 7892 38214
rect 7840 38150 7892 38156
rect 7656 36372 7708 36378
rect 7656 36314 7708 36320
rect 7656 36236 7708 36242
rect 7656 36178 7708 36184
rect 7392 35958 7512 35986
rect 7564 36032 7616 36038
rect 7564 35974 7616 35980
rect 7288 35760 7340 35766
rect 7288 35702 7340 35708
rect 7288 34944 7340 34950
rect 7288 34886 7340 34892
rect 7196 31204 7248 31210
rect 7196 31146 7248 31152
rect 7300 30938 7328 34886
rect 7392 34542 7420 35958
rect 7380 34536 7432 34542
rect 7380 34478 7432 34484
rect 7288 30932 7340 30938
rect 7288 30874 7340 30880
rect 7392 29594 7420 34478
rect 7472 33856 7524 33862
rect 7472 33798 7524 33804
rect 7484 31482 7512 33798
rect 7576 33114 7604 35974
rect 7668 33522 7696 36178
rect 7748 35148 7800 35154
rect 7748 35090 7800 35096
rect 7760 34746 7788 35090
rect 7748 34740 7800 34746
rect 7748 34682 7800 34688
rect 7760 33998 7788 34682
rect 7852 34202 7880 38150
rect 7950 38108 8258 38117
rect 7950 38106 7956 38108
rect 8012 38106 8036 38108
rect 8092 38106 8116 38108
rect 8172 38106 8196 38108
rect 8252 38106 8258 38108
rect 8012 38054 8014 38106
rect 8194 38054 8196 38106
rect 7950 38052 7956 38054
rect 8012 38052 8036 38054
rect 8092 38052 8116 38054
rect 8172 38052 8196 38054
rect 8252 38052 8258 38054
rect 7950 38043 8258 38052
rect 8208 37936 8260 37942
rect 8208 37878 8260 37884
rect 8220 37262 8248 37878
rect 8208 37256 8260 37262
rect 8208 37198 8260 37204
rect 7950 37020 8258 37029
rect 7950 37018 7956 37020
rect 8012 37018 8036 37020
rect 8092 37018 8116 37020
rect 8172 37018 8196 37020
rect 8252 37018 8258 37020
rect 8012 36966 8014 37018
rect 8194 36966 8196 37018
rect 7950 36964 7956 36966
rect 8012 36964 8036 36966
rect 8092 36964 8116 36966
rect 8172 36964 8196 36966
rect 8252 36964 8258 36966
rect 7950 36955 8258 36964
rect 7950 35932 8258 35941
rect 7950 35930 7956 35932
rect 8012 35930 8036 35932
rect 8092 35930 8116 35932
rect 8172 35930 8196 35932
rect 8252 35930 8258 35932
rect 8012 35878 8014 35930
rect 8194 35878 8196 35930
rect 7950 35876 7956 35878
rect 8012 35876 8036 35878
rect 8092 35876 8116 35878
rect 8172 35876 8196 35878
rect 8252 35876 8258 35878
rect 7950 35867 8258 35876
rect 8116 35760 8168 35766
rect 8116 35702 8168 35708
rect 8128 35222 8156 35702
rect 8116 35216 8168 35222
rect 8116 35158 8168 35164
rect 7950 34844 8258 34853
rect 7950 34842 7956 34844
rect 8012 34842 8036 34844
rect 8092 34842 8116 34844
rect 8172 34842 8196 34844
rect 8252 34842 8258 34844
rect 8012 34790 8014 34842
rect 8194 34790 8196 34842
rect 7950 34788 7956 34790
rect 8012 34788 8036 34790
rect 8092 34788 8116 34790
rect 8172 34788 8196 34790
rect 8252 34788 8258 34790
rect 7950 34779 8258 34788
rect 8312 34490 8340 40446
rect 8496 40390 8524 40462
rect 8484 40384 8536 40390
rect 8484 40326 8536 40332
rect 8392 40112 8444 40118
rect 8392 40054 8444 40060
rect 8404 39098 8432 40054
rect 8496 39642 8524 40326
rect 8588 40118 8616 40870
rect 8680 40730 8708 41550
rect 8864 41414 8892 45766
rect 8944 45620 8996 45626
rect 8944 45562 8996 45568
rect 8956 43246 8984 45562
rect 9312 45552 9364 45558
rect 9312 45494 9364 45500
rect 9220 44396 9272 44402
rect 9220 44338 9272 44344
rect 9232 44198 9260 44338
rect 9220 44192 9272 44198
rect 9220 44134 9272 44140
rect 9036 43784 9088 43790
rect 9036 43726 9088 43732
rect 8944 43240 8996 43246
rect 8944 43182 8996 43188
rect 8956 42906 8984 43182
rect 8944 42900 8996 42906
rect 8944 42842 8996 42848
rect 8956 41818 8984 42842
rect 8944 41812 8996 41818
rect 8944 41754 8996 41760
rect 8956 41682 8984 41754
rect 8944 41676 8996 41682
rect 8944 41618 8996 41624
rect 8864 41386 8984 41414
rect 8668 40724 8720 40730
rect 8668 40666 8720 40672
rect 8680 40458 8708 40666
rect 8760 40588 8812 40594
rect 8760 40530 8812 40536
rect 8668 40452 8720 40458
rect 8668 40394 8720 40400
rect 8576 40112 8628 40118
rect 8576 40054 8628 40060
rect 8576 39976 8628 39982
rect 8576 39918 8628 39924
rect 8668 39976 8720 39982
rect 8668 39918 8720 39924
rect 8588 39642 8616 39918
rect 8484 39636 8536 39642
rect 8484 39578 8536 39584
rect 8576 39636 8628 39642
rect 8576 39578 8628 39584
rect 8680 39574 8708 39918
rect 8668 39568 8720 39574
rect 8668 39510 8720 39516
rect 8576 39500 8628 39506
rect 8576 39442 8628 39448
rect 8392 39092 8444 39098
rect 8392 39034 8444 39040
rect 8588 37754 8616 39442
rect 8772 39438 8800 40530
rect 8852 40180 8904 40186
rect 8852 40122 8904 40128
rect 8760 39432 8812 39438
rect 8760 39374 8812 39380
rect 8668 39364 8720 39370
rect 8668 39306 8720 39312
rect 8680 37942 8708 39306
rect 8668 37936 8720 37942
rect 8668 37878 8720 37884
rect 8588 37726 8708 37754
rect 8576 37664 8628 37670
rect 8576 37606 8628 37612
rect 8588 37466 8616 37606
rect 8576 37460 8628 37466
rect 8576 37402 8628 37408
rect 8576 37324 8628 37330
rect 8576 37266 8628 37272
rect 8588 36582 8616 37266
rect 8576 36576 8628 36582
rect 8576 36518 8628 36524
rect 8392 35488 8444 35494
rect 8392 35430 8444 35436
rect 8404 35222 8432 35430
rect 8392 35216 8444 35222
rect 8392 35158 8444 35164
rect 8404 34746 8432 35158
rect 8484 35080 8536 35086
rect 8484 35022 8536 35028
rect 8392 34740 8444 34746
rect 8392 34682 8444 34688
rect 8496 34678 8524 35022
rect 8484 34672 8536 34678
rect 8484 34614 8536 34620
rect 8588 34626 8616 36518
rect 8680 34762 8708 37726
rect 8760 36236 8812 36242
rect 8760 36178 8812 36184
rect 8772 35290 8800 36178
rect 8864 35290 8892 40122
rect 8956 39030 8984 41386
rect 8944 39024 8996 39030
rect 8944 38966 8996 38972
rect 8944 38820 8996 38826
rect 8944 38762 8996 38768
rect 8956 36378 8984 38762
rect 9048 38010 9076 43726
rect 9128 41472 9180 41478
rect 9128 41414 9180 41420
rect 9140 39506 9168 41414
rect 9128 39500 9180 39506
rect 9128 39442 9180 39448
rect 9232 38486 9260 44134
rect 9324 43314 9352 45494
rect 9416 45082 9444 50866
rect 9496 46572 9548 46578
rect 9496 46514 9548 46520
rect 9404 45076 9456 45082
rect 9404 45018 9456 45024
rect 9312 43308 9364 43314
rect 9312 43250 9364 43256
rect 9508 42362 9536 46514
rect 9600 43382 9628 52906
rect 9692 51950 9720 53536
rect 9772 53100 9824 53106
rect 9772 53042 9824 53048
rect 9680 51944 9732 51950
rect 9680 51886 9732 51892
rect 9784 49910 9812 53042
rect 9864 52012 9916 52018
rect 9864 51954 9916 51960
rect 9772 49904 9824 49910
rect 9772 49846 9824 49852
rect 9680 46980 9732 46986
rect 9680 46922 9732 46928
rect 9588 43376 9640 43382
rect 9588 43318 9640 43324
rect 9600 42906 9628 43318
rect 9692 42906 9720 46922
rect 9876 45082 9904 51954
rect 9968 51610 9996 54130
rect 10232 54120 10284 54126
rect 10232 54062 10284 54068
rect 9956 51604 10008 51610
rect 9956 51546 10008 51552
rect 10244 45626 10272 54062
rect 10324 53576 10376 53582
rect 10324 53518 10376 53524
rect 10232 45620 10284 45626
rect 10232 45562 10284 45568
rect 9864 45076 9916 45082
rect 9864 45018 9916 45024
rect 10336 45014 10364 53518
rect 10428 53038 10456 55186
rect 10416 53032 10468 53038
rect 10416 52974 10468 52980
rect 10704 52562 10732 56200
rect 11072 53650 11100 56200
rect 11440 54262 11468 56200
rect 11428 54256 11480 54262
rect 11428 54198 11480 54204
rect 11704 53984 11756 53990
rect 11704 53926 11756 53932
rect 11060 53644 11112 53650
rect 11060 53586 11112 53592
rect 10968 53168 11020 53174
rect 10968 53110 11020 53116
rect 10692 52556 10744 52562
rect 10692 52498 10744 52504
rect 10784 52488 10836 52494
rect 10784 52430 10836 52436
rect 10796 50998 10824 52430
rect 10784 50992 10836 50998
rect 10784 50934 10836 50940
rect 10692 49224 10744 49230
rect 10692 49166 10744 49172
rect 10508 49088 10560 49094
rect 10508 49030 10560 49036
rect 10324 45008 10376 45014
rect 10324 44950 10376 44956
rect 9772 44736 9824 44742
rect 9770 44704 9772 44713
rect 9824 44704 9826 44713
rect 9770 44639 9826 44648
rect 10232 44396 10284 44402
rect 10232 44338 10284 44344
rect 10244 44305 10272 44338
rect 10230 44296 10286 44305
rect 10230 44231 10286 44240
rect 10416 44192 10468 44198
rect 10416 44134 10468 44140
rect 9956 43988 10008 43994
rect 9956 43930 10008 43936
rect 9588 42900 9640 42906
rect 9588 42842 9640 42848
rect 9680 42900 9732 42906
rect 9680 42842 9732 42848
rect 9496 42356 9548 42362
rect 9496 42298 9548 42304
rect 9496 41608 9548 41614
rect 9496 41550 9548 41556
rect 9404 40384 9456 40390
rect 9404 40326 9456 40332
rect 9312 39432 9364 39438
rect 9312 39374 9364 39380
rect 9220 38480 9272 38486
rect 9220 38422 9272 38428
rect 9036 38004 9088 38010
rect 9036 37946 9088 37952
rect 9324 37466 9352 39374
rect 9416 39370 9444 40326
rect 9508 40118 9536 41550
rect 9600 41414 9628 42842
rect 9772 42696 9824 42702
rect 9772 42638 9824 42644
rect 9784 42158 9812 42638
rect 9772 42152 9824 42158
rect 9772 42094 9824 42100
rect 9600 41386 9720 41414
rect 9692 40390 9720 41386
rect 9680 40384 9732 40390
rect 9680 40326 9732 40332
rect 9680 40180 9732 40186
rect 9680 40122 9732 40128
rect 9496 40112 9548 40118
rect 9496 40054 9548 40060
rect 9404 39364 9456 39370
rect 9404 39306 9456 39312
rect 9588 39024 9640 39030
rect 9588 38966 9640 38972
rect 9600 38894 9628 38966
rect 9588 38888 9640 38894
rect 9588 38830 9640 38836
rect 9600 38758 9628 38830
rect 9588 38752 9640 38758
rect 9588 38694 9640 38700
rect 9692 38418 9720 40122
rect 9680 38412 9732 38418
rect 9784 38400 9812 42094
rect 9864 38412 9916 38418
rect 9784 38372 9864 38400
rect 9680 38354 9732 38360
rect 9864 38354 9916 38360
rect 9864 38208 9916 38214
rect 9864 38150 9916 38156
rect 9496 38004 9548 38010
rect 9496 37946 9548 37952
rect 9404 37868 9456 37874
rect 9404 37810 9456 37816
rect 9312 37460 9364 37466
rect 9312 37402 9364 37408
rect 8944 36372 8996 36378
rect 8944 36314 8996 36320
rect 8760 35284 8812 35290
rect 8760 35226 8812 35232
rect 8852 35284 8904 35290
rect 8852 35226 8904 35232
rect 9324 35154 9352 37402
rect 9312 35148 9364 35154
rect 9312 35090 9364 35096
rect 8680 34734 8892 34762
rect 8588 34598 8708 34626
rect 8312 34462 8524 34490
rect 8392 34400 8444 34406
rect 8392 34342 8444 34348
rect 7840 34196 7892 34202
rect 7840 34138 7892 34144
rect 8300 34128 8352 34134
rect 8300 34070 8352 34076
rect 7748 33992 7800 33998
rect 7748 33934 7800 33940
rect 7760 33658 7788 33934
rect 7950 33756 8258 33765
rect 7950 33754 7956 33756
rect 8012 33754 8036 33756
rect 8092 33754 8116 33756
rect 8172 33754 8196 33756
rect 8252 33754 8258 33756
rect 8012 33702 8014 33754
rect 8194 33702 8196 33754
rect 7950 33700 7956 33702
rect 8012 33700 8036 33702
rect 8092 33700 8116 33702
rect 8172 33700 8196 33702
rect 8252 33700 8258 33702
rect 7950 33691 8258 33700
rect 7748 33652 7800 33658
rect 7748 33594 7800 33600
rect 7656 33516 7708 33522
rect 7656 33458 7708 33464
rect 7564 33108 7616 33114
rect 7564 33050 7616 33056
rect 7668 33046 7696 33458
rect 7840 33312 7892 33318
rect 7840 33254 7892 33260
rect 7656 33040 7708 33046
rect 7656 32982 7708 32988
rect 7748 32836 7800 32842
rect 7748 32778 7800 32784
rect 7656 32768 7708 32774
rect 7656 32710 7708 32716
rect 7668 32570 7696 32710
rect 7656 32564 7708 32570
rect 7656 32506 7708 32512
rect 7472 31476 7524 31482
rect 7472 31418 7524 31424
rect 7564 31272 7616 31278
rect 7564 31214 7616 31220
rect 7472 30592 7524 30598
rect 7472 30534 7524 30540
rect 6184 29572 6236 29578
rect 6184 29514 6236 29520
rect 7300 29566 7420 29594
rect 6196 26586 6224 29514
rect 7300 29510 7328 29566
rect 7288 29504 7340 29510
rect 7288 29446 7340 29452
rect 6460 29096 6512 29102
rect 6460 29038 6512 29044
rect 6472 28014 6500 29038
rect 7300 28490 7328 29446
rect 7288 28484 7340 28490
rect 7288 28426 7340 28432
rect 6828 28416 6880 28422
rect 6828 28358 6880 28364
rect 6840 28150 6868 28358
rect 6828 28144 6880 28150
rect 6828 28086 6880 28092
rect 6460 28008 6512 28014
rect 6460 27950 6512 27956
rect 6472 26926 6500 27950
rect 6736 27328 6788 27334
rect 6736 27270 6788 27276
rect 6460 26920 6512 26926
rect 6460 26862 6512 26868
rect 6184 26580 6236 26586
rect 6184 26522 6236 26528
rect 6092 24608 6144 24614
rect 6092 24550 6144 24556
rect 6104 24342 6132 24550
rect 6092 24336 6144 24342
rect 6092 24278 6144 24284
rect 6092 21888 6144 21894
rect 6092 21830 6144 21836
rect 6104 20874 6132 21830
rect 6092 20868 6144 20874
rect 6092 20810 6144 20816
rect 6104 20262 6132 20810
rect 6092 20256 6144 20262
rect 6092 20198 6144 20204
rect 6092 18760 6144 18766
rect 6092 18702 6144 18708
rect 6104 18222 6132 18702
rect 6092 18216 6144 18222
rect 6092 18158 6144 18164
rect 6104 17882 6132 18158
rect 6092 17876 6144 17882
rect 6092 17818 6144 17824
rect 6196 6914 6224 26522
rect 6472 26382 6500 26862
rect 6748 26450 6776 27270
rect 6828 26580 6880 26586
rect 6828 26522 6880 26528
rect 6840 26450 6868 26522
rect 6736 26444 6788 26450
rect 6736 26386 6788 26392
rect 6828 26444 6880 26450
rect 6828 26386 6880 26392
rect 6460 26376 6512 26382
rect 6460 26318 6512 26324
rect 6472 25888 6500 26318
rect 6552 25900 6604 25906
rect 6472 25860 6552 25888
rect 6552 25842 6604 25848
rect 6460 25220 6512 25226
rect 6460 25162 6512 25168
rect 6472 24410 6500 25162
rect 6460 24404 6512 24410
rect 6460 24346 6512 24352
rect 6564 23662 6592 25842
rect 6828 25832 6880 25838
rect 6828 25774 6880 25780
rect 6840 25294 6868 25774
rect 6828 25288 6880 25294
rect 6828 25230 6880 25236
rect 6828 24608 6880 24614
rect 6828 24550 6880 24556
rect 6736 24064 6788 24070
rect 6736 24006 6788 24012
rect 6552 23656 6604 23662
rect 6552 23598 6604 23604
rect 6368 22636 6420 22642
rect 6368 22578 6420 22584
rect 6276 21616 6328 21622
rect 6276 21558 6328 21564
rect 6104 6886 6224 6914
rect 6104 6730 6132 6886
rect 6092 6724 6144 6730
rect 6092 6666 6144 6672
rect 6288 5574 6316 21558
rect 6380 19174 6408 22578
rect 6748 21894 6776 24006
rect 6840 23798 6868 24550
rect 7104 24268 7156 24274
rect 7104 24210 7156 24216
rect 7116 23866 7144 24210
rect 7104 23860 7156 23866
rect 7104 23802 7156 23808
rect 6828 23792 6880 23798
rect 6828 23734 6880 23740
rect 7116 22642 7144 23802
rect 7196 23656 7248 23662
rect 7196 23598 7248 23604
rect 7104 22636 7156 22642
rect 7104 22578 7156 22584
rect 6736 21888 6788 21894
rect 6736 21830 6788 21836
rect 7208 21690 7236 23598
rect 7196 21684 7248 21690
rect 7196 21626 7248 21632
rect 6920 21548 6972 21554
rect 6920 21490 6972 21496
rect 6460 20460 6512 20466
rect 6460 20402 6512 20408
rect 6368 19168 6420 19174
rect 6368 19110 6420 19116
rect 6472 16810 6500 20402
rect 6736 20256 6788 20262
rect 6736 20198 6788 20204
rect 6748 19990 6776 20198
rect 6932 20058 6960 21490
rect 7104 21480 7156 21486
rect 7104 21422 7156 21428
rect 7012 21412 7064 21418
rect 7012 21354 7064 21360
rect 7024 20942 7052 21354
rect 7012 20936 7064 20942
rect 7012 20878 7064 20884
rect 6920 20052 6972 20058
rect 6920 19994 6972 20000
rect 6736 19984 6788 19990
rect 6736 19926 6788 19932
rect 6748 19854 6776 19926
rect 6736 19848 6788 19854
rect 6736 19790 6788 19796
rect 6748 19334 6776 19790
rect 7024 19718 7052 20878
rect 7116 20602 7144 21422
rect 7104 20596 7156 20602
rect 7104 20538 7156 20544
rect 7012 19712 7064 19718
rect 7012 19654 7064 19660
rect 6748 19306 6960 19334
rect 6828 19168 6880 19174
rect 6828 19110 6880 19116
rect 6840 18766 6868 19110
rect 6828 18760 6880 18766
rect 6828 18702 6880 18708
rect 6736 18692 6788 18698
rect 6736 18634 6788 18640
rect 6552 18216 6604 18222
rect 6552 18158 6604 18164
rect 6564 16998 6592 18158
rect 6748 17626 6776 18634
rect 6828 18624 6880 18630
rect 6828 18566 6880 18572
rect 6840 18358 6868 18566
rect 6932 18358 6960 19306
rect 7010 19272 7066 19281
rect 7010 19207 7066 19216
rect 6828 18352 6880 18358
rect 6828 18294 6880 18300
rect 6920 18352 6972 18358
rect 6920 18294 6972 18300
rect 6748 17598 6868 17626
rect 6932 17610 6960 18294
rect 6552 16992 6604 16998
rect 6552 16934 6604 16940
rect 6380 16782 6500 16810
rect 6380 16250 6408 16782
rect 6564 16538 6592 16934
rect 6644 16652 6696 16658
rect 6644 16594 6696 16600
rect 6656 16538 6684 16594
rect 6564 16510 6684 16538
rect 6656 16402 6684 16510
rect 6656 16374 6776 16402
rect 6368 16244 6420 16250
rect 6368 16186 6420 16192
rect 6748 15502 6776 16374
rect 6736 15496 6788 15502
rect 6736 15438 6788 15444
rect 6748 13870 6776 15438
rect 6736 13864 6788 13870
rect 6736 13806 6788 13812
rect 6840 8498 6868 17598
rect 6920 17604 6972 17610
rect 6920 17546 6972 17552
rect 6932 17338 6960 17546
rect 6920 17332 6972 17338
rect 6920 17274 6972 17280
rect 6932 16454 6960 17274
rect 6920 16448 6972 16454
rect 6920 16390 6972 16396
rect 6828 8492 6880 8498
rect 6828 8434 6880 8440
rect 6276 5568 6328 5574
rect 6276 5510 6328 5516
rect 6092 3936 6144 3942
rect 6092 3878 6144 3884
rect 6000 3732 6052 3738
rect 6000 3674 6052 3680
rect 6104 3534 6132 3878
rect 6092 3528 6144 3534
rect 6092 3470 6144 3476
rect 6460 3528 6512 3534
rect 6460 3470 6512 3476
rect 5908 3188 5960 3194
rect 5908 3130 5960 3136
rect 5816 2916 5868 2922
rect 5816 2858 5868 2864
rect 5724 2372 5776 2378
rect 5724 2314 5776 2320
rect 5736 800 5764 2314
rect 6104 800 6132 3470
rect 6472 2854 6500 3470
rect 6828 3392 6880 3398
rect 6828 3334 6880 3340
rect 6840 3058 6868 3334
rect 7024 3194 7052 19207
rect 7104 18420 7156 18426
rect 7104 18362 7156 18368
rect 7116 17882 7144 18362
rect 7104 17876 7156 17882
rect 7104 17818 7156 17824
rect 7104 13252 7156 13258
rect 7104 13194 7156 13200
rect 7116 9178 7144 13194
rect 7104 9172 7156 9178
rect 7104 9114 7156 9120
rect 7300 3194 7328 28426
rect 7484 25362 7512 30534
rect 7472 25356 7524 25362
rect 7472 25298 7524 25304
rect 7576 24750 7604 31214
rect 7760 28762 7788 32778
rect 7852 32502 7880 33254
rect 8312 32978 8340 34070
rect 8404 32978 8432 34342
rect 8496 33046 8524 34462
rect 8576 33924 8628 33930
rect 8576 33866 8628 33872
rect 8484 33040 8536 33046
rect 8484 32982 8536 32988
rect 8300 32972 8352 32978
rect 8300 32914 8352 32920
rect 8392 32972 8444 32978
rect 8392 32914 8444 32920
rect 7950 32668 8258 32677
rect 7950 32666 7956 32668
rect 8012 32666 8036 32668
rect 8092 32666 8116 32668
rect 8172 32666 8196 32668
rect 8252 32666 8258 32668
rect 8012 32614 8014 32666
rect 8194 32614 8196 32666
rect 7950 32612 7956 32614
rect 8012 32612 8036 32614
rect 8092 32612 8116 32614
rect 8172 32612 8196 32614
rect 8252 32612 8258 32614
rect 7950 32603 8258 32612
rect 7840 32496 7892 32502
rect 7840 32438 7892 32444
rect 8024 32496 8076 32502
rect 8024 32438 8076 32444
rect 8312 32450 8340 32914
rect 8588 32842 8616 33866
rect 8576 32836 8628 32842
rect 8576 32778 8628 32784
rect 8036 32366 8064 32438
rect 8312 32422 8432 32450
rect 8024 32360 8076 32366
rect 8024 32302 8076 32308
rect 8300 32360 8352 32366
rect 8300 32302 8352 32308
rect 7840 31952 7892 31958
rect 7840 31894 7892 31900
rect 7656 28756 7708 28762
rect 7656 28698 7708 28704
rect 7748 28756 7800 28762
rect 7748 28698 7800 28704
rect 7668 28422 7696 28698
rect 7852 28626 7880 31894
rect 8036 31890 8064 32302
rect 8024 31884 8076 31890
rect 8024 31826 8076 31832
rect 7950 31580 8258 31589
rect 7950 31578 7956 31580
rect 8012 31578 8036 31580
rect 8092 31578 8116 31580
rect 8172 31578 8196 31580
rect 8252 31578 8258 31580
rect 8012 31526 8014 31578
rect 8194 31526 8196 31578
rect 7950 31524 7956 31526
rect 8012 31524 8036 31526
rect 8092 31524 8116 31526
rect 8172 31524 8196 31526
rect 8252 31524 8258 31526
rect 7950 31515 8258 31524
rect 7932 31272 7984 31278
rect 7932 31214 7984 31220
rect 7944 30734 7972 31214
rect 7932 30728 7984 30734
rect 7932 30670 7984 30676
rect 8312 30666 8340 32302
rect 8404 32026 8432 32422
rect 8588 32026 8616 32778
rect 8680 32230 8708 34598
rect 8864 33658 8892 34734
rect 8852 33652 8904 33658
rect 8852 33594 8904 33600
rect 8668 32224 8720 32230
rect 8668 32166 8720 32172
rect 8392 32020 8444 32026
rect 8392 31962 8444 31968
rect 8576 32020 8628 32026
rect 8576 31962 8628 31968
rect 8680 30938 8708 32166
rect 8668 30932 8720 30938
rect 8668 30874 8720 30880
rect 8300 30660 8352 30666
rect 8300 30602 8352 30608
rect 7950 30492 8258 30501
rect 7950 30490 7956 30492
rect 8012 30490 8036 30492
rect 8092 30490 8116 30492
rect 8172 30490 8196 30492
rect 8252 30490 8258 30492
rect 8012 30438 8014 30490
rect 8194 30438 8196 30490
rect 7950 30436 7956 30438
rect 8012 30436 8036 30438
rect 8092 30436 8116 30438
rect 8172 30436 8196 30438
rect 8252 30436 8258 30438
rect 7950 30427 8258 30436
rect 8300 30048 8352 30054
rect 8300 29990 8352 29996
rect 7950 29404 8258 29413
rect 7950 29402 7956 29404
rect 8012 29402 8036 29404
rect 8092 29402 8116 29404
rect 8172 29402 8196 29404
rect 8252 29402 8258 29404
rect 8012 29350 8014 29402
rect 8194 29350 8196 29402
rect 7950 29348 7956 29350
rect 8012 29348 8036 29350
rect 8092 29348 8116 29350
rect 8172 29348 8196 29350
rect 8252 29348 8258 29350
rect 7950 29339 8258 29348
rect 8312 28966 8340 29990
rect 8576 29232 8628 29238
rect 8576 29174 8628 29180
rect 8300 28960 8352 28966
rect 8300 28902 8352 28908
rect 7748 28620 7800 28626
rect 7748 28562 7800 28568
rect 7840 28620 7892 28626
rect 7840 28562 7892 28568
rect 7656 28416 7708 28422
rect 7656 28358 7708 28364
rect 7760 26586 7788 28562
rect 7852 27674 7880 28562
rect 7950 28316 8258 28325
rect 7950 28314 7956 28316
rect 8012 28314 8036 28316
rect 8092 28314 8116 28316
rect 8172 28314 8196 28316
rect 8252 28314 8258 28316
rect 8012 28262 8014 28314
rect 8194 28262 8196 28314
rect 7950 28260 7956 28262
rect 8012 28260 8036 28262
rect 8092 28260 8116 28262
rect 8172 28260 8196 28262
rect 8252 28260 8258 28262
rect 7950 28251 8258 28260
rect 8588 28218 8616 29174
rect 8668 29164 8720 29170
rect 8668 29106 8720 29112
rect 8680 28966 8708 29106
rect 8760 29028 8812 29034
rect 8760 28970 8812 28976
rect 8668 28960 8720 28966
rect 8668 28902 8720 28908
rect 8680 28218 8708 28902
rect 8772 28558 8800 28970
rect 8760 28552 8812 28558
rect 8760 28494 8812 28500
rect 8576 28212 8628 28218
rect 8576 28154 8628 28160
rect 8668 28212 8720 28218
rect 8668 28154 8720 28160
rect 7840 27668 7892 27674
rect 7840 27610 7892 27616
rect 8300 27464 8352 27470
rect 8300 27406 8352 27412
rect 7950 27228 8258 27237
rect 7950 27226 7956 27228
rect 8012 27226 8036 27228
rect 8092 27226 8116 27228
rect 8172 27226 8196 27228
rect 8252 27226 8258 27228
rect 8012 27174 8014 27226
rect 8194 27174 8196 27226
rect 7950 27172 7956 27174
rect 8012 27172 8036 27174
rect 8092 27172 8116 27174
rect 8172 27172 8196 27174
rect 8252 27172 8258 27174
rect 7950 27163 8258 27172
rect 7840 27124 7892 27130
rect 7840 27066 7892 27072
rect 7748 26580 7800 26586
rect 7748 26522 7800 26528
rect 7760 25974 7788 26522
rect 7748 25968 7800 25974
rect 7748 25910 7800 25916
rect 7760 24954 7788 25910
rect 7852 25430 7880 27066
rect 8312 26858 8340 27406
rect 8588 27130 8616 28154
rect 8680 27130 8708 28154
rect 8772 27538 8800 28494
rect 8760 27532 8812 27538
rect 8760 27474 8812 27480
rect 8576 27124 8628 27130
rect 8576 27066 8628 27072
rect 8668 27124 8720 27130
rect 8668 27066 8720 27072
rect 8576 26920 8628 26926
rect 8576 26862 8628 26868
rect 8300 26852 8352 26858
rect 8300 26794 8352 26800
rect 7950 26140 8258 26149
rect 7950 26138 7956 26140
rect 8012 26138 8036 26140
rect 8092 26138 8116 26140
rect 8172 26138 8196 26140
rect 8252 26138 8258 26140
rect 8012 26086 8014 26138
rect 8194 26086 8196 26138
rect 7950 26084 7956 26086
rect 8012 26084 8036 26086
rect 8092 26084 8116 26086
rect 8172 26084 8196 26086
rect 8252 26084 8258 26086
rect 7950 26075 8258 26084
rect 8484 26036 8536 26042
rect 8484 25978 8536 25984
rect 7840 25424 7892 25430
rect 7840 25366 7892 25372
rect 7950 25052 8258 25061
rect 7950 25050 7956 25052
rect 8012 25050 8036 25052
rect 8092 25050 8116 25052
rect 8172 25050 8196 25052
rect 8252 25050 8258 25052
rect 8012 24998 8014 25050
rect 8194 24998 8196 25050
rect 7950 24996 7956 24998
rect 8012 24996 8036 24998
rect 8092 24996 8116 24998
rect 8172 24996 8196 24998
rect 8252 24996 8258 24998
rect 7950 24987 8258 24996
rect 7748 24948 7800 24954
rect 7748 24890 7800 24896
rect 7748 24812 7800 24818
rect 7748 24754 7800 24760
rect 7564 24744 7616 24750
rect 7564 24686 7616 24692
rect 7656 24676 7708 24682
rect 7656 24618 7708 24624
rect 7472 24404 7524 24410
rect 7472 24346 7524 24352
rect 7484 21026 7512 24346
rect 7564 22976 7616 22982
rect 7564 22918 7616 22924
rect 7576 21146 7604 22918
rect 7668 22030 7696 24618
rect 7760 23322 7788 24754
rect 8496 24342 8524 25978
rect 8588 24410 8616 26862
rect 8680 26586 8708 27066
rect 8864 26926 8892 33594
rect 9416 33114 9444 37810
rect 9508 36582 9536 37946
rect 9588 37732 9640 37738
rect 9588 37674 9640 37680
rect 9496 36576 9548 36582
rect 9496 36518 9548 36524
rect 9496 35216 9548 35222
rect 9496 35158 9548 35164
rect 9404 33108 9456 33114
rect 9404 33050 9456 33056
rect 9404 32428 9456 32434
rect 9404 32370 9456 32376
rect 9416 31890 9444 32370
rect 9508 31890 9536 35158
rect 9600 34746 9628 37674
rect 9876 37398 9904 38150
rect 9864 37392 9916 37398
rect 9864 37334 9916 37340
rect 9680 36712 9732 36718
rect 9680 36654 9732 36660
rect 9588 34740 9640 34746
rect 9588 34682 9640 34688
rect 9600 33998 9628 34682
rect 9588 33992 9640 33998
rect 9588 33934 9640 33940
rect 9692 32570 9720 36654
rect 9968 36378 9996 43930
rect 10428 43450 10456 44134
rect 10520 43994 10548 49030
rect 10600 46572 10652 46578
rect 10600 46514 10652 46520
rect 10508 43988 10560 43994
rect 10508 43930 10560 43936
rect 10416 43444 10468 43450
rect 10416 43386 10468 43392
rect 10520 43330 10548 43930
rect 10232 43308 10284 43314
rect 10232 43250 10284 43256
rect 10428 43302 10548 43330
rect 10140 42220 10192 42226
rect 10140 42162 10192 42168
rect 10048 39296 10100 39302
rect 10048 39238 10100 39244
rect 10060 38350 10088 39238
rect 10152 38826 10180 42162
rect 10244 42090 10272 43250
rect 10324 42152 10376 42158
rect 10324 42094 10376 42100
rect 10232 42084 10284 42090
rect 10232 42026 10284 42032
rect 10244 41414 10272 42026
rect 10336 41750 10364 42094
rect 10324 41744 10376 41750
rect 10324 41686 10376 41692
rect 10244 41386 10364 41414
rect 10232 40724 10284 40730
rect 10232 40666 10284 40672
rect 10244 40458 10272 40666
rect 10232 40452 10284 40458
rect 10232 40394 10284 40400
rect 10140 38820 10192 38826
rect 10140 38762 10192 38768
rect 10048 38344 10100 38350
rect 10048 38286 10100 38292
rect 10336 37330 10364 41386
rect 10428 37466 10456 43302
rect 10508 42220 10560 42226
rect 10508 42162 10560 42168
rect 10520 38554 10548 42162
rect 10612 41478 10640 46514
rect 10704 46170 10732 49166
rect 10876 46504 10928 46510
rect 10876 46446 10928 46452
rect 10692 46164 10744 46170
rect 10692 46106 10744 46112
rect 10888 45286 10916 46446
rect 10876 45280 10928 45286
rect 10876 45222 10928 45228
rect 10980 44538 11008 53110
rect 11716 48278 11744 53926
rect 11808 53038 11836 56200
rect 12176 53650 12204 56200
rect 12348 54188 12400 54194
rect 12348 54130 12400 54136
rect 12164 53644 12216 53650
rect 12164 53586 12216 53592
rect 11888 53100 11940 53106
rect 11888 53042 11940 53048
rect 11796 53032 11848 53038
rect 11796 52974 11848 52980
rect 11900 52154 11928 53042
rect 12360 52154 12388 54130
rect 12544 54126 12572 56200
rect 12912 54262 12940 56200
rect 13280 55214 13308 56200
rect 13280 55186 13400 55214
rect 12900 54256 12952 54262
rect 12900 54198 12952 54204
rect 12532 54120 12584 54126
rect 12532 54062 12584 54068
rect 12950 53884 13258 53893
rect 12950 53882 12956 53884
rect 13012 53882 13036 53884
rect 13092 53882 13116 53884
rect 13172 53882 13196 53884
rect 13252 53882 13258 53884
rect 13012 53830 13014 53882
rect 13194 53830 13196 53882
rect 12950 53828 12956 53830
rect 13012 53828 13036 53830
rect 13092 53828 13116 53830
rect 13172 53828 13196 53830
rect 13252 53828 13258 53830
rect 12950 53819 13258 53828
rect 12624 53576 12676 53582
rect 12624 53518 12676 53524
rect 12636 52698 12664 53518
rect 12950 52796 13258 52805
rect 12950 52794 12956 52796
rect 13012 52794 13036 52796
rect 13092 52794 13116 52796
rect 13172 52794 13196 52796
rect 13252 52794 13258 52796
rect 13012 52742 13014 52794
rect 13194 52742 13196 52794
rect 12950 52740 12956 52742
rect 13012 52740 13036 52742
rect 13092 52740 13116 52742
rect 13172 52740 13196 52742
rect 13252 52740 13258 52742
rect 12950 52731 13258 52740
rect 12624 52692 12676 52698
rect 12624 52634 12676 52640
rect 12808 52488 12860 52494
rect 12808 52430 12860 52436
rect 11888 52148 11940 52154
rect 11888 52090 11940 52096
rect 12348 52148 12400 52154
rect 12348 52090 12400 52096
rect 11888 52012 11940 52018
rect 11888 51954 11940 51960
rect 11980 52012 12032 52018
rect 11980 51954 12032 51960
rect 11704 48272 11756 48278
rect 11704 48214 11756 48220
rect 11704 47660 11756 47666
rect 11704 47602 11756 47608
rect 11428 47456 11480 47462
rect 11428 47398 11480 47404
rect 11440 46986 11468 47398
rect 11428 46980 11480 46986
rect 11428 46922 11480 46928
rect 11152 46912 11204 46918
rect 11152 46854 11204 46860
rect 11336 46912 11388 46918
rect 11336 46854 11388 46860
rect 11164 46714 11192 46854
rect 11152 46708 11204 46714
rect 11152 46650 11204 46656
rect 11348 46034 11376 46854
rect 11336 46028 11388 46034
rect 11336 45970 11388 45976
rect 11152 45824 11204 45830
rect 11152 45766 11204 45772
rect 11060 45348 11112 45354
rect 11060 45290 11112 45296
rect 10968 44532 11020 44538
rect 10968 44474 11020 44480
rect 10876 43852 10928 43858
rect 10876 43794 10928 43800
rect 10888 42770 10916 43794
rect 10876 42764 10928 42770
rect 10876 42706 10928 42712
rect 11072 42362 11100 45290
rect 11164 44538 11192 45766
rect 11440 45558 11468 46922
rect 11520 45960 11572 45966
rect 11520 45902 11572 45908
rect 11428 45552 11480 45558
rect 11428 45494 11480 45500
rect 11440 44946 11468 45494
rect 11428 44940 11480 44946
rect 11428 44882 11480 44888
rect 11152 44532 11204 44538
rect 11152 44474 11204 44480
rect 11440 43994 11468 44882
rect 11428 43988 11480 43994
rect 11428 43930 11480 43936
rect 11244 42900 11296 42906
rect 11244 42842 11296 42848
rect 11060 42356 11112 42362
rect 11060 42298 11112 42304
rect 10784 42016 10836 42022
rect 10784 41958 10836 41964
rect 10796 41682 10824 41958
rect 10784 41676 10836 41682
rect 10784 41618 10836 41624
rect 10876 41676 10928 41682
rect 10876 41618 10928 41624
rect 10600 41472 10652 41478
rect 10600 41414 10652 41420
rect 10692 41472 10744 41478
rect 10692 41414 10744 41420
rect 10600 40112 10652 40118
rect 10600 40054 10652 40060
rect 10508 38548 10560 38554
rect 10508 38490 10560 38496
rect 10612 38010 10640 40054
rect 10704 39098 10732 41414
rect 10796 40118 10824 41618
rect 10888 41274 10916 41618
rect 11072 41274 11100 42298
rect 11152 41540 11204 41546
rect 11152 41482 11204 41488
rect 11164 41290 11192 41482
rect 11256 41414 11284 42842
rect 11532 41818 11560 45902
rect 11612 44736 11664 44742
rect 11610 44704 11612 44713
rect 11664 44704 11666 44713
rect 11610 44639 11666 44648
rect 11610 44296 11666 44305
rect 11610 44231 11612 44240
rect 11664 44231 11666 44240
rect 11612 44202 11664 44208
rect 11716 42362 11744 47602
rect 11900 46714 11928 51954
rect 11992 49434 12020 51954
rect 12820 49434 12848 52430
rect 13372 52426 13400 55186
rect 13648 53174 13676 56200
rect 14016 53582 14044 56200
rect 14004 53576 14056 53582
rect 14004 53518 14056 53524
rect 13636 53168 13688 53174
rect 13636 53110 13688 53116
rect 13648 52698 13676 53110
rect 14384 53106 14412 56200
rect 14752 54330 14780 56200
rect 14740 54324 14792 54330
rect 14740 54266 14792 54272
rect 15120 54176 15148 56200
rect 15200 54188 15252 54194
rect 15120 54148 15200 54176
rect 15200 54130 15252 54136
rect 15488 53582 15516 56200
rect 15752 53984 15804 53990
rect 15750 53952 15752 53961
rect 15804 53952 15806 53961
rect 15750 53887 15806 53896
rect 15476 53576 15528 53582
rect 15476 53518 15528 53524
rect 14464 53440 14516 53446
rect 14464 53382 14516 53388
rect 15752 53440 15804 53446
rect 15752 53382 15804 53388
rect 14372 53100 14424 53106
rect 14372 53042 14424 53048
rect 14004 52964 14056 52970
rect 14004 52906 14056 52912
rect 13636 52692 13688 52698
rect 13636 52634 13688 52640
rect 14016 52601 14044 52906
rect 13634 52592 13690 52601
rect 13634 52527 13636 52536
rect 13688 52527 13690 52536
rect 14002 52592 14058 52601
rect 14002 52527 14058 52536
rect 13636 52498 13688 52504
rect 13360 52420 13412 52426
rect 13360 52362 13412 52368
rect 13372 52154 13400 52362
rect 13360 52148 13412 52154
rect 13360 52090 13412 52096
rect 12950 51708 13258 51717
rect 12950 51706 12956 51708
rect 13012 51706 13036 51708
rect 13092 51706 13116 51708
rect 13172 51706 13196 51708
rect 13252 51706 13258 51708
rect 13012 51654 13014 51706
rect 13194 51654 13196 51706
rect 12950 51652 12956 51654
rect 13012 51652 13036 51654
rect 13092 51652 13116 51654
rect 13172 51652 13196 51654
rect 13252 51652 13258 51654
rect 12950 51643 13258 51652
rect 12950 50620 13258 50629
rect 12950 50618 12956 50620
rect 13012 50618 13036 50620
rect 13092 50618 13116 50620
rect 13172 50618 13196 50620
rect 13252 50618 13258 50620
rect 13012 50566 13014 50618
rect 13194 50566 13196 50618
rect 12950 50564 12956 50566
rect 13012 50564 13036 50566
rect 13092 50564 13116 50566
rect 13172 50564 13196 50566
rect 13252 50564 13258 50566
rect 12950 50555 13258 50564
rect 12950 49532 13258 49541
rect 12950 49530 12956 49532
rect 13012 49530 13036 49532
rect 13092 49530 13116 49532
rect 13172 49530 13196 49532
rect 13252 49530 13258 49532
rect 13012 49478 13014 49530
rect 13194 49478 13196 49530
rect 12950 49476 12956 49478
rect 13012 49476 13036 49478
rect 13092 49476 13116 49478
rect 13172 49476 13196 49478
rect 13252 49476 13258 49478
rect 12950 49467 13258 49476
rect 11980 49428 12032 49434
rect 11980 49370 12032 49376
rect 12808 49428 12860 49434
rect 12808 49370 12860 49376
rect 13452 49224 13504 49230
rect 13452 49166 13504 49172
rect 12950 48444 13258 48453
rect 12950 48442 12956 48444
rect 13012 48442 13036 48444
rect 13092 48442 13116 48444
rect 13172 48442 13196 48444
rect 13252 48442 13258 48444
rect 13012 48390 13014 48442
rect 13194 48390 13196 48442
rect 12950 48388 12956 48390
rect 13012 48388 13036 48390
rect 13092 48388 13116 48390
rect 13172 48388 13196 48390
rect 13252 48388 13258 48390
rect 12950 48379 13258 48388
rect 12716 48272 12768 48278
rect 12716 48214 12768 48220
rect 12164 47116 12216 47122
rect 12164 47058 12216 47064
rect 11888 46708 11940 46714
rect 11888 46650 11940 46656
rect 12176 46510 12204 47058
rect 12440 46912 12492 46918
rect 12440 46854 12492 46860
rect 12164 46504 12216 46510
rect 12164 46446 12216 46452
rect 12176 46034 12204 46446
rect 12164 46028 12216 46034
rect 12164 45970 12216 45976
rect 11796 45484 11848 45490
rect 11796 45426 11848 45432
rect 11808 45393 11836 45426
rect 11794 45384 11850 45393
rect 11794 45319 11850 45328
rect 12072 45280 12124 45286
rect 12072 45222 12124 45228
rect 12084 44266 12112 45222
rect 12176 44470 12204 45970
rect 12452 45898 12480 46854
rect 12440 45892 12492 45898
rect 12440 45834 12492 45840
rect 12440 44532 12492 44538
rect 12440 44474 12492 44480
rect 12164 44464 12216 44470
rect 12164 44406 12216 44412
rect 12072 44260 12124 44266
rect 12072 44202 12124 44208
rect 11704 42356 11756 42362
rect 11704 42298 11756 42304
rect 11520 41812 11572 41818
rect 11520 41754 11572 41760
rect 12084 41682 12112 44202
rect 12176 42770 12204 44406
rect 12164 42764 12216 42770
rect 12164 42706 12216 42712
rect 12348 42764 12400 42770
rect 12348 42706 12400 42712
rect 12176 42650 12204 42706
rect 12176 42622 12296 42650
rect 12164 42288 12216 42294
rect 12164 42230 12216 42236
rect 12072 41676 12124 41682
rect 12072 41618 12124 41624
rect 11428 41608 11480 41614
rect 11428 41550 11480 41556
rect 11256 41386 11376 41414
rect 10876 41268 10928 41274
rect 10876 41210 10928 41216
rect 11060 41268 11112 41274
rect 11164 41262 11284 41290
rect 11060 41210 11112 41216
rect 10876 41132 10928 41138
rect 10876 41074 10928 41080
rect 11060 41132 11112 41138
rect 11060 41074 11112 41080
rect 10888 40934 10916 41074
rect 10876 40928 10928 40934
rect 10876 40870 10928 40876
rect 10888 40662 10916 40870
rect 11072 40730 11100 41074
rect 11060 40724 11112 40730
rect 11060 40666 11112 40672
rect 10876 40656 10928 40662
rect 10876 40598 10928 40604
rect 10784 40112 10836 40118
rect 10784 40054 10836 40060
rect 10692 39092 10744 39098
rect 10692 39034 10744 39040
rect 10968 39024 11020 39030
rect 10968 38966 11020 38972
rect 10876 38888 10928 38894
rect 10876 38830 10928 38836
rect 10692 38208 10744 38214
rect 10692 38150 10744 38156
rect 10600 38004 10652 38010
rect 10600 37946 10652 37952
rect 10704 37942 10732 38150
rect 10508 37936 10560 37942
rect 10508 37878 10560 37884
rect 10692 37936 10744 37942
rect 10692 37878 10744 37884
rect 10416 37460 10468 37466
rect 10416 37402 10468 37408
rect 10324 37324 10376 37330
rect 10324 37266 10376 37272
rect 10520 37194 10548 37878
rect 10598 37360 10654 37369
rect 10704 37346 10732 37878
rect 10704 37318 10824 37346
rect 10598 37295 10600 37304
rect 10652 37295 10654 37304
rect 10600 37266 10652 37272
rect 10508 37188 10560 37194
rect 10428 37148 10508 37176
rect 10138 36816 10194 36825
rect 10138 36751 10194 36760
rect 9956 36372 10008 36378
rect 9956 36314 10008 36320
rect 9772 35624 9824 35630
rect 9772 35566 9824 35572
rect 9784 34202 9812 35566
rect 9864 35488 9916 35494
rect 9864 35430 9916 35436
rect 9876 35086 9904 35430
rect 9864 35080 9916 35086
rect 9864 35022 9916 35028
rect 9876 34746 9904 35022
rect 9864 34740 9916 34746
rect 9864 34682 9916 34688
rect 9772 34196 9824 34202
rect 9772 34138 9824 34144
rect 9772 33448 9824 33454
rect 9772 33390 9824 33396
rect 9784 32910 9812 33390
rect 9956 33040 10008 33046
rect 9956 32982 10008 32988
rect 9772 32904 9824 32910
rect 9772 32846 9824 32852
rect 9772 32768 9824 32774
rect 9772 32710 9824 32716
rect 9680 32564 9732 32570
rect 9680 32506 9732 32512
rect 9588 32496 9640 32502
rect 9588 32438 9640 32444
rect 9600 32230 9628 32438
rect 9588 32224 9640 32230
rect 9588 32166 9640 32172
rect 9404 31884 9456 31890
rect 9404 31826 9456 31832
rect 9496 31884 9548 31890
rect 9496 31826 9548 31832
rect 9508 31754 9536 31826
rect 9416 31726 9536 31754
rect 9416 31346 9444 31726
rect 9404 31340 9456 31346
rect 9404 31282 9456 31288
rect 9692 29714 9720 32506
rect 9680 29708 9732 29714
rect 9680 29650 9732 29656
rect 9784 29306 9812 32710
rect 9864 32224 9916 32230
rect 9864 32166 9916 32172
rect 9876 31890 9904 32166
rect 9968 32026 9996 32982
rect 9956 32020 10008 32026
rect 9956 31962 10008 31968
rect 9864 31884 9916 31890
rect 9864 31826 9916 31832
rect 9968 31754 9996 31962
rect 9876 31726 9996 31754
rect 8944 29300 8996 29306
rect 8944 29242 8996 29248
rect 9220 29300 9272 29306
rect 9220 29242 9272 29248
rect 9772 29300 9824 29306
rect 9772 29242 9824 29248
rect 8852 26920 8904 26926
rect 8852 26862 8904 26868
rect 8668 26580 8720 26586
rect 8668 26522 8720 26528
rect 8680 26382 8708 26522
rect 8668 26376 8720 26382
rect 8668 26318 8720 26324
rect 8680 26042 8708 26318
rect 8668 26036 8720 26042
rect 8668 25978 8720 25984
rect 8668 24812 8720 24818
rect 8668 24754 8720 24760
rect 8576 24404 8628 24410
rect 8576 24346 8628 24352
rect 8484 24336 8536 24342
rect 8484 24278 8536 24284
rect 7950 23964 8258 23973
rect 7950 23962 7956 23964
rect 8012 23962 8036 23964
rect 8092 23962 8116 23964
rect 8172 23962 8196 23964
rect 8252 23962 8258 23964
rect 8012 23910 8014 23962
rect 8194 23910 8196 23962
rect 7950 23908 7956 23910
rect 8012 23908 8036 23910
rect 8092 23908 8116 23910
rect 8172 23908 8196 23910
rect 8252 23908 8258 23910
rect 7950 23899 8258 23908
rect 8496 23866 8524 24278
rect 8680 24274 8708 24754
rect 8760 24744 8812 24750
rect 8760 24686 8812 24692
rect 8668 24268 8720 24274
rect 8668 24210 8720 24216
rect 8484 23860 8536 23866
rect 8484 23802 8536 23808
rect 7840 23520 7892 23526
rect 7840 23462 7892 23468
rect 7748 23316 7800 23322
rect 7748 23258 7800 23264
rect 7760 22778 7788 23258
rect 7748 22772 7800 22778
rect 7748 22714 7800 22720
rect 7852 22642 7880 23462
rect 8496 23322 8524 23802
rect 8484 23316 8536 23322
rect 8484 23258 8536 23264
rect 8496 23050 8524 23258
rect 8484 23044 8536 23050
rect 8484 22986 8536 22992
rect 7950 22876 8258 22885
rect 7950 22874 7956 22876
rect 8012 22874 8036 22876
rect 8092 22874 8116 22876
rect 8172 22874 8196 22876
rect 8252 22874 8258 22876
rect 8012 22822 8014 22874
rect 8194 22822 8196 22874
rect 7950 22820 7956 22822
rect 8012 22820 8036 22822
rect 8092 22820 8116 22822
rect 8172 22820 8196 22822
rect 8252 22820 8258 22822
rect 7950 22811 8258 22820
rect 8116 22772 8168 22778
rect 8116 22714 8168 22720
rect 7840 22636 7892 22642
rect 7840 22578 7892 22584
rect 7748 22432 7800 22438
rect 7748 22374 7800 22380
rect 7656 22024 7708 22030
rect 7656 21966 7708 21972
rect 7760 21622 7788 22374
rect 7748 21616 7800 21622
rect 7748 21558 7800 21564
rect 7852 21554 7880 22578
rect 8128 22098 8156 22714
rect 8116 22092 8168 22098
rect 8116 22034 8168 22040
rect 8128 21876 8156 22034
rect 8772 22030 8800 24686
rect 8852 23044 8904 23050
rect 8852 22986 8904 22992
rect 8864 22166 8892 22986
rect 8852 22160 8904 22166
rect 8852 22102 8904 22108
rect 8392 22024 8444 22030
rect 8392 21966 8444 21972
rect 8760 22024 8812 22030
rect 8760 21966 8812 21972
rect 8404 21894 8432 21966
rect 8392 21888 8444 21894
rect 8128 21848 8340 21876
rect 7950 21788 8258 21797
rect 7950 21786 7956 21788
rect 8012 21786 8036 21788
rect 8092 21786 8116 21788
rect 8172 21786 8196 21788
rect 8252 21786 8258 21788
rect 8012 21734 8014 21786
rect 8194 21734 8196 21786
rect 7950 21732 7956 21734
rect 8012 21732 8036 21734
rect 8092 21732 8116 21734
rect 8172 21732 8196 21734
rect 8252 21732 8258 21734
rect 7950 21723 8258 21732
rect 8312 21672 8340 21848
rect 8392 21830 8444 21836
rect 8220 21644 8340 21672
rect 7840 21548 7892 21554
rect 7840 21490 7892 21496
rect 7564 21140 7616 21146
rect 7564 21082 7616 21088
rect 7484 20998 7696 21026
rect 8220 21010 8248 21644
rect 7564 19984 7616 19990
rect 7564 19926 7616 19932
rect 7380 18216 7432 18222
rect 7380 18158 7432 18164
rect 7392 3738 7420 18158
rect 7472 18080 7524 18086
rect 7472 18022 7524 18028
rect 7484 17338 7512 18022
rect 7576 17746 7604 19926
rect 7564 17740 7616 17746
rect 7564 17682 7616 17688
rect 7472 17332 7524 17338
rect 7472 17274 7524 17280
rect 7668 16574 7696 20998
rect 8208 21004 8260 21010
rect 8208 20946 8260 20952
rect 7950 20700 8258 20709
rect 7950 20698 7956 20700
rect 8012 20698 8036 20700
rect 8092 20698 8116 20700
rect 8172 20698 8196 20700
rect 8252 20698 8258 20700
rect 8012 20646 8014 20698
rect 8194 20646 8196 20698
rect 7950 20644 7956 20646
rect 8012 20644 8036 20646
rect 8092 20644 8116 20646
rect 8172 20644 8196 20646
rect 8252 20644 8258 20646
rect 7950 20635 8258 20644
rect 7748 20256 7800 20262
rect 7748 20198 7800 20204
rect 7760 19922 7788 20198
rect 7748 19916 7800 19922
rect 7748 19858 7800 19864
rect 7950 19612 8258 19621
rect 7950 19610 7956 19612
rect 8012 19610 8036 19612
rect 8092 19610 8116 19612
rect 8172 19610 8196 19612
rect 8252 19610 8258 19612
rect 8012 19558 8014 19610
rect 8194 19558 8196 19610
rect 7950 19556 7956 19558
rect 8012 19556 8036 19558
rect 8092 19556 8116 19558
rect 8172 19556 8196 19558
rect 8252 19556 8258 19558
rect 7950 19547 8258 19556
rect 7950 18524 8258 18533
rect 7950 18522 7956 18524
rect 8012 18522 8036 18524
rect 8092 18522 8116 18524
rect 8172 18522 8196 18524
rect 8252 18522 8258 18524
rect 8012 18470 8014 18522
rect 8194 18470 8196 18522
rect 7950 18468 7956 18470
rect 8012 18468 8036 18470
rect 8092 18468 8116 18470
rect 8172 18468 8196 18470
rect 8252 18468 8258 18470
rect 7950 18459 8258 18468
rect 7748 17740 7800 17746
rect 7748 17682 7800 17688
rect 7760 17270 7788 17682
rect 7950 17436 8258 17445
rect 7950 17434 7956 17436
rect 8012 17434 8036 17436
rect 8092 17434 8116 17436
rect 8172 17434 8196 17436
rect 8252 17434 8258 17436
rect 8012 17382 8014 17434
rect 8194 17382 8196 17434
rect 7950 17380 7956 17382
rect 8012 17380 8036 17382
rect 8092 17380 8116 17382
rect 8172 17380 8196 17382
rect 8252 17380 8258 17382
rect 7950 17371 8258 17380
rect 7748 17264 7800 17270
rect 7748 17206 7800 17212
rect 7760 16658 7788 17206
rect 7840 17060 7892 17066
rect 7840 17002 7892 17008
rect 7748 16652 7800 16658
rect 7748 16594 7800 16600
rect 7576 16546 7696 16574
rect 7472 9512 7524 9518
rect 7472 9454 7524 9460
rect 7484 8974 7512 9454
rect 7472 8968 7524 8974
rect 7472 8910 7524 8916
rect 7380 3732 7432 3738
rect 7380 3674 7432 3680
rect 7012 3188 7064 3194
rect 7012 3130 7064 3136
rect 7288 3188 7340 3194
rect 7288 3130 7340 3136
rect 6828 3052 6880 3058
rect 6828 2994 6880 3000
rect 6460 2848 6512 2854
rect 6460 2790 6512 2796
rect 6472 800 6500 2790
rect 6840 800 6868 2994
rect 7576 2582 7604 16546
rect 7748 15972 7800 15978
rect 7748 15914 7800 15920
rect 7656 15360 7708 15366
rect 7656 15302 7708 15308
rect 7668 15094 7696 15302
rect 7656 15088 7708 15094
rect 7656 15030 7708 15036
rect 7656 9580 7708 9586
rect 7656 9522 7708 9528
rect 7668 2650 7696 9522
rect 7760 2990 7788 15914
rect 7852 15162 7880 17002
rect 7932 16788 7984 16794
rect 7932 16730 7984 16736
rect 7944 16522 7972 16730
rect 8404 16574 8432 21830
rect 8864 21622 8892 22102
rect 8852 21616 8904 21622
rect 8852 21558 8904 21564
rect 8484 21344 8536 21350
rect 8484 21286 8536 21292
rect 8496 19854 8524 21286
rect 8484 19848 8536 19854
rect 8484 19790 8536 19796
rect 8864 19446 8892 21558
rect 8956 20602 8984 29242
rect 9232 29170 9260 29242
rect 9220 29164 9272 29170
rect 9220 29106 9272 29112
rect 9680 29028 9732 29034
rect 9680 28970 9732 28976
rect 9128 28552 9180 28558
rect 9180 28512 9260 28540
rect 9128 28494 9180 28500
rect 9232 28014 9260 28512
rect 9404 28484 9456 28490
rect 9404 28426 9456 28432
rect 9416 28218 9444 28426
rect 9588 28416 9640 28422
rect 9588 28358 9640 28364
rect 9404 28212 9456 28218
rect 9404 28154 9456 28160
rect 9220 28008 9272 28014
rect 9220 27950 9272 27956
rect 9128 27396 9180 27402
rect 9128 27338 9180 27344
rect 9140 27130 9168 27338
rect 9128 27124 9180 27130
rect 9128 27066 9180 27072
rect 9232 25362 9260 27950
rect 9496 27328 9548 27334
rect 9496 27270 9548 27276
rect 9508 27130 9536 27270
rect 9496 27124 9548 27130
rect 9496 27066 9548 27072
rect 9312 26376 9364 26382
rect 9312 26318 9364 26324
rect 9324 25702 9352 26318
rect 9312 25696 9364 25702
rect 9312 25638 9364 25644
rect 9220 25356 9272 25362
rect 9220 25298 9272 25304
rect 9324 24886 9352 25638
rect 9312 24880 9364 24886
rect 9312 24822 9364 24828
rect 9404 24744 9456 24750
rect 9404 24686 9456 24692
rect 9128 24064 9180 24070
rect 9128 24006 9180 24012
rect 9036 23520 9088 23526
rect 9036 23462 9088 23468
rect 8944 20596 8996 20602
rect 8944 20538 8996 20544
rect 8668 19440 8720 19446
rect 8668 19382 8720 19388
rect 8852 19440 8904 19446
rect 8852 19382 8904 19388
rect 8576 19168 8628 19174
rect 8576 19110 8628 19116
rect 8588 18970 8616 19110
rect 8576 18964 8628 18970
rect 8576 18906 8628 18912
rect 8484 16992 8536 16998
rect 8484 16934 8536 16940
rect 8496 16794 8524 16934
rect 8484 16788 8536 16794
rect 8484 16730 8536 16736
rect 8312 16546 8432 16574
rect 8588 16574 8616 18906
rect 8680 18834 8708 19382
rect 8668 18828 8720 18834
rect 8668 18770 8720 18776
rect 8956 16658 8984 20538
rect 9048 18222 9076 23462
rect 9140 21146 9168 24006
rect 9312 23792 9364 23798
rect 9312 23734 9364 23740
rect 9220 22500 9272 22506
rect 9220 22442 9272 22448
rect 9128 21140 9180 21146
rect 9128 21082 9180 21088
rect 9232 20618 9260 22442
rect 9140 20590 9260 20618
rect 9324 20602 9352 23734
rect 9416 22098 9444 24686
rect 9600 24342 9628 28358
rect 9692 25106 9720 28970
rect 9876 26908 9904 31726
rect 9956 30592 10008 30598
rect 9956 30534 10008 30540
rect 9968 29714 9996 30534
rect 9956 29708 10008 29714
rect 9956 29650 10008 29656
rect 10152 29034 10180 36751
rect 10324 36372 10376 36378
rect 10324 36314 10376 36320
rect 10232 36032 10284 36038
rect 10232 35974 10284 35980
rect 10244 34202 10272 35974
rect 10232 34196 10284 34202
rect 10232 34138 10284 34144
rect 10232 32428 10284 32434
rect 10232 32370 10284 32376
rect 10244 32298 10272 32370
rect 10232 32292 10284 32298
rect 10232 32234 10284 32240
rect 10336 30274 10364 36314
rect 10244 30246 10364 30274
rect 10140 29028 10192 29034
rect 10140 28970 10192 28976
rect 9876 26880 10180 26908
rect 10048 26784 10100 26790
rect 10048 26726 10100 26732
rect 9772 26240 9824 26246
rect 9772 26182 9824 26188
rect 9784 25226 9812 26182
rect 9864 25356 9916 25362
rect 9864 25298 9916 25304
rect 9772 25220 9824 25226
rect 9772 25162 9824 25168
rect 9692 25078 9812 25106
rect 9588 24336 9640 24342
rect 9588 24278 9640 24284
rect 9600 23866 9628 24278
rect 9680 24132 9732 24138
rect 9680 24074 9732 24080
rect 9692 23866 9720 24074
rect 9588 23860 9640 23866
rect 9588 23802 9640 23808
rect 9680 23860 9732 23866
rect 9680 23802 9732 23808
rect 9588 23724 9640 23730
rect 9588 23666 9640 23672
rect 9600 23118 9628 23666
rect 9784 23526 9812 25078
rect 9876 24290 9904 25298
rect 9956 24948 10008 24954
rect 9956 24890 10008 24896
rect 9968 24410 9996 24890
rect 9956 24404 10008 24410
rect 9956 24346 10008 24352
rect 9876 24274 9996 24290
rect 9876 24268 10008 24274
rect 9876 24262 9956 24268
rect 9956 24210 10008 24216
rect 9864 23656 9916 23662
rect 9864 23598 9916 23604
rect 9772 23520 9824 23526
rect 9772 23462 9824 23468
rect 9588 23112 9640 23118
rect 9588 23054 9640 23060
rect 9772 22772 9824 22778
rect 9772 22714 9824 22720
rect 9404 22092 9456 22098
rect 9404 22034 9456 22040
rect 9416 21078 9444 22034
rect 9588 21888 9640 21894
rect 9588 21830 9640 21836
rect 9496 21412 9548 21418
rect 9496 21354 9548 21360
rect 9404 21072 9456 21078
rect 9404 21014 9456 21020
rect 9416 20942 9444 21014
rect 9404 20936 9456 20942
rect 9404 20878 9456 20884
rect 9508 20754 9536 21354
rect 9416 20726 9536 20754
rect 9312 20596 9364 20602
rect 9036 18216 9088 18222
rect 9036 18158 9088 18164
rect 9036 18080 9088 18086
rect 9036 18022 9088 18028
rect 9048 17678 9076 18022
rect 9036 17672 9088 17678
rect 9036 17614 9088 17620
rect 9140 17202 9168 20590
rect 9312 20538 9364 20544
rect 9416 20534 9444 20726
rect 9496 20596 9548 20602
rect 9496 20538 9548 20544
rect 9404 20528 9456 20534
rect 9404 20470 9456 20476
rect 9220 20460 9272 20466
rect 9220 20402 9272 20408
rect 9232 17338 9260 20402
rect 9312 20324 9364 20330
rect 9312 20266 9364 20272
rect 9324 17626 9352 20266
rect 9404 19916 9456 19922
rect 9404 19858 9456 19864
rect 9416 19258 9444 19858
rect 9508 19854 9536 20538
rect 9496 19848 9548 19854
rect 9496 19790 9548 19796
rect 9508 19334 9536 19790
rect 9600 19530 9628 21830
rect 9600 19514 9720 19530
rect 9600 19508 9732 19514
rect 9600 19502 9680 19508
rect 9680 19450 9732 19456
rect 9508 19306 9628 19334
rect 9416 19230 9536 19258
rect 9404 18284 9456 18290
rect 9404 18226 9456 18232
rect 9416 17746 9444 18226
rect 9508 18222 9536 19230
rect 9496 18216 9548 18222
rect 9496 18158 9548 18164
rect 9404 17740 9456 17746
rect 9404 17682 9456 17688
rect 9324 17598 9444 17626
rect 9312 17536 9364 17542
rect 9312 17478 9364 17484
rect 9220 17332 9272 17338
rect 9220 17274 9272 17280
rect 9128 17196 9180 17202
rect 9128 17138 9180 17144
rect 9324 17134 9352 17478
rect 9312 17128 9364 17134
rect 9048 17076 9312 17082
rect 9048 17070 9364 17076
rect 9048 17054 9352 17070
rect 8944 16652 8996 16658
rect 8944 16594 8996 16600
rect 8588 16546 8708 16574
rect 7932 16516 7984 16522
rect 7932 16458 7984 16464
rect 7950 16348 8258 16357
rect 7950 16346 7956 16348
rect 8012 16346 8036 16348
rect 8092 16346 8116 16348
rect 8172 16346 8196 16348
rect 8252 16346 8258 16348
rect 8012 16294 8014 16346
rect 8194 16294 8196 16346
rect 7950 16292 7956 16294
rect 8012 16292 8036 16294
rect 8092 16292 8116 16294
rect 8172 16292 8196 16294
rect 8252 16292 8258 16294
rect 7950 16283 8258 16292
rect 8208 16108 8260 16114
rect 8208 16050 8260 16056
rect 8220 15706 8248 16050
rect 8208 15700 8260 15706
rect 8208 15642 8260 15648
rect 7950 15260 8258 15269
rect 7950 15258 7956 15260
rect 8012 15258 8036 15260
rect 8092 15258 8116 15260
rect 8172 15258 8196 15260
rect 8252 15258 8258 15260
rect 8012 15206 8014 15258
rect 8194 15206 8196 15258
rect 7950 15204 7956 15206
rect 8012 15204 8036 15206
rect 8092 15204 8116 15206
rect 8172 15204 8196 15206
rect 8252 15204 8258 15206
rect 7950 15195 8258 15204
rect 7840 15156 7892 15162
rect 7840 15098 7892 15104
rect 7950 14172 8258 14181
rect 7950 14170 7956 14172
rect 8012 14170 8036 14172
rect 8092 14170 8116 14172
rect 8172 14170 8196 14172
rect 8252 14170 8258 14172
rect 8012 14118 8014 14170
rect 8194 14118 8196 14170
rect 7950 14116 7956 14118
rect 8012 14116 8036 14118
rect 8092 14116 8116 14118
rect 8172 14116 8196 14118
rect 8252 14116 8258 14118
rect 7950 14107 8258 14116
rect 7950 13084 8258 13093
rect 7950 13082 7956 13084
rect 8012 13082 8036 13084
rect 8092 13082 8116 13084
rect 8172 13082 8196 13084
rect 8252 13082 8258 13084
rect 8012 13030 8014 13082
rect 8194 13030 8196 13082
rect 7950 13028 7956 13030
rect 8012 13028 8036 13030
rect 8092 13028 8116 13030
rect 8172 13028 8196 13030
rect 8252 13028 8258 13030
rect 7950 13019 8258 13028
rect 7950 11996 8258 12005
rect 7950 11994 7956 11996
rect 8012 11994 8036 11996
rect 8092 11994 8116 11996
rect 8172 11994 8196 11996
rect 8252 11994 8258 11996
rect 8012 11942 8014 11994
rect 8194 11942 8196 11994
rect 7950 11940 7956 11942
rect 8012 11940 8036 11942
rect 8092 11940 8116 11942
rect 8172 11940 8196 11942
rect 8252 11940 8258 11942
rect 7950 11931 8258 11940
rect 7950 10908 8258 10917
rect 7950 10906 7956 10908
rect 8012 10906 8036 10908
rect 8092 10906 8116 10908
rect 8172 10906 8196 10908
rect 8252 10906 8258 10908
rect 8012 10854 8014 10906
rect 8194 10854 8196 10906
rect 7950 10852 7956 10854
rect 8012 10852 8036 10854
rect 8092 10852 8116 10854
rect 8172 10852 8196 10854
rect 8252 10852 8258 10854
rect 7950 10843 8258 10852
rect 7950 9820 8258 9829
rect 7950 9818 7956 9820
rect 8012 9818 8036 9820
rect 8092 9818 8116 9820
rect 8172 9818 8196 9820
rect 8252 9818 8258 9820
rect 8012 9766 8014 9818
rect 8194 9766 8196 9818
rect 7950 9764 7956 9766
rect 8012 9764 8036 9766
rect 8092 9764 8116 9766
rect 8172 9764 8196 9766
rect 8252 9764 8258 9766
rect 7950 9755 8258 9764
rect 7950 8732 8258 8741
rect 7950 8730 7956 8732
rect 8012 8730 8036 8732
rect 8092 8730 8116 8732
rect 8172 8730 8196 8732
rect 8252 8730 8258 8732
rect 8012 8678 8014 8730
rect 8194 8678 8196 8730
rect 7950 8676 7956 8678
rect 8012 8676 8036 8678
rect 8092 8676 8116 8678
rect 8172 8676 8196 8678
rect 8252 8676 8258 8678
rect 7950 8667 8258 8676
rect 7950 7644 8258 7653
rect 7950 7642 7956 7644
rect 8012 7642 8036 7644
rect 8092 7642 8116 7644
rect 8172 7642 8196 7644
rect 8252 7642 8258 7644
rect 8012 7590 8014 7642
rect 8194 7590 8196 7642
rect 7950 7588 7956 7590
rect 8012 7588 8036 7590
rect 8092 7588 8116 7590
rect 8172 7588 8196 7590
rect 8252 7588 8258 7590
rect 7950 7579 8258 7588
rect 7950 6556 8258 6565
rect 7950 6554 7956 6556
rect 8012 6554 8036 6556
rect 8092 6554 8116 6556
rect 8172 6554 8196 6556
rect 8252 6554 8258 6556
rect 8012 6502 8014 6554
rect 8194 6502 8196 6554
rect 7950 6500 7956 6502
rect 8012 6500 8036 6502
rect 8092 6500 8116 6502
rect 8172 6500 8196 6502
rect 8252 6500 8258 6502
rect 7950 6491 8258 6500
rect 7950 5468 8258 5477
rect 7950 5466 7956 5468
rect 8012 5466 8036 5468
rect 8092 5466 8116 5468
rect 8172 5466 8196 5468
rect 8252 5466 8258 5468
rect 8012 5414 8014 5466
rect 8194 5414 8196 5466
rect 7950 5412 7956 5414
rect 8012 5412 8036 5414
rect 8092 5412 8116 5414
rect 8172 5412 8196 5414
rect 8252 5412 8258 5414
rect 7950 5403 8258 5412
rect 7950 4380 8258 4389
rect 7950 4378 7956 4380
rect 8012 4378 8036 4380
rect 8092 4378 8116 4380
rect 8172 4378 8196 4380
rect 8252 4378 8258 4380
rect 8012 4326 8014 4378
rect 8194 4326 8196 4378
rect 7950 4324 7956 4326
rect 8012 4324 8036 4326
rect 8092 4324 8116 4326
rect 8172 4324 8196 4326
rect 8252 4324 8258 4326
rect 7950 4315 8258 4324
rect 8312 4282 8340 16546
rect 8484 16448 8536 16454
rect 8484 16390 8536 16396
rect 8392 15904 8444 15910
rect 8392 15846 8444 15852
rect 8404 15094 8432 15846
rect 8496 15434 8524 16390
rect 8576 15564 8628 15570
rect 8576 15506 8628 15512
rect 8484 15428 8536 15434
rect 8484 15370 8536 15376
rect 8392 15088 8444 15094
rect 8392 15030 8444 15036
rect 8496 14958 8524 15370
rect 8484 14952 8536 14958
rect 8484 14894 8536 14900
rect 8392 14816 8444 14822
rect 8392 14758 8444 14764
rect 8404 13734 8432 14758
rect 8588 14618 8616 15506
rect 8576 14612 8628 14618
rect 8576 14554 8628 14560
rect 8680 14278 8708 16546
rect 9048 15502 9076 17054
rect 9416 16980 9444 17598
rect 9232 16952 9444 16980
rect 9232 16590 9260 16952
rect 9600 16810 9628 19306
rect 9680 18624 9732 18630
rect 9680 18566 9732 18572
rect 9324 16782 9628 16810
rect 9220 16584 9272 16590
rect 9324 16574 9352 16782
rect 9588 16652 9640 16658
rect 9588 16594 9640 16600
rect 9324 16546 9444 16574
rect 9220 16526 9272 16532
rect 9128 16448 9180 16454
rect 9128 16390 9180 16396
rect 9140 16250 9168 16390
rect 9128 16244 9180 16250
rect 9128 16186 9180 16192
rect 9036 15496 9088 15502
rect 9036 15438 9088 15444
rect 8760 15428 8812 15434
rect 8760 15370 8812 15376
rect 8668 14272 8720 14278
rect 8668 14214 8720 14220
rect 8484 13864 8536 13870
rect 8484 13806 8536 13812
rect 8392 13728 8444 13734
rect 8392 13670 8444 13676
rect 8496 13530 8524 13806
rect 8484 13524 8536 13530
rect 8484 13466 8536 13472
rect 8772 12850 8800 15370
rect 8852 13728 8904 13734
rect 8852 13670 8904 13676
rect 8760 12844 8812 12850
rect 8760 12786 8812 12792
rect 8864 12782 8892 13670
rect 8852 12776 8904 12782
rect 8852 12718 8904 12724
rect 9048 9042 9076 15438
rect 9128 15360 9180 15366
rect 9128 15302 9180 15308
rect 9140 12918 9168 15302
rect 9128 12912 9180 12918
rect 9128 12854 9180 12860
rect 9036 9036 9088 9042
rect 9036 8978 9088 8984
rect 9312 5704 9364 5710
rect 9312 5646 9364 5652
rect 8300 4276 8352 4282
rect 8300 4218 8352 4224
rect 8482 4176 8538 4185
rect 8482 4111 8538 4120
rect 8300 3596 8352 3602
rect 8300 3538 8352 3544
rect 7840 3392 7892 3398
rect 7840 3334 7892 3340
rect 7748 2984 7800 2990
rect 7748 2926 7800 2932
rect 7656 2644 7708 2650
rect 7656 2586 7708 2592
rect 7564 2576 7616 2582
rect 7564 2518 7616 2524
rect 7196 2440 7248 2446
rect 7196 2382 7248 2388
rect 7564 2440 7616 2446
rect 7564 2382 7616 2388
rect 7208 800 7236 2382
rect 7576 800 7604 2382
rect 7852 1986 7880 3334
rect 7950 3292 8258 3301
rect 7950 3290 7956 3292
rect 8012 3290 8036 3292
rect 8092 3290 8116 3292
rect 8172 3290 8196 3292
rect 8252 3290 8258 3292
rect 8012 3238 8014 3290
rect 8194 3238 8196 3290
rect 7950 3236 7956 3238
rect 8012 3236 8036 3238
rect 8092 3236 8116 3238
rect 8172 3236 8196 3238
rect 8252 3236 8258 3238
rect 7950 3227 8258 3236
rect 8208 3052 8260 3058
rect 8312 3040 8340 3538
rect 8496 3194 8524 4111
rect 9036 4004 9088 4010
rect 9036 3946 9088 3952
rect 8668 3392 8720 3398
rect 8668 3334 8720 3340
rect 8484 3188 8536 3194
rect 8484 3130 8536 3136
rect 8680 3058 8708 3334
rect 8260 3012 8340 3040
rect 8208 2994 8260 3000
rect 7950 2204 8258 2213
rect 7950 2202 7956 2204
rect 8012 2202 8036 2204
rect 8092 2202 8116 2204
rect 8172 2202 8196 2204
rect 8252 2202 8258 2204
rect 8012 2150 8014 2202
rect 8194 2150 8196 2202
rect 7950 2148 7956 2150
rect 8012 2148 8036 2150
rect 8092 2148 8116 2150
rect 8172 2148 8196 2150
rect 8252 2148 8258 2150
rect 7950 2139 8258 2148
rect 7852 1958 7972 1986
rect 7944 800 7972 1958
rect 8312 800 8340 3012
rect 8668 3052 8720 3058
rect 8668 2994 8720 3000
rect 8680 800 8708 2994
rect 9048 2990 9076 3946
rect 9324 3058 9352 5646
rect 9416 5642 9444 16546
rect 9600 16538 9628 16594
rect 9508 16510 9628 16538
rect 9508 12442 9536 16510
rect 9588 16448 9640 16454
rect 9588 16390 9640 16396
rect 9600 16250 9628 16390
rect 9588 16244 9640 16250
rect 9588 16186 9640 16192
rect 9692 14346 9720 18566
rect 9680 14340 9732 14346
rect 9680 14282 9732 14288
rect 9588 12776 9640 12782
rect 9588 12718 9640 12724
rect 9496 12436 9548 12442
rect 9496 12378 9548 12384
rect 9600 12306 9628 12718
rect 9588 12300 9640 12306
rect 9588 12242 9640 12248
rect 9496 8900 9548 8906
rect 9496 8842 9548 8848
rect 9404 5636 9456 5642
rect 9404 5578 9456 5584
rect 9404 3936 9456 3942
rect 9404 3878 9456 3884
rect 9416 3534 9444 3878
rect 9508 3738 9536 8842
rect 9784 6322 9812 22714
rect 9876 21434 9904 23598
rect 9968 23186 9996 24210
rect 9956 23180 10008 23186
rect 9956 23122 10008 23128
rect 9956 21480 10008 21486
rect 9876 21428 9956 21434
rect 9876 21422 10008 21428
rect 9876 21406 9996 21422
rect 9876 20398 9904 21406
rect 9864 20392 9916 20398
rect 9864 20334 9916 20340
rect 9876 19174 9904 20334
rect 9864 19168 9916 19174
rect 9864 19110 9916 19116
rect 9876 18222 9904 19110
rect 10060 18426 10088 26726
rect 10152 20058 10180 26880
rect 10244 26586 10272 30246
rect 10324 30184 10376 30190
rect 10428 30172 10456 37148
rect 10508 37130 10560 37136
rect 10692 37188 10744 37194
rect 10692 37130 10744 37136
rect 10704 34066 10732 37130
rect 10796 36854 10824 37318
rect 10784 36848 10836 36854
rect 10784 36790 10836 36796
rect 10692 34060 10744 34066
rect 10692 34002 10744 34008
rect 10508 33856 10560 33862
rect 10508 33798 10560 33804
rect 10520 30938 10548 33798
rect 10888 33114 10916 38830
rect 10980 38418 11008 38966
rect 10968 38412 11020 38418
rect 10968 38354 11020 38360
rect 10968 38208 11020 38214
rect 10968 38150 11020 38156
rect 10980 38010 11008 38150
rect 10968 38004 11020 38010
rect 10968 37946 11020 37952
rect 10968 37460 11020 37466
rect 10968 37402 11020 37408
rect 10980 37330 11008 37402
rect 10968 37324 11020 37330
rect 10968 37266 11020 37272
rect 11072 36922 11100 40666
rect 11256 38400 11284 41262
rect 11348 40050 11376 41386
rect 11336 40044 11388 40050
rect 11336 39986 11388 39992
rect 11164 38372 11284 38400
rect 11164 37262 11192 38372
rect 11244 38276 11296 38282
rect 11244 38218 11296 38224
rect 11152 37256 11204 37262
rect 11152 37198 11204 37204
rect 11152 37120 11204 37126
rect 11152 37062 11204 37068
rect 11060 36916 11112 36922
rect 11060 36858 11112 36864
rect 11072 36378 11100 36858
rect 11060 36372 11112 36378
rect 11060 36314 11112 36320
rect 11072 36174 11100 36314
rect 11060 36168 11112 36174
rect 11060 36110 11112 36116
rect 11060 35284 11112 35290
rect 11060 35226 11112 35232
rect 11072 34746 11100 35226
rect 11060 34740 11112 34746
rect 11060 34682 11112 34688
rect 11060 34468 11112 34474
rect 11060 34410 11112 34416
rect 10968 33652 11020 33658
rect 10968 33594 11020 33600
rect 10876 33108 10928 33114
rect 10876 33050 10928 33056
rect 10980 32774 11008 33594
rect 10968 32768 11020 32774
rect 10968 32710 11020 32716
rect 10692 32428 10744 32434
rect 10692 32370 10744 32376
rect 10508 30932 10560 30938
rect 10508 30874 10560 30880
rect 10376 30144 10456 30172
rect 10324 30126 10376 30132
rect 10232 26580 10284 26586
rect 10232 26522 10284 26528
rect 10244 24834 10272 26522
rect 10336 25378 10364 30126
rect 10508 29708 10560 29714
rect 10508 29650 10560 29656
rect 10520 28014 10548 29650
rect 10704 29102 10732 32370
rect 11072 31754 11100 34410
rect 10980 31726 11100 31754
rect 10980 31278 11008 31726
rect 11060 31408 11112 31414
rect 11060 31350 11112 31356
rect 10968 31272 11020 31278
rect 10968 31214 11020 31220
rect 10876 30864 10928 30870
rect 10876 30806 10928 30812
rect 10888 30326 10916 30806
rect 10876 30320 10928 30326
rect 10876 30262 10928 30268
rect 10692 29096 10744 29102
rect 10692 29038 10744 29044
rect 10784 29028 10836 29034
rect 10784 28970 10836 28976
rect 10508 28008 10560 28014
rect 10508 27950 10560 27956
rect 10692 26852 10744 26858
rect 10692 26794 10744 26800
rect 10508 25900 10560 25906
rect 10508 25842 10560 25848
rect 10520 25498 10548 25842
rect 10704 25838 10732 26794
rect 10796 26042 10824 28970
rect 10888 28762 10916 30262
rect 10980 30190 11008 31214
rect 10968 30184 11020 30190
rect 10968 30126 11020 30132
rect 11072 29646 11100 31350
rect 11060 29640 11112 29646
rect 11060 29582 11112 29588
rect 11072 29306 11100 29582
rect 11060 29300 11112 29306
rect 11060 29242 11112 29248
rect 11072 28994 11100 29242
rect 10980 28966 11100 28994
rect 10968 28960 11020 28966
rect 10968 28902 11020 28908
rect 10876 28756 10928 28762
rect 10876 28698 10928 28704
rect 10888 26926 10916 28698
rect 10980 28490 11008 28902
rect 10968 28484 11020 28490
rect 10968 28426 11020 28432
rect 10980 28150 11008 28426
rect 11060 28416 11112 28422
rect 11060 28358 11112 28364
rect 10968 28144 11020 28150
rect 10968 28086 11020 28092
rect 10980 27674 11008 28086
rect 11072 27878 11100 28358
rect 11060 27872 11112 27878
rect 11060 27814 11112 27820
rect 10968 27668 11020 27674
rect 10968 27610 11020 27616
rect 10968 26988 11020 26994
rect 10968 26930 11020 26936
rect 10876 26920 10928 26926
rect 10876 26862 10928 26868
rect 10784 26036 10836 26042
rect 10784 25978 10836 25984
rect 10692 25832 10744 25838
rect 10692 25774 10744 25780
rect 10692 25696 10744 25702
rect 10692 25638 10744 25644
rect 10508 25492 10560 25498
rect 10508 25434 10560 25440
rect 10600 25492 10652 25498
rect 10600 25434 10652 25440
rect 10336 25350 10548 25378
rect 10244 24806 10456 24834
rect 10324 24744 10376 24750
rect 10324 24686 10376 24692
rect 10232 23044 10284 23050
rect 10232 22986 10284 22992
rect 10244 22710 10272 22986
rect 10232 22704 10284 22710
rect 10232 22646 10284 22652
rect 10232 20800 10284 20806
rect 10232 20742 10284 20748
rect 10140 20052 10192 20058
rect 10140 19994 10192 20000
rect 10244 19990 10272 20742
rect 10232 19984 10284 19990
rect 10232 19926 10284 19932
rect 10336 19802 10364 24686
rect 10428 22710 10456 24806
rect 10416 22704 10468 22710
rect 10416 22646 10468 22652
rect 10416 22432 10468 22438
rect 10416 22374 10468 22380
rect 10428 19854 10456 22374
rect 10520 22094 10548 25350
rect 10612 23662 10640 25434
rect 10600 23656 10652 23662
rect 10600 23598 10652 23604
rect 10704 22642 10732 25638
rect 10980 25498 11008 26930
rect 11072 26314 11100 27814
rect 11164 27062 11192 37062
rect 11256 36650 11284 38218
rect 11440 38010 11468 41550
rect 11796 41472 11848 41478
rect 11796 41414 11848 41420
rect 11808 40730 11836 41414
rect 11980 41132 12032 41138
rect 11980 41074 12032 41080
rect 11796 40724 11848 40730
rect 11796 40666 11848 40672
rect 11520 39840 11572 39846
rect 11520 39782 11572 39788
rect 11428 38004 11480 38010
rect 11428 37946 11480 37952
rect 11336 37868 11388 37874
rect 11336 37810 11388 37816
rect 11244 36644 11296 36650
rect 11244 36586 11296 36592
rect 11242 36408 11298 36417
rect 11242 36343 11244 36352
rect 11296 36343 11298 36352
rect 11244 36314 11296 36320
rect 11348 35290 11376 37810
rect 11440 37806 11468 37946
rect 11532 37942 11560 39782
rect 11888 39636 11940 39642
rect 11888 39578 11940 39584
rect 11704 38956 11756 38962
rect 11704 38898 11756 38904
rect 11716 38010 11744 38898
rect 11704 38004 11756 38010
rect 11704 37946 11756 37952
rect 11520 37936 11572 37942
rect 11520 37878 11572 37884
rect 11428 37800 11480 37806
rect 11428 37742 11480 37748
rect 11532 37738 11560 37878
rect 11520 37732 11572 37738
rect 11520 37674 11572 37680
rect 11704 37732 11756 37738
rect 11704 37674 11756 37680
rect 11716 37262 11744 37674
rect 11704 37256 11756 37262
rect 11704 37198 11756 37204
rect 11704 36100 11756 36106
rect 11704 36042 11756 36048
rect 11716 35698 11744 36042
rect 11704 35692 11756 35698
rect 11704 35634 11756 35640
rect 11336 35284 11388 35290
rect 11336 35226 11388 35232
rect 11716 35222 11744 35634
rect 11704 35216 11756 35222
rect 11704 35158 11756 35164
rect 11244 34944 11296 34950
rect 11244 34886 11296 34892
rect 11256 32570 11284 34886
rect 11716 34066 11744 35158
rect 11704 34060 11756 34066
rect 11704 34002 11756 34008
rect 11900 33114 11928 39578
rect 11992 39506 12020 41074
rect 12072 40384 12124 40390
rect 12072 40326 12124 40332
rect 12084 40186 12112 40326
rect 12072 40180 12124 40186
rect 12072 40122 12124 40128
rect 11980 39500 12032 39506
rect 11980 39442 12032 39448
rect 11992 38418 12020 39442
rect 12176 39098 12204 42230
rect 12268 41138 12296 42622
rect 12360 42158 12388 42706
rect 12348 42152 12400 42158
rect 12348 42094 12400 42100
rect 12256 41132 12308 41138
rect 12256 41074 12308 41080
rect 12348 40928 12400 40934
rect 12348 40870 12400 40876
rect 12360 39438 12388 40870
rect 12348 39432 12400 39438
rect 12348 39374 12400 39380
rect 12164 39092 12216 39098
rect 12164 39034 12216 39040
rect 12164 38752 12216 38758
rect 12164 38694 12216 38700
rect 11980 38412 12032 38418
rect 11980 38354 12032 38360
rect 11980 35080 12032 35086
rect 11980 35022 12032 35028
rect 11888 33108 11940 33114
rect 11888 33050 11940 33056
rect 11334 33008 11390 33017
rect 11334 32943 11336 32952
rect 11388 32943 11390 32952
rect 11336 32914 11388 32920
rect 11348 32774 11376 32914
rect 11992 32910 12020 35022
rect 12072 34944 12124 34950
rect 12072 34886 12124 34892
rect 12084 34474 12112 34886
rect 12072 34468 12124 34474
rect 12072 34410 12124 34416
rect 11980 32904 12032 32910
rect 11980 32846 12032 32852
rect 11336 32768 11388 32774
rect 11336 32710 11388 32716
rect 11244 32564 11296 32570
rect 11244 32506 11296 32512
rect 11992 32026 12020 32846
rect 11980 32020 12032 32026
rect 11980 31962 12032 31968
rect 11612 31680 11664 31686
rect 11612 31622 11664 31628
rect 11624 31414 11652 31622
rect 11612 31408 11664 31414
rect 11612 31350 11664 31356
rect 11624 31142 11652 31350
rect 11612 31136 11664 31142
rect 11612 31078 11664 31084
rect 11978 30832 12034 30841
rect 11978 30767 11980 30776
rect 12032 30767 12034 30776
rect 11980 30738 12032 30744
rect 11992 30598 12020 30738
rect 11980 30592 12032 30598
rect 11980 30534 12032 30540
rect 11428 29504 11480 29510
rect 11428 29446 11480 29452
rect 11336 29232 11388 29238
rect 11336 29174 11388 29180
rect 11152 27056 11204 27062
rect 11152 26998 11204 27004
rect 11244 26784 11296 26790
rect 11244 26726 11296 26732
rect 11060 26308 11112 26314
rect 11060 26250 11112 26256
rect 11152 26240 11204 26246
rect 11152 26182 11204 26188
rect 11164 26042 11192 26182
rect 11152 26036 11204 26042
rect 11152 25978 11204 25984
rect 11152 25900 11204 25906
rect 11152 25842 11204 25848
rect 11164 25702 11192 25842
rect 11152 25696 11204 25702
rect 11152 25638 11204 25644
rect 10968 25492 11020 25498
rect 10968 25434 11020 25440
rect 11164 25430 11192 25638
rect 11152 25424 11204 25430
rect 11152 25366 11204 25372
rect 10784 24608 10836 24614
rect 10784 24550 10836 24556
rect 10692 22636 10744 22642
rect 10692 22578 10744 22584
rect 10692 22094 10744 22098
rect 10520 22092 10744 22094
rect 10520 22066 10692 22092
rect 10692 22034 10744 22040
rect 10704 21690 10732 22034
rect 10796 21690 10824 24550
rect 11256 24274 11284 26726
rect 11348 24410 11376 29174
rect 11440 28150 11468 29446
rect 11612 28960 11664 28966
rect 11612 28902 11664 28908
rect 11428 28144 11480 28150
rect 11428 28086 11480 28092
rect 11440 26450 11468 28086
rect 11624 27946 11652 28902
rect 11704 28076 11756 28082
rect 11704 28018 11756 28024
rect 11612 27940 11664 27946
rect 11612 27882 11664 27888
rect 11428 26444 11480 26450
rect 11428 26386 11480 26392
rect 11716 25906 11744 28018
rect 12072 27532 12124 27538
rect 12072 27474 12124 27480
rect 12084 26994 12112 27474
rect 12072 26988 12124 26994
rect 12072 26930 12124 26936
rect 11796 26512 11848 26518
rect 11796 26454 11848 26460
rect 11808 26042 11836 26454
rect 12072 26308 12124 26314
rect 12072 26250 12124 26256
rect 11796 26036 11848 26042
rect 11796 25978 11848 25984
rect 12084 25974 12112 26250
rect 12072 25968 12124 25974
rect 12072 25910 12124 25916
rect 11704 25900 11756 25906
rect 11704 25842 11756 25848
rect 12084 25158 12112 25910
rect 12072 25152 12124 25158
rect 12072 25094 12124 25100
rect 11428 24948 11480 24954
rect 11428 24890 11480 24896
rect 12072 24948 12124 24954
rect 12176 24936 12204 38694
rect 12256 37664 12308 37670
rect 12256 37606 12308 37612
rect 12268 37466 12296 37606
rect 12256 37460 12308 37466
rect 12256 37402 12308 37408
rect 12268 32842 12296 37402
rect 12452 36786 12480 44474
rect 12532 41608 12584 41614
rect 12532 41550 12584 41556
rect 12544 39642 12572 41550
rect 12624 40656 12676 40662
rect 12624 40598 12676 40604
rect 12532 39636 12584 39642
rect 12532 39578 12584 39584
rect 12544 38894 12572 39578
rect 12636 39098 12664 40598
rect 12728 40526 12756 48214
rect 12950 47356 13258 47365
rect 12950 47354 12956 47356
rect 13012 47354 13036 47356
rect 13092 47354 13116 47356
rect 13172 47354 13196 47356
rect 13252 47354 13258 47356
rect 13012 47302 13014 47354
rect 13194 47302 13196 47354
rect 12950 47300 12956 47302
rect 13012 47300 13036 47302
rect 13092 47300 13116 47302
rect 13172 47300 13196 47302
rect 13252 47300 13258 47302
rect 12950 47291 13258 47300
rect 12950 46268 13258 46277
rect 12950 46266 12956 46268
rect 13012 46266 13036 46268
rect 13092 46266 13116 46268
rect 13172 46266 13196 46268
rect 13252 46266 13258 46268
rect 13012 46214 13014 46266
rect 13194 46214 13196 46266
rect 12950 46212 12956 46214
rect 13012 46212 13036 46214
rect 13092 46212 13116 46214
rect 13172 46212 13196 46214
rect 13252 46212 13258 46214
rect 12950 46203 13258 46212
rect 13176 45824 13228 45830
rect 13176 45766 13228 45772
rect 13188 45558 13216 45766
rect 13176 45552 13228 45558
rect 13176 45494 13228 45500
rect 13464 45354 13492 49166
rect 14188 46912 14240 46918
rect 14188 46854 14240 46860
rect 14200 46646 14228 46854
rect 14188 46640 14240 46646
rect 14188 46582 14240 46588
rect 14096 46368 14148 46374
rect 14096 46310 14148 46316
rect 13728 45824 13780 45830
rect 13728 45766 13780 45772
rect 13636 45552 13688 45558
rect 13636 45494 13688 45500
rect 13544 45484 13596 45490
rect 13544 45426 13596 45432
rect 13452 45348 13504 45354
rect 13452 45290 13504 45296
rect 12950 45180 13258 45189
rect 12950 45178 12956 45180
rect 13012 45178 13036 45180
rect 13092 45178 13116 45180
rect 13172 45178 13196 45180
rect 13252 45178 13258 45180
rect 13012 45126 13014 45178
rect 13194 45126 13196 45178
rect 12950 45124 12956 45126
rect 13012 45124 13036 45126
rect 13092 45124 13116 45126
rect 13172 45124 13196 45126
rect 13252 45124 13258 45126
rect 12950 45115 13258 45124
rect 12808 44736 12860 44742
rect 12808 44678 12860 44684
rect 12820 43382 12848 44678
rect 12950 44092 13258 44101
rect 12950 44090 12956 44092
rect 13012 44090 13036 44092
rect 13092 44090 13116 44092
rect 13172 44090 13196 44092
rect 13252 44090 13258 44092
rect 13012 44038 13014 44090
rect 13194 44038 13196 44090
rect 12950 44036 12956 44038
rect 13012 44036 13036 44038
rect 13092 44036 13116 44038
rect 13172 44036 13196 44038
rect 13252 44036 13258 44038
rect 12950 44027 13258 44036
rect 12808 43376 12860 43382
rect 12808 43318 12860 43324
rect 12950 43004 13258 43013
rect 12950 43002 12956 43004
rect 13012 43002 13036 43004
rect 13092 43002 13116 43004
rect 13172 43002 13196 43004
rect 13252 43002 13258 43004
rect 13012 42950 13014 43002
rect 13194 42950 13196 43002
rect 12950 42948 12956 42950
rect 13012 42948 13036 42950
rect 13092 42948 13116 42950
rect 13172 42948 13196 42950
rect 13252 42948 13258 42950
rect 12950 42939 13258 42948
rect 13556 42362 13584 45426
rect 13544 42356 13596 42362
rect 13544 42298 13596 42304
rect 13452 42288 13504 42294
rect 13452 42230 13504 42236
rect 12950 41916 13258 41925
rect 12950 41914 12956 41916
rect 13012 41914 13036 41916
rect 13092 41914 13116 41916
rect 13172 41914 13196 41916
rect 13252 41914 13258 41916
rect 13012 41862 13014 41914
rect 13194 41862 13196 41914
rect 12950 41860 12956 41862
rect 13012 41860 13036 41862
rect 13092 41860 13116 41862
rect 13172 41860 13196 41862
rect 13252 41860 13258 41862
rect 12950 41851 13258 41860
rect 12808 41744 12860 41750
rect 12808 41686 12860 41692
rect 12716 40520 12768 40526
rect 12716 40462 12768 40468
rect 12716 40044 12768 40050
rect 12716 39986 12768 39992
rect 12728 39506 12756 39986
rect 12716 39500 12768 39506
rect 12716 39442 12768 39448
rect 12624 39092 12676 39098
rect 12624 39034 12676 39040
rect 12716 38956 12768 38962
rect 12716 38898 12768 38904
rect 12532 38888 12584 38894
rect 12532 38830 12584 38836
rect 12624 38412 12676 38418
rect 12624 38354 12676 38360
rect 12636 38321 12664 38354
rect 12622 38312 12678 38321
rect 12622 38247 12678 38256
rect 12728 37754 12756 38898
rect 12636 37726 12756 37754
rect 12532 37664 12584 37670
rect 12532 37606 12584 37612
rect 12440 36780 12492 36786
rect 12440 36722 12492 36728
rect 12440 36576 12492 36582
rect 12440 36518 12492 36524
rect 12348 35488 12400 35494
rect 12348 35430 12400 35436
rect 12360 35018 12388 35430
rect 12348 35012 12400 35018
rect 12348 34954 12400 34960
rect 12452 33862 12480 36518
rect 12544 36242 12572 37606
rect 12532 36236 12584 36242
rect 12532 36178 12584 36184
rect 12636 36122 12664 37726
rect 12716 37664 12768 37670
rect 12716 37606 12768 37612
rect 12728 37126 12756 37606
rect 12820 37194 12848 41686
rect 13360 41472 13412 41478
rect 13360 41414 13412 41420
rect 13372 41070 13400 41414
rect 13360 41064 13412 41070
rect 13360 41006 13412 41012
rect 12950 40828 13258 40837
rect 12950 40826 12956 40828
rect 13012 40826 13036 40828
rect 13092 40826 13116 40828
rect 13172 40826 13196 40828
rect 13252 40826 13258 40828
rect 13012 40774 13014 40826
rect 13194 40774 13196 40826
rect 12950 40772 12956 40774
rect 13012 40772 13036 40774
rect 13092 40772 13116 40774
rect 13172 40772 13196 40774
rect 13252 40772 13258 40774
rect 12950 40763 13258 40772
rect 12900 40588 12952 40594
rect 12900 40530 12952 40536
rect 13360 40588 13412 40594
rect 13360 40530 13412 40536
rect 12912 40390 12940 40530
rect 12900 40384 12952 40390
rect 12900 40326 12952 40332
rect 12950 39740 13258 39749
rect 12950 39738 12956 39740
rect 13012 39738 13036 39740
rect 13092 39738 13116 39740
rect 13172 39738 13196 39740
rect 13252 39738 13258 39740
rect 13012 39686 13014 39738
rect 13194 39686 13196 39738
rect 12950 39684 12956 39686
rect 13012 39684 13036 39686
rect 13092 39684 13116 39686
rect 13172 39684 13196 39686
rect 13252 39684 13258 39686
rect 12950 39675 13258 39684
rect 13372 39642 13400 40530
rect 13360 39636 13412 39642
rect 13360 39578 13412 39584
rect 12992 39296 13044 39302
rect 12992 39238 13044 39244
rect 13084 39296 13136 39302
rect 13084 39238 13136 39244
rect 13004 38894 13032 39238
rect 13096 38962 13124 39238
rect 13084 38956 13136 38962
rect 13084 38898 13136 38904
rect 12992 38888 13044 38894
rect 12992 38830 13044 38836
rect 12950 38652 13258 38661
rect 12950 38650 12956 38652
rect 13012 38650 13036 38652
rect 13092 38650 13116 38652
rect 13172 38650 13196 38652
rect 13252 38650 13258 38652
rect 13012 38598 13014 38650
rect 13194 38598 13196 38650
rect 12950 38596 12956 38598
rect 13012 38596 13036 38598
rect 13092 38596 13116 38598
rect 13172 38596 13196 38598
rect 13252 38596 13258 38598
rect 12950 38587 13258 38596
rect 13360 38480 13412 38486
rect 13360 38422 13412 38428
rect 12950 37564 13258 37573
rect 12950 37562 12956 37564
rect 13012 37562 13036 37564
rect 13092 37562 13116 37564
rect 13172 37562 13196 37564
rect 13252 37562 13258 37564
rect 13012 37510 13014 37562
rect 13194 37510 13196 37562
rect 12950 37508 12956 37510
rect 13012 37508 13036 37510
rect 13092 37508 13116 37510
rect 13172 37508 13196 37510
rect 13252 37508 13258 37510
rect 12950 37499 13258 37508
rect 13084 37460 13136 37466
rect 13372 37448 13400 38422
rect 13084 37402 13136 37408
rect 13280 37420 13400 37448
rect 13096 37330 13124 37402
rect 13084 37324 13136 37330
rect 13084 37266 13136 37272
rect 12808 37188 12860 37194
rect 12808 37130 12860 37136
rect 13084 37188 13136 37194
rect 13084 37130 13136 37136
rect 12716 37120 12768 37126
rect 12716 37062 12768 37068
rect 12544 36094 12664 36122
rect 12544 35601 12572 36094
rect 12624 36032 12676 36038
rect 12624 35974 12676 35980
rect 12530 35592 12586 35601
rect 12530 35527 12586 35536
rect 12532 35488 12584 35494
rect 12532 35430 12584 35436
rect 12544 34610 12572 35430
rect 12532 34604 12584 34610
rect 12532 34546 12584 34552
rect 12440 33856 12492 33862
rect 12440 33798 12492 33804
rect 12636 33658 12664 35974
rect 12728 35222 12756 37062
rect 13096 36922 13124 37130
rect 13084 36916 13136 36922
rect 13084 36858 13136 36864
rect 13280 36718 13308 37420
rect 13358 37360 13414 37369
rect 13358 37295 13360 37304
rect 13412 37295 13414 37304
rect 13360 37266 13412 37272
rect 13360 36780 13412 36786
rect 13360 36722 13412 36728
rect 12808 36712 12860 36718
rect 12808 36654 12860 36660
rect 13268 36712 13320 36718
rect 13268 36654 13320 36660
rect 12716 35216 12768 35222
rect 12716 35158 12768 35164
rect 12716 34740 12768 34746
rect 12716 34682 12768 34688
rect 12624 33652 12676 33658
rect 12624 33594 12676 33600
rect 12532 33516 12584 33522
rect 12532 33458 12584 33464
rect 12544 33318 12572 33458
rect 12532 33312 12584 33318
rect 12530 33280 12532 33289
rect 12584 33280 12586 33289
rect 12530 33215 12586 33224
rect 12256 32836 12308 32842
rect 12256 32778 12308 32784
rect 12440 32360 12492 32366
rect 12440 32302 12492 32308
rect 12452 31822 12480 32302
rect 12440 31816 12492 31822
rect 12440 31758 12492 31764
rect 12624 31272 12676 31278
rect 12624 31214 12676 31220
rect 12440 31204 12492 31210
rect 12440 31146 12492 31152
rect 12452 30734 12480 31146
rect 12440 30728 12492 30734
rect 12440 30670 12492 30676
rect 12636 30326 12664 31214
rect 12624 30320 12676 30326
rect 12624 30262 12676 30268
rect 12728 30190 12756 34682
rect 12820 31890 12848 36654
rect 12950 36476 13258 36485
rect 12950 36474 12956 36476
rect 13012 36474 13036 36476
rect 13092 36474 13116 36476
rect 13172 36474 13196 36476
rect 13252 36474 13258 36476
rect 13012 36422 13014 36474
rect 13194 36422 13196 36474
rect 12950 36420 12956 36422
rect 13012 36420 13036 36422
rect 13092 36420 13116 36422
rect 13172 36420 13196 36422
rect 13252 36420 13258 36422
rect 12950 36411 13258 36420
rect 13372 36242 13400 36722
rect 13464 36378 13492 42230
rect 13544 40452 13596 40458
rect 13544 40394 13596 40400
rect 13452 36372 13504 36378
rect 13452 36314 13504 36320
rect 13360 36236 13412 36242
rect 13360 36178 13412 36184
rect 13360 35828 13412 35834
rect 13360 35770 13412 35776
rect 12950 35388 13258 35397
rect 12950 35386 12956 35388
rect 13012 35386 13036 35388
rect 13092 35386 13116 35388
rect 13172 35386 13196 35388
rect 13252 35386 13258 35388
rect 13012 35334 13014 35386
rect 13194 35334 13196 35386
rect 12950 35332 12956 35334
rect 13012 35332 13036 35334
rect 13092 35332 13116 35334
rect 13172 35332 13196 35334
rect 13252 35332 13258 35334
rect 12950 35323 13258 35332
rect 12950 34300 13258 34309
rect 12950 34298 12956 34300
rect 13012 34298 13036 34300
rect 13092 34298 13116 34300
rect 13172 34298 13196 34300
rect 13252 34298 13258 34300
rect 13012 34246 13014 34298
rect 13194 34246 13196 34298
rect 12950 34244 12956 34246
rect 13012 34244 13036 34246
rect 13092 34244 13116 34246
rect 13172 34244 13196 34246
rect 13252 34244 13258 34246
rect 12950 34235 13258 34244
rect 13372 33454 13400 35770
rect 13452 35760 13504 35766
rect 13452 35702 13504 35708
rect 13464 35018 13492 35702
rect 13452 35012 13504 35018
rect 13452 34954 13504 34960
rect 13464 33998 13492 34954
rect 13556 34746 13584 40394
rect 13648 39574 13676 45494
rect 13740 44538 13768 45766
rect 14108 45422 14136 46310
rect 14200 46170 14228 46582
rect 14280 46504 14332 46510
rect 14280 46446 14332 46452
rect 14188 46164 14240 46170
rect 14188 46106 14240 46112
rect 14200 45898 14228 46106
rect 14188 45892 14240 45898
rect 14188 45834 14240 45840
rect 13820 45416 13872 45422
rect 13820 45358 13872 45364
rect 14096 45416 14148 45422
rect 14096 45358 14148 45364
rect 13832 44878 13860 45358
rect 14096 44940 14148 44946
rect 14096 44882 14148 44888
rect 13820 44872 13872 44878
rect 13820 44814 13872 44820
rect 13728 44532 13780 44538
rect 13728 44474 13780 44480
rect 13740 43450 13768 44474
rect 14108 44334 14136 44882
rect 14188 44804 14240 44810
rect 14188 44746 14240 44752
rect 14096 44328 14148 44334
rect 14096 44270 14148 44276
rect 13820 43784 13872 43790
rect 13820 43726 13872 43732
rect 13728 43444 13780 43450
rect 13728 43386 13780 43392
rect 13832 42770 13860 43726
rect 14108 43382 14136 44270
rect 14096 43376 14148 43382
rect 14016 43336 14096 43364
rect 14016 42838 14044 43336
rect 14096 43318 14148 43324
rect 14200 43194 14228 44746
rect 14292 44282 14320 46446
rect 14372 45416 14424 45422
rect 14372 45358 14424 45364
rect 14384 44946 14412 45358
rect 14372 44940 14424 44946
rect 14372 44882 14424 44888
rect 14476 44520 14504 53382
rect 14648 52896 14700 52902
rect 14648 52838 14700 52844
rect 14556 46504 14608 46510
rect 14556 46446 14608 46452
rect 14568 45558 14596 46446
rect 14556 45552 14608 45558
rect 14556 45494 14608 45500
rect 14476 44492 14596 44520
rect 14292 44254 14504 44282
rect 14476 44198 14504 44254
rect 14372 44192 14424 44198
rect 14372 44134 14424 44140
rect 14464 44192 14516 44198
rect 14464 44134 14516 44140
rect 14096 43172 14148 43178
rect 14200 43166 14320 43194
rect 14096 43114 14148 43120
rect 14004 42832 14056 42838
rect 14004 42774 14056 42780
rect 13820 42764 13872 42770
rect 13820 42706 13872 42712
rect 14108 42650 14136 43114
rect 14108 42622 14228 42650
rect 14200 41478 14228 42622
rect 14188 41472 14240 41478
rect 14188 41414 14240 41420
rect 13820 40928 13872 40934
rect 13820 40870 13872 40876
rect 13728 40520 13780 40526
rect 13728 40462 13780 40468
rect 13636 39568 13688 39574
rect 13636 39510 13688 39516
rect 13636 39432 13688 39438
rect 13636 39374 13688 39380
rect 13648 38282 13676 39374
rect 13636 38276 13688 38282
rect 13636 38218 13688 38224
rect 13648 38010 13676 38218
rect 13636 38004 13688 38010
rect 13636 37946 13688 37952
rect 13636 37800 13688 37806
rect 13636 37742 13688 37748
rect 13648 35834 13676 37742
rect 13636 35828 13688 35834
rect 13636 35770 13688 35776
rect 13740 35578 13768 40462
rect 13832 40458 13860 40870
rect 13820 40452 13872 40458
rect 13820 40394 13872 40400
rect 14200 39642 14228 41414
rect 13820 39636 13872 39642
rect 13820 39578 13872 39584
rect 14188 39636 14240 39642
rect 14188 39578 14240 39584
rect 13832 39302 13860 39578
rect 13912 39500 13964 39506
rect 13912 39442 13964 39448
rect 13820 39296 13872 39302
rect 13820 39238 13872 39244
rect 13832 38826 13860 39238
rect 13820 38820 13872 38826
rect 13820 38762 13872 38768
rect 13820 37460 13872 37466
rect 13820 37402 13872 37408
rect 13832 36718 13860 37402
rect 13820 36712 13872 36718
rect 13820 36654 13872 36660
rect 13820 36032 13872 36038
rect 13818 36000 13820 36009
rect 13872 36000 13874 36009
rect 13818 35935 13874 35944
rect 13924 35834 13952 39442
rect 14004 39296 14056 39302
rect 14004 39238 14056 39244
rect 14016 38758 14044 39238
rect 14004 38752 14056 38758
rect 14004 38694 14056 38700
rect 14096 38752 14148 38758
rect 14096 38694 14148 38700
rect 14188 38752 14240 38758
rect 14188 38694 14240 38700
rect 14108 38554 14136 38694
rect 14096 38548 14148 38554
rect 14096 38490 14148 38496
rect 14004 38004 14056 38010
rect 14004 37946 14056 37952
rect 13912 35828 13964 35834
rect 13912 35770 13964 35776
rect 14016 35766 14044 37946
rect 14200 37262 14228 38694
rect 14292 37670 14320 43166
rect 14384 42294 14412 44134
rect 14372 42288 14424 42294
rect 14372 42230 14424 42236
rect 14464 41540 14516 41546
rect 14464 41482 14516 41488
rect 14372 40044 14424 40050
rect 14372 39986 14424 39992
rect 14384 39438 14412 39986
rect 14372 39432 14424 39438
rect 14372 39374 14424 39380
rect 14280 37664 14332 37670
rect 14280 37606 14332 37612
rect 14188 37256 14240 37262
rect 14188 37198 14240 37204
rect 14476 37126 14504 41482
rect 14280 37120 14332 37126
rect 14280 37062 14332 37068
rect 14464 37120 14516 37126
rect 14464 37062 14516 37068
rect 14292 36922 14320 37062
rect 14280 36916 14332 36922
rect 14280 36858 14332 36864
rect 14096 36780 14148 36786
rect 14096 36722 14148 36728
rect 14004 35760 14056 35766
rect 14004 35702 14056 35708
rect 14108 35612 14136 36722
rect 14372 36576 14424 36582
rect 14372 36518 14424 36524
rect 14464 36576 14516 36582
rect 14464 36518 14516 36524
rect 14384 36038 14412 36518
rect 14372 36032 14424 36038
rect 14372 35974 14424 35980
rect 13648 35562 13768 35578
rect 13636 35556 13768 35562
rect 13688 35550 13768 35556
rect 13924 35584 14136 35612
rect 13636 35498 13688 35504
rect 13634 35456 13690 35465
rect 13634 35391 13690 35400
rect 13544 34740 13596 34746
rect 13544 34682 13596 34688
rect 13544 34604 13596 34610
rect 13544 34546 13596 34552
rect 13452 33992 13504 33998
rect 13452 33934 13504 33940
rect 13464 33590 13492 33934
rect 13452 33584 13504 33590
rect 13452 33526 13504 33532
rect 13360 33448 13412 33454
rect 13360 33390 13412 33396
rect 13452 33448 13504 33454
rect 13452 33390 13504 33396
rect 12950 33212 13258 33221
rect 12950 33210 12956 33212
rect 13012 33210 13036 33212
rect 13092 33210 13116 33212
rect 13172 33210 13196 33212
rect 13252 33210 13258 33212
rect 13012 33158 13014 33210
rect 13194 33158 13196 33210
rect 12950 33156 12956 33158
rect 13012 33156 13036 33158
rect 13092 33156 13116 33158
rect 13172 33156 13196 33158
rect 13252 33156 13258 33158
rect 12950 33147 13258 33156
rect 13266 32600 13322 32609
rect 13266 32535 13322 32544
rect 13280 32230 13308 32535
rect 13268 32224 13320 32230
rect 13268 32166 13320 32172
rect 12950 32124 13258 32133
rect 12950 32122 12956 32124
rect 13012 32122 13036 32124
rect 13092 32122 13116 32124
rect 13172 32122 13196 32124
rect 13252 32122 13258 32124
rect 13012 32070 13014 32122
rect 13194 32070 13196 32122
rect 12950 32068 12956 32070
rect 13012 32068 13036 32070
rect 13092 32068 13116 32070
rect 13172 32068 13196 32070
rect 13252 32068 13258 32070
rect 12950 32059 13258 32068
rect 13464 31890 13492 33390
rect 12808 31884 12860 31890
rect 12808 31826 12860 31832
rect 13452 31884 13504 31890
rect 13452 31826 13504 31832
rect 12808 31408 12860 31414
rect 12808 31350 12860 31356
rect 12716 30184 12768 30190
rect 12716 30126 12768 30132
rect 12716 30048 12768 30054
rect 12716 29990 12768 29996
rect 12256 29504 12308 29510
rect 12256 29446 12308 29452
rect 12268 29238 12296 29446
rect 12256 29232 12308 29238
rect 12256 29174 12308 29180
rect 12624 29028 12676 29034
rect 12624 28970 12676 28976
rect 12348 28484 12400 28490
rect 12348 28426 12400 28432
rect 12256 27328 12308 27334
rect 12256 27270 12308 27276
rect 12124 24908 12204 24936
rect 12072 24890 12124 24896
rect 11440 24857 11468 24890
rect 11426 24848 11482 24857
rect 11426 24783 11482 24792
rect 11336 24404 11388 24410
rect 11336 24346 11388 24352
rect 11244 24268 11296 24274
rect 11244 24210 11296 24216
rect 11704 23724 11756 23730
rect 11704 23666 11756 23672
rect 11060 23656 11112 23662
rect 11060 23598 11112 23604
rect 11072 23066 11100 23598
rect 11520 23316 11572 23322
rect 11520 23258 11572 23264
rect 10888 23038 11100 23066
rect 10692 21684 10744 21690
rect 10692 21626 10744 21632
rect 10784 21684 10836 21690
rect 10784 21626 10836 21632
rect 10888 21570 10916 23038
rect 11532 22982 11560 23258
rect 11520 22976 11572 22982
rect 11520 22918 11572 22924
rect 10968 22568 11020 22574
rect 10968 22510 11020 22516
rect 10980 21622 11008 22510
rect 11152 21888 11204 21894
rect 11152 21830 11204 21836
rect 10796 21542 10916 21570
rect 10968 21616 11020 21622
rect 10968 21558 11020 21564
rect 10244 19774 10364 19802
rect 10416 19848 10468 19854
rect 10416 19790 10468 19796
rect 10140 19712 10192 19718
rect 10140 19654 10192 19660
rect 10152 19378 10180 19654
rect 10140 19372 10192 19378
rect 10140 19314 10192 19320
rect 10152 18630 10180 19314
rect 10244 19242 10272 19774
rect 10324 19712 10376 19718
rect 10324 19654 10376 19660
rect 10232 19236 10284 19242
rect 10232 19178 10284 19184
rect 10140 18624 10192 18630
rect 10140 18566 10192 18572
rect 10048 18420 10100 18426
rect 10048 18362 10100 18368
rect 9864 18216 9916 18222
rect 9864 18158 9916 18164
rect 9864 17604 9916 17610
rect 9864 17546 9916 17552
rect 9876 16726 9904 17546
rect 9864 16720 9916 16726
rect 9864 16662 9916 16668
rect 9956 16652 10008 16658
rect 9956 16594 10008 16600
rect 9968 14414 9996 16594
rect 9956 14408 10008 14414
rect 9956 14350 10008 14356
rect 9968 14074 9996 14350
rect 9956 14068 10008 14074
rect 9956 14010 10008 14016
rect 9864 12164 9916 12170
rect 9864 12106 9916 12112
rect 9876 11898 9904 12106
rect 9864 11892 9916 11898
rect 9864 11834 9916 11840
rect 10060 10742 10088 18362
rect 10244 18358 10272 19178
rect 10336 18426 10364 19654
rect 10508 19508 10560 19514
rect 10508 19450 10560 19456
rect 10520 19394 10548 19450
rect 10428 19366 10548 19394
rect 10796 19394 10824 21542
rect 10876 20052 10928 20058
rect 10876 19994 10928 20000
rect 10888 19514 10916 19994
rect 11060 19916 11112 19922
rect 11060 19858 11112 19864
rect 10876 19508 10928 19514
rect 10876 19450 10928 19456
rect 10796 19378 10916 19394
rect 10796 19372 10928 19378
rect 10796 19366 10876 19372
rect 10324 18420 10376 18426
rect 10324 18362 10376 18368
rect 10232 18352 10284 18358
rect 10232 18294 10284 18300
rect 10140 17332 10192 17338
rect 10140 17274 10192 17280
rect 10152 15706 10180 17274
rect 10244 17218 10272 18294
rect 10244 17190 10364 17218
rect 10336 17134 10364 17190
rect 10324 17128 10376 17134
rect 10324 17070 10376 17076
rect 10324 16448 10376 16454
rect 10324 16390 10376 16396
rect 10336 16182 10364 16390
rect 10324 16176 10376 16182
rect 10324 16118 10376 16124
rect 10140 15700 10192 15706
rect 10140 15642 10192 15648
rect 10152 15434 10180 15642
rect 10140 15428 10192 15434
rect 10140 15370 10192 15376
rect 10324 12776 10376 12782
rect 10324 12718 10376 12724
rect 10336 12170 10364 12718
rect 10324 12164 10376 12170
rect 10324 12106 10376 12112
rect 10336 11694 10364 12106
rect 10428 11830 10456 19366
rect 10876 19314 10928 19320
rect 10692 18896 10744 18902
rect 10692 18838 10744 18844
rect 10508 17536 10560 17542
rect 10508 17478 10560 17484
rect 10520 17338 10548 17478
rect 10508 17332 10560 17338
rect 10508 17274 10560 17280
rect 10508 17060 10560 17066
rect 10508 17002 10560 17008
rect 10520 13394 10548 17002
rect 10704 16590 10732 18838
rect 10888 18766 10916 19314
rect 11072 18970 11100 19858
rect 11060 18964 11112 18970
rect 11060 18906 11112 18912
rect 10968 18828 11020 18834
rect 10968 18770 11020 18776
rect 10876 18760 10928 18766
rect 10876 18702 10928 18708
rect 10980 17898 11008 18770
rect 10980 17870 11100 17898
rect 11072 17746 11100 17870
rect 11060 17740 11112 17746
rect 11060 17682 11112 17688
rect 11072 17270 11100 17682
rect 11060 17264 11112 17270
rect 11060 17206 11112 17212
rect 10784 17128 10836 17134
rect 10784 17070 10836 17076
rect 10692 16584 10744 16590
rect 10692 16526 10744 16532
rect 10796 15434 10824 17070
rect 11060 16448 11112 16454
rect 11060 16390 11112 16396
rect 10876 16040 10928 16046
rect 10876 15982 10928 15988
rect 10888 15570 10916 15982
rect 10876 15564 10928 15570
rect 10876 15506 10928 15512
rect 10784 15428 10836 15434
rect 10784 15370 10836 15376
rect 10796 15094 10824 15370
rect 10784 15088 10836 15094
rect 10784 15030 10836 15036
rect 10888 14482 10916 15506
rect 11072 14618 11100 16390
rect 11164 16250 11192 21830
rect 11244 20936 11296 20942
rect 11244 20878 11296 20884
rect 11256 20058 11284 20878
rect 11244 20052 11296 20058
rect 11244 19994 11296 20000
rect 11244 18624 11296 18630
rect 11244 18566 11296 18572
rect 11256 16454 11284 18566
rect 11532 17882 11560 22918
rect 11716 22710 11744 23666
rect 12164 23656 12216 23662
rect 12084 23604 12164 23610
rect 12084 23598 12216 23604
rect 11980 23588 12032 23594
rect 11980 23530 12032 23536
rect 12084 23582 12204 23598
rect 11796 23248 11848 23254
rect 11794 23216 11796 23225
rect 11848 23216 11850 23225
rect 11794 23151 11850 23160
rect 11808 22778 11836 23151
rect 11992 22982 12020 23530
rect 11980 22976 12032 22982
rect 11980 22918 12032 22924
rect 11796 22772 11848 22778
rect 12084 22760 12112 23582
rect 12164 23520 12216 23526
rect 12164 23462 12216 23468
rect 11796 22714 11848 22720
rect 11992 22732 12112 22760
rect 11704 22704 11756 22710
rect 11704 22646 11756 22652
rect 11992 22506 12020 22732
rect 12072 22636 12124 22642
rect 12072 22578 12124 22584
rect 11980 22500 12032 22506
rect 11980 22442 12032 22448
rect 11704 22092 11756 22098
rect 11704 22034 11756 22040
rect 11612 21888 11664 21894
rect 11612 21830 11664 21836
rect 11624 21486 11652 21830
rect 11716 21690 11744 22034
rect 11704 21684 11756 21690
rect 11704 21626 11756 21632
rect 11612 21480 11664 21486
rect 11612 21422 11664 21428
rect 11796 21004 11848 21010
rect 11796 20946 11848 20952
rect 11808 19922 11836 20946
rect 12084 20262 12112 22578
rect 12176 20942 12204 23462
rect 12268 22710 12296 27270
rect 12360 26450 12388 28426
rect 12440 27328 12492 27334
rect 12440 27270 12492 27276
rect 12348 26444 12400 26450
rect 12348 26386 12400 26392
rect 12348 25696 12400 25702
rect 12348 25638 12400 25644
rect 12360 24206 12388 25638
rect 12452 25430 12480 27270
rect 12440 25424 12492 25430
rect 12440 25366 12492 25372
rect 12532 25356 12584 25362
rect 12532 25298 12584 25304
rect 12440 25152 12492 25158
rect 12544 25140 12572 25298
rect 12492 25112 12572 25140
rect 12440 25094 12492 25100
rect 12440 24880 12492 24886
rect 12440 24822 12492 24828
rect 12452 24410 12480 24822
rect 12440 24404 12492 24410
rect 12440 24346 12492 24352
rect 12440 24268 12492 24274
rect 12440 24210 12492 24216
rect 12348 24200 12400 24206
rect 12348 24142 12400 24148
rect 12452 23746 12480 24210
rect 12360 23718 12480 23746
rect 12360 23050 12388 23718
rect 12348 23044 12400 23050
rect 12348 22986 12400 22992
rect 12544 22778 12572 25112
rect 12532 22772 12584 22778
rect 12532 22714 12584 22720
rect 12256 22704 12308 22710
rect 12256 22646 12308 22652
rect 12636 22642 12664 28970
rect 12728 24954 12756 29990
rect 12820 28558 12848 31350
rect 12950 31036 13258 31045
rect 12950 31034 12956 31036
rect 13012 31034 13036 31036
rect 13092 31034 13116 31036
rect 13172 31034 13196 31036
rect 13252 31034 13258 31036
rect 13012 30982 13014 31034
rect 13194 30982 13196 31034
rect 12950 30980 12956 30982
rect 13012 30980 13036 30982
rect 13092 30980 13116 30982
rect 13172 30980 13196 30982
rect 13252 30980 13258 30982
rect 12950 30971 13258 30980
rect 12992 30728 13044 30734
rect 13044 30676 13124 30682
rect 12992 30670 13124 30676
rect 13004 30654 13124 30670
rect 13096 30190 13124 30654
rect 13084 30184 13136 30190
rect 13084 30126 13136 30132
rect 12950 29948 13258 29957
rect 12950 29946 12956 29948
rect 13012 29946 13036 29948
rect 13092 29946 13116 29948
rect 13172 29946 13196 29948
rect 13252 29946 13258 29948
rect 13012 29894 13014 29946
rect 13194 29894 13196 29946
rect 12950 29892 12956 29894
rect 13012 29892 13036 29894
rect 13092 29892 13116 29894
rect 13172 29892 13196 29894
rect 13252 29892 13258 29894
rect 12950 29883 13258 29892
rect 13360 29164 13412 29170
rect 13360 29106 13412 29112
rect 12950 28860 13258 28869
rect 12950 28858 12956 28860
rect 13012 28858 13036 28860
rect 13092 28858 13116 28860
rect 13172 28858 13196 28860
rect 13252 28858 13258 28860
rect 13012 28806 13014 28858
rect 13194 28806 13196 28858
rect 12950 28804 12956 28806
rect 13012 28804 13036 28806
rect 13092 28804 13116 28806
rect 13172 28804 13196 28806
rect 13252 28804 13258 28806
rect 12950 28795 13258 28804
rect 13372 28762 13400 29106
rect 13360 28756 13412 28762
rect 13360 28698 13412 28704
rect 13452 28688 13504 28694
rect 13452 28630 13504 28636
rect 12808 28552 12860 28558
rect 12808 28494 12860 28500
rect 12808 28008 12860 28014
rect 12808 27950 12860 27956
rect 13360 28008 13412 28014
rect 13360 27950 13412 27956
rect 12820 26994 12848 27950
rect 12950 27772 13258 27781
rect 12950 27770 12956 27772
rect 13012 27770 13036 27772
rect 13092 27770 13116 27772
rect 13172 27770 13196 27772
rect 13252 27770 13258 27772
rect 13012 27718 13014 27770
rect 13194 27718 13196 27770
rect 12950 27716 12956 27718
rect 13012 27716 13036 27718
rect 13092 27716 13116 27718
rect 13172 27716 13196 27718
rect 13252 27716 13258 27718
rect 12950 27707 13258 27716
rect 13268 27328 13320 27334
rect 13268 27270 13320 27276
rect 12808 26988 12860 26994
rect 12808 26930 12860 26936
rect 12716 24948 12768 24954
rect 12716 24890 12768 24896
rect 12820 23186 12848 26930
rect 13280 26790 13308 27270
rect 13268 26784 13320 26790
rect 13268 26726 13320 26732
rect 12950 26684 13258 26693
rect 12950 26682 12956 26684
rect 13012 26682 13036 26684
rect 13092 26682 13116 26684
rect 13172 26682 13196 26684
rect 13252 26682 13258 26684
rect 13012 26630 13014 26682
rect 13194 26630 13196 26682
rect 12950 26628 12956 26630
rect 13012 26628 13036 26630
rect 13092 26628 13116 26630
rect 13172 26628 13196 26630
rect 13252 26628 13258 26630
rect 12950 26619 13258 26628
rect 13372 26382 13400 27950
rect 13360 26376 13412 26382
rect 13360 26318 13412 26324
rect 13360 26240 13412 26246
rect 13360 26182 13412 26188
rect 12950 25596 13258 25605
rect 12950 25594 12956 25596
rect 13012 25594 13036 25596
rect 13092 25594 13116 25596
rect 13172 25594 13196 25596
rect 13252 25594 13258 25596
rect 13012 25542 13014 25594
rect 13194 25542 13196 25594
rect 12950 25540 12956 25542
rect 13012 25540 13036 25542
rect 13092 25540 13116 25542
rect 13172 25540 13196 25542
rect 13252 25540 13258 25542
rect 12950 25531 13258 25540
rect 13372 25498 13400 26182
rect 13360 25492 13412 25498
rect 13360 25434 13412 25440
rect 13268 25424 13320 25430
rect 13320 25372 13400 25378
rect 13268 25366 13400 25372
rect 13280 25350 13400 25366
rect 12950 24508 13258 24517
rect 12950 24506 12956 24508
rect 13012 24506 13036 24508
rect 13092 24506 13116 24508
rect 13172 24506 13196 24508
rect 13252 24506 13258 24508
rect 13012 24454 13014 24506
rect 13194 24454 13196 24506
rect 12950 24452 12956 24454
rect 13012 24452 13036 24454
rect 13092 24452 13116 24454
rect 13172 24452 13196 24454
rect 13252 24452 13258 24454
rect 12950 24443 13258 24452
rect 12992 24404 13044 24410
rect 12992 24346 13044 24352
rect 13004 24138 13032 24346
rect 12992 24132 13044 24138
rect 12992 24074 13044 24080
rect 13004 23730 13032 24074
rect 13372 24070 13400 25350
rect 13464 24750 13492 28630
rect 13556 27418 13584 34546
rect 13648 33454 13676 35391
rect 13728 33992 13780 33998
rect 13728 33934 13780 33940
rect 13740 33522 13768 33934
rect 13728 33516 13780 33522
rect 13728 33458 13780 33464
rect 13636 33448 13688 33454
rect 13636 33390 13688 33396
rect 13636 33312 13688 33318
rect 13636 33254 13688 33260
rect 13648 31482 13676 33254
rect 13636 31476 13688 31482
rect 13636 31418 13688 31424
rect 13740 30326 13768 33458
rect 13728 30320 13780 30326
rect 13728 30262 13780 30268
rect 13820 28620 13872 28626
rect 13820 28562 13872 28568
rect 13832 28506 13860 28562
rect 13648 28478 13860 28506
rect 13924 28506 13952 35584
rect 14188 35488 14240 35494
rect 14188 35430 14240 35436
rect 14200 35222 14228 35430
rect 14188 35216 14240 35222
rect 14188 35158 14240 35164
rect 14280 35080 14332 35086
rect 14280 35022 14332 35028
rect 14292 34134 14320 35022
rect 14280 34128 14332 34134
rect 14280 34070 14332 34076
rect 14384 33946 14412 35974
rect 14108 33918 14412 33946
rect 14004 32224 14056 32230
rect 14004 32166 14056 32172
rect 14016 30734 14044 32166
rect 14108 31958 14136 33918
rect 14280 33856 14332 33862
rect 14280 33798 14332 33804
rect 14292 32774 14320 33798
rect 14476 32978 14504 36518
rect 14464 32972 14516 32978
rect 14464 32914 14516 32920
rect 14372 32904 14424 32910
rect 14372 32846 14424 32852
rect 14280 32768 14332 32774
rect 14280 32710 14332 32716
rect 14188 32428 14240 32434
rect 14188 32370 14240 32376
rect 14200 32230 14228 32370
rect 14188 32224 14240 32230
rect 14188 32166 14240 32172
rect 14096 31952 14148 31958
rect 14096 31894 14148 31900
rect 14096 31136 14148 31142
rect 14292 31124 14320 32710
rect 14384 31142 14412 32846
rect 14096 31078 14148 31084
rect 14200 31096 14320 31124
rect 14372 31136 14424 31142
rect 14004 30728 14056 30734
rect 14004 30670 14056 30676
rect 14004 30592 14056 30598
rect 14004 30534 14056 30540
rect 14016 28642 14044 30534
rect 14108 29102 14136 31078
rect 14096 29096 14148 29102
rect 14096 29038 14148 29044
rect 14016 28614 14136 28642
rect 13924 28478 14044 28506
rect 13648 28218 13676 28478
rect 13728 28416 13780 28422
rect 13728 28358 13780 28364
rect 13912 28416 13964 28422
rect 13912 28358 13964 28364
rect 13636 28212 13688 28218
rect 13636 28154 13688 28160
rect 13556 27390 13676 27418
rect 13544 27328 13596 27334
rect 13544 27270 13596 27276
rect 13556 27062 13584 27270
rect 13544 27056 13596 27062
rect 13544 26998 13596 27004
rect 13544 26376 13596 26382
rect 13544 26318 13596 26324
rect 13556 25362 13584 26318
rect 13544 25356 13596 25362
rect 13544 25298 13596 25304
rect 13544 25220 13596 25226
rect 13544 25162 13596 25168
rect 13452 24744 13504 24750
rect 13452 24686 13504 24692
rect 13360 24064 13412 24070
rect 13360 24006 13412 24012
rect 13452 24064 13504 24070
rect 13452 24006 13504 24012
rect 12992 23724 13044 23730
rect 12992 23666 13044 23672
rect 12950 23420 13258 23429
rect 12950 23418 12956 23420
rect 13012 23418 13036 23420
rect 13092 23418 13116 23420
rect 13172 23418 13196 23420
rect 13252 23418 13258 23420
rect 13012 23366 13014 23418
rect 13194 23366 13196 23418
rect 12950 23364 12956 23366
rect 13012 23364 13036 23366
rect 13092 23364 13116 23366
rect 13172 23364 13196 23366
rect 13252 23364 13258 23366
rect 12950 23355 13258 23364
rect 12808 23180 12860 23186
rect 12808 23122 12860 23128
rect 12624 22636 12676 22642
rect 12624 22578 12676 22584
rect 12624 22432 12676 22438
rect 12624 22374 12676 22380
rect 12532 22092 12584 22098
rect 12532 22034 12584 22040
rect 12256 22024 12308 22030
rect 12256 21966 12308 21972
rect 12268 21418 12296 21966
rect 12438 21584 12494 21593
rect 12348 21548 12400 21554
rect 12438 21519 12494 21528
rect 12348 21490 12400 21496
rect 12256 21412 12308 21418
rect 12256 21354 12308 21360
rect 12164 20936 12216 20942
rect 12164 20878 12216 20884
rect 12256 20392 12308 20398
rect 12256 20334 12308 20340
rect 12072 20256 12124 20262
rect 12072 20198 12124 20204
rect 11796 19916 11848 19922
rect 11796 19858 11848 19864
rect 12164 19712 12216 19718
rect 12164 19654 12216 19660
rect 12072 19372 12124 19378
rect 12072 19314 12124 19320
rect 11612 19304 11664 19310
rect 11612 19246 11664 19252
rect 11624 18154 11652 19246
rect 11704 19168 11756 19174
rect 11704 19110 11756 19116
rect 11980 19168 12032 19174
rect 11980 19110 12032 19116
rect 11612 18148 11664 18154
rect 11612 18090 11664 18096
rect 11520 17876 11572 17882
rect 11520 17818 11572 17824
rect 11532 17202 11560 17818
rect 11520 17196 11572 17202
rect 11520 17138 11572 17144
rect 11532 16794 11560 17138
rect 11520 16788 11572 16794
rect 11520 16730 11572 16736
rect 11520 16584 11572 16590
rect 11624 16574 11652 18090
rect 11716 17338 11744 19110
rect 11888 18828 11940 18834
rect 11888 18770 11940 18776
rect 11704 17332 11756 17338
rect 11704 17274 11756 17280
rect 11796 17264 11848 17270
rect 11796 17206 11848 17212
rect 11572 16546 11652 16574
rect 11520 16526 11572 16532
rect 11244 16448 11296 16454
rect 11244 16390 11296 16396
rect 11152 16244 11204 16250
rect 11152 16186 11204 16192
rect 11256 15434 11284 16390
rect 11244 15428 11296 15434
rect 11244 15370 11296 15376
rect 11256 15026 11284 15370
rect 11532 15366 11560 16526
rect 11808 16046 11836 17206
rect 11900 16250 11928 18770
rect 11992 18766 12020 19110
rect 11980 18760 12032 18766
rect 11980 18702 12032 18708
rect 11980 18284 12032 18290
rect 11980 18226 12032 18232
rect 11888 16244 11940 16250
rect 11888 16186 11940 16192
rect 11796 16040 11848 16046
rect 11796 15982 11848 15988
rect 11704 15972 11756 15978
rect 11704 15914 11756 15920
rect 11520 15360 11572 15366
rect 11520 15302 11572 15308
rect 11244 15020 11296 15026
rect 11244 14962 11296 14968
rect 11256 14634 11284 14962
rect 11060 14612 11112 14618
rect 11256 14606 11376 14634
rect 11060 14554 11112 14560
rect 11348 14482 11376 14606
rect 10876 14476 10928 14482
rect 10876 14418 10928 14424
rect 11336 14476 11388 14482
rect 11336 14418 11388 14424
rect 10508 13388 10560 13394
rect 10508 13330 10560 13336
rect 10888 12306 10916 14418
rect 11348 14074 11376 14418
rect 11612 14272 11664 14278
rect 11612 14214 11664 14220
rect 11336 14068 11388 14074
rect 11336 14010 11388 14016
rect 10968 13388 11020 13394
rect 10968 13330 11020 13336
rect 10980 12986 11008 13330
rect 10968 12980 11020 12986
rect 10968 12922 11020 12928
rect 10876 12300 10928 12306
rect 10876 12242 10928 12248
rect 10416 11824 10468 11830
rect 10416 11766 10468 11772
rect 10980 11762 11008 12922
rect 10968 11756 11020 11762
rect 10968 11698 11020 11704
rect 10324 11688 10376 11694
rect 10324 11630 10376 11636
rect 10048 10736 10100 10742
rect 10048 10678 10100 10684
rect 10048 9648 10100 9654
rect 10048 9590 10100 9596
rect 9772 6316 9824 6322
rect 9772 6258 9824 6264
rect 9772 3936 9824 3942
rect 9772 3878 9824 3884
rect 9496 3732 9548 3738
rect 9496 3674 9548 3680
rect 9784 3534 9812 3878
rect 10060 3738 10088 9590
rect 10336 8566 10364 11630
rect 11624 11626 11652 14214
rect 11716 14074 11744 15914
rect 11992 15162 12020 18226
rect 12084 17338 12112 19314
rect 12072 17332 12124 17338
rect 12072 17274 12124 17280
rect 12072 16584 12124 16590
rect 12072 16526 12124 16532
rect 12084 16182 12112 16526
rect 12072 16176 12124 16182
rect 12072 16118 12124 16124
rect 12176 15706 12204 19654
rect 12268 18834 12296 20334
rect 12360 19446 12388 21490
rect 12348 19440 12400 19446
rect 12348 19382 12400 19388
rect 12256 18828 12308 18834
rect 12256 18770 12308 18776
rect 12348 18352 12400 18358
rect 12346 18320 12348 18329
rect 12400 18320 12402 18329
rect 12346 18255 12402 18264
rect 12452 16946 12480 21519
rect 12544 18630 12572 22034
rect 12636 19378 12664 22374
rect 12950 22332 13258 22341
rect 12950 22330 12956 22332
rect 13012 22330 13036 22332
rect 13092 22330 13116 22332
rect 13172 22330 13196 22332
rect 13252 22330 13258 22332
rect 13012 22278 13014 22330
rect 13194 22278 13196 22330
rect 12950 22276 12956 22278
rect 13012 22276 13036 22278
rect 13092 22276 13116 22278
rect 13172 22276 13196 22278
rect 13252 22276 13258 22278
rect 12950 22267 13258 22276
rect 12808 21888 12860 21894
rect 12808 21830 12860 21836
rect 12820 21690 12848 21830
rect 12808 21684 12860 21690
rect 12808 21626 12860 21632
rect 12716 21616 12768 21622
rect 12716 21558 12768 21564
rect 12728 19514 12756 21558
rect 12950 21244 13258 21253
rect 12950 21242 12956 21244
rect 13012 21242 13036 21244
rect 13092 21242 13116 21244
rect 13172 21242 13196 21244
rect 13252 21242 13258 21244
rect 13012 21190 13014 21242
rect 13194 21190 13196 21242
rect 12950 21188 12956 21190
rect 13012 21188 13036 21190
rect 13092 21188 13116 21190
rect 13172 21188 13196 21190
rect 13252 21188 13258 21190
rect 12950 21179 13258 21188
rect 12950 20156 13258 20165
rect 12950 20154 12956 20156
rect 13012 20154 13036 20156
rect 13092 20154 13116 20156
rect 13172 20154 13196 20156
rect 13252 20154 13258 20156
rect 13012 20102 13014 20154
rect 13194 20102 13196 20154
rect 12950 20100 12956 20102
rect 13012 20100 13036 20102
rect 13092 20100 13116 20102
rect 13172 20100 13196 20102
rect 13252 20100 13258 20102
rect 12950 20091 13258 20100
rect 12808 19780 12860 19786
rect 12808 19722 12860 19728
rect 12716 19508 12768 19514
rect 12716 19450 12768 19456
rect 12624 19372 12676 19378
rect 12624 19314 12676 19320
rect 12532 18624 12584 18630
rect 12532 18566 12584 18572
rect 12452 16918 12572 16946
rect 12438 16824 12494 16833
rect 12438 16759 12494 16768
rect 12164 15700 12216 15706
rect 12164 15642 12216 15648
rect 12348 15360 12400 15366
rect 12348 15302 12400 15308
rect 11980 15156 12032 15162
rect 11980 15098 12032 15104
rect 12360 14958 12388 15302
rect 12348 14952 12400 14958
rect 12348 14894 12400 14900
rect 12452 14634 12480 16759
rect 12360 14606 12480 14634
rect 11796 14544 11848 14550
rect 11796 14486 11848 14492
rect 11704 14068 11756 14074
rect 11704 14010 11756 14016
rect 11704 13796 11756 13802
rect 11704 13738 11756 13744
rect 11716 12850 11744 13738
rect 11704 12844 11756 12850
rect 11704 12786 11756 12792
rect 11716 12442 11744 12786
rect 11704 12436 11756 12442
rect 11704 12378 11756 12384
rect 11808 12322 11836 14486
rect 12360 13954 12388 14606
rect 12544 14074 12572 16918
rect 12532 14068 12584 14074
rect 12532 14010 12584 14016
rect 12360 13926 12572 13954
rect 12348 13184 12400 13190
rect 12348 13126 12400 13132
rect 11888 12708 11940 12714
rect 11888 12650 11940 12656
rect 11716 12294 11836 12322
rect 11612 11620 11664 11626
rect 11612 11562 11664 11568
rect 10324 8560 10376 8566
rect 10324 8502 10376 8508
rect 11058 7984 11114 7993
rect 11058 7919 11114 7928
rect 10600 5840 10652 5846
rect 10600 5782 10652 5788
rect 10508 3936 10560 3942
rect 10508 3878 10560 3884
rect 10048 3732 10100 3738
rect 10048 3674 10100 3680
rect 9404 3528 9456 3534
rect 9404 3470 9456 3476
rect 9772 3528 9824 3534
rect 9772 3470 9824 3476
rect 9312 3052 9364 3058
rect 9312 2994 9364 3000
rect 9036 2984 9088 2990
rect 9036 2926 9088 2932
rect 9048 800 9076 2926
rect 9416 800 9444 3470
rect 9784 800 9812 3470
rect 10520 2990 10548 3878
rect 10612 3058 10640 5782
rect 10876 3528 10928 3534
rect 10876 3470 10928 3476
rect 10600 3052 10652 3058
rect 10600 2994 10652 3000
rect 10508 2984 10560 2990
rect 10508 2926 10560 2932
rect 10140 2440 10192 2446
rect 10140 2382 10192 2388
rect 10152 800 10180 2382
rect 10520 800 10548 2926
rect 10888 800 10916 3470
rect 11072 2650 11100 7919
rect 11612 4072 11664 4078
rect 11612 4014 11664 4020
rect 11244 3392 11296 3398
rect 11244 3334 11296 3340
rect 11256 3058 11284 3334
rect 11244 3052 11296 3058
rect 11244 2994 11296 3000
rect 11060 2644 11112 2650
rect 11060 2586 11112 2592
rect 11256 800 11284 2994
rect 11624 800 11652 4014
rect 11716 2446 11744 12294
rect 11796 12232 11848 12238
rect 11796 12174 11848 12180
rect 11808 11762 11836 12174
rect 11796 11756 11848 11762
rect 11796 11698 11848 11704
rect 11796 11620 11848 11626
rect 11796 11562 11848 11568
rect 11808 6458 11836 11562
rect 11796 6452 11848 6458
rect 11796 6394 11848 6400
rect 11900 5846 11928 12650
rect 12072 12640 12124 12646
rect 12072 12582 12124 12588
rect 12084 12306 12112 12582
rect 12072 12300 12124 12306
rect 12072 12242 12124 12248
rect 11980 11552 12032 11558
rect 11980 11494 12032 11500
rect 11888 5840 11940 5846
rect 11888 5782 11940 5788
rect 11992 4146 12020 11494
rect 12360 11218 12388 13126
rect 12348 11212 12400 11218
rect 12348 11154 12400 11160
rect 12544 10690 12572 13926
rect 12452 10662 12572 10690
rect 12452 9586 12480 10662
rect 12532 10532 12584 10538
rect 12532 10474 12584 10480
rect 12440 9580 12492 9586
rect 12440 9522 12492 9528
rect 11980 4140 12032 4146
rect 11980 4082 12032 4088
rect 11886 3224 11942 3233
rect 11886 3159 11888 3168
rect 11940 3159 11942 3168
rect 11888 3130 11940 3136
rect 11980 2508 12032 2514
rect 11980 2450 12032 2456
rect 11704 2440 11756 2446
rect 11704 2382 11756 2388
rect 11992 800 12020 2450
rect 12544 2446 12572 10474
rect 12636 10062 12664 19314
rect 12820 18970 12848 19722
rect 12950 19068 13258 19077
rect 12950 19066 12956 19068
rect 13012 19066 13036 19068
rect 13092 19066 13116 19068
rect 13172 19066 13196 19068
rect 13252 19066 13258 19068
rect 13012 19014 13014 19066
rect 13194 19014 13196 19066
rect 12950 19012 12956 19014
rect 13012 19012 13036 19014
rect 13092 19012 13116 19014
rect 13172 19012 13196 19014
rect 13252 19012 13258 19014
rect 12950 19003 13258 19012
rect 12808 18964 12860 18970
rect 12808 18906 12860 18912
rect 13176 18624 13228 18630
rect 13176 18566 13228 18572
rect 13188 18426 13216 18566
rect 13176 18420 13228 18426
rect 13176 18362 13228 18368
rect 12950 17980 13258 17989
rect 12950 17978 12956 17980
rect 13012 17978 13036 17980
rect 13092 17978 13116 17980
rect 13172 17978 13196 17980
rect 13252 17978 13258 17980
rect 13012 17926 13014 17978
rect 13194 17926 13196 17978
rect 12950 17924 12956 17926
rect 13012 17924 13036 17926
rect 13092 17924 13116 17926
rect 13172 17924 13196 17926
rect 13252 17924 13258 17926
rect 12950 17915 13258 17924
rect 12808 17128 12860 17134
rect 12808 17070 12860 17076
rect 12820 16833 12848 17070
rect 12950 16892 13258 16901
rect 12950 16890 12956 16892
rect 13012 16890 13036 16892
rect 13092 16890 13116 16892
rect 13172 16890 13196 16892
rect 13252 16890 13258 16892
rect 13012 16838 13014 16890
rect 13194 16838 13196 16890
rect 12950 16836 12956 16838
rect 13012 16836 13036 16838
rect 13092 16836 13116 16838
rect 13172 16836 13196 16838
rect 13252 16836 13258 16838
rect 12806 16824 12862 16833
rect 12950 16827 13258 16836
rect 12806 16759 12808 16768
rect 12860 16759 12862 16768
rect 12808 16730 12860 16736
rect 12950 15804 13258 15813
rect 12950 15802 12956 15804
rect 13012 15802 13036 15804
rect 13092 15802 13116 15804
rect 13172 15802 13196 15804
rect 13252 15802 13258 15804
rect 13012 15750 13014 15802
rect 13194 15750 13196 15802
rect 12950 15748 12956 15750
rect 13012 15748 13036 15750
rect 13092 15748 13116 15750
rect 13172 15748 13196 15750
rect 13252 15748 13258 15750
rect 12950 15739 13258 15748
rect 13268 15428 13320 15434
rect 13268 15370 13320 15376
rect 13280 15162 13308 15370
rect 13268 15156 13320 15162
rect 13268 15098 13320 15104
rect 12808 15020 12860 15026
rect 12808 14962 12860 14968
rect 12716 14340 12768 14346
rect 12716 14282 12768 14288
rect 12624 10056 12676 10062
rect 12624 9998 12676 10004
rect 12728 6914 12756 14282
rect 12820 12986 12848 14962
rect 12950 14716 13258 14725
rect 12950 14714 12956 14716
rect 13012 14714 13036 14716
rect 13092 14714 13116 14716
rect 13172 14714 13196 14716
rect 13252 14714 13258 14716
rect 13012 14662 13014 14714
rect 13194 14662 13196 14714
rect 12950 14660 12956 14662
rect 13012 14660 13036 14662
rect 13092 14660 13116 14662
rect 13172 14660 13196 14662
rect 13252 14660 13258 14662
rect 12950 14651 13258 14660
rect 13372 14074 13400 24006
rect 13464 23866 13492 24006
rect 13452 23860 13504 23866
rect 13452 23802 13504 23808
rect 13556 20602 13584 25162
rect 13648 21593 13676 27390
rect 13740 25226 13768 28358
rect 13820 27464 13872 27470
rect 13820 27406 13872 27412
rect 13832 26450 13860 27406
rect 13820 26444 13872 26450
rect 13820 26386 13872 26392
rect 13924 26042 13952 28358
rect 13912 26036 13964 26042
rect 13912 25978 13964 25984
rect 13912 25288 13964 25294
rect 13912 25230 13964 25236
rect 13728 25220 13780 25226
rect 13728 25162 13780 25168
rect 13728 24064 13780 24070
rect 13728 24006 13780 24012
rect 13740 23769 13768 24006
rect 13726 23760 13782 23769
rect 13726 23695 13782 23704
rect 13728 23588 13780 23594
rect 13728 23530 13780 23536
rect 13634 21584 13690 21593
rect 13634 21519 13690 21528
rect 13636 21480 13688 21486
rect 13636 21422 13688 21428
rect 13648 21146 13676 21422
rect 13636 21140 13688 21146
rect 13636 21082 13688 21088
rect 13740 20602 13768 23530
rect 13820 22976 13872 22982
rect 13820 22918 13872 22924
rect 13832 22166 13860 22918
rect 13924 22778 13952 25230
rect 14016 23866 14044 28478
rect 14108 27538 14136 28614
rect 14096 27532 14148 27538
rect 14096 27474 14148 27480
rect 14096 26784 14148 26790
rect 14096 26726 14148 26732
rect 14108 26450 14136 26726
rect 14096 26444 14148 26450
rect 14096 26386 14148 26392
rect 14096 25696 14148 25702
rect 14096 25638 14148 25644
rect 14108 25498 14136 25638
rect 14096 25492 14148 25498
rect 14096 25434 14148 25440
rect 14096 24336 14148 24342
rect 14096 24278 14148 24284
rect 14108 24206 14136 24278
rect 14096 24200 14148 24206
rect 14096 24142 14148 24148
rect 14004 23860 14056 23866
rect 14004 23802 14056 23808
rect 13912 22772 13964 22778
rect 13912 22714 13964 22720
rect 13820 22160 13872 22166
rect 13820 22102 13872 22108
rect 13924 22098 13952 22714
rect 14096 22568 14148 22574
rect 14096 22510 14148 22516
rect 13912 22092 13964 22098
rect 13912 22034 13964 22040
rect 14108 21894 14136 22510
rect 14200 22098 14228 31096
rect 14372 31078 14424 31084
rect 14280 30728 14332 30734
rect 14280 30670 14332 30676
rect 14188 22092 14240 22098
rect 14188 22034 14240 22040
rect 14096 21888 14148 21894
rect 14096 21830 14148 21836
rect 14096 21548 14148 21554
rect 14096 21490 14148 21496
rect 13912 21480 13964 21486
rect 13912 21422 13964 21428
rect 13820 21412 13872 21418
rect 13820 21354 13872 21360
rect 13832 20942 13860 21354
rect 13924 21350 13952 21422
rect 13912 21344 13964 21350
rect 13912 21286 13964 21292
rect 13820 20936 13872 20942
rect 13820 20878 13872 20884
rect 13544 20596 13596 20602
rect 13544 20538 13596 20544
rect 13728 20596 13780 20602
rect 13728 20538 13780 20544
rect 13452 19236 13504 19242
rect 13452 19178 13504 19184
rect 13464 18222 13492 19178
rect 13556 18970 13584 20538
rect 13740 19854 13768 20538
rect 13832 20534 13860 20878
rect 13820 20528 13872 20534
rect 13820 20470 13872 20476
rect 13728 19848 13780 19854
rect 13728 19790 13780 19796
rect 13636 19712 13688 19718
rect 13636 19654 13688 19660
rect 13544 18964 13596 18970
rect 13544 18906 13596 18912
rect 13542 18864 13598 18873
rect 13542 18799 13544 18808
rect 13596 18799 13598 18808
rect 13544 18770 13596 18776
rect 13556 18426 13584 18770
rect 13544 18420 13596 18426
rect 13544 18362 13596 18368
rect 13452 18216 13504 18222
rect 13452 18158 13504 18164
rect 13464 15094 13492 18158
rect 13648 17746 13676 19654
rect 13728 19304 13780 19310
rect 13726 19272 13728 19281
rect 13780 19272 13782 19281
rect 13726 19207 13782 19216
rect 13728 19168 13780 19174
rect 13728 19110 13780 19116
rect 13740 18834 13768 19110
rect 13728 18828 13780 18834
rect 13728 18770 13780 18776
rect 13636 17740 13688 17746
rect 13636 17682 13688 17688
rect 13636 17536 13688 17542
rect 13636 17478 13688 17484
rect 13648 16454 13676 17478
rect 13636 16448 13688 16454
rect 13636 16390 13688 16396
rect 13544 16244 13596 16250
rect 13544 16186 13596 16192
rect 13556 15910 13584 16186
rect 13648 16114 13676 16390
rect 13636 16108 13688 16114
rect 13636 16050 13688 16056
rect 13544 15904 13596 15910
rect 13544 15846 13596 15852
rect 13452 15088 13504 15094
rect 13452 15030 13504 15036
rect 13556 14482 13584 15846
rect 13740 15570 13768 18770
rect 13820 18216 13872 18222
rect 13820 18158 13872 18164
rect 13832 17542 13860 18158
rect 13820 17536 13872 17542
rect 13820 17478 13872 17484
rect 13832 16998 13860 17478
rect 13820 16992 13872 16998
rect 13820 16934 13872 16940
rect 13728 15564 13780 15570
rect 13728 15506 13780 15512
rect 13636 15496 13688 15502
rect 13636 15438 13688 15444
rect 13648 14890 13676 15438
rect 13728 15156 13780 15162
rect 13728 15098 13780 15104
rect 13636 14884 13688 14890
rect 13636 14826 13688 14832
rect 13544 14476 13596 14482
rect 13544 14418 13596 14424
rect 13452 14272 13504 14278
rect 13452 14214 13504 14220
rect 12900 14068 12952 14074
rect 12900 14010 12952 14016
rect 13360 14068 13412 14074
rect 13360 14010 13412 14016
rect 12912 13938 12940 14010
rect 12900 13932 12952 13938
rect 12900 13874 12952 13880
rect 12950 13628 13258 13637
rect 12950 13626 12956 13628
rect 13012 13626 13036 13628
rect 13092 13626 13116 13628
rect 13172 13626 13196 13628
rect 13252 13626 13258 13628
rect 13012 13574 13014 13626
rect 13194 13574 13196 13626
rect 12950 13572 12956 13574
rect 13012 13572 13036 13574
rect 13092 13572 13116 13574
rect 13172 13572 13196 13574
rect 13252 13572 13258 13574
rect 12950 13563 13258 13572
rect 13372 13258 13400 14010
rect 13360 13252 13412 13258
rect 13360 13194 13412 13200
rect 13358 13152 13414 13161
rect 13358 13087 13414 13096
rect 12808 12980 12860 12986
rect 12808 12922 12860 12928
rect 12950 12540 13258 12549
rect 12950 12538 12956 12540
rect 13012 12538 13036 12540
rect 13092 12538 13116 12540
rect 13172 12538 13196 12540
rect 13252 12538 13258 12540
rect 13012 12486 13014 12538
rect 13194 12486 13196 12538
rect 12950 12484 12956 12486
rect 13012 12484 13036 12486
rect 13092 12484 13116 12486
rect 13172 12484 13196 12486
rect 13252 12484 13258 12486
rect 12950 12475 13258 12484
rect 12950 11452 13258 11461
rect 12950 11450 12956 11452
rect 13012 11450 13036 11452
rect 13092 11450 13116 11452
rect 13172 11450 13196 11452
rect 13252 11450 13258 11452
rect 13012 11398 13014 11450
rect 13194 11398 13196 11450
rect 12950 11396 12956 11398
rect 13012 11396 13036 11398
rect 13092 11396 13116 11398
rect 13172 11396 13196 11398
rect 13252 11396 13258 11398
rect 12950 11387 13258 11396
rect 12950 10364 13258 10373
rect 12950 10362 12956 10364
rect 13012 10362 13036 10364
rect 13092 10362 13116 10364
rect 13172 10362 13196 10364
rect 13252 10362 13258 10364
rect 13012 10310 13014 10362
rect 13194 10310 13196 10362
rect 12950 10308 12956 10310
rect 13012 10308 13036 10310
rect 13092 10308 13116 10310
rect 13172 10308 13196 10310
rect 13252 10308 13258 10310
rect 12950 10299 13258 10308
rect 12950 9276 13258 9285
rect 12950 9274 12956 9276
rect 13012 9274 13036 9276
rect 13092 9274 13116 9276
rect 13172 9274 13196 9276
rect 13252 9274 13258 9276
rect 13012 9222 13014 9274
rect 13194 9222 13196 9274
rect 12950 9220 12956 9222
rect 13012 9220 13036 9222
rect 13092 9220 13116 9222
rect 13172 9220 13196 9222
rect 13252 9220 13258 9222
rect 12950 9211 13258 9220
rect 12950 8188 13258 8197
rect 12950 8186 12956 8188
rect 13012 8186 13036 8188
rect 13092 8186 13116 8188
rect 13172 8186 13196 8188
rect 13252 8186 13258 8188
rect 13012 8134 13014 8186
rect 13194 8134 13196 8186
rect 12950 8132 12956 8134
rect 13012 8132 13036 8134
rect 13092 8132 13116 8134
rect 13172 8132 13196 8134
rect 13252 8132 13258 8134
rect 12950 8123 13258 8132
rect 12950 7100 13258 7109
rect 12950 7098 12956 7100
rect 13012 7098 13036 7100
rect 13092 7098 13116 7100
rect 13172 7098 13196 7100
rect 13252 7098 13258 7100
rect 13012 7046 13014 7098
rect 13194 7046 13196 7098
rect 12950 7044 12956 7046
rect 13012 7044 13036 7046
rect 13092 7044 13116 7046
rect 13172 7044 13196 7046
rect 13252 7044 13258 7046
rect 12950 7035 13258 7044
rect 13372 6914 13400 13087
rect 13464 12442 13492 14214
rect 13556 13394 13584 14418
rect 13648 14346 13676 14826
rect 13636 14340 13688 14346
rect 13636 14282 13688 14288
rect 13544 13388 13596 13394
rect 13544 13330 13596 13336
rect 13636 13184 13688 13190
rect 13556 13144 13636 13172
rect 13452 12436 13504 12442
rect 13452 12378 13504 12384
rect 12728 6886 12848 6914
rect 13372 6886 13492 6914
rect 12624 5568 12676 5574
rect 12624 5510 12676 5516
rect 12636 3058 12664 5510
rect 12716 3596 12768 3602
rect 12716 3538 12768 3544
rect 12624 3052 12676 3058
rect 12624 2994 12676 3000
rect 12532 2440 12584 2446
rect 12532 2382 12584 2388
rect 12348 2372 12400 2378
rect 12348 2314 12400 2320
rect 12360 800 12388 2314
rect 12728 800 12756 3538
rect 12820 2582 12848 6886
rect 12950 6012 13258 6021
rect 12950 6010 12956 6012
rect 13012 6010 13036 6012
rect 13092 6010 13116 6012
rect 13172 6010 13196 6012
rect 13252 6010 13258 6012
rect 13012 5958 13014 6010
rect 13194 5958 13196 6010
rect 12950 5956 12956 5958
rect 13012 5956 13036 5958
rect 13092 5956 13116 5958
rect 13172 5956 13196 5958
rect 13252 5956 13258 5958
rect 12950 5947 13258 5956
rect 13464 5710 13492 6886
rect 13452 5704 13504 5710
rect 13452 5646 13504 5652
rect 12950 4924 13258 4933
rect 12950 4922 12956 4924
rect 13012 4922 13036 4924
rect 13092 4922 13116 4924
rect 13172 4922 13196 4924
rect 13252 4922 13258 4924
rect 13012 4870 13014 4922
rect 13194 4870 13196 4922
rect 12950 4868 12956 4870
rect 13012 4868 13036 4870
rect 13092 4868 13116 4870
rect 13172 4868 13196 4870
rect 13252 4868 13258 4870
rect 12950 4859 13258 4868
rect 13556 4146 13584 13144
rect 13636 13126 13688 13132
rect 13740 12714 13768 15098
rect 13832 14550 13860 16934
rect 13820 14544 13872 14550
rect 13820 14486 13872 14492
rect 13820 14272 13872 14278
rect 13820 14214 13872 14220
rect 13728 12708 13780 12714
rect 13728 12650 13780 12656
rect 13832 12434 13860 14214
rect 13648 12406 13860 12434
rect 13544 4140 13596 4146
rect 13544 4082 13596 4088
rect 13452 4072 13504 4078
rect 13452 4014 13504 4020
rect 12950 3836 13258 3845
rect 12950 3834 12956 3836
rect 13012 3834 13036 3836
rect 13092 3834 13116 3836
rect 13172 3834 13196 3836
rect 13252 3834 13258 3836
rect 13012 3782 13014 3834
rect 13194 3782 13196 3834
rect 12950 3780 12956 3782
rect 13012 3780 13036 3782
rect 13092 3780 13116 3782
rect 13172 3780 13196 3782
rect 13252 3780 13258 3782
rect 12950 3771 13258 3780
rect 13360 2984 13412 2990
rect 13360 2926 13412 2932
rect 12950 2748 13258 2757
rect 12950 2746 12956 2748
rect 13012 2746 13036 2748
rect 13092 2746 13116 2748
rect 13172 2746 13196 2748
rect 13252 2746 13258 2748
rect 13012 2694 13014 2746
rect 13194 2694 13196 2746
rect 12950 2692 12956 2694
rect 13012 2692 13036 2694
rect 13092 2692 13116 2694
rect 13172 2692 13196 2694
rect 13252 2692 13258 2694
rect 12950 2683 13258 2692
rect 12808 2576 12860 2582
rect 12808 2518 12860 2524
rect 13096 870 13216 898
rect 13096 800 13124 870
rect 1674 0 1730 800
rect 2042 0 2098 800
rect 2410 0 2466 800
rect 2778 0 2834 800
rect 3146 0 3202 800
rect 3514 0 3570 800
rect 3882 0 3938 800
rect 4250 0 4306 800
rect 4618 0 4674 800
rect 4986 0 5042 800
rect 5354 0 5410 800
rect 5722 0 5778 800
rect 6090 0 6146 800
rect 6458 0 6514 800
rect 6826 0 6882 800
rect 7194 0 7250 800
rect 7562 0 7618 800
rect 7930 0 7986 800
rect 8298 0 8354 800
rect 8666 0 8722 800
rect 9034 0 9090 800
rect 9402 0 9458 800
rect 9770 0 9826 800
rect 10138 0 10194 800
rect 10506 0 10562 800
rect 10874 0 10930 800
rect 11242 0 11298 800
rect 11610 0 11666 800
rect 11978 0 12034 800
rect 12346 0 12402 800
rect 12714 0 12770 800
rect 13082 0 13138 800
rect 13188 762 13216 870
rect 13372 762 13400 2926
rect 13464 800 13492 4014
rect 13648 3534 13676 12406
rect 13728 12096 13780 12102
rect 13728 12038 13780 12044
rect 13740 11830 13768 12038
rect 13728 11824 13780 11830
rect 13728 11766 13780 11772
rect 13924 8906 13952 21286
rect 14004 20868 14056 20874
rect 14004 20810 14056 20816
rect 14016 20534 14044 20810
rect 14004 20528 14056 20534
rect 14004 20470 14056 20476
rect 14016 19990 14044 20470
rect 14004 19984 14056 19990
rect 14004 19926 14056 19932
rect 14004 19440 14056 19446
rect 14004 19382 14056 19388
rect 14016 19174 14044 19382
rect 14004 19168 14056 19174
rect 14004 19110 14056 19116
rect 14004 18692 14056 18698
rect 14004 18634 14056 18640
rect 14016 18426 14044 18634
rect 14004 18420 14056 18426
rect 14004 18362 14056 18368
rect 14108 17202 14136 21490
rect 14200 21350 14228 22034
rect 14292 21486 14320 30670
rect 14568 30054 14596 44492
rect 14660 43450 14688 52838
rect 15764 52601 15792 53382
rect 15856 53106 15884 56200
rect 16224 54330 16252 56200
rect 16212 54324 16264 54330
rect 16212 54266 16264 54272
rect 16212 54052 16264 54058
rect 16212 53994 16264 54000
rect 16120 53984 16172 53990
rect 16120 53926 16172 53932
rect 15844 53100 15896 53106
rect 15844 53042 15896 53048
rect 15936 52896 15988 52902
rect 15936 52838 15988 52844
rect 15750 52592 15806 52601
rect 15750 52527 15806 52536
rect 15948 47802 15976 52838
rect 16028 48000 16080 48006
rect 16028 47942 16080 47948
rect 15936 47796 15988 47802
rect 15936 47738 15988 47744
rect 16040 46986 16068 47942
rect 16028 46980 16080 46986
rect 16028 46922 16080 46928
rect 16132 45554 16160 53926
rect 15948 45526 16160 45554
rect 15292 45280 15344 45286
rect 15292 45222 15344 45228
rect 14832 44192 14884 44198
rect 14832 44134 14884 44140
rect 14648 43444 14700 43450
rect 14648 43386 14700 43392
rect 14648 43240 14700 43246
rect 14648 43182 14700 43188
rect 14660 42770 14688 43182
rect 14740 43172 14792 43178
rect 14740 43114 14792 43120
rect 14648 42764 14700 42770
rect 14648 42706 14700 42712
rect 14752 40186 14780 43114
rect 14844 42158 14872 44134
rect 15016 43648 15068 43654
rect 15016 43590 15068 43596
rect 14924 43104 14976 43110
rect 14924 43046 14976 43052
rect 14832 42152 14884 42158
rect 14832 42094 14884 42100
rect 14740 40180 14792 40186
rect 14740 40122 14792 40128
rect 14648 39840 14700 39846
rect 14648 39782 14700 39788
rect 14660 39030 14688 39782
rect 14648 39024 14700 39030
rect 14648 38966 14700 38972
rect 14752 38962 14780 40122
rect 14832 39296 14884 39302
rect 14832 39238 14884 39244
rect 14740 38956 14792 38962
rect 14740 38898 14792 38904
rect 14844 38418 14872 39238
rect 14832 38412 14884 38418
rect 14832 38354 14884 38360
rect 14936 36922 14964 43046
rect 15028 42634 15056 43590
rect 15016 42628 15068 42634
rect 15016 42570 15068 42576
rect 15304 42362 15332 45222
rect 15384 44804 15436 44810
rect 15384 44746 15436 44752
rect 15396 43926 15424 44746
rect 15384 43920 15436 43926
rect 15384 43862 15436 43868
rect 15292 42356 15344 42362
rect 15292 42298 15344 42304
rect 15108 42084 15160 42090
rect 15108 42026 15160 42032
rect 15016 40384 15068 40390
rect 15016 40326 15068 40332
rect 14924 36916 14976 36922
rect 14924 36858 14976 36864
rect 14832 36780 14884 36786
rect 14832 36722 14884 36728
rect 14844 36582 14872 36722
rect 14832 36576 14884 36582
rect 14832 36518 14884 36524
rect 15028 36310 15056 40326
rect 15120 40186 15148 42026
rect 15292 41472 15344 41478
rect 15292 41414 15344 41420
rect 15200 41132 15252 41138
rect 15200 41074 15252 41080
rect 15108 40180 15160 40186
rect 15108 40122 15160 40128
rect 15212 40050 15240 41074
rect 15304 40526 15332 41414
rect 15292 40520 15344 40526
rect 15292 40462 15344 40468
rect 15292 40112 15344 40118
rect 15292 40054 15344 40060
rect 15200 40044 15252 40050
rect 15200 39986 15252 39992
rect 15200 39296 15252 39302
rect 15200 39238 15252 39244
rect 15108 38888 15160 38894
rect 15108 38830 15160 38836
rect 15120 38554 15148 38830
rect 15108 38548 15160 38554
rect 15108 38490 15160 38496
rect 15106 38448 15162 38457
rect 15106 38383 15162 38392
rect 15120 37874 15148 38383
rect 15108 37868 15160 37874
rect 15108 37810 15160 37816
rect 15212 36378 15240 39238
rect 15304 37806 15332 40054
rect 15396 39506 15424 43862
rect 15844 43716 15896 43722
rect 15844 43658 15896 43664
rect 15856 40730 15884 43658
rect 15948 43314 15976 45526
rect 16224 44198 16252 53994
rect 16592 53786 16620 56200
rect 16960 54194 16988 56200
rect 16948 54188 17000 54194
rect 16948 54130 17000 54136
rect 17040 53984 17092 53990
rect 17040 53926 17092 53932
rect 16580 53780 16632 53786
rect 16580 53722 16632 53728
rect 16592 53582 16620 53722
rect 16580 53576 16632 53582
rect 16580 53518 16632 53524
rect 16856 53440 16908 53446
rect 16856 53382 16908 53388
rect 16868 52601 16896 53382
rect 16854 52592 16910 52601
rect 16854 52527 16910 52536
rect 16580 47456 16632 47462
rect 16580 47398 16632 47404
rect 16396 46912 16448 46918
rect 16396 46854 16448 46860
rect 16408 46646 16436 46854
rect 16396 46640 16448 46646
rect 16396 46582 16448 46588
rect 16408 46016 16436 46582
rect 16488 46504 16540 46510
rect 16488 46446 16540 46452
rect 16500 46170 16528 46446
rect 16488 46164 16540 46170
rect 16488 46106 16540 46112
rect 16488 46028 16540 46034
rect 16408 45988 16488 46016
rect 16488 45970 16540 45976
rect 16500 45558 16528 45970
rect 16592 45778 16620 47398
rect 16764 47116 16816 47122
rect 16764 47058 16816 47064
rect 16776 46578 16804 47058
rect 16948 46708 17000 46714
rect 16948 46650 17000 46656
rect 16764 46572 16816 46578
rect 16764 46514 16816 46520
rect 16776 46034 16804 46514
rect 16764 46028 16816 46034
rect 16764 45970 16816 45976
rect 16776 45914 16804 45970
rect 16776 45886 16896 45914
rect 16764 45824 16816 45830
rect 16592 45750 16712 45778
rect 16764 45766 16816 45772
rect 16488 45552 16540 45558
rect 16488 45494 16540 45500
rect 16500 45286 16528 45494
rect 16304 45280 16356 45286
rect 16304 45222 16356 45228
rect 16488 45280 16540 45286
rect 16488 45222 16540 45228
rect 16212 44192 16264 44198
rect 16212 44134 16264 44140
rect 16316 43790 16344 45222
rect 16500 44878 16528 45222
rect 16488 44872 16540 44878
rect 16488 44814 16540 44820
rect 16500 44538 16528 44814
rect 16488 44532 16540 44538
rect 16488 44474 16540 44480
rect 16304 43784 16356 43790
rect 16304 43726 16356 43732
rect 16028 43648 16080 43654
rect 16028 43590 16080 43596
rect 15936 43308 15988 43314
rect 15936 43250 15988 43256
rect 15948 43110 15976 43250
rect 15936 43104 15988 43110
rect 15936 43046 15988 43052
rect 15844 40724 15896 40730
rect 15844 40666 15896 40672
rect 15752 40520 15804 40526
rect 15752 40462 15804 40468
rect 15384 39500 15436 39506
rect 15384 39442 15436 39448
rect 15568 39500 15620 39506
rect 15568 39442 15620 39448
rect 15476 39024 15528 39030
rect 15476 38966 15528 38972
rect 15384 38888 15436 38894
rect 15384 38830 15436 38836
rect 15396 38758 15424 38830
rect 15384 38752 15436 38758
rect 15384 38694 15436 38700
rect 15384 38208 15436 38214
rect 15384 38150 15436 38156
rect 15396 38010 15424 38150
rect 15384 38004 15436 38010
rect 15384 37946 15436 37952
rect 15292 37800 15344 37806
rect 15292 37742 15344 37748
rect 15200 36372 15252 36378
rect 15200 36314 15252 36320
rect 15016 36304 15068 36310
rect 15016 36246 15068 36252
rect 14740 35624 14792 35630
rect 14740 35566 14792 35572
rect 15016 35624 15068 35630
rect 15016 35566 15068 35572
rect 14752 35290 14780 35566
rect 14740 35284 14792 35290
rect 14740 35226 14792 35232
rect 14924 34944 14976 34950
rect 14924 34886 14976 34892
rect 14832 34128 14884 34134
rect 14832 34070 14884 34076
rect 14844 32978 14872 34070
rect 14832 32972 14884 32978
rect 14832 32914 14884 32920
rect 14830 32872 14886 32881
rect 14830 32807 14886 32816
rect 14648 32768 14700 32774
rect 14648 32710 14700 32716
rect 14740 32768 14792 32774
rect 14740 32710 14792 32716
rect 14660 32026 14688 32710
rect 14752 32230 14780 32710
rect 14844 32230 14872 32807
rect 14740 32224 14792 32230
rect 14740 32166 14792 32172
rect 14832 32224 14884 32230
rect 14832 32166 14884 32172
rect 14648 32020 14700 32026
rect 14648 31962 14700 31968
rect 14556 30048 14608 30054
rect 14556 29990 14608 29996
rect 14464 28416 14516 28422
rect 14464 28358 14516 28364
rect 14476 27962 14504 28358
rect 14384 27946 14504 27962
rect 14384 27940 14516 27946
rect 14384 27934 14464 27940
rect 14280 21480 14332 21486
rect 14280 21422 14332 21428
rect 14188 21344 14240 21350
rect 14188 21286 14240 21292
rect 14096 17196 14148 17202
rect 14096 17138 14148 17144
rect 14108 16640 14136 17138
rect 14016 16612 14136 16640
rect 14016 15162 14044 16612
rect 14096 15632 14148 15638
rect 14096 15574 14148 15580
rect 14108 15162 14136 15574
rect 14004 15156 14056 15162
rect 14004 15098 14056 15104
rect 14096 15156 14148 15162
rect 14096 15098 14148 15104
rect 14200 15042 14228 21286
rect 14280 20800 14332 20806
rect 14280 20742 14332 20748
rect 14292 18970 14320 20742
rect 14384 18986 14412 27934
rect 14464 27882 14516 27888
rect 14568 27690 14596 29990
rect 14740 29096 14792 29102
rect 14740 29038 14792 29044
rect 14752 28218 14780 29038
rect 14740 28212 14792 28218
rect 14740 28154 14792 28160
rect 14476 27662 14596 27690
rect 14476 27402 14504 27662
rect 14556 27600 14608 27606
rect 14556 27542 14608 27548
rect 14464 27396 14516 27402
rect 14464 27338 14516 27344
rect 14464 23860 14516 23866
rect 14464 23802 14516 23808
rect 14476 19122 14504 23802
rect 14568 23186 14596 27542
rect 14752 27470 14780 28154
rect 14740 27464 14792 27470
rect 14740 27406 14792 27412
rect 14648 26852 14700 26858
rect 14648 26794 14700 26800
rect 14556 23180 14608 23186
rect 14556 23122 14608 23128
rect 14556 22976 14608 22982
rect 14660 22964 14688 26794
rect 14844 26738 14872 32166
rect 14936 31210 14964 34886
rect 15028 32298 15056 35566
rect 15200 34740 15252 34746
rect 15200 34682 15252 34688
rect 15016 32292 15068 32298
rect 15016 32234 15068 32240
rect 14924 31204 14976 31210
rect 14924 31146 14976 31152
rect 15028 31142 15056 32234
rect 15016 31136 15068 31142
rect 15016 31078 15068 31084
rect 15212 29306 15240 34682
rect 15304 34406 15332 37742
rect 15384 37664 15436 37670
rect 15384 37606 15436 37612
rect 15396 37262 15424 37606
rect 15384 37256 15436 37262
rect 15384 37198 15436 37204
rect 15396 35034 15424 37198
rect 15488 35698 15516 38966
rect 15580 36242 15608 39442
rect 15764 38894 15792 40462
rect 15752 38888 15804 38894
rect 15752 38830 15804 38836
rect 15660 38820 15712 38826
rect 15660 38762 15712 38768
rect 15568 36236 15620 36242
rect 15568 36178 15620 36184
rect 15672 36174 15700 38762
rect 15764 37806 15792 38830
rect 15948 38758 15976 43046
rect 16040 41070 16068 43590
rect 16120 43172 16172 43178
rect 16120 43114 16172 43120
rect 16132 42702 16160 43114
rect 16120 42696 16172 42702
rect 16120 42638 16172 42644
rect 16316 41682 16344 43726
rect 16396 43104 16448 43110
rect 16396 43046 16448 43052
rect 16408 42906 16436 43046
rect 16396 42900 16448 42906
rect 16396 42842 16448 42848
rect 16580 42832 16632 42838
rect 16580 42774 16632 42780
rect 16488 42696 16540 42702
rect 16488 42638 16540 42644
rect 16304 41676 16356 41682
rect 16304 41618 16356 41624
rect 16120 41540 16172 41546
rect 16120 41482 16172 41488
rect 16132 41206 16160 41482
rect 16120 41200 16172 41206
rect 16120 41142 16172 41148
rect 16028 41064 16080 41070
rect 16028 41006 16080 41012
rect 16120 39976 16172 39982
rect 16120 39918 16172 39924
rect 16132 39098 16160 39918
rect 16120 39092 16172 39098
rect 16120 39034 16172 39040
rect 15936 38752 15988 38758
rect 15934 38720 15936 38729
rect 15988 38720 15990 38729
rect 15934 38655 15990 38664
rect 15844 38344 15896 38350
rect 15844 38286 15896 38292
rect 15752 37800 15804 37806
rect 15752 37742 15804 37748
rect 15660 36168 15712 36174
rect 15660 36110 15712 36116
rect 15476 35692 15528 35698
rect 15476 35634 15528 35640
rect 15488 35154 15516 35634
rect 15660 35488 15712 35494
rect 15660 35430 15712 35436
rect 15476 35148 15528 35154
rect 15476 35090 15528 35096
rect 15396 35006 15516 35034
rect 15292 34400 15344 34406
rect 15292 34342 15344 34348
rect 15292 31816 15344 31822
rect 15292 31758 15344 31764
rect 15304 31686 15332 31758
rect 15292 31680 15344 31686
rect 15292 31622 15344 31628
rect 15384 30592 15436 30598
rect 15382 30560 15384 30569
rect 15436 30560 15438 30569
rect 15382 30495 15438 30504
rect 15292 29504 15344 29510
rect 15292 29446 15344 29452
rect 15304 29345 15332 29446
rect 15290 29336 15346 29345
rect 15200 29300 15252 29306
rect 15290 29271 15346 29280
rect 15200 29242 15252 29248
rect 15488 29152 15516 35006
rect 15672 34678 15700 35430
rect 15764 35290 15792 37742
rect 15752 35284 15804 35290
rect 15752 35226 15804 35232
rect 15752 35012 15804 35018
rect 15752 34954 15804 34960
rect 15764 34746 15792 34954
rect 15752 34740 15804 34746
rect 15752 34682 15804 34688
rect 15660 34672 15712 34678
rect 15660 34614 15712 34620
rect 15752 34468 15804 34474
rect 15752 34410 15804 34416
rect 15764 33318 15792 34410
rect 15752 33312 15804 33318
rect 15752 33254 15804 33260
rect 15750 31784 15806 31793
rect 15568 31748 15620 31754
rect 15568 31690 15620 31696
rect 15660 31748 15712 31754
rect 15750 31719 15806 31728
rect 15660 31690 15712 31696
rect 15580 31482 15608 31690
rect 15568 31476 15620 31482
rect 15568 31418 15620 31424
rect 15568 31272 15620 31278
rect 15672 31260 15700 31690
rect 15620 31232 15700 31260
rect 15568 31214 15620 31220
rect 15568 30592 15620 30598
rect 15568 30534 15620 30540
rect 15580 30190 15608 30534
rect 15672 30394 15700 31232
rect 15764 30938 15792 31719
rect 15752 30932 15804 30938
rect 15752 30874 15804 30880
rect 15660 30388 15712 30394
rect 15660 30330 15712 30336
rect 15568 30184 15620 30190
rect 15568 30126 15620 30132
rect 15856 29850 15884 38286
rect 16212 37868 16264 37874
rect 16212 37810 16264 37816
rect 16028 37732 16080 37738
rect 16028 37674 16080 37680
rect 15936 37120 15988 37126
rect 15936 37062 15988 37068
rect 15948 35834 15976 37062
rect 15936 35828 15988 35834
rect 15936 35770 15988 35776
rect 16040 34542 16068 37674
rect 16120 37120 16172 37126
rect 16120 37062 16172 37068
rect 16028 34536 16080 34542
rect 16028 34478 16080 34484
rect 16132 34456 16160 37062
rect 16224 36378 16252 37810
rect 16316 37466 16344 41618
rect 16396 41472 16448 41478
rect 16396 41414 16448 41420
rect 16304 37460 16356 37466
rect 16304 37402 16356 37408
rect 16408 37330 16436 41414
rect 16500 41138 16528 42638
rect 16488 41132 16540 41138
rect 16488 41074 16540 41080
rect 16488 40996 16540 41002
rect 16488 40938 16540 40944
rect 16500 40050 16528 40938
rect 16592 40934 16620 42774
rect 16684 41614 16712 45750
rect 16776 44810 16804 45766
rect 16868 44946 16896 45886
rect 16960 45490 16988 46650
rect 16948 45484 17000 45490
rect 16948 45426 17000 45432
rect 16856 44940 16908 44946
rect 16856 44882 16908 44888
rect 16764 44804 16816 44810
rect 16764 44746 16816 44752
rect 16868 44402 16896 44882
rect 16856 44396 16908 44402
rect 16856 44338 16908 44344
rect 16764 44192 16816 44198
rect 16764 44134 16816 44140
rect 16672 41608 16724 41614
rect 16672 41550 16724 41556
rect 16580 40928 16632 40934
rect 16580 40870 16632 40876
rect 16580 40656 16632 40662
rect 16578 40624 16580 40633
rect 16632 40624 16634 40633
rect 16578 40559 16634 40568
rect 16580 40112 16632 40118
rect 16580 40054 16632 40060
rect 16488 40044 16540 40050
rect 16488 39986 16540 39992
rect 16500 37398 16528 39986
rect 16592 38554 16620 40054
rect 16672 39976 16724 39982
rect 16672 39918 16724 39924
rect 16684 38962 16712 39918
rect 16672 38956 16724 38962
rect 16672 38898 16724 38904
rect 16580 38548 16632 38554
rect 16580 38490 16632 38496
rect 16580 38208 16632 38214
rect 16580 38150 16632 38156
rect 16592 38010 16620 38150
rect 16580 38004 16632 38010
rect 16580 37946 16632 37952
rect 16488 37392 16540 37398
rect 16488 37334 16540 37340
rect 16396 37324 16448 37330
rect 16396 37266 16448 37272
rect 16670 36816 16726 36825
rect 16670 36751 16672 36760
rect 16724 36751 16726 36760
rect 16672 36722 16724 36728
rect 16212 36372 16264 36378
rect 16212 36314 16264 36320
rect 16672 36032 16724 36038
rect 16672 35974 16724 35980
rect 16488 35692 16540 35698
rect 16488 35634 16540 35640
rect 16132 34428 16252 34456
rect 15936 33924 15988 33930
rect 15936 33866 15988 33872
rect 15948 33114 15976 33866
rect 16120 33448 16172 33454
rect 16120 33390 16172 33396
rect 16028 33312 16080 33318
rect 16028 33254 16080 33260
rect 15936 33108 15988 33114
rect 15936 33050 15988 33056
rect 15936 32428 15988 32434
rect 15936 32370 15988 32376
rect 15948 32026 15976 32370
rect 15936 32020 15988 32026
rect 15936 31962 15988 31968
rect 16040 31754 16068 33254
rect 16132 32570 16160 33390
rect 16120 32564 16172 32570
rect 16120 32506 16172 32512
rect 16028 31748 16080 31754
rect 16028 31690 16080 31696
rect 16224 31634 16252 34428
rect 16396 34400 16448 34406
rect 16396 34342 16448 34348
rect 16408 34202 16436 34342
rect 16304 34196 16356 34202
rect 16304 34138 16356 34144
rect 16396 34196 16448 34202
rect 16396 34138 16448 34144
rect 16316 33810 16344 34138
rect 16316 33782 16436 33810
rect 16304 32904 16356 32910
rect 16304 32846 16356 32852
rect 15948 31606 16252 31634
rect 15948 30938 15976 31606
rect 16316 31396 16344 32846
rect 16408 31482 16436 33782
rect 16500 31686 16528 35634
rect 16684 35494 16712 35974
rect 16672 35488 16724 35494
rect 16672 35430 16724 35436
rect 16580 34944 16632 34950
rect 16580 34886 16632 34892
rect 16592 34066 16620 34886
rect 16580 34060 16632 34066
rect 16580 34002 16632 34008
rect 16592 33930 16620 34002
rect 16580 33924 16632 33930
rect 16580 33866 16632 33872
rect 16592 33318 16620 33866
rect 16580 33312 16632 33318
rect 16580 33254 16632 33260
rect 16580 33108 16632 33114
rect 16580 33050 16632 33056
rect 16592 32366 16620 33050
rect 16672 32836 16724 32842
rect 16672 32778 16724 32784
rect 16684 32502 16712 32778
rect 16672 32496 16724 32502
rect 16672 32438 16724 32444
rect 16580 32360 16632 32366
rect 16580 32302 16632 32308
rect 16488 31680 16540 31686
rect 16488 31622 16540 31628
rect 16580 31680 16632 31686
rect 16776 31634 16804 44134
rect 16868 43382 16896 44338
rect 16856 43376 16908 43382
rect 16856 43318 16908 43324
rect 16868 42770 16896 43318
rect 16948 43104 17000 43110
rect 16948 43046 17000 43052
rect 16856 42764 16908 42770
rect 16856 42706 16908 42712
rect 16868 41138 16896 42706
rect 16960 42362 16988 43046
rect 16948 42356 17000 42362
rect 16948 42298 17000 42304
rect 16856 41132 16908 41138
rect 16856 41074 16908 41080
rect 16946 40488 17002 40497
rect 16946 40423 17002 40432
rect 16856 40384 16908 40390
rect 16856 40326 16908 40332
rect 16868 39642 16896 40326
rect 16856 39636 16908 39642
rect 16856 39578 16908 39584
rect 16854 37768 16910 37777
rect 16854 37703 16910 37712
rect 16868 34610 16896 37703
rect 16960 36242 16988 40423
rect 17052 36378 17080 53926
rect 17328 53582 17356 56200
rect 17696 54262 17724 56200
rect 18064 56114 18092 56200
rect 18156 56114 18184 56222
rect 18064 56086 18184 56114
rect 17950 54428 18258 54437
rect 17950 54426 17956 54428
rect 18012 54426 18036 54428
rect 18092 54426 18116 54428
rect 18172 54426 18196 54428
rect 18252 54426 18258 54428
rect 18012 54374 18014 54426
rect 18194 54374 18196 54426
rect 17950 54372 17956 54374
rect 18012 54372 18036 54374
rect 18092 54372 18116 54374
rect 18172 54372 18196 54374
rect 18252 54372 18258 54374
rect 17950 54363 18258 54372
rect 17684 54256 17736 54262
rect 17684 54198 17736 54204
rect 18340 53582 18368 56222
rect 18418 56200 18474 57000
rect 18786 56200 18842 57000
rect 19154 56200 19210 57000
rect 19522 56200 19578 57000
rect 19890 56200 19946 57000
rect 20258 56200 20314 57000
rect 20626 56200 20682 57000
rect 20994 56200 21050 57000
rect 21362 56200 21418 57000
rect 21730 56200 21786 57000
rect 22098 56200 22154 57000
rect 22466 56200 22522 57000
rect 22834 56200 22890 57000
rect 23202 56200 23258 57000
rect 23570 56200 23626 57000
rect 24490 56264 24546 56273
rect 18432 54126 18460 56200
rect 18420 54120 18472 54126
rect 18420 54062 18472 54068
rect 18420 53984 18472 53990
rect 18420 53926 18472 53932
rect 17316 53576 17368 53582
rect 17316 53518 17368 53524
rect 18328 53576 18380 53582
rect 18328 53518 18380 53524
rect 17328 53242 17356 53518
rect 17408 53440 17460 53446
rect 17408 53382 17460 53388
rect 17316 53236 17368 53242
rect 17316 53178 17368 53184
rect 17420 47802 17448 53382
rect 17950 53340 18258 53349
rect 17950 53338 17956 53340
rect 18012 53338 18036 53340
rect 18092 53338 18116 53340
rect 18172 53338 18196 53340
rect 18252 53338 18258 53340
rect 18012 53286 18014 53338
rect 18194 53286 18196 53338
rect 17950 53284 17956 53286
rect 18012 53284 18036 53286
rect 18092 53284 18116 53286
rect 18172 53284 18196 53286
rect 18252 53284 18258 53286
rect 17950 53275 18258 53284
rect 17950 52252 18258 52261
rect 17950 52250 17956 52252
rect 18012 52250 18036 52252
rect 18092 52250 18116 52252
rect 18172 52250 18196 52252
rect 18252 52250 18258 52252
rect 18012 52198 18014 52250
rect 18194 52198 18196 52250
rect 17950 52196 17956 52198
rect 18012 52196 18036 52198
rect 18092 52196 18116 52198
rect 18172 52196 18196 52198
rect 18252 52196 18258 52198
rect 17950 52187 18258 52196
rect 17950 51164 18258 51173
rect 17950 51162 17956 51164
rect 18012 51162 18036 51164
rect 18092 51162 18116 51164
rect 18172 51162 18196 51164
rect 18252 51162 18258 51164
rect 18012 51110 18014 51162
rect 18194 51110 18196 51162
rect 17950 51108 17956 51110
rect 18012 51108 18036 51110
rect 18092 51108 18116 51110
rect 18172 51108 18196 51110
rect 18252 51108 18258 51110
rect 17950 51099 18258 51108
rect 17950 50076 18258 50085
rect 17950 50074 17956 50076
rect 18012 50074 18036 50076
rect 18092 50074 18116 50076
rect 18172 50074 18196 50076
rect 18252 50074 18258 50076
rect 18012 50022 18014 50074
rect 18194 50022 18196 50074
rect 17950 50020 17956 50022
rect 18012 50020 18036 50022
rect 18092 50020 18116 50022
rect 18172 50020 18196 50022
rect 18252 50020 18258 50022
rect 17950 50011 18258 50020
rect 17950 48988 18258 48997
rect 17950 48986 17956 48988
rect 18012 48986 18036 48988
rect 18092 48986 18116 48988
rect 18172 48986 18196 48988
rect 18252 48986 18258 48988
rect 18012 48934 18014 48986
rect 18194 48934 18196 48986
rect 17950 48932 17956 48934
rect 18012 48932 18036 48934
rect 18092 48932 18116 48934
rect 18172 48932 18196 48934
rect 18252 48932 18258 48934
rect 17950 48923 18258 48932
rect 18432 48278 18460 53926
rect 18512 53508 18564 53514
rect 18512 53450 18564 53456
rect 18420 48272 18472 48278
rect 18420 48214 18472 48220
rect 17950 47900 18258 47909
rect 17950 47898 17956 47900
rect 18012 47898 18036 47900
rect 18092 47898 18116 47900
rect 18172 47898 18196 47900
rect 18252 47898 18258 47900
rect 18012 47846 18014 47898
rect 18194 47846 18196 47898
rect 17950 47844 17956 47846
rect 18012 47844 18036 47846
rect 18092 47844 18116 47846
rect 18172 47844 18196 47846
rect 18252 47844 18258 47846
rect 17950 47835 18258 47844
rect 17408 47796 17460 47802
rect 17408 47738 17460 47744
rect 18432 47666 18460 48214
rect 18524 47802 18552 53450
rect 18800 53106 18828 56200
rect 18880 54256 18932 54262
rect 18880 54198 18932 54204
rect 18892 53786 18920 54198
rect 18880 53780 18932 53786
rect 18880 53722 18932 53728
rect 19168 53582 19196 56200
rect 19536 54194 19564 56200
rect 19524 54188 19576 54194
rect 19524 54130 19576 54136
rect 19708 54120 19760 54126
rect 19708 54062 19760 54068
rect 19340 54052 19392 54058
rect 19340 53994 19392 54000
rect 19156 53576 19208 53582
rect 19156 53518 19208 53524
rect 19168 53242 19196 53518
rect 19156 53236 19208 53242
rect 19156 53178 19208 53184
rect 18788 53100 18840 53106
rect 18788 53042 18840 53048
rect 18604 52896 18656 52902
rect 18604 52838 18656 52844
rect 18512 47796 18564 47802
rect 18512 47738 18564 47744
rect 18420 47660 18472 47666
rect 18420 47602 18472 47608
rect 18512 47660 18564 47666
rect 18512 47602 18564 47608
rect 17408 47592 17460 47598
rect 17408 47534 17460 47540
rect 17420 46714 17448 47534
rect 17500 47456 17552 47462
rect 17500 47398 17552 47404
rect 17408 46708 17460 46714
rect 17408 46650 17460 46656
rect 17316 44804 17368 44810
rect 17316 44746 17368 44752
rect 17224 43648 17276 43654
rect 17224 43590 17276 43596
rect 17132 42628 17184 42634
rect 17132 42570 17184 42576
rect 17144 41274 17172 42570
rect 17132 41268 17184 41274
rect 17132 41210 17184 41216
rect 17144 38350 17172 41210
rect 17236 40594 17264 43590
rect 17328 40594 17356 44746
rect 17512 43858 17540 47398
rect 18328 47184 18380 47190
rect 18328 47126 18380 47132
rect 17592 47116 17644 47122
rect 17592 47058 17644 47064
rect 17604 43858 17632 47058
rect 17776 46912 17828 46918
rect 17776 46854 17828 46860
rect 17788 46714 17816 46854
rect 17950 46812 18258 46821
rect 17950 46810 17956 46812
rect 18012 46810 18036 46812
rect 18092 46810 18116 46812
rect 18172 46810 18196 46812
rect 18252 46810 18258 46812
rect 18012 46758 18014 46810
rect 18194 46758 18196 46810
rect 17950 46756 17956 46758
rect 18012 46756 18036 46758
rect 18092 46756 18116 46758
rect 18172 46756 18196 46758
rect 18252 46756 18258 46758
rect 17950 46747 18258 46756
rect 17776 46708 17828 46714
rect 17776 46650 17828 46656
rect 17950 45724 18258 45733
rect 17950 45722 17956 45724
rect 18012 45722 18036 45724
rect 18092 45722 18116 45724
rect 18172 45722 18196 45724
rect 18252 45722 18258 45724
rect 18012 45670 18014 45722
rect 18194 45670 18196 45722
rect 17950 45668 17956 45670
rect 18012 45668 18036 45670
rect 18092 45668 18116 45670
rect 18172 45668 18196 45670
rect 18252 45668 18258 45670
rect 17950 45659 18258 45668
rect 17950 44636 18258 44645
rect 17950 44634 17956 44636
rect 18012 44634 18036 44636
rect 18092 44634 18116 44636
rect 18172 44634 18196 44636
rect 18252 44634 18258 44636
rect 18012 44582 18014 44634
rect 18194 44582 18196 44634
rect 17950 44580 17956 44582
rect 18012 44580 18036 44582
rect 18092 44580 18116 44582
rect 18172 44580 18196 44582
rect 18252 44580 18258 44582
rect 17950 44571 18258 44580
rect 17684 43920 17736 43926
rect 17684 43862 17736 43868
rect 17500 43852 17552 43858
rect 17500 43794 17552 43800
rect 17592 43852 17644 43858
rect 17592 43794 17644 43800
rect 17408 43784 17460 43790
rect 17408 43726 17460 43732
rect 17224 40588 17276 40594
rect 17224 40530 17276 40536
rect 17316 40588 17368 40594
rect 17316 40530 17368 40536
rect 17224 39296 17276 39302
rect 17224 39238 17276 39244
rect 17236 39030 17264 39238
rect 17224 39024 17276 39030
rect 17224 38966 17276 38972
rect 17132 38344 17184 38350
rect 17132 38286 17184 38292
rect 17130 37632 17186 37641
rect 17130 37567 17186 37576
rect 17144 36922 17172 37567
rect 17316 37120 17368 37126
rect 17316 37062 17368 37068
rect 17132 36916 17184 36922
rect 17132 36858 17184 36864
rect 17224 36848 17276 36854
rect 17224 36790 17276 36796
rect 17040 36372 17092 36378
rect 17040 36314 17092 36320
rect 16948 36236 17000 36242
rect 16948 36178 17000 36184
rect 16856 34604 16908 34610
rect 16856 34546 16908 34552
rect 17040 33108 17092 33114
rect 17040 33050 17092 33056
rect 17052 32978 17080 33050
rect 17236 32978 17264 36790
rect 17328 36650 17356 37062
rect 17316 36644 17368 36650
rect 17316 36586 17368 36592
rect 17316 35556 17368 35562
rect 17316 35498 17368 35504
rect 17328 35290 17356 35498
rect 17316 35284 17368 35290
rect 17316 35226 17368 35232
rect 17420 34082 17448 43726
rect 17696 43450 17724 43862
rect 17950 43548 18258 43557
rect 17950 43546 17956 43548
rect 18012 43546 18036 43548
rect 18092 43546 18116 43548
rect 18172 43546 18196 43548
rect 18252 43546 18258 43548
rect 18012 43494 18014 43546
rect 18194 43494 18196 43546
rect 17950 43492 17956 43494
rect 18012 43492 18036 43494
rect 18092 43492 18116 43494
rect 18172 43492 18196 43494
rect 18252 43492 18258 43494
rect 17950 43483 18258 43492
rect 17684 43444 17736 43450
rect 17684 43386 17736 43392
rect 18236 43308 18288 43314
rect 18236 43250 18288 43256
rect 17592 42764 17644 42770
rect 17592 42706 17644 42712
rect 17500 42220 17552 42226
rect 17500 42162 17552 42168
rect 17512 41750 17540 42162
rect 17500 41744 17552 41750
rect 17500 41686 17552 41692
rect 17604 41614 17632 42706
rect 18248 42702 18276 43250
rect 18236 42696 18288 42702
rect 18236 42638 18288 42644
rect 17950 42460 18258 42469
rect 17950 42458 17956 42460
rect 18012 42458 18036 42460
rect 18092 42458 18116 42460
rect 18172 42458 18196 42460
rect 18252 42458 18258 42460
rect 18012 42406 18014 42458
rect 18194 42406 18196 42458
rect 17950 42404 17956 42406
rect 18012 42404 18036 42406
rect 18092 42404 18116 42406
rect 18172 42404 18196 42406
rect 18252 42404 18258 42406
rect 17950 42395 18258 42404
rect 17776 42016 17828 42022
rect 17776 41958 17828 41964
rect 17592 41608 17644 41614
rect 17592 41550 17644 41556
rect 17592 40656 17644 40662
rect 17592 40598 17644 40604
rect 17500 38412 17552 38418
rect 17500 38354 17552 38360
rect 17512 38282 17540 38354
rect 17500 38276 17552 38282
rect 17500 38218 17552 38224
rect 17512 38010 17540 38218
rect 17500 38004 17552 38010
rect 17500 37946 17552 37952
rect 17604 36530 17632 40598
rect 17788 39982 17816 41958
rect 18340 41682 18368 47126
rect 18524 47054 18552 47602
rect 18616 47122 18644 52838
rect 18788 49088 18840 49094
rect 18788 49030 18840 49036
rect 18696 48136 18748 48142
rect 18696 48078 18748 48084
rect 18708 47598 18736 48078
rect 18696 47592 18748 47598
rect 18696 47534 18748 47540
rect 18604 47116 18656 47122
rect 18604 47058 18656 47064
rect 18512 47048 18564 47054
rect 18510 47016 18512 47025
rect 18564 47016 18566 47025
rect 18420 46980 18472 46986
rect 18510 46951 18566 46960
rect 18420 46922 18472 46928
rect 18432 46034 18460 46922
rect 18708 46714 18736 47534
rect 18696 46708 18748 46714
rect 18696 46650 18748 46656
rect 18800 46594 18828 49030
rect 19064 47796 19116 47802
rect 19064 47738 19116 47744
rect 18972 47728 19024 47734
rect 18972 47670 19024 47676
rect 18616 46566 18828 46594
rect 18420 46028 18472 46034
rect 18420 45970 18472 45976
rect 18512 45416 18564 45422
rect 18512 45358 18564 45364
rect 18524 44538 18552 45358
rect 18512 44532 18564 44538
rect 18512 44474 18564 44480
rect 18512 44328 18564 44334
rect 18512 44270 18564 44276
rect 18328 41676 18380 41682
rect 18328 41618 18380 41624
rect 18524 41614 18552 44270
rect 18616 42362 18644 46566
rect 18880 46504 18932 46510
rect 18880 46446 18932 46452
rect 18788 46368 18840 46374
rect 18788 46310 18840 46316
rect 18800 45898 18828 46310
rect 18788 45892 18840 45898
rect 18788 45834 18840 45840
rect 18696 45824 18748 45830
rect 18696 45766 18748 45772
rect 18708 44334 18736 45766
rect 18800 44742 18828 45834
rect 18892 45082 18920 46446
rect 18880 45076 18932 45082
rect 18880 45018 18932 45024
rect 18880 44872 18932 44878
rect 18880 44814 18932 44820
rect 18788 44736 18840 44742
rect 18788 44678 18840 44684
rect 18800 44470 18828 44678
rect 18788 44464 18840 44470
rect 18788 44406 18840 44412
rect 18696 44328 18748 44334
rect 18696 44270 18748 44276
rect 18800 43654 18828 44406
rect 18892 44198 18920 44814
rect 18880 44192 18932 44198
rect 18880 44134 18932 44140
rect 18788 43648 18840 43654
rect 18788 43590 18840 43596
rect 18788 42696 18840 42702
rect 18788 42638 18840 42644
rect 18604 42356 18656 42362
rect 18604 42298 18656 42304
rect 18512 41608 18564 41614
rect 18512 41550 18564 41556
rect 18328 41540 18380 41546
rect 18328 41482 18380 41488
rect 17950 41372 18258 41381
rect 17950 41370 17956 41372
rect 18012 41370 18036 41372
rect 18092 41370 18116 41372
rect 18172 41370 18196 41372
rect 18252 41370 18258 41372
rect 18012 41318 18014 41370
rect 18194 41318 18196 41370
rect 17950 41316 17956 41318
rect 18012 41316 18036 41318
rect 18092 41316 18116 41318
rect 18172 41316 18196 41318
rect 18252 41316 18258 41318
rect 17950 41307 18258 41316
rect 17868 40928 17920 40934
rect 17868 40870 17920 40876
rect 17880 40526 17908 40870
rect 17868 40520 17920 40526
rect 17868 40462 17920 40468
rect 17950 40284 18258 40293
rect 17950 40282 17956 40284
rect 18012 40282 18036 40284
rect 18092 40282 18116 40284
rect 18172 40282 18196 40284
rect 18252 40282 18258 40284
rect 18012 40230 18014 40282
rect 18194 40230 18196 40282
rect 17950 40228 17956 40230
rect 18012 40228 18036 40230
rect 18092 40228 18116 40230
rect 18172 40228 18196 40230
rect 18252 40228 18258 40230
rect 17950 40219 18258 40228
rect 18236 40180 18288 40186
rect 18236 40122 18288 40128
rect 18248 40089 18276 40122
rect 18234 40080 18290 40089
rect 18234 40015 18290 40024
rect 17776 39976 17828 39982
rect 17776 39918 17828 39924
rect 17950 39196 18258 39205
rect 17950 39194 17956 39196
rect 18012 39194 18036 39196
rect 18092 39194 18116 39196
rect 18172 39194 18196 39196
rect 18252 39194 18258 39196
rect 18012 39142 18014 39194
rect 18194 39142 18196 39194
rect 17950 39140 17956 39142
rect 18012 39140 18036 39142
rect 18092 39140 18116 39142
rect 18172 39140 18196 39142
rect 18252 39140 18258 39142
rect 17950 39131 18258 39140
rect 17950 38108 18258 38117
rect 17950 38106 17956 38108
rect 18012 38106 18036 38108
rect 18092 38106 18116 38108
rect 18172 38106 18196 38108
rect 18252 38106 18258 38108
rect 18012 38054 18014 38106
rect 18194 38054 18196 38106
rect 17950 38052 17956 38054
rect 18012 38052 18036 38054
rect 18092 38052 18116 38054
rect 18172 38052 18196 38054
rect 18252 38052 18258 38054
rect 17950 38043 18258 38052
rect 17868 37664 17920 37670
rect 17868 37606 17920 37612
rect 17880 37330 17908 37606
rect 17868 37324 17920 37330
rect 17868 37266 17920 37272
rect 17776 37188 17828 37194
rect 17776 37130 17828 37136
rect 17328 34054 17448 34082
rect 17512 36502 17632 36530
rect 17040 32972 17092 32978
rect 17040 32914 17092 32920
rect 17224 32972 17276 32978
rect 17224 32914 17276 32920
rect 17052 32858 17080 32914
rect 17052 32830 17172 32858
rect 16948 32768 17000 32774
rect 16948 32710 17000 32716
rect 16960 32298 16988 32710
rect 17040 32496 17092 32502
rect 17040 32438 17092 32444
rect 16948 32292 17000 32298
rect 16948 32234 17000 32240
rect 16856 32224 16908 32230
rect 16856 32166 16908 32172
rect 16632 31628 16804 31634
rect 16580 31622 16804 31628
rect 16396 31476 16448 31482
rect 16396 31418 16448 31424
rect 16132 31368 16344 31396
rect 15936 30932 15988 30938
rect 15936 30874 15988 30880
rect 15844 29844 15896 29850
rect 15844 29786 15896 29792
rect 15568 29776 15620 29782
rect 15568 29718 15620 29724
rect 15396 29124 15516 29152
rect 15016 28960 15068 28966
rect 15016 28902 15068 28908
rect 14752 26710 14872 26738
rect 14752 23866 14780 26710
rect 14832 26580 14884 26586
rect 14832 26522 14884 26528
rect 14844 25294 14872 26522
rect 14832 25288 14884 25294
rect 14832 25230 14884 25236
rect 14924 25152 14976 25158
rect 14924 25094 14976 25100
rect 14832 24200 14884 24206
rect 14832 24142 14884 24148
rect 14740 23860 14792 23866
rect 14740 23802 14792 23808
rect 14608 22936 14688 22964
rect 14556 22918 14608 22924
rect 14660 22642 14688 22936
rect 14648 22636 14700 22642
rect 14648 22578 14700 22584
rect 14556 22432 14608 22438
rect 14556 22374 14608 22380
rect 14568 21010 14596 22374
rect 14648 22228 14700 22234
rect 14648 22170 14700 22176
rect 14556 21004 14608 21010
rect 14556 20946 14608 20952
rect 14476 19094 14596 19122
rect 14280 18964 14332 18970
rect 14384 18958 14504 18986
rect 14280 18906 14332 18912
rect 14372 18896 14424 18902
rect 14372 18838 14424 18844
rect 14280 17060 14332 17066
rect 14280 17002 14332 17008
rect 14292 15201 14320 17002
rect 14278 15192 14334 15201
rect 14278 15127 14334 15136
rect 14108 15014 14228 15042
rect 14004 13388 14056 13394
rect 14004 13330 14056 13336
rect 14016 12986 14044 13330
rect 14004 12980 14056 12986
rect 14004 12922 14056 12928
rect 14108 9654 14136 15014
rect 14280 13320 14332 13326
rect 14280 13262 14332 13268
rect 14188 12776 14240 12782
rect 14188 12718 14240 12724
rect 14200 12374 14228 12718
rect 14188 12368 14240 12374
rect 14188 12310 14240 12316
rect 14292 12306 14320 13262
rect 14280 12300 14332 12306
rect 14280 12242 14332 12248
rect 14384 12238 14412 18838
rect 14476 17066 14504 18958
rect 14464 17060 14516 17066
rect 14464 17002 14516 17008
rect 14568 16522 14596 19094
rect 14660 18222 14688 22170
rect 14752 22094 14780 23802
rect 14844 23186 14872 24142
rect 14832 23180 14884 23186
rect 14832 23122 14884 23128
rect 14752 22066 14872 22094
rect 14740 19168 14792 19174
rect 14740 19110 14792 19116
rect 14752 18630 14780 19110
rect 14740 18624 14792 18630
rect 14738 18592 14740 18601
rect 14792 18592 14794 18601
rect 14738 18527 14794 18536
rect 14648 18216 14700 18222
rect 14648 18158 14700 18164
rect 14556 16516 14608 16522
rect 14556 16458 14608 16464
rect 14648 15360 14700 15366
rect 14568 15320 14648 15348
rect 14372 12232 14424 12238
rect 14372 12174 14424 12180
rect 14280 12096 14332 12102
rect 14280 12038 14332 12044
rect 14096 9648 14148 9654
rect 14096 9590 14148 9596
rect 13912 8900 13964 8906
rect 13912 8842 13964 8848
rect 13636 3528 13688 3534
rect 13636 3470 13688 3476
rect 14292 3058 14320 12038
rect 14568 5574 14596 15320
rect 14648 15302 14700 15308
rect 14740 14952 14792 14958
rect 14740 14894 14792 14900
rect 14648 13864 14700 13870
rect 14648 13806 14700 13812
rect 14556 5568 14608 5574
rect 14556 5510 14608 5516
rect 14280 3052 14332 3058
rect 14280 2994 14332 3000
rect 14188 2984 14240 2990
rect 14188 2926 14240 2932
rect 13820 2372 13872 2378
rect 13820 2314 13872 2320
rect 13832 800 13860 2314
rect 14200 800 14228 2926
rect 14556 2508 14608 2514
rect 14556 2450 14608 2456
rect 14568 800 14596 2450
rect 14660 2446 14688 13806
rect 14752 11898 14780 14894
rect 14844 14618 14872 22066
rect 14936 17678 14964 25094
rect 15028 23866 15056 28902
rect 15292 28552 15344 28558
rect 15292 28494 15344 28500
rect 15108 27124 15160 27130
rect 15108 27066 15160 27072
rect 15120 25362 15148 27066
rect 15108 25356 15160 25362
rect 15108 25298 15160 25304
rect 15200 24608 15252 24614
rect 15200 24550 15252 24556
rect 15016 23860 15068 23866
rect 15016 23802 15068 23808
rect 15108 22092 15160 22098
rect 15108 22034 15160 22040
rect 15016 22024 15068 22030
rect 15016 21966 15068 21972
rect 15028 21894 15056 21966
rect 15016 21888 15068 21894
rect 15016 21830 15068 21836
rect 15120 21350 15148 22034
rect 15108 21344 15160 21350
rect 15108 21286 15160 21292
rect 15016 21004 15068 21010
rect 15016 20946 15068 20952
rect 15028 20874 15056 20946
rect 15016 20868 15068 20874
rect 15016 20810 15068 20816
rect 15212 19922 15240 24550
rect 15304 21298 15332 28494
rect 15396 28257 15424 29124
rect 15476 29028 15528 29034
rect 15476 28970 15528 28976
rect 15382 28248 15438 28257
rect 15382 28183 15438 28192
rect 15384 28076 15436 28082
rect 15384 28018 15436 28024
rect 15396 27130 15424 28018
rect 15384 27124 15436 27130
rect 15384 27066 15436 27072
rect 15488 25294 15516 28970
rect 15580 26314 15608 29718
rect 15660 29708 15712 29714
rect 15660 29650 15712 29656
rect 15672 29238 15700 29650
rect 15660 29232 15712 29238
rect 15660 29174 15712 29180
rect 15660 28212 15712 28218
rect 15660 28154 15712 28160
rect 15568 26308 15620 26314
rect 15568 26250 15620 26256
rect 15476 25288 15528 25294
rect 15476 25230 15528 25236
rect 15384 24812 15436 24818
rect 15384 24754 15436 24760
rect 15396 23866 15424 24754
rect 15384 23860 15436 23866
rect 15384 23802 15436 23808
rect 15672 23746 15700 28154
rect 15752 24744 15804 24750
rect 15752 24686 15804 24692
rect 15764 23866 15792 24686
rect 15752 23860 15804 23866
rect 15752 23802 15804 23808
rect 15672 23718 15792 23746
rect 15764 23225 15792 23718
rect 15856 23322 15884 29786
rect 16132 28558 16160 31368
rect 16304 31272 16356 31278
rect 16304 31214 16356 31220
rect 16212 30660 16264 30666
rect 16212 30602 16264 30608
rect 16224 29850 16252 30602
rect 16316 30054 16344 31214
rect 16500 30802 16528 31622
rect 16592 31606 16804 31622
rect 16488 30796 16540 30802
rect 16488 30738 16540 30744
rect 16776 30376 16804 31606
rect 16500 30348 16804 30376
rect 16304 30048 16356 30054
rect 16304 29990 16356 29996
rect 16212 29844 16264 29850
rect 16212 29786 16264 29792
rect 16316 28626 16344 29990
rect 16396 29776 16448 29782
rect 16396 29718 16448 29724
rect 16304 28620 16356 28626
rect 16304 28562 16356 28568
rect 16120 28552 16172 28558
rect 16120 28494 16172 28500
rect 16212 28416 16264 28422
rect 16212 28358 16264 28364
rect 16120 28008 16172 28014
rect 16120 27950 16172 27956
rect 15936 27872 15988 27878
rect 15936 27814 15988 27820
rect 16028 27872 16080 27878
rect 16028 27814 16080 27820
rect 15948 27402 15976 27814
rect 16040 27674 16068 27814
rect 16028 27668 16080 27674
rect 16028 27610 16080 27616
rect 16132 27554 16160 27950
rect 16040 27526 16160 27554
rect 15936 27396 15988 27402
rect 15936 27338 15988 27344
rect 15948 26790 15976 27338
rect 15936 26784 15988 26790
rect 15936 26726 15988 26732
rect 15948 25906 15976 26726
rect 15936 25900 15988 25906
rect 15936 25842 15988 25848
rect 15844 23316 15896 23322
rect 15844 23258 15896 23264
rect 15750 23216 15806 23225
rect 15750 23151 15806 23160
rect 15568 22976 15620 22982
rect 15568 22918 15620 22924
rect 15304 21270 15516 21298
rect 15200 19916 15252 19922
rect 15200 19858 15252 19864
rect 15016 19236 15068 19242
rect 15016 19178 15068 19184
rect 15108 19236 15160 19242
rect 15108 19178 15160 19184
rect 15028 18630 15056 19178
rect 15120 18766 15148 19178
rect 15108 18760 15160 18766
rect 15108 18702 15160 18708
rect 15016 18624 15068 18630
rect 15016 18566 15068 18572
rect 15108 18216 15160 18222
rect 15108 18158 15160 18164
rect 15120 17898 15148 18158
rect 15488 17898 15516 21270
rect 15580 21010 15608 22918
rect 15660 21888 15712 21894
rect 15660 21830 15712 21836
rect 15672 21350 15700 21830
rect 15660 21344 15712 21350
rect 15660 21286 15712 21292
rect 15568 21004 15620 21010
rect 15568 20946 15620 20952
rect 15120 17870 15240 17898
rect 14924 17672 14976 17678
rect 14924 17614 14976 17620
rect 15212 16726 15240 17870
rect 15304 17870 15516 17898
rect 15200 16720 15252 16726
rect 15200 16662 15252 16668
rect 14924 16652 14976 16658
rect 14924 16594 14976 16600
rect 14832 14612 14884 14618
rect 14832 14554 14884 14560
rect 14844 14346 14872 14554
rect 14832 14340 14884 14346
rect 14832 14282 14884 14288
rect 14936 14226 14964 16594
rect 15212 16590 15240 16662
rect 15200 16584 15252 16590
rect 15200 16526 15252 16532
rect 15108 16448 15160 16454
rect 15108 16390 15160 16396
rect 15014 15736 15070 15745
rect 15014 15671 15016 15680
rect 15068 15671 15070 15680
rect 15016 15642 15068 15648
rect 15028 15502 15056 15642
rect 15016 15496 15068 15502
rect 15016 15438 15068 15444
rect 15120 14414 15148 16390
rect 15304 15706 15332 17870
rect 15476 17536 15528 17542
rect 15476 17478 15528 17484
rect 15568 17536 15620 17542
rect 15568 17478 15620 17484
rect 15384 17332 15436 17338
rect 15384 17274 15436 17280
rect 15292 15700 15344 15706
rect 15292 15642 15344 15648
rect 15200 15496 15252 15502
rect 15200 15438 15252 15444
rect 15212 14414 15240 15438
rect 15304 15162 15332 15642
rect 15292 15156 15344 15162
rect 15292 15098 15344 15104
rect 15108 14408 15160 14414
rect 15108 14350 15160 14356
rect 15200 14408 15252 14414
rect 15200 14350 15252 14356
rect 14844 14198 14964 14226
rect 14740 11892 14792 11898
rect 14740 11834 14792 11840
rect 14752 11150 14780 11834
rect 14740 11144 14792 11150
rect 14740 11086 14792 11092
rect 14844 10962 14872 14198
rect 14922 14104 14978 14113
rect 14922 14039 14924 14048
rect 14976 14039 14978 14048
rect 14924 14010 14976 14016
rect 14936 13938 14964 14010
rect 14924 13932 14976 13938
rect 14924 13874 14976 13880
rect 14924 13184 14976 13190
rect 14924 13126 14976 13132
rect 14936 11694 14964 13126
rect 15212 12986 15240 14350
rect 15396 13326 15424 17274
rect 15384 13320 15436 13326
rect 15384 13262 15436 13268
rect 15200 12980 15252 12986
rect 15200 12922 15252 12928
rect 15292 12912 15344 12918
rect 15488 12866 15516 17478
rect 15580 15434 15608 17478
rect 15764 17354 15792 23151
rect 15856 22778 15884 23258
rect 15844 22772 15896 22778
rect 15844 22714 15896 22720
rect 16040 22094 16068 27526
rect 16120 26920 16172 26926
rect 16120 26862 16172 26868
rect 16132 26790 16160 26862
rect 16120 26784 16172 26790
rect 16118 26752 16120 26761
rect 16172 26752 16174 26761
rect 16118 26687 16174 26696
rect 16120 26376 16172 26382
rect 16120 26318 16172 26324
rect 16132 24410 16160 26318
rect 16120 24404 16172 24410
rect 16120 24346 16172 24352
rect 16132 23662 16160 24346
rect 16120 23656 16172 23662
rect 16120 23598 16172 23604
rect 16120 22432 16172 22438
rect 16120 22374 16172 22380
rect 16132 22273 16160 22374
rect 16118 22264 16174 22273
rect 16118 22199 16174 22208
rect 16040 22066 16160 22094
rect 15936 21888 15988 21894
rect 15936 21830 15988 21836
rect 15842 21176 15898 21185
rect 15842 21111 15844 21120
rect 15896 21111 15898 21120
rect 15844 21082 15896 21088
rect 15844 20800 15896 20806
rect 15844 20742 15896 20748
rect 15672 17338 15792 17354
rect 15660 17332 15792 17338
rect 15712 17326 15792 17332
rect 15660 17274 15712 17280
rect 15752 17264 15804 17270
rect 15856 17252 15884 20742
rect 15948 20505 15976 21830
rect 16028 21140 16080 21146
rect 16028 21082 16080 21088
rect 15934 20496 15990 20505
rect 16040 20466 16068 21082
rect 15934 20431 15990 20440
rect 16028 20460 16080 20466
rect 16028 20402 16080 20408
rect 16028 19780 16080 19786
rect 16028 19722 16080 19728
rect 16040 19310 16068 19722
rect 15936 19304 15988 19310
rect 15936 19246 15988 19252
rect 16028 19304 16080 19310
rect 16028 19246 16080 19252
rect 15948 18970 15976 19246
rect 15936 18964 15988 18970
rect 15936 18906 15988 18912
rect 16040 18698 16068 19246
rect 16028 18692 16080 18698
rect 16028 18634 16080 18640
rect 15804 17224 15884 17252
rect 15752 17206 15804 17212
rect 15660 17128 15712 17134
rect 15660 17070 15712 17076
rect 15568 15428 15620 15434
rect 15568 15370 15620 15376
rect 15672 15026 15700 17070
rect 15764 16658 15792 17206
rect 15752 16652 15804 16658
rect 15752 16594 15804 16600
rect 16028 16584 16080 16590
rect 16028 16526 16080 16532
rect 15844 15428 15896 15434
rect 15844 15370 15896 15376
rect 15936 15428 15988 15434
rect 15936 15370 15988 15376
rect 15660 15020 15712 15026
rect 15660 14962 15712 14968
rect 15672 14618 15700 14962
rect 15660 14612 15712 14618
rect 15660 14554 15712 14560
rect 15568 14340 15620 14346
rect 15568 14282 15620 14288
rect 15580 14074 15608 14282
rect 15568 14068 15620 14074
rect 15568 14010 15620 14016
rect 15660 14000 15712 14006
rect 15660 13942 15712 13948
rect 15568 13864 15620 13870
rect 15568 13806 15620 13812
rect 15292 12854 15344 12860
rect 15200 12640 15252 12646
rect 15200 12582 15252 12588
rect 15016 12300 15068 12306
rect 15016 12242 15068 12248
rect 15028 11762 15056 12242
rect 15016 11756 15068 11762
rect 15016 11698 15068 11704
rect 14924 11688 14976 11694
rect 14924 11630 14976 11636
rect 14752 10934 14872 10962
rect 14752 3466 14780 10934
rect 14832 9988 14884 9994
rect 14832 9930 14884 9936
rect 14740 3460 14792 3466
rect 14740 3402 14792 3408
rect 14844 2582 14872 9930
rect 15212 7478 15240 12582
rect 15304 12170 15332 12854
rect 15396 12838 15516 12866
rect 15396 12646 15424 12838
rect 15476 12776 15528 12782
rect 15476 12718 15528 12724
rect 15384 12640 15436 12646
rect 15384 12582 15436 12588
rect 15292 12164 15344 12170
rect 15292 12106 15344 12112
rect 15488 11354 15516 12718
rect 15580 12102 15608 13806
rect 15568 12096 15620 12102
rect 15568 12038 15620 12044
rect 15476 11348 15528 11354
rect 15476 11290 15528 11296
rect 15200 7472 15252 7478
rect 15200 7414 15252 7420
rect 15580 6798 15608 12038
rect 15672 11830 15700 13942
rect 15752 12368 15804 12374
rect 15752 12310 15804 12316
rect 15764 12102 15792 12310
rect 15752 12096 15804 12102
rect 15752 12038 15804 12044
rect 15660 11824 15712 11830
rect 15660 11766 15712 11772
rect 15568 6792 15620 6798
rect 15568 6734 15620 6740
rect 15108 4208 15160 4214
rect 15108 4150 15160 4156
rect 14924 3596 14976 3602
rect 14924 3538 14976 3544
rect 14832 2576 14884 2582
rect 14832 2518 14884 2524
rect 14648 2440 14700 2446
rect 14648 2382 14700 2388
rect 14936 800 14964 3538
rect 15120 3534 15148 4150
rect 15108 3528 15160 3534
rect 15108 3470 15160 3476
rect 15660 2984 15712 2990
rect 15660 2926 15712 2932
rect 15292 2508 15344 2514
rect 15292 2450 15344 2456
rect 15304 800 15332 2450
rect 15672 800 15700 2926
rect 15764 2650 15792 12038
rect 15856 7410 15884 15370
rect 15948 15162 15976 15370
rect 15936 15156 15988 15162
rect 15936 15098 15988 15104
rect 16040 15042 16068 16526
rect 16132 16454 16160 22066
rect 16224 20942 16252 28358
rect 16408 27690 16436 29718
rect 16500 28490 16528 30348
rect 16672 29640 16724 29646
rect 16672 29582 16724 29588
rect 16488 28484 16540 28490
rect 16488 28426 16540 28432
rect 16408 27662 16528 27690
rect 16396 27532 16448 27538
rect 16396 27474 16448 27480
rect 16304 27124 16356 27130
rect 16304 27066 16356 27072
rect 16316 26450 16344 27066
rect 16304 26444 16356 26450
rect 16304 26386 16356 26392
rect 16316 25974 16344 26386
rect 16304 25968 16356 25974
rect 16304 25910 16356 25916
rect 16408 25702 16436 27474
rect 16396 25696 16448 25702
rect 16396 25638 16448 25644
rect 16408 24818 16436 25638
rect 16396 24812 16448 24818
rect 16396 24754 16448 24760
rect 16408 24274 16436 24754
rect 16396 24268 16448 24274
rect 16396 24210 16448 24216
rect 16500 24154 16528 27662
rect 16684 26450 16712 29582
rect 16764 29504 16816 29510
rect 16762 29472 16764 29481
rect 16816 29472 16818 29481
rect 16762 29407 16818 29416
rect 16868 28490 16896 32166
rect 16948 31952 17000 31958
rect 16948 31894 17000 31900
rect 16960 29306 16988 31894
rect 17052 31278 17080 32438
rect 17144 31754 17172 32830
rect 17144 31726 17264 31754
rect 17132 31340 17184 31346
rect 17132 31282 17184 31288
rect 17040 31272 17092 31278
rect 17040 31214 17092 31220
rect 17040 29504 17092 29510
rect 17040 29446 17092 29452
rect 16948 29300 17000 29306
rect 16948 29242 17000 29248
rect 17052 28558 17080 29446
rect 17040 28552 17092 28558
rect 17040 28494 17092 28500
rect 16856 28484 16908 28490
rect 16856 28426 16908 28432
rect 16856 26784 16908 26790
rect 16856 26726 16908 26732
rect 16672 26444 16724 26450
rect 16672 26386 16724 26392
rect 16672 26308 16724 26314
rect 16672 26250 16724 26256
rect 16580 25900 16632 25906
rect 16580 25842 16632 25848
rect 16592 25702 16620 25842
rect 16580 25696 16632 25702
rect 16580 25638 16632 25644
rect 16316 24126 16528 24154
rect 16592 24138 16620 25638
rect 16580 24132 16632 24138
rect 16212 20936 16264 20942
rect 16212 20878 16264 20884
rect 16316 17338 16344 24126
rect 16580 24074 16632 24080
rect 16592 23050 16620 24074
rect 16580 23044 16632 23050
rect 16580 22986 16632 22992
rect 16488 22092 16540 22098
rect 16488 22034 16540 22040
rect 16500 21146 16528 22034
rect 16580 22024 16632 22030
rect 16580 21966 16632 21972
rect 16592 21894 16620 21966
rect 16580 21888 16632 21894
rect 16580 21830 16632 21836
rect 16684 21350 16712 26250
rect 16764 26240 16816 26246
rect 16764 26182 16816 26188
rect 16776 26042 16804 26182
rect 16764 26036 16816 26042
rect 16764 25978 16816 25984
rect 16764 25152 16816 25158
rect 16764 25094 16816 25100
rect 16776 24750 16804 25094
rect 16764 24744 16816 24750
rect 16764 24686 16816 24692
rect 16868 24426 16896 26726
rect 17144 25770 17172 31282
rect 17236 27418 17264 31726
rect 17328 29646 17356 34054
rect 17408 32972 17460 32978
rect 17408 32914 17460 32920
rect 17420 30666 17448 32914
rect 17512 32502 17540 36502
rect 17592 36372 17644 36378
rect 17592 36314 17644 36320
rect 17500 32496 17552 32502
rect 17500 32438 17552 32444
rect 17604 31754 17632 36314
rect 17682 33144 17738 33153
rect 17682 33079 17684 33088
rect 17736 33079 17738 33088
rect 17684 33050 17736 33056
rect 17788 32570 17816 37130
rect 17950 37020 18258 37029
rect 17950 37018 17956 37020
rect 18012 37018 18036 37020
rect 18092 37018 18116 37020
rect 18172 37018 18196 37020
rect 18252 37018 18258 37020
rect 18012 36966 18014 37018
rect 18194 36966 18196 37018
rect 17950 36964 17956 36966
rect 18012 36964 18036 36966
rect 18092 36964 18116 36966
rect 18172 36964 18196 36966
rect 18252 36964 18258 36966
rect 17950 36955 18258 36964
rect 18340 36689 18368 41482
rect 18420 41472 18472 41478
rect 18420 41414 18472 41420
rect 18432 39982 18460 41414
rect 18420 39976 18472 39982
rect 18420 39918 18472 39924
rect 18524 38486 18552 41550
rect 18616 41414 18644 42298
rect 18800 42226 18828 42638
rect 18788 42220 18840 42226
rect 18788 42162 18840 42168
rect 18616 41386 18736 41414
rect 18604 41064 18656 41070
rect 18604 41006 18656 41012
rect 18616 40730 18644 41006
rect 18604 40724 18656 40730
rect 18604 40666 18656 40672
rect 18604 39500 18656 39506
rect 18604 39442 18656 39448
rect 18616 39098 18644 39442
rect 18604 39092 18656 39098
rect 18604 39034 18656 39040
rect 18512 38480 18564 38486
rect 18512 38422 18564 38428
rect 18420 38412 18472 38418
rect 18420 38354 18472 38360
rect 18432 38214 18460 38354
rect 18420 38208 18472 38214
rect 18420 38150 18472 38156
rect 18420 37732 18472 37738
rect 18420 37674 18472 37680
rect 18326 36680 18382 36689
rect 18326 36615 18382 36624
rect 18328 36576 18380 36582
rect 18328 36518 18380 36524
rect 17950 35932 18258 35941
rect 17950 35930 17956 35932
rect 18012 35930 18036 35932
rect 18092 35930 18116 35932
rect 18172 35930 18196 35932
rect 18252 35930 18258 35932
rect 18012 35878 18014 35930
rect 18194 35878 18196 35930
rect 17950 35876 17956 35878
rect 18012 35876 18036 35878
rect 18092 35876 18116 35878
rect 18172 35876 18196 35878
rect 18252 35876 18258 35878
rect 17950 35867 18258 35876
rect 18052 35760 18104 35766
rect 18052 35702 18104 35708
rect 18064 35154 18092 35702
rect 18340 35630 18368 36518
rect 18328 35624 18380 35630
rect 18432 35612 18460 37674
rect 18512 37120 18564 37126
rect 18512 37062 18564 37068
rect 18524 36922 18552 37062
rect 18512 36916 18564 36922
rect 18512 36858 18564 36864
rect 18616 36786 18644 39034
rect 18708 38554 18736 41386
rect 18788 40928 18840 40934
rect 18788 40870 18840 40876
rect 18800 39506 18828 40870
rect 18892 39982 18920 44134
rect 18984 41478 19012 47670
rect 18972 41472 19024 41478
rect 18972 41414 19024 41420
rect 18972 41200 19024 41206
rect 18972 41142 19024 41148
rect 18984 40934 19012 41142
rect 18972 40928 19024 40934
rect 18972 40870 19024 40876
rect 18880 39976 18932 39982
rect 18880 39918 18932 39924
rect 18788 39500 18840 39506
rect 18788 39442 18840 39448
rect 18984 39030 19012 40870
rect 18972 39024 19024 39030
rect 18972 38966 19024 38972
rect 18696 38548 18748 38554
rect 18696 38490 18748 38496
rect 18708 38010 18736 38490
rect 18788 38276 18840 38282
rect 18788 38218 18840 38224
rect 18696 38004 18748 38010
rect 18696 37946 18748 37952
rect 18696 37664 18748 37670
rect 18696 37606 18748 37612
rect 18708 37466 18736 37606
rect 18696 37460 18748 37466
rect 18696 37402 18748 37408
rect 18800 37346 18828 38218
rect 19076 38214 19104 47738
rect 19248 45416 19300 45422
rect 19352 45370 19380 53994
rect 19432 53984 19484 53990
rect 19432 53926 19484 53932
rect 19444 47734 19472 53926
rect 19616 53440 19668 53446
rect 19616 53382 19668 53388
rect 19432 47728 19484 47734
rect 19432 47670 19484 47676
rect 19628 46714 19656 53382
rect 19720 53242 19748 54062
rect 19904 53582 19932 56200
rect 19892 53576 19944 53582
rect 19892 53518 19944 53524
rect 19708 53236 19760 53242
rect 19708 53178 19760 53184
rect 20272 53106 20300 56200
rect 20640 55214 20668 56200
rect 20640 55186 20760 55214
rect 20732 54194 20760 55186
rect 20720 54188 20772 54194
rect 20720 54130 20772 54136
rect 20628 53508 20680 53514
rect 20628 53450 20680 53456
rect 20260 53100 20312 53106
rect 20260 53042 20312 53048
rect 20352 52896 20404 52902
rect 20352 52838 20404 52844
rect 19984 47048 20036 47054
rect 19984 46990 20036 46996
rect 19616 46708 19668 46714
rect 19616 46650 19668 46656
rect 19628 46617 19656 46650
rect 19614 46608 19670 46617
rect 19614 46543 19670 46552
rect 19800 46368 19852 46374
rect 19800 46310 19852 46316
rect 19524 45960 19576 45966
rect 19576 45920 19656 45948
rect 19524 45902 19576 45908
rect 19300 45364 19380 45370
rect 19248 45358 19380 45364
rect 19260 45342 19380 45358
rect 19352 44742 19380 45342
rect 19628 45286 19656 45920
rect 19616 45280 19668 45286
rect 19616 45222 19668 45228
rect 19628 44742 19656 45222
rect 19340 44736 19392 44742
rect 19338 44704 19340 44713
rect 19616 44736 19668 44742
rect 19392 44704 19394 44713
rect 19616 44678 19668 44684
rect 19338 44639 19394 44648
rect 19524 44192 19576 44198
rect 19524 44134 19576 44140
rect 19248 43648 19300 43654
rect 19248 43590 19300 43596
rect 19340 43648 19392 43654
rect 19340 43590 19392 43596
rect 19260 43382 19288 43590
rect 19248 43376 19300 43382
rect 19248 43318 19300 43324
rect 19260 42906 19288 43318
rect 19248 42900 19300 42906
rect 19248 42842 19300 42848
rect 19156 41472 19208 41478
rect 19156 41414 19208 41420
rect 19168 39574 19196 41414
rect 19260 41206 19288 42842
rect 19352 42294 19380 43590
rect 19536 43246 19564 44134
rect 19524 43240 19576 43246
rect 19524 43182 19576 43188
rect 19524 43104 19576 43110
rect 19524 43046 19576 43052
rect 19340 42288 19392 42294
rect 19340 42230 19392 42236
rect 19432 42152 19484 42158
rect 19432 42094 19484 42100
rect 19248 41200 19300 41206
rect 19248 41142 19300 41148
rect 19340 40928 19392 40934
rect 19340 40870 19392 40876
rect 19352 40186 19380 40870
rect 19340 40180 19392 40186
rect 19340 40122 19392 40128
rect 19248 39840 19300 39846
rect 19248 39782 19300 39788
rect 19156 39568 19208 39574
rect 19156 39510 19208 39516
rect 18880 38208 18932 38214
rect 18880 38150 18932 38156
rect 19064 38208 19116 38214
rect 19064 38150 19116 38156
rect 18892 37874 18920 38150
rect 18880 37868 18932 37874
rect 18880 37810 18932 37816
rect 18708 37318 18828 37346
rect 18708 36922 18736 37318
rect 18788 37256 18840 37262
rect 18788 37198 18840 37204
rect 18696 36916 18748 36922
rect 18696 36858 18748 36864
rect 18800 36786 18828 37198
rect 18604 36780 18656 36786
rect 18604 36722 18656 36728
rect 18788 36780 18840 36786
rect 18788 36722 18840 36728
rect 18696 35760 18748 35766
rect 18696 35702 18748 35708
rect 18604 35624 18656 35630
rect 18432 35584 18604 35612
rect 18328 35566 18380 35572
rect 18604 35566 18656 35572
rect 18052 35148 18104 35154
rect 18052 35090 18104 35096
rect 18328 35148 18380 35154
rect 18328 35090 18380 35096
rect 17950 34844 18258 34853
rect 17950 34842 17956 34844
rect 18012 34842 18036 34844
rect 18092 34842 18116 34844
rect 18172 34842 18196 34844
rect 18252 34842 18258 34844
rect 18012 34790 18014 34842
rect 18194 34790 18196 34842
rect 17950 34788 17956 34790
rect 18012 34788 18036 34790
rect 18092 34788 18116 34790
rect 18172 34788 18196 34790
rect 18252 34788 18258 34790
rect 17950 34779 18258 34788
rect 17868 34468 17920 34474
rect 17868 34410 17920 34416
rect 17776 32564 17828 32570
rect 17776 32506 17828 32512
rect 17776 32292 17828 32298
rect 17776 32234 17828 32240
rect 17684 32224 17736 32230
rect 17684 32166 17736 32172
rect 17696 31890 17724 32166
rect 17684 31884 17736 31890
rect 17684 31826 17736 31832
rect 17604 31726 17724 31754
rect 17408 30660 17460 30666
rect 17460 30620 17632 30648
rect 17408 30602 17460 30608
rect 17316 29640 17368 29646
rect 17500 29640 17552 29646
rect 17316 29582 17368 29588
rect 17420 29588 17500 29594
rect 17420 29582 17552 29588
rect 17420 29566 17540 29582
rect 17314 29336 17370 29345
rect 17314 29271 17316 29280
rect 17368 29271 17370 29280
rect 17316 29242 17368 29248
rect 17328 28422 17356 29242
rect 17420 29102 17448 29566
rect 17500 29504 17552 29510
rect 17500 29446 17552 29452
rect 17512 29306 17540 29446
rect 17500 29300 17552 29306
rect 17500 29242 17552 29248
rect 17604 29102 17632 30620
rect 17696 29594 17724 31726
rect 17788 30802 17816 32234
rect 17880 31906 17908 34410
rect 17950 33756 18258 33765
rect 17950 33754 17956 33756
rect 18012 33754 18036 33756
rect 18092 33754 18116 33756
rect 18172 33754 18196 33756
rect 18252 33754 18258 33756
rect 18012 33702 18014 33754
rect 18194 33702 18196 33754
rect 17950 33700 17956 33702
rect 18012 33700 18036 33702
rect 18092 33700 18116 33702
rect 18172 33700 18196 33702
rect 18252 33700 18258 33702
rect 17950 33691 18258 33700
rect 18340 33522 18368 35090
rect 18512 34944 18564 34950
rect 18512 34886 18564 34892
rect 18420 34400 18472 34406
rect 18420 34342 18472 34348
rect 18328 33516 18380 33522
rect 18328 33458 18380 33464
rect 17950 32668 18258 32677
rect 17950 32666 17956 32668
rect 18012 32666 18036 32668
rect 18092 32666 18116 32668
rect 18172 32666 18196 32668
rect 18252 32666 18258 32668
rect 18012 32614 18014 32666
rect 18194 32614 18196 32666
rect 17950 32612 17956 32614
rect 18012 32612 18036 32614
rect 18092 32612 18116 32614
rect 18172 32612 18196 32614
rect 18252 32612 18258 32614
rect 17950 32603 18258 32612
rect 17880 31890 18092 31906
rect 17880 31884 18104 31890
rect 17880 31878 18052 31884
rect 17776 30796 17828 30802
rect 17776 30738 17828 30744
rect 17788 29714 17816 30738
rect 17776 29708 17828 29714
rect 17776 29650 17828 29656
rect 17696 29566 17816 29594
rect 17684 29164 17736 29170
rect 17684 29106 17736 29112
rect 17408 29096 17460 29102
rect 17592 29096 17644 29102
rect 17460 29056 17540 29084
rect 17408 29038 17460 29044
rect 17316 28416 17368 28422
rect 17314 28384 17316 28393
rect 17368 28384 17370 28393
rect 17314 28319 17370 28328
rect 17236 27390 17448 27418
rect 17316 27328 17368 27334
rect 17316 27270 17368 27276
rect 17328 27062 17356 27270
rect 17316 27056 17368 27062
rect 17316 26998 17368 27004
rect 17224 26988 17276 26994
rect 17224 26930 17276 26936
rect 17236 26586 17264 26930
rect 17316 26920 17368 26926
rect 17314 26888 17316 26897
rect 17368 26888 17370 26897
rect 17314 26823 17370 26832
rect 17224 26580 17276 26586
rect 17224 26522 17276 26528
rect 17132 25764 17184 25770
rect 17132 25706 17184 25712
rect 17144 25362 17172 25706
rect 17420 25684 17448 27390
rect 17328 25656 17448 25684
rect 17132 25356 17184 25362
rect 17132 25298 17184 25304
rect 17132 24812 17184 24818
rect 17132 24754 17184 24760
rect 16776 24398 16896 24426
rect 16776 22030 16804 24398
rect 16856 23520 16908 23526
rect 16856 23462 16908 23468
rect 16764 22024 16816 22030
rect 16764 21966 16816 21972
rect 16764 21888 16816 21894
rect 16764 21830 16816 21836
rect 16580 21344 16632 21350
rect 16580 21286 16632 21292
rect 16672 21344 16724 21350
rect 16672 21286 16724 21292
rect 16592 21146 16620 21286
rect 16670 21176 16726 21185
rect 16488 21140 16540 21146
rect 16488 21082 16540 21088
rect 16580 21140 16632 21146
rect 16670 21111 16726 21120
rect 16580 21082 16632 21088
rect 16580 20052 16632 20058
rect 16580 19994 16632 20000
rect 16304 17332 16356 17338
rect 16304 17274 16356 17280
rect 16316 16794 16344 17274
rect 16488 16992 16540 16998
rect 16488 16934 16540 16940
rect 16304 16788 16356 16794
rect 16304 16730 16356 16736
rect 16120 16448 16172 16454
rect 16120 16390 16172 16396
rect 16210 16280 16266 16289
rect 16210 16215 16212 16224
rect 16264 16215 16266 16224
rect 16212 16186 16264 16192
rect 16304 15972 16356 15978
rect 16304 15914 16356 15920
rect 15948 15014 16068 15042
rect 15948 12434 15976 15014
rect 16120 14952 16172 14958
rect 16120 14894 16172 14900
rect 16132 13274 16160 14894
rect 16212 14884 16264 14890
rect 16212 14826 16264 14832
rect 16224 13394 16252 14826
rect 16316 14226 16344 15914
rect 16500 15162 16528 16934
rect 16488 15156 16540 15162
rect 16488 15098 16540 15104
rect 16316 14198 16436 14226
rect 16212 13388 16264 13394
rect 16212 13330 16264 13336
rect 16132 13246 16252 13274
rect 16120 12640 16172 12646
rect 16120 12582 16172 12588
rect 15948 12406 16068 12434
rect 16040 12306 16068 12406
rect 16132 12322 16160 12582
rect 16224 12442 16252 13246
rect 16304 13252 16356 13258
rect 16304 13194 16356 13200
rect 16212 12436 16264 12442
rect 16212 12378 16264 12384
rect 16028 12300 16080 12306
rect 16132 12294 16252 12322
rect 16028 12242 16080 12248
rect 16224 12170 16252 12294
rect 16212 12164 16264 12170
rect 16212 12106 16264 12112
rect 16224 11830 16252 12106
rect 16212 11824 16264 11830
rect 16212 11766 16264 11772
rect 16028 11280 16080 11286
rect 16026 11248 16028 11257
rect 16080 11248 16082 11257
rect 16026 11183 16082 11192
rect 16040 11150 16068 11183
rect 16028 11144 16080 11150
rect 16028 11086 16080 11092
rect 15844 7404 15896 7410
rect 15844 7346 15896 7352
rect 16212 7336 16264 7342
rect 16212 7278 16264 7284
rect 16224 4146 16252 7278
rect 16120 4140 16172 4146
rect 16120 4082 16172 4088
rect 16212 4140 16264 4146
rect 16212 4082 16264 4088
rect 16132 3670 16160 4082
rect 16120 3664 16172 3670
rect 16120 3606 16172 3612
rect 16028 3596 16080 3602
rect 16028 3538 16080 3544
rect 15752 2644 15804 2650
rect 15752 2586 15804 2592
rect 16040 800 16068 3538
rect 16316 3534 16344 13194
rect 16408 6914 16436 14198
rect 16592 13938 16620 19994
rect 16684 16250 16712 21111
rect 16776 17678 16804 21830
rect 16868 19854 16896 23462
rect 17040 23248 17092 23254
rect 17040 23190 17092 23196
rect 17052 22094 17080 23190
rect 17144 23186 17172 24754
rect 17224 24608 17276 24614
rect 17224 24550 17276 24556
rect 17236 23866 17264 24550
rect 17224 23860 17276 23866
rect 17224 23802 17276 23808
rect 17328 23730 17356 25656
rect 17512 25362 17540 29056
rect 17592 29038 17644 29044
rect 17592 28688 17644 28694
rect 17592 28630 17644 28636
rect 17500 25356 17552 25362
rect 17500 25298 17552 25304
rect 17408 25152 17460 25158
rect 17408 25094 17460 25100
rect 17316 23724 17368 23730
rect 17316 23666 17368 23672
rect 17132 23180 17184 23186
rect 17132 23122 17184 23128
rect 17144 22710 17172 23122
rect 17132 22704 17184 22710
rect 17132 22646 17184 22652
rect 17052 22066 17172 22094
rect 16856 19848 16908 19854
rect 16856 19790 16908 19796
rect 17144 19378 17172 22066
rect 17132 19372 17184 19378
rect 17132 19314 17184 19320
rect 16948 19304 17000 19310
rect 16948 19246 17000 19252
rect 16856 18828 16908 18834
rect 16856 18770 16908 18776
rect 16868 17678 16896 18770
rect 16764 17672 16816 17678
rect 16764 17614 16816 17620
rect 16856 17672 16908 17678
rect 16856 17614 16908 17620
rect 16868 16998 16896 17614
rect 16856 16992 16908 16998
rect 16856 16934 16908 16940
rect 16672 16244 16724 16250
rect 16672 16186 16724 16192
rect 16684 15094 16712 16186
rect 16672 15088 16724 15094
rect 16672 15030 16724 15036
rect 16764 14816 16816 14822
rect 16764 14758 16816 14764
rect 16580 13932 16632 13938
rect 16580 13874 16632 13880
rect 16776 11234 16804 14758
rect 16856 13184 16908 13190
rect 16856 13126 16908 13132
rect 16868 12918 16896 13126
rect 16856 12912 16908 12918
rect 16856 12854 16908 12860
rect 16960 12434 16988 19246
rect 17040 15904 17092 15910
rect 17040 15846 17092 15852
rect 17052 15502 17080 15846
rect 17040 15496 17092 15502
rect 17040 15438 17092 15444
rect 17052 14346 17080 15438
rect 17328 14414 17356 23666
rect 17420 18698 17448 25094
rect 17512 24886 17540 25298
rect 17604 25158 17632 28630
rect 17696 28422 17724 29106
rect 17684 28416 17736 28422
rect 17682 28384 17684 28393
rect 17736 28384 17738 28393
rect 17682 28319 17738 28328
rect 17682 28248 17738 28257
rect 17682 28183 17684 28192
rect 17736 28183 17738 28192
rect 17684 28154 17736 28160
rect 17788 27946 17816 29566
rect 17776 27940 17828 27946
rect 17776 27882 17828 27888
rect 17880 27554 17908 31878
rect 18052 31826 18104 31832
rect 18328 31680 18380 31686
rect 18328 31622 18380 31628
rect 17950 31580 18258 31589
rect 17950 31578 17956 31580
rect 18012 31578 18036 31580
rect 18092 31578 18116 31580
rect 18172 31578 18196 31580
rect 18252 31578 18258 31580
rect 18012 31526 18014 31578
rect 18194 31526 18196 31578
rect 17950 31524 17956 31526
rect 18012 31524 18036 31526
rect 18092 31524 18116 31526
rect 18172 31524 18196 31526
rect 18252 31524 18258 31526
rect 17950 31515 18258 31524
rect 18340 30598 18368 31622
rect 18328 30592 18380 30598
rect 18328 30534 18380 30540
rect 17950 30492 18258 30501
rect 17950 30490 17956 30492
rect 18012 30490 18036 30492
rect 18092 30490 18116 30492
rect 18172 30490 18196 30492
rect 18252 30490 18258 30492
rect 18012 30438 18014 30490
rect 18194 30438 18196 30490
rect 17950 30436 17956 30438
rect 18012 30436 18036 30438
rect 18092 30436 18116 30438
rect 18172 30436 18196 30438
rect 18252 30436 18258 30438
rect 17950 30427 18258 30436
rect 18340 30394 18368 30534
rect 18328 30388 18380 30394
rect 18328 30330 18380 30336
rect 18328 30048 18380 30054
rect 18328 29990 18380 29996
rect 18340 29714 18368 29990
rect 18328 29708 18380 29714
rect 18328 29650 18380 29656
rect 17950 29404 18258 29413
rect 17950 29402 17956 29404
rect 18012 29402 18036 29404
rect 18092 29402 18116 29404
rect 18172 29402 18196 29404
rect 18252 29402 18258 29404
rect 18012 29350 18014 29402
rect 18194 29350 18196 29402
rect 17950 29348 17956 29350
rect 18012 29348 18036 29350
rect 18092 29348 18116 29350
rect 18172 29348 18196 29350
rect 18252 29348 18258 29350
rect 17950 29339 18258 29348
rect 18432 29306 18460 34342
rect 18524 34202 18552 34886
rect 18512 34196 18564 34202
rect 18512 34138 18564 34144
rect 18512 32224 18564 32230
rect 18512 32166 18564 32172
rect 18420 29300 18472 29306
rect 18420 29242 18472 29248
rect 17960 29164 18012 29170
rect 17960 29106 18012 29112
rect 17972 28966 18000 29106
rect 18420 29028 18472 29034
rect 18420 28970 18472 28976
rect 17960 28960 18012 28966
rect 17960 28902 18012 28908
rect 17972 28762 18000 28902
rect 17960 28756 18012 28762
rect 17960 28698 18012 28704
rect 17950 28316 18258 28325
rect 17950 28314 17956 28316
rect 18012 28314 18036 28316
rect 18092 28314 18116 28316
rect 18172 28314 18196 28316
rect 18252 28314 18258 28316
rect 18012 28262 18014 28314
rect 18194 28262 18196 28314
rect 17950 28260 17956 28262
rect 18012 28260 18036 28262
rect 18092 28260 18116 28262
rect 18172 28260 18196 28262
rect 18252 28260 18258 28262
rect 17950 28251 18258 28260
rect 17960 27940 18012 27946
rect 17960 27882 18012 27888
rect 17972 27606 18000 27882
rect 18328 27872 18380 27878
rect 18328 27814 18380 27820
rect 17788 27526 17908 27554
rect 17960 27600 18012 27606
rect 17960 27542 18012 27548
rect 17684 27328 17736 27334
rect 17684 27270 17736 27276
rect 17592 25152 17644 25158
rect 17592 25094 17644 25100
rect 17500 24880 17552 24886
rect 17500 24822 17552 24828
rect 17512 23594 17540 24822
rect 17696 23866 17724 27270
rect 17788 27130 17816 27526
rect 17868 27464 17920 27470
rect 17868 27406 17920 27412
rect 17776 27124 17828 27130
rect 17776 27066 17828 27072
rect 17776 25696 17828 25702
rect 17776 25638 17828 25644
rect 17684 23860 17736 23866
rect 17684 23802 17736 23808
rect 17500 23588 17552 23594
rect 17500 23530 17552 23536
rect 17512 22574 17540 23530
rect 17500 22568 17552 22574
rect 17500 22510 17552 22516
rect 17592 22500 17644 22506
rect 17592 22442 17644 22448
rect 17500 21888 17552 21894
rect 17500 21830 17552 21836
rect 17512 21690 17540 21830
rect 17604 21690 17632 22442
rect 17788 22098 17816 25638
rect 17880 24732 17908 27406
rect 17950 27228 18258 27237
rect 17950 27226 17956 27228
rect 18012 27226 18036 27228
rect 18092 27226 18116 27228
rect 18172 27226 18196 27228
rect 18252 27226 18258 27228
rect 18012 27174 18014 27226
rect 18194 27174 18196 27226
rect 17950 27172 17956 27174
rect 18012 27172 18036 27174
rect 18092 27172 18116 27174
rect 18172 27172 18196 27174
rect 18252 27172 18258 27174
rect 17950 27163 18258 27172
rect 17960 26988 18012 26994
rect 17960 26930 18012 26936
rect 17972 26586 18000 26930
rect 18052 26784 18104 26790
rect 18052 26726 18104 26732
rect 17960 26580 18012 26586
rect 17960 26522 18012 26528
rect 18064 26450 18092 26726
rect 18052 26444 18104 26450
rect 18052 26386 18104 26392
rect 17950 26140 18258 26149
rect 17950 26138 17956 26140
rect 18012 26138 18036 26140
rect 18092 26138 18116 26140
rect 18172 26138 18196 26140
rect 18252 26138 18258 26140
rect 18012 26086 18014 26138
rect 18194 26086 18196 26138
rect 17950 26084 17956 26086
rect 18012 26084 18036 26086
rect 18092 26084 18116 26086
rect 18172 26084 18196 26086
rect 18252 26084 18258 26086
rect 17950 26075 18258 26084
rect 18340 26042 18368 27814
rect 18432 27470 18460 28970
rect 18420 27464 18472 27470
rect 18420 27406 18472 27412
rect 18524 26976 18552 32166
rect 18616 32026 18644 35566
rect 18708 34066 18736 35702
rect 18800 34746 18828 36722
rect 18788 34740 18840 34746
rect 18788 34682 18840 34688
rect 18696 34060 18748 34066
rect 18696 34002 18748 34008
rect 18708 33590 18736 34002
rect 18696 33584 18748 33590
rect 18696 33526 18748 33532
rect 18696 33040 18748 33046
rect 18696 32982 18748 32988
rect 18604 32020 18656 32026
rect 18604 31962 18656 31968
rect 18602 31920 18658 31929
rect 18602 31855 18604 31864
rect 18656 31855 18658 31864
rect 18604 31826 18656 31832
rect 18432 26948 18552 26976
rect 18328 26036 18380 26042
rect 18328 25978 18380 25984
rect 18432 25974 18460 26948
rect 18616 26874 18644 31826
rect 18708 30394 18736 32982
rect 18788 32428 18840 32434
rect 18788 32370 18840 32376
rect 18800 30784 18828 32370
rect 18892 31754 18920 37810
rect 19168 37754 19196 39510
rect 18984 37726 19196 37754
rect 18984 37505 19012 37726
rect 19064 37664 19116 37670
rect 19260 37641 19288 39782
rect 19444 39098 19472 42094
rect 19432 39092 19484 39098
rect 19432 39034 19484 39040
rect 19536 38962 19564 43046
rect 19628 42702 19656 44678
rect 19616 42696 19668 42702
rect 19616 42638 19668 42644
rect 19616 41472 19668 41478
rect 19616 41414 19668 41420
rect 19524 38956 19576 38962
rect 19524 38898 19576 38904
rect 19628 38010 19656 41414
rect 19812 41274 19840 46310
rect 19892 45824 19944 45830
rect 19892 45766 19944 45772
rect 19904 44402 19932 45766
rect 19996 45626 20024 46990
rect 20364 46714 20392 52838
rect 20444 47048 20496 47054
rect 20444 46990 20496 46996
rect 20352 46708 20404 46714
rect 20352 46650 20404 46656
rect 20352 46504 20404 46510
rect 20456 46492 20484 46990
rect 20640 46753 20668 53450
rect 20732 53174 20760 54130
rect 21008 53582 21036 56200
rect 21376 54194 21404 56200
rect 21364 54188 21416 54194
rect 21364 54130 21416 54136
rect 21088 53984 21140 53990
rect 21088 53926 21140 53932
rect 20996 53576 21048 53582
rect 20996 53518 21048 53524
rect 20904 53440 20956 53446
rect 20904 53382 20956 53388
rect 20720 53168 20772 53174
rect 20720 53110 20772 53116
rect 20626 46744 20682 46753
rect 20682 46714 20760 46730
rect 20682 46708 20772 46714
rect 20682 46702 20720 46708
rect 20626 46679 20682 46688
rect 20720 46650 20772 46656
rect 20404 46464 20484 46492
rect 20352 46446 20404 46452
rect 19984 45620 20036 45626
rect 19984 45562 20036 45568
rect 20260 45280 20312 45286
rect 20260 45222 20312 45228
rect 19892 44396 19944 44402
rect 19892 44338 19944 44344
rect 20076 44396 20128 44402
rect 20076 44338 20128 44344
rect 19800 41268 19852 41274
rect 19800 41210 19852 41216
rect 19904 41070 19932 44338
rect 20088 43110 20116 44338
rect 20168 43308 20220 43314
rect 20168 43250 20220 43256
rect 20076 43104 20128 43110
rect 20076 43046 20128 43052
rect 19984 41472 20036 41478
rect 19984 41414 20036 41420
rect 19892 41064 19944 41070
rect 19812 41024 19892 41052
rect 19708 40452 19760 40458
rect 19708 40394 19760 40400
rect 19616 38004 19668 38010
rect 19616 37946 19668 37952
rect 19340 37868 19392 37874
rect 19340 37810 19392 37816
rect 19064 37606 19116 37612
rect 19246 37632 19302 37641
rect 18970 37496 19026 37505
rect 19076 37482 19104 37606
rect 19246 37567 19302 37576
rect 19076 37466 19288 37482
rect 19352 37466 19380 37810
rect 19076 37460 19300 37466
rect 19076 37454 19248 37460
rect 18970 37431 19026 37440
rect 19248 37402 19300 37408
rect 19340 37460 19392 37466
rect 19340 37402 19392 37408
rect 19352 37369 19380 37402
rect 19062 37360 19118 37369
rect 19338 37360 19394 37369
rect 19062 37295 19118 37304
rect 19156 37324 19208 37330
rect 18972 37188 19024 37194
rect 18972 37130 19024 37136
rect 18984 34746 19012 37130
rect 18972 34740 19024 34746
rect 18972 34682 19024 34688
rect 18892 31726 19012 31754
rect 18800 30756 18920 30784
rect 18788 30660 18840 30666
rect 18788 30602 18840 30608
rect 18696 30388 18748 30394
rect 18696 30330 18748 30336
rect 18800 30326 18828 30602
rect 18788 30320 18840 30326
rect 18788 30262 18840 30268
rect 18696 30048 18748 30054
rect 18694 30016 18696 30025
rect 18748 30016 18750 30025
rect 18694 29951 18750 29960
rect 18892 28694 18920 30756
rect 18880 28688 18932 28694
rect 18880 28630 18932 28636
rect 18788 27940 18840 27946
rect 18788 27882 18840 27888
rect 18524 26846 18644 26874
rect 18420 25968 18472 25974
rect 18420 25910 18472 25916
rect 18420 25492 18472 25498
rect 18420 25434 18472 25440
rect 17950 25052 18258 25061
rect 17950 25050 17956 25052
rect 18012 25050 18036 25052
rect 18092 25050 18116 25052
rect 18172 25050 18196 25052
rect 18252 25050 18258 25052
rect 18012 24998 18014 25050
rect 18194 24998 18196 25050
rect 17950 24996 17956 24998
rect 18012 24996 18036 24998
rect 18092 24996 18116 24998
rect 18172 24996 18196 24998
rect 18252 24996 18258 24998
rect 17950 24987 18258 24996
rect 18328 24948 18380 24954
rect 18328 24890 18380 24896
rect 18052 24880 18104 24886
rect 18052 24822 18104 24828
rect 17960 24744 18012 24750
rect 17880 24704 17960 24732
rect 17880 24206 17908 24704
rect 17960 24686 18012 24692
rect 17972 24614 18000 24686
rect 17960 24608 18012 24614
rect 17960 24550 18012 24556
rect 17868 24200 17920 24206
rect 17868 24142 17920 24148
rect 18064 24070 18092 24822
rect 17868 24064 17920 24070
rect 17868 24006 17920 24012
rect 18052 24064 18104 24070
rect 18052 24006 18104 24012
rect 17880 23662 17908 24006
rect 17950 23964 18258 23973
rect 17950 23962 17956 23964
rect 18012 23962 18036 23964
rect 18092 23962 18116 23964
rect 18172 23962 18196 23964
rect 18252 23962 18258 23964
rect 18012 23910 18014 23962
rect 18194 23910 18196 23962
rect 17950 23908 17956 23910
rect 18012 23908 18036 23910
rect 18092 23908 18116 23910
rect 18172 23908 18196 23910
rect 18252 23908 18258 23910
rect 17950 23899 18258 23908
rect 18340 23730 18368 24890
rect 18328 23724 18380 23730
rect 18328 23666 18380 23672
rect 17868 23656 17920 23662
rect 17868 23598 17920 23604
rect 17880 23050 17908 23598
rect 17868 23044 17920 23050
rect 17868 22986 17920 22992
rect 17950 22876 18258 22885
rect 17950 22874 17956 22876
rect 18012 22874 18036 22876
rect 18092 22874 18116 22876
rect 18172 22874 18196 22876
rect 18252 22874 18258 22876
rect 18012 22822 18014 22874
rect 18194 22822 18196 22874
rect 17950 22820 17956 22822
rect 18012 22820 18036 22822
rect 18092 22820 18116 22822
rect 18172 22820 18196 22822
rect 18252 22820 18258 22822
rect 17950 22811 18258 22820
rect 18328 22704 18380 22710
rect 18328 22646 18380 22652
rect 17776 22092 17828 22098
rect 17776 22034 17828 22040
rect 17868 21888 17920 21894
rect 17788 21836 17868 21842
rect 17788 21830 17920 21836
rect 17788 21814 17908 21830
rect 17500 21684 17552 21690
rect 17500 21626 17552 21632
rect 17592 21684 17644 21690
rect 17592 21626 17644 21632
rect 17788 21536 17816 21814
rect 17950 21788 18258 21797
rect 17950 21786 17956 21788
rect 18012 21786 18036 21788
rect 18092 21786 18116 21788
rect 18172 21786 18196 21788
rect 18252 21786 18258 21788
rect 18012 21734 18014 21786
rect 18194 21734 18196 21786
rect 17950 21732 17956 21734
rect 18012 21732 18036 21734
rect 18092 21732 18116 21734
rect 18172 21732 18196 21734
rect 18252 21732 18258 21734
rect 17950 21723 18258 21732
rect 17868 21616 17920 21622
rect 17868 21558 17920 21564
rect 17696 21508 17816 21536
rect 17696 20942 17724 21508
rect 17880 21350 17908 21558
rect 18340 21486 18368 22646
rect 18052 21480 18104 21486
rect 18052 21422 18104 21428
rect 18328 21480 18380 21486
rect 18328 21422 18380 21428
rect 17776 21344 17828 21350
rect 17776 21286 17828 21292
rect 17868 21344 17920 21350
rect 17868 21286 17920 21292
rect 17788 21010 17816 21286
rect 18064 21010 18092 21422
rect 17776 21004 17828 21010
rect 17776 20946 17828 20952
rect 18052 21004 18104 21010
rect 18052 20946 18104 20952
rect 18432 20942 18460 25434
rect 18524 21978 18552 26846
rect 18604 26580 18656 26586
rect 18604 26522 18656 26528
rect 18696 26580 18748 26586
rect 18696 26522 18748 26528
rect 18616 25226 18644 26522
rect 18708 26314 18736 26522
rect 18696 26308 18748 26314
rect 18696 26250 18748 26256
rect 18604 25220 18656 25226
rect 18604 25162 18656 25168
rect 18696 24676 18748 24682
rect 18696 24618 18748 24624
rect 18604 23724 18656 23730
rect 18604 23666 18656 23672
rect 18616 22098 18644 23666
rect 18604 22092 18656 22098
rect 18604 22034 18656 22040
rect 18524 21950 18644 21978
rect 17684 20936 17736 20942
rect 17684 20878 17736 20884
rect 18420 20936 18472 20942
rect 18420 20878 18472 20884
rect 17950 20700 18258 20709
rect 17950 20698 17956 20700
rect 18012 20698 18036 20700
rect 18092 20698 18116 20700
rect 18172 20698 18196 20700
rect 18252 20698 18258 20700
rect 18012 20646 18014 20698
rect 18194 20646 18196 20698
rect 17950 20644 17956 20646
rect 18012 20644 18036 20646
rect 18092 20644 18116 20646
rect 18172 20644 18196 20646
rect 18252 20644 18258 20646
rect 17950 20635 18258 20644
rect 17868 20256 17920 20262
rect 17868 20198 17920 20204
rect 18052 20256 18104 20262
rect 18052 20198 18104 20204
rect 17500 19168 17552 19174
rect 17500 19110 17552 19116
rect 17408 18692 17460 18698
rect 17408 18634 17460 18640
rect 17408 15972 17460 15978
rect 17408 15914 17460 15920
rect 17420 15502 17448 15914
rect 17408 15496 17460 15502
rect 17408 15438 17460 15444
rect 17316 14408 17368 14414
rect 17316 14350 17368 14356
rect 17040 14340 17092 14346
rect 17040 14282 17092 14288
rect 17328 14006 17356 14350
rect 17316 14000 17368 14006
rect 17316 13942 17368 13948
rect 17040 13932 17092 13938
rect 17040 13874 17092 13880
rect 17052 13394 17080 13874
rect 17040 13388 17092 13394
rect 17040 13330 17092 13336
rect 17052 12782 17080 13330
rect 17040 12776 17092 12782
rect 17040 12718 17092 12724
rect 16960 12406 17080 12434
rect 16856 12096 16908 12102
rect 16856 12038 16908 12044
rect 16868 11558 16896 12038
rect 16856 11552 16908 11558
rect 16856 11494 16908 11500
rect 16684 11206 16804 11234
rect 16408 6886 16528 6914
rect 16500 4214 16528 6886
rect 16488 4208 16540 4214
rect 16488 4150 16540 4156
rect 16684 4146 16712 11206
rect 16764 11076 16816 11082
rect 16764 11018 16816 11024
rect 16672 4140 16724 4146
rect 16672 4082 16724 4088
rect 16396 4072 16448 4078
rect 16396 4014 16448 4020
rect 16304 3528 16356 3534
rect 16304 3470 16356 3476
rect 16408 800 16436 4014
rect 16776 3058 16804 11018
rect 16948 9920 17000 9926
rect 16948 9862 17000 9868
rect 16764 3052 16816 3058
rect 16764 2994 16816 3000
rect 16960 2446 16988 9862
rect 17052 8566 17080 12406
rect 17420 12102 17448 15438
rect 17512 14618 17540 19110
rect 17590 18728 17646 18737
rect 17590 18663 17646 18672
rect 17604 18630 17632 18663
rect 17592 18624 17644 18630
rect 17592 18566 17644 18572
rect 17592 16652 17644 16658
rect 17592 16594 17644 16600
rect 17500 14612 17552 14618
rect 17500 14554 17552 14560
rect 17500 14340 17552 14346
rect 17500 14282 17552 14288
rect 17512 13734 17540 14282
rect 17500 13728 17552 13734
rect 17500 13670 17552 13676
rect 17512 12646 17540 13670
rect 17500 12640 17552 12646
rect 17500 12582 17552 12588
rect 17604 12434 17632 16594
rect 17776 16584 17828 16590
rect 17776 16526 17828 16532
rect 17788 15910 17816 16526
rect 17776 15904 17828 15910
rect 17776 15846 17828 15852
rect 17684 14272 17736 14278
rect 17684 14214 17736 14220
rect 17512 12406 17632 12434
rect 17408 12096 17460 12102
rect 17408 12038 17460 12044
rect 17512 9654 17540 12406
rect 17592 12096 17644 12102
rect 17592 12038 17644 12044
rect 17604 11898 17632 12038
rect 17592 11892 17644 11898
rect 17592 11834 17644 11840
rect 17696 10554 17724 14214
rect 17776 13456 17828 13462
rect 17776 13398 17828 13404
rect 17788 11286 17816 13398
rect 17776 11280 17828 11286
rect 17776 11222 17828 11228
rect 17604 10526 17724 10554
rect 17500 9648 17552 9654
rect 17500 9590 17552 9596
rect 17408 9444 17460 9450
rect 17408 9386 17460 9392
rect 17040 8560 17092 8566
rect 17040 8502 17092 8508
rect 17132 2916 17184 2922
rect 17132 2858 17184 2864
rect 16948 2440 17000 2446
rect 16948 2382 17000 2388
rect 16764 2372 16816 2378
rect 16764 2314 16816 2320
rect 16776 800 16804 2314
rect 17144 800 17172 2858
rect 17420 2650 17448 9386
rect 17500 4072 17552 4078
rect 17500 4014 17552 4020
rect 17408 2644 17460 2650
rect 17408 2586 17460 2592
rect 17512 800 17540 4014
rect 17604 3534 17632 10526
rect 17684 7268 17736 7274
rect 17684 7210 17736 7216
rect 17696 4622 17724 7210
rect 17776 5228 17828 5234
rect 17776 5170 17828 5176
rect 17788 4758 17816 5170
rect 17776 4752 17828 4758
rect 17776 4694 17828 4700
rect 17684 4616 17736 4622
rect 17684 4558 17736 4564
rect 17776 3596 17828 3602
rect 17776 3538 17828 3544
rect 17592 3528 17644 3534
rect 17592 3470 17644 3476
rect 17788 1714 17816 3538
rect 17880 3058 17908 20198
rect 18064 20058 18092 20198
rect 18052 20052 18104 20058
rect 18052 19994 18104 20000
rect 18512 19712 18564 19718
rect 18512 19654 18564 19660
rect 17950 19612 18258 19621
rect 17950 19610 17956 19612
rect 18012 19610 18036 19612
rect 18092 19610 18116 19612
rect 18172 19610 18196 19612
rect 18252 19610 18258 19612
rect 18012 19558 18014 19610
rect 18194 19558 18196 19610
rect 17950 19556 17956 19558
rect 18012 19556 18036 19558
rect 18092 19556 18116 19558
rect 18172 19556 18196 19558
rect 18252 19556 18258 19558
rect 17950 19547 18258 19556
rect 18326 18728 18382 18737
rect 18326 18663 18382 18672
rect 17950 18524 18258 18533
rect 17950 18522 17956 18524
rect 18012 18522 18036 18524
rect 18092 18522 18116 18524
rect 18172 18522 18196 18524
rect 18252 18522 18258 18524
rect 18012 18470 18014 18522
rect 18194 18470 18196 18522
rect 17950 18468 17956 18470
rect 18012 18468 18036 18470
rect 18092 18468 18116 18470
rect 18172 18468 18196 18470
rect 18252 18468 18258 18470
rect 17950 18459 18258 18468
rect 18340 18426 18368 18663
rect 18328 18420 18380 18426
rect 18328 18362 18380 18368
rect 18144 18216 18196 18222
rect 18144 18158 18196 18164
rect 18156 17882 18184 18158
rect 18144 17876 18196 17882
rect 18144 17818 18196 17824
rect 17950 17436 18258 17445
rect 17950 17434 17956 17436
rect 18012 17434 18036 17436
rect 18092 17434 18116 17436
rect 18172 17434 18196 17436
rect 18252 17434 18258 17436
rect 18012 17382 18014 17434
rect 18194 17382 18196 17434
rect 17950 17380 17956 17382
rect 18012 17380 18036 17382
rect 18092 17380 18116 17382
rect 18172 17380 18196 17382
rect 18252 17380 18258 17382
rect 17950 17371 18258 17380
rect 18236 17196 18288 17202
rect 18236 17138 18288 17144
rect 18248 16658 18276 17138
rect 18236 16652 18288 16658
rect 18236 16594 18288 16600
rect 18328 16584 18380 16590
rect 18328 16526 18380 16532
rect 17950 16348 18258 16357
rect 17950 16346 17956 16348
rect 18012 16346 18036 16348
rect 18092 16346 18116 16348
rect 18172 16346 18196 16348
rect 18252 16346 18258 16348
rect 18012 16294 18014 16346
rect 18194 16294 18196 16346
rect 17950 16292 17956 16294
rect 18012 16292 18036 16294
rect 18092 16292 18116 16294
rect 18172 16292 18196 16294
rect 18252 16292 18258 16294
rect 17950 16283 18258 16292
rect 18236 15904 18288 15910
rect 18236 15846 18288 15852
rect 18248 15570 18276 15846
rect 18340 15706 18368 16526
rect 18420 16448 18472 16454
rect 18420 16390 18472 16396
rect 18432 15706 18460 16390
rect 18328 15700 18380 15706
rect 18328 15642 18380 15648
rect 18420 15700 18472 15706
rect 18420 15642 18472 15648
rect 18236 15564 18288 15570
rect 18236 15506 18288 15512
rect 18248 15366 18276 15506
rect 18236 15360 18288 15366
rect 18236 15302 18288 15308
rect 17950 15260 18258 15269
rect 17950 15258 17956 15260
rect 18012 15258 18036 15260
rect 18092 15258 18116 15260
rect 18172 15258 18196 15260
rect 18252 15258 18258 15260
rect 18012 15206 18014 15258
rect 18194 15206 18196 15258
rect 17950 15204 17956 15206
rect 18012 15204 18036 15206
rect 18092 15204 18116 15206
rect 18172 15204 18196 15206
rect 18252 15204 18258 15206
rect 17950 15195 18258 15204
rect 18340 15144 18368 15642
rect 18248 15116 18368 15144
rect 17960 15020 18012 15026
rect 17960 14962 18012 14968
rect 17972 14482 18000 14962
rect 18248 14958 18276 15116
rect 18236 14952 18288 14958
rect 18236 14894 18288 14900
rect 18328 14952 18380 14958
rect 18328 14894 18380 14900
rect 17960 14476 18012 14482
rect 17960 14418 18012 14424
rect 17950 14172 18258 14181
rect 17950 14170 17956 14172
rect 18012 14170 18036 14172
rect 18092 14170 18116 14172
rect 18172 14170 18196 14172
rect 18252 14170 18258 14172
rect 18012 14118 18014 14170
rect 18194 14118 18196 14170
rect 17950 14116 17956 14118
rect 18012 14116 18036 14118
rect 18092 14116 18116 14118
rect 18172 14116 18196 14118
rect 18252 14116 18258 14118
rect 17950 14107 18258 14116
rect 18144 13864 18196 13870
rect 18144 13806 18196 13812
rect 18156 13394 18184 13806
rect 18144 13388 18196 13394
rect 18144 13330 18196 13336
rect 17950 13084 18258 13093
rect 17950 13082 17956 13084
rect 18012 13082 18036 13084
rect 18092 13082 18116 13084
rect 18172 13082 18196 13084
rect 18252 13082 18258 13084
rect 18012 13030 18014 13082
rect 18194 13030 18196 13082
rect 17950 13028 17956 13030
rect 18012 13028 18036 13030
rect 18092 13028 18116 13030
rect 18172 13028 18196 13030
rect 18252 13028 18258 13030
rect 17950 13019 18258 13028
rect 18340 12986 18368 14894
rect 18418 14512 18474 14521
rect 18418 14447 18474 14456
rect 18432 14414 18460 14447
rect 18420 14408 18472 14414
rect 18420 14350 18472 14356
rect 18420 13252 18472 13258
rect 18420 13194 18472 13200
rect 18328 12980 18380 12986
rect 18328 12922 18380 12928
rect 17950 11996 18258 12005
rect 17950 11994 17956 11996
rect 18012 11994 18036 11996
rect 18092 11994 18116 11996
rect 18172 11994 18196 11996
rect 18252 11994 18258 11996
rect 18012 11942 18014 11994
rect 18194 11942 18196 11994
rect 17950 11940 17956 11942
rect 18012 11940 18036 11942
rect 18092 11940 18116 11942
rect 18172 11940 18196 11942
rect 18252 11940 18258 11942
rect 17950 11931 18258 11940
rect 18340 11830 18368 12922
rect 18432 12374 18460 13194
rect 18420 12368 18472 12374
rect 18420 12310 18472 12316
rect 18328 11824 18380 11830
rect 18328 11766 18380 11772
rect 18328 11552 18380 11558
rect 18328 11494 18380 11500
rect 17950 10908 18258 10917
rect 17950 10906 17956 10908
rect 18012 10906 18036 10908
rect 18092 10906 18116 10908
rect 18172 10906 18196 10908
rect 18252 10906 18258 10908
rect 18012 10854 18014 10906
rect 18194 10854 18196 10906
rect 17950 10852 17956 10854
rect 18012 10852 18036 10854
rect 18092 10852 18116 10854
rect 18172 10852 18196 10854
rect 18252 10852 18258 10854
rect 17950 10843 18258 10852
rect 18340 10674 18368 11494
rect 18328 10668 18380 10674
rect 18328 10610 18380 10616
rect 18524 10062 18552 19654
rect 18616 18766 18644 21950
rect 18708 19378 18736 24618
rect 18800 23730 18828 27882
rect 18892 27130 18920 28630
rect 18880 27124 18932 27130
rect 18880 27066 18932 27072
rect 18880 25832 18932 25838
rect 18880 25774 18932 25780
rect 18788 23724 18840 23730
rect 18788 23666 18840 23672
rect 18892 23322 18920 25774
rect 18880 23316 18932 23322
rect 18880 23258 18932 23264
rect 18892 22642 18920 23258
rect 18880 22636 18932 22642
rect 18880 22578 18932 22584
rect 18892 21010 18920 22578
rect 18880 21004 18932 21010
rect 18880 20946 18932 20952
rect 18984 20058 19012 31726
rect 19076 20602 19104 37295
rect 19338 37295 19394 37304
rect 19156 37266 19208 37272
rect 19168 36854 19196 37266
rect 19294 37256 19346 37262
rect 19294 37198 19346 37204
rect 19306 37074 19334 37198
rect 19260 37046 19334 37074
rect 19156 36848 19208 36854
rect 19156 36790 19208 36796
rect 19260 36786 19288 37046
rect 19248 36780 19300 36786
rect 19248 36722 19300 36728
rect 19616 36780 19668 36786
rect 19616 36722 19668 36728
rect 19154 36680 19210 36689
rect 19154 36615 19210 36624
rect 19168 28762 19196 36615
rect 19628 36582 19656 36722
rect 19616 36576 19668 36582
rect 19616 36518 19668 36524
rect 19628 36145 19656 36518
rect 19614 36136 19670 36145
rect 19614 36071 19670 36080
rect 19524 35488 19576 35494
rect 19524 35430 19576 35436
rect 19248 35216 19300 35222
rect 19248 35158 19300 35164
rect 19260 32450 19288 35158
rect 19536 34678 19564 35430
rect 19524 34672 19576 34678
rect 19524 34614 19576 34620
rect 19720 32570 19748 40394
rect 19812 36718 19840 41024
rect 19892 41006 19944 41012
rect 19996 40186 20024 41414
rect 19984 40180 20036 40186
rect 19984 40122 20036 40128
rect 20088 39982 20116 43046
rect 20180 42634 20208 43250
rect 20168 42628 20220 42634
rect 20168 42570 20220 42576
rect 20168 41676 20220 41682
rect 20168 41618 20220 41624
rect 20180 40497 20208 41618
rect 20272 41614 20300 45222
rect 20364 45082 20392 46446
rect 20916 45558 20944 53382
rect 21008 53242 21036 53518
rect 20996 53236 21048 53242
rect 20996 53178 21048 53184
rect 20904 45552 20956 45558
rect 20904 45494 20956 45500
rect 20352 45076 20404 45082
rect 20352 45018 20404 45024
rect 20812 44192 20864 44198
rect 20812 44134 20864 44140
rect 20628 43784 20680 43790
rect 20628 43726 20680 43732
rect 20536 43648 20588 43654
rect 20536 43590 20588 43596
rect 20548 43314 20576 43590
rect 20536 43308 20588 43314
rect 20536 43250 20588 43256
rect 20640 42566 20668 43726
rect 20628 42560 20680 42566
rect 20628 42502 20680 42508
rect 20534 42120 20590 42129
rect 20534 42055 20590 42064
rect 20352 41744 20404 41750
rect 20352 41686 20404 41692
rect 20260 41608 20312 41614
rect 20260 41550 20312 41556
rect 20166 40488 20222 40497
rect 20166 40423 20222 40432
rect 20076 39976 20128 39982
rect 20076 39918 20128 39924
rect 19984 39364 20036 39370
rect 19984 39306 20036 39312
rect 19892 39024 19944 39030
rect 19892 38966 19944 38972
rect 19800 36712 19852 36718
rect 19800 36654 19852 36660
rect 19798 33552 19854 33561
rect 19798 33487 19854 33496
rect 19812 33454 19840 33487
rect 19800 33448 19852 33454
rect 19800 33390 19852 33396
rect 19432 32564 19484 32570
rect 19432 32506 19484 32512
rect 19708 32564 19760 32570
rect 19708 32506 19760 32512
rect 19260 32422 19380 32450
rect 19352 32366 19380 32422
rect 19248 32360 19300 32366
rect 19248 32302 19300 32308
rect 19340 32360 19392 32366
rect 19340 32302 19392 32308
rect 19260 32026 19288 32302
rect 19248 32020 19300 32026
rect 19248 31962 19300 31968
rect 19156 28756 19208 28762
rect 19156 28698 19208 28704
rect 19156 28008 19208 28014
rect 19156 27950 19208 27956
rect 19168 27674 19196 27950
rect 19260 27878 19288 31962
rect 19444 31890 19472 32506
rect 19800 32496 19852 32502
rect 19800 32438 19852 32444
rect 19524 32224 19576 32230
rect 19524 32166 19576 32172
rect 19432 31884 19484 31890
rect 19432 31826 19484 31832
rect 19536 31754 19564 32166
rect 19616 31952 19668 31958
rect 19616 31894 19668 31900
rect 19352 31726 19564 31754
rect 19248 27872 19300 27878
rect 19248 27814 19300 27820
rect 19156 27668 19208 27674
rect 19156 27610 19208 27616
rect 19352 27402 19380 31726
rect 19524 31136 19576 31142
rect 19524 31078 19576 31084
rect 19432 30388 19484 30394
rect 19432 30330 19484 30336
rect 19340 27396 19392 27402
rect 19340 27338 19392 27344
rect 19444 26994 19472 30330
rect 19432 26988 19484 26994
rect 19432 26930 19484 26936
rect 19156 26376 19208 26382
rect 19156 26318 19208 26324
rect 19168 25906 19196 26318
rect 19432 26240 19484 26246
rect 19432 26182 19484 26188
rect 19156 25900 19208 25906
rect 19156 25842 19208 25848
rect 19248 25696 19300 25702
rect 19248 25638 19300 25644
rect 19156 24200 19208 24206
rect 19156 24142 19208 24148
rect 19168 23798 19196 24142
rect 19156 23792 19208 23798
rect 19156 23734 19208 23740
rect 19156 23520 19208 23526
rect 19156 23462 19208 23468
rect 19168 21622 19196 23462
rect 19156 21616 19208 21622
rect 19156 21558 19208 21564
rect 19156 21072 19208 21078
rect 19156 21014 19208 21020
rect 19064 20596 19116 20602
rect 19064 20538 19116 20544
rect 19168 20466 19196 21014
rect 19260 20602 19288 25638
rect 19444 24954 19472 26182
rect 19432 24948 19484 24954
rect 19432 24890 19484 24896
rect 19340 23180 19392 23186
rect 19340 23122 19392 23128
rect 19352 22098 19380 23122
rect 19340 22092 19392 22098
rect 19340 22034 19392 22040
rect 19248 20596 19300 20602
rect 19248 20538 19300 20544
rect 19156 20460 19208 20466
rect 19156 20402 19208 20408
rect 18972 20052 19024 20058
rect 18972 19994 19024 20000
rect 18984 19922 19012 19994
rect 19064 19984 19116 19990
rect 19064 19926 19116 19932
rect 18972 19916 19024 19922
rect 18972 19858 19024 19864
rect 18696 19372 18748 19378
rect 18696 19314 18748 19320
rect 18604 18760 18656 18766
rect 18604 18702 18656 18708
rect 18878 18728 18934 18737
rect 18878 18663 18934 18672
rect 18972 18692 19024 18698
rect 18696 18080 18748 18086
rect 18696 18022 18748 18028
rect 18708 17610 18736 18022
rect 18696 17604 18748 17610
rect 18696 17546 18748 17552
rect 18604 17128 18656 17134
rect 18604 17070 18656 17076
rect 18616 16590 18644 17070
rect 18604 16584 18656 16590
rect 18604 16526 18656 16532
rect 18708 14958 18736 17546
rect 18788 16720 18840 16726
rect 18788 16662 18840 16668
rect 18800 16250 18828 16662
rect 18788 16244 18840 16250
rect 18788 16186 18840 16192
rect 18892 15688 18920 18663
rect 18972 18634 19024 18640
rect 18800 15660 18920 15688
rect 18696 14952 18748 14958
rect 18696 14894 18748 14900
rect 18800 14770 18828 15660
rect 18880 15564 18932 15570
rect 18880 15506 18932 15512
rect 18616 14742 18828 14770
rect 18616 11218 18644 14742
rect 18788 14340 18840 14346
rect 18788 14282 18840 14288
rect 18696 13388 18748 13394
rect 18696 13330 18748 13336
rect 18708 12238 18736 13330
rect 18696 12232 18748 12238
rect 18696 12174 18748 12180
rect 18604 11212 18656 11218
rect 18604 11154 18656 11160
rect 18696 11076 18748 11082
rect 18696 11018 18748 11024
rect 18512 10056 18564 10062
rect 18512 9998 18564 10004
rect 17950 9820 18258 9829
rect 17950 9818 17956 9820
rect 18012 9818 18036 9820
rect 18092 9818 18116 9820
rect 18172 9818 18196 9820
rect 18252 9818 18258 9820
rect 18012 9766 18014 9818
rect 18194 9766 18196 9818
rect 17950 9764 17956 9766
rect 18012 9764 18036 9766
rect 18092 9764 18116 9766
rect 18172 9764 18196 9766
rect 18252 9764 18258 9766
rect 17950 9755 18258 9764
rect 17950 8732 18258 8741
rect 17950 8730 17956 8732
rect 18012 8730 18036 8732
rect 18092 8730 18116 8732
rect 18172 8730 18196 8732
rect 18252 8730 18258 8732
rect 18012 8678 18014 8730
rect 18194 8678 18196 8730
rect 17950 8676 17956 8678
rect 18012 8676 18036 8678
rect 18092 8676 18116 8678
rect 18172 8676 18196 8678
rect 18252 8676 18258 8678
rect 17950 8667 18258 8676
rect 17950 7644 18258 7653
rect 17950 7642 17956 7644
rect 18012 7642 18036 7644
rect 18092 7642 18116 7644
rect 18172 7642 18196 7644
rect 18252 7642 18258 7644
rect 18012 7590 18014 7642
rect 18194 7590 18196 7642
rect 17950 7588 17956 7590
rect 18012 7588 18036 7590
rect 18092 7588 18116 7590
rect 18172 7588 18196 7590
rect 18252 7588 18258 7590
rect 17950 7579 18258 7588
rect 17950 6556 18258 6565
rect 17950 6554 17956 6556
rect 18012 6554 18036 6556
rect 18092 6554 18116 6556
rect 18172 6554 18196 6556
rect 18252 6554 18258 6556
rect 18012 6502 18014 6554
rect 18194 6502 18196 6554
rect 17950 6500 17956 6502
rect 18012 6500 18036 6502
rect 18092 6500 18116 6502
rect 18172 6500 18196 6502
rect 18252 6500 18258 6502
rect 17950 6491 18258 6500
rect 17950 5468 18258 5477
rect 17950 5466 17956 5468
rect 18012 5466 18036 5468
rect 18092 5466 18116 5468
rect 18172 5466 18196 5468
rect 18252 5466 18258 5468
rect 18012 5414 18014 5466
rect 18194 5414 18196 5466
rect 17950 5412 17956 5414
rect 18012 5412 18036 5414
rect 18092 5412 18116 5414
rect 18172 5412 18196 5414
rect 18252 5412 18258 5414
rect 17950 5403 18258 5412
rect 18708 4622 18736 11018
rect 18800 10606 18828 14282
rect 18892 13938 18920 15506
rect 18880 13932 18932 13938
rect 18880 13874 18932 13880
rect 18892 12986 18920 13874
rect 18880 12980 18932 12986
rect 18880 12922 18932 12928
rect 18880 12096 18932 12102
rect 18880 12038 18932 12044
rect 18892 11694 18920 12038
rect 18880 11688 18932 11694
rect 18880 11630 18932 11636
rect 18788 10600 18840 10606
rect 18788 10542 18840 10548
rect 18984 6914 19012 18634
rect 19076 13954 19104 19926
rect 19536 19854 19564 31078
rect 19628 26042 19656 31894
rect 19812 31482 19840 32438
rect 19800 31476 19852 31482
rect 19800 31418 19852 31424
rect 19708 31408 19760 31414
rect 19708 31350 19760 31356
rect 19720 30734 19748 31350
rect 19800 30932 19852 30938
rect 19800 30874 19852 30880
rect 19708 30728 19760 30734
rect 19708 30670 19760 30676
rect 19812 30258 19840 30874
rect 19904 30682 19932 38966
rect 19996 36650 20024 39306
rect 20076 39296 20128 39302
rect 20076 39238 20128 39244
rect 19984 36644 20036 36650
rect 19984 36586 20036 36592
rect 20088 36417 20116 39238
rect 20168 38276 20220 38282
rect 20168 38218 20220 38224
rect 20074 36408 20130 36417
rect 20074 36343 20130 36352
rect 19984 36032 20036 36038
rect 19984 35974 20036 35980
rect 19996 31482 20024 35974
rect 20180 35154 20208 38218
rect 20260 37664 20312 37670
rect 20260 37606 20312 37612
rect 20168 35148 20220 35154
rect 20168 35090 20220 35096
rect 20076 34604 20128 34610
rect 20076 34546 20128 34552
rect 20088 33454 20116 34546
rect 20168 33856 20220 33862
rect 20168 33798 20220 33804
rect 20180 33590 20208 33798
rect 20168 33584 20220 33590
rect 20168 33526 20220 33532
rect 20076 33448 20128 33454
rect 20076 33390 20128 33396
rect 19984 31476 20036 31482
rect 19984 31418 20036 31424
rect 20088 31278 20116 33390
rect 20168 33380 20220 33386
rect 20168 33322 20220 33328
rect 20180 31822 20208 33322
rect 20272 32570 20300 37606
rect 20364 35834 20392 41686
rect 20444 40928 20496 40934
rect 20444 40870 20496 40876
rect 20456 39438 20484 40870
rect 20548 40458 20576 42055
rect 20640 41682 20668 42502
rect 20628 41676 20680 41682
rect 20628 41618 20680 41624
rect 20628 41540 20680 41546
rect 20628 41482 20680 41488
rect 20720 41540 20772 41546
rect 20720 41482 20772 41488
rect 20640 40526 20668 41482
rect 20628 40520 20680 40526
rect 20628 40462 20680 40468
rect 20536 40452 20588 40458
rect 20536 40394 20588 40400
rect 20444 39432 20496 39438
rect 20444 39374 20496 39380
rect 20628 39432 20680 39438
rect 20628 39374 20680 39380
rect 20536 38820 20588 38826
rect 20536 38762 20588 38768
rect 20444 37868 20496 37874
rect 20444 37810 20496 37816
rect 20456 36786 20484 37810
rect 20548 37262 20576 38762
rect 20536 37256 20588 37262
rect 20536 37198 20588 37204
rect 20640 36922 20668 39374
rect 20732 37738 20760 41482
rect 20720 37732 20772 37738
rect 20720 37674 20772 37680
rect 20628 36916 20680 36922
rect 20628 36858 20680 36864
rect 20444 36780 20496 36786
rect 20444 36722 20496 36728
rect 20444 36576 20496 36582
rect 20444 36518 20496 36524
rect 20352 35828 20404 35834
rect 20352 35770 20404 35776
rect 20456 33946 20484 36518
rect 20720 35488 20772 35494
rect 20720 35430 20772 35436
rect 20628 34400 20680 34406
rect 20628 34342 20680 34348
rect 20364 33918 20484 33946
rect 20536 33924 20588 33930
rect 20260 32564 20312 32570
rect 20260 32506 20312 32512
rect 20364 32502 20392 33918
rect 20536 33866 20588 33872
rect 20444 33856 20496 33862
rect 20444 33798 20496 33804
rect 20456 33658 20484 33798
rect 20548 33658 20576 33866
rect 20444 33652 20496 33658
rect 20444 33594 20496 33600
rect 20536 33652 20588 33658
rect 20536 33594 20588 33600
rect 20352 32496 20404 32502
rect 20352 32438 20404 32444
rect 20444 32360 20496 32366
rect 20444 32302 20496 32308
rect 20352 31884 20404 31890
rect 20352 31826 20404 31832
rect 20168 31816 20220 31822
rect 20168 31758 20220 31764
rect 20260 31680 20312 31686
rect 20260 31622 20312 31628
rect 20168 31476 20220 31482
rect 20168 31418 20220 31424
rect 20076 31272 20128 31278
rect 20076 31214 20128 31220
rect 20180 30802 20208 31418
rect 20168 30796 20220 30802
rect 20168 30738 20220 30744
rect 19904 30654 20116 30682
rect 19892 30592 19944 30598
rect 19890 30560 19892 30569
rect 19944 30560 19946 30569
rect 19890 30495 19946 30504
rect 19892 30388 19944 30394
rect 19892 30330 19944 30336
rect 19800 30252 19852 30258
rect 19800 30194 19852 30200
rect 19800 30116 19852 30122
rect 19800 30058 19852 30064
rect 19812 30025 19840 30058
rect 19798 30016 19854 30025
rect 19798 29951 19854 29960
rect 19904 29782 19932 30330
rect 20088 29782 20116 30654
rect 20168 30660 20220 30666
rect 20168 30602 20220 30608
rect 20180 30122 20208 30602
rect 20168 30116 20220 30122
rect 20168 30058 20220 30064
rect 19892 29776 19944 29782
rect 19892 29718 19944 29724
rect 20076 29776 20128 29782
rect 20076 29718 20128 29724
rect 19800 29504 19852 29510
rect 19852 29464 19932 29492
rect 19800 29446 19852 29452
rect 19800 29164 19852 29170
rect 19800 29106 19852 29112
rect 19812 29073 19840 29106
rect 19798 29064 19854 29073
rect 19798 28999 19854 29008
rect 19800 28008 19852 28014
rect 19800 27950 19852 27956
rect 19708 27328 19760 27334
rect 19708 27270 19760 27276
rect 19720 26042 19748 27270
rect 19812 27062 19840 27950
rect 19800 27056 19852 27062
rect 19800 26998 19852 27004
rect 19800 26920 19852 26926
rect 19800 26862 19852 26868
rect 19812 26382 19840 26862
rect 19800 26376 19852 26382
rect 19800 26318 19852 26324
rect 19800 26240 19852 26246
rect 19800 26182 19852 26188
rect 19616 26036 19668 26042
rect 19616 25978 19668 25984
rect 19708 26036 19760 26042
rect 19708 25978 19760 25984
rect 19616 25900 19668 25906
rect 19616 25842 19668 25848
rect 19524 19848 19576 19854
rect 19524 19790 19576 19796
rect 19248 19168 19300 19174
rect 19248 19110 19300 19116
rect 19156 18692 19208 18698
rect 19156 18634 19208 18640
rect 19168 16250 19196 18634
rect 19156 16244 19208 16250
rect 19156 16186 19208 16192
rect 19156 14952 19208 14958
rect 19156 14894 19208 14900
rect 19168 14074 19196 14894
rect 19156 14068 19208 14074
rect 19156 14010 19208 14016
rect 19076 13926 19196 13954
rect 19064 13864 19116 13870
rect 19064 13806 19116 13812
rect 19076 9654 19104 13806
rect 19168 11778 19196 13926
rect 19260 13870 19288 19110
rect 19524 18624 19576 18630
rect 19524 18566 19576 18572
rect 19432 17196 19484 17202
rect 19432 17138 19484 17144
rect 19444 16794 19472 17138
rect 19536 17082 19564 18566
rect 19628 17270 19656 25842
rect 19708 25288 19760 25294
rect 19708 25230 19760 25236
rect 19720 23662 19748 25230
rect 19708 23656 19760 23662
rect 19708 23598 19760 23604
rect 19720 23186 19748 23598
rect 19708 23180 19760 23186
rect 19708 23122 19760 23128
rect 19812 21146 19840 26182
rect 19904 24818 19932 29464
rect 20088 29306 20116 29718
rect 20272 29578 20300 31622
rect 20260 29572 20312 29578
rect 20260 29514 20312 29520
rect 20076 29300 20128 29306
rect 20076 29242 20128 29248
rect 20260 29096 20312 29102
rect 20180 29056 20260 29084
rect 19984 27532 20036 27538
rect 19984 27474 20036 27480
rect 19892 24812 19944 24818
rect 19892 24754 19944 24760
rect 19892 24132 19944 24138
rect 19892 24074 19944 24080
rect 19904 23866 19932 24074
rect 19892 23860 19944 23866
rect 19892 23802 19944 23808
rect 19996 23798 20024 27474
rect 19984 23792 20036 23798
rect 19984 23734 20036 23740
rect 19996 23338 20024 23734
rect 19996 23322 20116 23338
rect 19996 23316 20128 23322
rect 19996 23310 20076 23316
rect 20076 23258 20128 23264
rect 20180 23202 20208 29056
rect 20260 29038 20312 29044
rect 20364 27538 20392 31826
rect 20456 31686 20484 32302
rect 20444 31680 20496 31686
rect 20444 31622 20496 31628
rect 20444 31340 20496 31346
rect 20444 31282 20496 31288
rect 20352 27532 20404 27538
rect 20352 27474 20404 27480
rect 20456 27418 20484 31282
rect 20640 29646 20668 34342
rect 20732 33998 20760 35430
rect 20720 33992 20772 33998
rect 20720 33934 20772 33940
rect 20732 32978 20760 33934
rect 20720 32972 20772 32978
rect 20720 32914 20772 32920
rect 20720 32292 20772 32298
rect 20720 32234 20772 32240
rect 20732 32026 20760 32234
rect 20720 32020 20772 32026
rect 20720 31962 20772 31968
rect 20720 30864 20772 30870
rect 20720 30806 20772 30812
rect 20628 29640 20680 29646
rect 20628 29582 20680 29588
rect 20732 29238 20760 30806
rect 20720 29232 20772 29238
rect 20720 29174 20772 29180
rect 20824 29170 20852 44134
rect 20904 43648 20956 43654
rect 20904 43590 20956 43596
rect 20916 42634 20944 43590
rect 21100 43217 21128 53926
rect 21744 53582 21772 56200
rect 21916 53712 21968 53718
rect 21916 53654 21968 53660
rect 21732 53576 21784 53582
rect 21732 53518 21784 53524
rect 21744 53242 21772 53518
rect 21732 53236 21784 53242
rect 21732 53178 21784 53184
rect 21456 50448 21508 50454
rect 21456 50390 21508 50396
rect 21180 46912 21232 46918
rect 21180 46854 21232 46860
rect 21192 46034 21220 46854
rect 21180 46028 21232 46034
rect 21180 45970 21232 45976
rect 21272 45416 21324 45422
rect 21272 45358 21324 45364
rect 21284 43790 21312 45358
rect 21180 43784 21232 43790
rect 21180 43726 21232 43732
rect 21272 43784 21324 43790
rect 21272 43726 21324 43732
rect 21086 43208 21142 43217
rect 21086 43143 21142 43152
rect 20904 42628 20956 42634
rect 20904 42570 20956 42576
rect 20916 42294 20944 42570
rect 20904 42288 20956 42294
rect 20904 42230 20956 42236
rect 20916 42022 20944 42230
rect 21192 42090 21220 43726
rect 21180 42084 21232 42090
rect 21180 42026 21232 42032
rect 20904 42016 20956 42022
rect 20904 41958 20956 41964
rect 20904 41268 20956 41274
rect 20904 41210 20956 41216
rect 20916 41138 20944 41210
rect 20904 41132 20956 41138
rect 20904 41074 20956 41080
rect 20916 38978 20944 41074
rect 20996 41064 21048 41070
rect 20996 41006 21048 41012
rect 21008 39098 21036 41006
rect 21088 39568 21140 39574
rect 21088 39510 21140 39516
rect 21100 39098 21128 39510
rect 20996 39092 21048 39098
rect 20996 39034 21048 39040
rect 21088 39092 21140 39098
rect 21088 39034 21140 39040
rect 20916 38950 21036 38978
rect 20904 37460 20956 37466
rect 20904 37402 20956 37408
rect 20916 37262 20944 37402
rect 20904 37256 20956 37262
rect 20904 37198 20956 37204
rect 21008 36038 21036 38950
rect 21192 37806 21220 42026
rect 21284 39982 21312 43726
rect 21468 41002 21496 50390
rect 21640 49836 21692 49842
rect 21640 49778 21692 49784
rect 21548 44940 21600 44946
rect 21548 44882 21600 44888
rect 21560 43994 21588 44882
rect 21548 43988 21600 43994
rect 21548 43930 21600 43936
rect 21652 43926 21680 49778
rect 21824 46028 21876 46034
rect 21824 45970 21876 45976
rect 21732 45824 21784 45830
rect 21732 45766 21784 45772
rect 21744 45626 21772 45766
rect 21732 45620 21784 45626
rect 21732 45562 21784 45568
rect 21744 45286 21772 45562
rect 21732 45280 21784 45286
rect 21732 45222 21784 45228
rect 21744 45082 21772 45222
rect 21732 45076 21784 45082
rect 21732 45018 21784 45024
rect 21744 44810 21772 45018
rect 21732 44804 21784 44810
rect 21732 44746 21784 44752
rect 21640 43920 21692 43926
rect 21640 43862 21692 43868
rect 21548 42560 21600 42566
rect 21548 42502 21600 42508
rect 21456 40996 21508 41002
rect 21456 40938 21508 40944
rect 21560 40594 21588 42502
rect 21652 41188 21680 43862
rect 21836 42650 21864 45970
rect 21928 44198 21956 53654
rect 22112 53582 22140 56200
rect 22480 54194 22508 56200
rect 22468 54188 22520 54194
rect 22468 54130 22520 54136
rect 22480 54074 22508 54130
rect 22284 54052 22336 54058
rect 22480 54046 22600 54074
rect 22284 53994 22336 54000
rect 22192 53984 22244 53990
rect 22192 53926 22244 53932
rect 22100 53576 22152 53582
rect 22100 53518 22152 53524
rect 22112 53242 22140 53518
rect 22100 53236 22152 53242
rect 22100 53178 22152 53184
rect 22204 46170 22232 53926
rect 22192 46164 22244 46170
rect 22192 46106 22244 46112
rect 22204 45966 22232 46106
rect 22192 45960 22244 45966
rect 22006 45928 22062 45937
rect 22062 45908 22192 45914
rect 22062 45902 22244 45908
rect 22062 45886 22232 45902
rect 22006 45863 22062 45872
rect 22296 45642 22324 53994
rect 22376 53984 22428 53990
rect 22374 53952 22376 53961
rect 22428 53952 22430 53961
rect 22374 53887 22430 53896
rect 22376 53712 22428 53718
rect 22376 53654 22428 53660
rect 22204 45614 22324 45642
rect 22204 45506 22232 45614
rect 22020 45478 22232 45506
rect 22284 45552 22336 45558
rect 22284 45494 22336 45500
rect 21916 44192 21968 44198
rect 21916 44134 21968 44140
rect 21928 43722 21956 44134
rect 21916 43716 21968 43722
rect 21916 43658 21968 43664
rect 21916 43308 21968 43314
rect 21916 43250 21968 43256
rect 21928 43217 21956 43250
rect 21914 43208 21970 43217
rect 21914 43143 21970 43152
rect 22020 43058 22048 45478
rect 22296 44878 22324 45494
rect 22284 44872 22336 44878
rect 22284 44814 22336 44820
rect 22296 44742 22324 44814
rect 22284 44736 22336 44742
rect 22284 44678 22336 44684
rect 22296 44334 22324 44678
rect 22284 44328 22336 44334
rect 22284 44270 22336 44276
rect 22192 43648 22244 43654
rect 22192 43590 22244 43596
rect 22020 43030 22140 43058
rect 22006 42800 22062 42809
rect 22006 42735 22008 42744
rect 22060 42735 22062 42744
rect 22008 42706 22060 42712
rect 21836 42622 21956 42650
rect 21732 41472 21784 41478
rect 21732 41414 21784 41420
rect 21744 41256 21772 41414
rect 21824 41268 21876 41274
rect 21744 41228 21824 41256
rect 21824 41210 21876 41216
rect 21652 41160 21772 41188
rect 21744 41052 21772 41160
rect 21652 41024 21772 41052
rect 21456 40588 21508 40594
rect 21456 40530 21508 40536
rect 21548 40588 21600 40594
rect 21548 40530 21600 40536
rect 21364 40384 21416 40390
rect 21364 40326 21416 40332
rect 21272 39976 21324 39982
rect 21272 39918 21324 39924
rect 21376 39370 21404 40326
rect 21364 39364 21416 39370
rect 21364 39306 21416 39312
rect 21272 38888 21324 38894
rect 21272 38830 21324 38836
rect 21180 37800 21232 37806
rect 21180 37742 21232 37748
rect 21088 36780 21140 36786
rect 21088 36722 21140 36728
rect 21100 36582 21128 36722
rect 21088 36576 21140 36582
rect 21086 36544 21088 36553
rect 21140 36544 21142 36553
rect 21086 36479 21142 36488
rect 21284 36258 21312 38830
rect 21364 38752 21416 38758
rect 21364 38694 21416 38700
rect 21100 36230 21312 36258
rect 21376 36242 21404 38694
rect 21468 37874 21496 40530
rect 21548 38548 21600 38554
rect 21548 38490 21600 38496
rect 21560 38418 21588 38490
rect 21548 38412 21600 38418
rect 21548 38354 21600 38360
rect 21456 37868 21508 37874
rect 21456 37810 21508 37816
rect 21454 36408 21510 36417
rect 21454 36343 21510 36352
rect 21364 36236 21416 36242
rect 20996 36032 21048 36038
rect 20996 35974 21048 35980
rect 20996 35488 21048 35494
rect 20996 35430 21048 35436
rect 21008 35290 21036 35430
rect 20996 35284 21048 35290
rect 20996 35226 21048 35232
rect 21008 35018 21036 35226
rect 20996 35012 21048 35018
rect 20996 34954 21048 34960
rect 20904 34536 20956 34542
rect 20904 34478 20956 34484
rect 20916 33658 20944 34478
rect 21008 34134 21036 34954
rect 21100 34950 21128 36230
rect 21364 36178 21416 36184
rect 21272 36168 21324 36174
rect 21272 36110 21324 36116
rect 21180 36100 21232 36106
rect 21180 36042 21232 36048
rect 21088 34944 21140 34950
rect 21088 34886 21140 34892
rect 21088 34400 21140 34406
rect 21088 34342 21140 34348
rect 20996 34128 21048 34134
rect 20996 34070 21048 34076
rect 20904 33652 20956 33658
rect 20904 33594 20956 33600
rect 21008 33386 21036 34070
rect 20996 33380 21048 33386
rect 20996 33322 21048 33328
rect 20904 32768 20956 32774
rect 20904 32710 20956 32716
rect 20916 31890 20944 32710
rect 20996 32224 21048 32230
rect 20996 32166 21048 32172
rect 20904 31884 20956 31890
rect 20904 31826 20956 31832
rect 21008 31754 21036 32166
rect 20996 31748 21048 31754
rect 20996 31690 21048 31696
rect 21100 31498 21128 34342
rect 20916 31470 21128 31498
rect 20916 30190 20944 31470
rect 21192 30569 21220 36042
rect 21284 34950 21312 36110
rect 21272 34944 21324 34950
rect 21272 34886 21324 34892
rect 21284 34066 21312 34886
rect 21272 34060 21324 34066
rect 21272 34002 21324 34008
rect 21284 33522 21312 34002
rect 21468 33590 21496 36343
rect 21560 34678 21588 38354
rect 21652 37466 21680 41024
rect 21928 40934 21956 42622
rect 22008 42560 22060 42566
rect 22008 42502 22060 42508
rect 22020 42362 22048 42502
rect 22008 42356 22060 42362
rect 22008 42298 22060 42304
rect 22112 42242 22140 43030
rect 22204 42673 22232 43590
rect 22296 43382 22324 44270
rect 22388 43450 22416 53654
rect 22468 53440 22520 53446
rect 22468 53382 22520 53388
rect 22480 46714 22508 53382
rect 22572 53242 22600 54046
rect 22848 53582 22876 56200
rect 23216 55214 23244 56200
rect 23584 55214 23612 56200
rect 24490 56199 24546 56208
rect 23216 55186 23336 55214
rect 23584 55186 23704 55214
rect 22950 53884 23258 53893
rect 22950 53882 22956 53884
rect 23012 53882 23036 53884
rect 23092 53882 23116 53884
rect 23172 53882 23196 53884
rect 23252 53882 23258 53884
rect 23012 53830 23014 53882
rect 23194 53830 23196 53882
rect 22950 53828 22956 53830
rect 23012 53828 23036 53830
rect 23092 53828 23116 53830
rect 23172 53828 23196 53830
rect 23252 53828 23258 53830
rect 22950 53819 23258 53828
rect 22836 53576 22888 53582
rect 22836 53518 22888 53524
rect 23308 53242 23336 55186
rect 23572 53984 23624 53990
rect 23572 53926 23624 53932
rect 22560 53236 22612 53242
rect 22560 53178 22612 53184
rect 23296 53236 23348 53242
rect 23296 53178 23348 53184
rect 22560 52896 22612 52902
rect 22560 52838 22612 52844
rect 22468 46708 22520 46714
rect 22468 46650 22520 46656
rect 22468 46504 22520 46510
rect 22468 46446 22520 46452
rect 22376 43444 22428 43450
rect 22376 43386 22428 43392
rect 22284 43376 22336 43382
rect 22284 43318 22336 43324
rect 22376 42832 22428 42838
rect 22376 42774 22428 42780
rect 22190 42664 22246 42673
rect 22190 42599 22246 42608
rect 22282 42392 22338 42401
rect 22192 42356 22244 42362
rect 22282 42327 22338 42336
rect 22192 42298 22244 42304
rect 22020 42214 22140 42242
rect 21732 40928 21784 40934
rect 21732 40870 21784 40876
rect 21916 40928 21968 40934
rect 21916 40870 21968 40876
rect 21744 39574 21772 40870
rect 22020 40746 22048 42214
rect 22100 42084 22152 42090
rect 22100 42026 22152 42032
rect 22112 41585 22140 42026
rect 22098 41576 22154 41585
rect 22098 41511 22154 41520
rect 22098 41304 22154 41313
rect 22098 41239 22154 41248
rect 22112 41138 22140 41239
rect 22100 41132 22152 41138
rect 22100 41074 22152 41080
rect 21836 40718 22048 40746
rect 22204 40730 22232 42298
rect 22192 40724 22244 40730
rect 21836 40390 21864 40718
rect 22192 40666 22244 40672
rect 22008 40656 22060 40662
rect 22008 40598 22060 40604
rect 22100 40656 22152 40662
rect 22100 40598 22152 40604
rect 22020 40526 22048 40598
rect 22008 40520 22060 40526
rect 22008 40462 22060 40468
rect 21824 40384 21876 40390
rect 22112 40338 22140 40598
rect 21824 40326 21876 40332
rect 22020 40310 22140 40338
rect 21824 39976 21876 39982
rect 21824 39918 21876 39924
rect 21732 39568 21784 39574
rect 21732 39510 21784 39516
rect 21640 37460 21692 37466
rect 21640 37402 21692 37408
rect 21640 36916 21692 36922
rect 21640 36858 21692 36864
rect 21548 34672 21600 34678
rect 21548 34614 21600 34620
rect 21560 34202 21588 34614
rect 21652 34542 21680 36858
rect 21744 36718 21772 39510
rect 21836 39506 21864 39918
rect 21916 39840 21968 39846
rect 21916 39782 21968 39788
rect 21824 39500 21876 39506
rect 21824 39442 21876 39448
rect 21928 37942 21956 39782
rect 22020 38826 22048 40310
rect 22098 40216 22154 40225
rect 22098 40151 22100 40160
rect 22152 40151 22154 40160
rect 22100 40122 22152 40128
rect 22008 38820 22060 38826
rect 22008 38762 22060 38768
rect 22112 38486 22140 40122
rect 22100 38480 22152 38486
rect 22100 38422 22152 38428
rect 22008 38276 22060 38282
rect 22008 38218 22060 38224
rect 22020 38010 22048 38218
rect 22112 38010 22140 38422
rect 22296 38418 22324 42327
rect 22388 41682 22416 42774
rect 22480 42226 22508 46446
rect 22572 43858 22600 52838
rect 22950 52796 23258 52805
rect 22950 52794 22956 52796
rect 23012 52794 23036 52796
rect 23092 52794 23116 52796
rect 23172 52794 23196 52796
rect 23252 52794 23258 52796
rect 23012 52742 23014 52794
rect 23194 52742 23196 52794
rect 22950 52740 22956 52742
rect 23012 52740 23036 52742
rect 23092 52740 23116 52742
rect 23172 52740 23196 52742
rect 23252 52740 23258 52742
rect 22950 52731 23258 52740
rect 22950 51708 23258 51717
rect 22950 51706 22956 51708
rect 23012 51706 23036 51708
rect 23092 51706 23116 51708
rect 23172 51706 23196 51708
rect 23252 51706 23258 51708
rect 23012 51654 23014 51706
rect 23194 51654 23196 51706
rect 22950 51652 22956 51654
rect 23012 51652 23036 51654
rect 23092 51652 23116 51654
rect 23172 51652 23196 51654
rect 23252 51652 23258 51654
rect 22950 51643 23258 51652
rect 22950 50620 23258 50629
rect 22950 50618 22956 50620
rect 23012 50618 23036 50620
rect 23092 50618 23116 50620
rect 23172 50618 23196 50620
rect 23252 50618 23258 50620
rect 23012 50566 23014 50618
rect 23194 50566 23196 50618
rect 22950 50564 22956 50566
rect 23012 50564 23036 50566
rect 23092 50564 23116 50566
rect 23172 50564 23196 50566
rect 23252 50564 23258 50566
rect 22950 50555 23258 50564
rect 22950 49532 23258 49541
rect 22950 49530 22956 49532
rect 23012 49530 23036 49532
rect 23092 49530 23116 49532
rect 23172 49530 23196 49532
rect 23252 49530 23258 49532
rect 23012 49478 23014 49530
rect 23194 49478 23196 49530
rect 22950 49476 22956 49478
rect 23012 49476 23036 49478
rect 23092 49476 23116 49478
rect 23172 49476 23196 49478
rect 23252 49476 23258 49478
rect 22950 49467 23258 49476
rect 22950 48444 23258 48453
rect 22950 48442 22956 48444
rect 23012 48442 23036 48444
rect 23092 48442 23116 48444
rect 23172 48442 23196 48444
rect 23252 48442 23258 48444
rect 23012 48390 23014 48442
rect 23194 48390 23196 48442
rect 22950 48388 22956 48390
rect 23012 48388 23036 48390
rect 23092 48388 23116 48390
rect 23172 48388 23196 48390
rect 23252 48388 23258 48390
rect 22950 48379 23258 48388
rect 23296 47592 23348 47598
rect 23296 47534 23348 47540
rect 22950 47356 23258 47365
rect 22950 47354 22956 47356
rect 23012 47354 23036 47356
rect 23092 47354 23116 47356
rect 23172 47354 23196 47356
rect 23252 47354 23258 47356
rect 23012 47302 23014 47354
rect 23194 47302 23196 47354
rect 22950 47300 22956 47302
rect 23012 47300 23036 47302
rect 23092 47300 23116 47302
rect 23172 47300 23196 47302
rect 23252 47300 23258 47302
rect 22950 47291 23258 47300
rect 22744 46368 22796 46374
rect 22744 46310 22796 46316
rect 22652 44328 22704 44334
rect 22652 44270 22704 44276
rect 22560 43852 22612 43858
rect 22560 43794 22612 43800
rect 22560 43240 22612 43246
rect 22560 43182 22612 43188
rect 22468 42220 22520 42226
rect 22468 42162 22520 42168
rect 22468 42016 22520 42022
rect 22468 41958 22520 41964
rect 22480 41818 22508 41958
rect 22468 41812 22520 41818
rect 22468 41754 22520 41760
rect 22376 41676 22428 41682
rect 22376 41618 22428 41624
rect 22376 40384 22428 40390
rect 22376 40326 22428 40332
rect 22388 40186 22416 40326
rect 22376 40180 22428 40186
rect 22376 40122 22428 40128
rect 22468 40112 22520 40118
rect 22468 40054 22520 40060
rect 22376 39976 22428 39982
rect 22376 39918 22428 39924
rect 22388 38894 22416 39918
rect 22376 38888 22428 38894
rect 22376 38830 22428 38836
rect 22284 38412 22336 38418
rect 22284 38354 22336 38360
rect 22388 38282 22416 38830
rect 22376 38276 22428 38282
rect 22376 38218 22428 38224
rect 22480 38162 22508 40054
rect 22296 38134 22508 38162
rect 22008 38004 22060 38010
rect 22008 37946 22060 37952
rect 22100 38004 22152 38010
rect 22100 37946 22152 37952
rect 21916 37936 21968 37942
rect 21916 37878 21968 37884
rect 22112 37777 22140 37946
rect 22098 37768 22154 37777
rect 22098 37703 22154 37712
rect 22192 37732 22244 37738
rect 22192 37674 22244 37680
rect 21916 37664 21968 37670
rect 21916 37606 21968 37612
rect 21928 37262 21956 37606
rect 22100 37460 22152 37466
rect 22100 37402 22152 37408
rect 22112 37262 22140 37402
rect 21916 37256 21968 37262
rect 21916 37198 21968 37204
rect 22100 37256 22152 37262
rect 22100 37198 22152 37204
rect 21824 37120 21876 37126
rect 21824 37062 21876 37068
rect 21732 36712 21784 36718
rect 21732 36654 21784 36660
rect 21640 34536 21692 34542
rect 21640 34478 21692 34484
rect 21548 34196 21600 34202
rect 21548 34138 21600 34144
rect 21456 33584 21508 33590
rect 21456 33526 21508 33532
rect 21272 33516 21324 33522
rect 21272 33458 21324 33464
rect 21270 33416 21326 33425
rect 21270 33351 21326 33360
rect 21284 32026 21312 33351
rect 21640 33312 21692 33318
rect 21640 33254 21692 33260
rect 21456 32904 21508 32910
rect 21456 32846 21508 32852
rect 21364 32836 21416 32842
rect 21364 32778 21416 32784
rect 21376 32502 21404 32778
rect 21364 32496 21416 32502
rect 21364 32438 21416 32444
rect 21272 32020 21324 32026
rect 21272 31962 21324 31968
rect 21272 31748 21324 31754
rect 21272 31690 21324 31696
rect 21178 30560 21234 30569
rect 21178 30495 21234 30504
rect 20904 30184 20956 30190
rect 20904 30126 20956 30132
rect 20916 29866 20944 30126
rect 20916 29838 21036 29866
rect 20904 29708 20956 29714
rect 20904 29650 20956 29656
rect 20812 29164 20864 29170
rect 20812 29106 20864 29112
rect 20536 29096 20588 29102
rect 20536 29038 20588 29044
rect 20364 27390 20484 27418
rect 20364 24682 20392 27390
rect 20444 27328 20496 27334
rect 20444 27270 20496 27276
rect 20456 27169 20484 27270
rect 20442 27160 20498 27169
rect 20442 27095 20444 27104
rect 20496 27095 20498 27104
rect 20444 27066 20496 27072
rect 20456 26382 20484 27066
rect 20444 26376 20496 26382
rect 20444 26318 20496 26324
rect 20352 24676 20404 24682
rect 20352 24618 20404 24624
rect 20364 24274 20392 24618
rect 20548 24274 20576 29038
rect 20720 28416 20772 28422
rect 20720 28358 20772 28364
rect 20732 28121 20760 28358
rect 20718 28112 20774 28121
rect 20718 28047 20774 28056
rect 20916 28014 20944 29650
rect 21008 28082 21036 29838
rect 21192 28994 21220 30495
rect 21284 30138 21312 31690
rect 21376 30394 21404 32438
rect 21364 30388 21416 30394
rect 21364 30330 21416 30336
rect 21284 30110 21404 30138
rect 21272 29096 21324 29102
rect 21272 29038 21324 29044
rect 21100 28966 21220 28994
rect 20996 28076 21048 28082
rect 20996 28018 21048 28024
rect 20904 28008 20956 28014
rect 20904 27950 20956 27956
rect 20628 27328 20680 27334
rect 20628 27270 20680 27276
rect 20640 26586 20668 27270
rect 20916 26994 20944 27950
rect 21100 27538 21128 28966
rect 21284 28558 21312 29038
rect 21272 28552 21324 28558
rect 21272 28494 21324 28500
rect 21088 27532 21140 27538
rect 21088 27474 21140 27480
rect 20904 26988 20956 26994
rect 20904 26930 20956 26936
rect 20720 26784 20772 26790
rect 20720 26726 20772 26732
rect 20628 26580 20680 26586
rect 20628 26522 20680 26528
rect 20628 25832 20680 25838
rect 20628 25774 20680 25780
rect 20352 24268 20404 24274
rect 20352 24210 20404 24216
rect 20536 24268 20588 24274
rect 20536 24210 20588 24216
rect 20260 23860 20312 23866
rect 20260 23802 20312 23808
rect 19904 23174 20208 23202
rect 19904 21350 19932 23174
rect 20076 22432 20128 22438
rect 20076 22374 20128 22380
rect 19984 22160 20036 22166
rect 19984 22102 20036 22108
rect 19996 21690 20024 22102
rect 19984 21684 20036 21690
rect 19984 21626 20036 21632
rect 20088 21486 20116 22374
rect 20076 21480 20128 21486
rect 20076 21422 20128 21428
rect 19892 21344 19944 21350
rect 19892 21286 19944 21292
rect 19800 21140 19852 21146
rect 19800 21082 19852 21088
rect 19708 17740 19760 17746
rect 19708 17682 19760 17688
rect 19720 17338 19748 17682
rect 19708 17332 19760 17338
rect 19708 17274 19760 17280
rect 19616 17264 19668 17270
rect 19616 17206 19668 17212
rect 19536 17054 19748 17082
rect 19432 16788 19484 16794
rect 19432 16730 19484 16736
rect 19444 14906 19472 16730
rect 19524 16448 19576 16454
rect 19524 16390 19576 16396
rect 19536 16250 19564 16390
rect 19524 16244 19576 16250
rect 19524 16186 19576 16192
rect 19352 14878 19472 14906
rect 19248 13864 19300 13870
rect 19248 13806 19300 13812
rect 19352 13326 19380 14878
rect 19432 14816 19484 14822
rect 19432 14758 19484 14764
rect 19524 14816 19576 14822
rect 19524 14758 19576 14764
rect 19444 13870 19472 14758
rect 19432 13864 19484 13870
rect 19432 13806 19484 13812
rect 19340 13320 19392 13326
rect 19340 13262 19392 13268
rect 19536 12170 19564 14758
rect 19616 13524 19668 13530
rect 19616 13466 19668 13472
rect 19524 12164 19576 12170
rect 19524 12106 19576 12112
rect 19168 11750 19288 11778
rect 19156 10600 19208 10606
rect 19156 10542 19208 10548
rect 19064 9648 19116 9654
rect 19064 9590 19116 9596
rect 18984 6886 19104 6914
rect 19076 5234 19104 6886
rect 19064 5228 19116 5234
rect 19064 5170 19116 5176
rect 18696 4616 18748 4622
rect 18696 4558 18748 4564
rect 17950 4380 18258 4389
rect 17950 4378 17956 4380
rect 18012 4378 18036 4380
rect 18092 4378 18116 4380
rect 18172 4378 18196 4380
rect 18252 4378 18258 4380
rect 18012 4326 18014 4378
rect 18194 4326 18196 4378
rect 17950 4324 17956 4326
rect 18012 4324 18036 4326
rect 18092 4324 18116 4326
rect 18172 4324 18196 4326
rect 18252 4324 18258 4326
rect 17950 4315 18258 4324
rect 19168 3670 19196 10542
rect 19260 4146 19288 11750
rect 19524 11008 19576 11014
rect 19524 10950 19576 10956
rect 19536 10810 19564 10950
rect 19628 10810 19656 13466
rect 19720 13394 19748 17054
rect 19812 14958 19840 21082
rect 19904 17490 19932 21286
rect 20272 20874 20300 23802
rect 20548 23662 20576 24210
rect 20640 23866 20668 25774
rect 20732 25362 20760 26726
rect 20810 26616 20866 26625
rect 20810 26551 20812 26560
rect 20864 26551 20866 26560
rect 20812 26522 20864 26528
rect 20824 26382 20852 26522
rect 20916 26450 20944 26930
rect 21272 26852 21324 26858
rect 21272 26794 21324 26800
rect 20904 26444 20956 26450
rect 20904 26386 20956 26392
rect 20812 26376 20864 26382
rect 20812 26318 20864 26324
rect 20720 25356 20772 25362
rect 20720 25298 20772 25304
rect 20628 23860 20680 23866
rect 20628 23802 20680 23808
rect 20536 23656 20588 23662
rect 20536 23598 20588 23604
rect 20720 23520 20772 23526
rect 20772 23480 20852 23508
rect 20720 23462 20772 23468
rect 20824 23118 20852 23480
rect 21088 23180 21140 23186
rect 21088 23122 21140 23128
rect 20812 23112 20864 23118
rect 20812 23054 20864 23060
rect 20720 22976 20772 22982
rect 20720 22918 20772 22924
rect 20536 22636 20588 22642
rect 20536 22578 20588 22584
rect 20548 21962 20576 22578
rect 20536 21956 20588 21962
rect 20536 21898 20588 21904
rect 20260 20868 20312 20874
rect 20260 20810 20312 20816
rect 20444 20800 20496 20806
rect 20444 20742 20496 20748
rect 20456 19854 20484 20742
rect 20444 19848 20496 19854
rect 20444 19790 20496 19796
rect 20260 19780 20312 19786
rect 20260 19722 20312 19728
rect 19984 18624 20036 18630
rect 19984 18566 20036 18572
rect 19996 17610 20024 18566
rect 19984 17604 20036 17610
rect 19984 17546 20036 17552
rect 19904 17462 20024 17490
rect 19892 16516 19944 16522
rect 19892 16458 19944 16464
rect 19904 15570 19932 16458
rect 19892 15564 19944 15570
rect 19892 15506 19944 15512
rect 19800 14952 19852 14958
rect 19800 14894 19852 14900
rect 19904 14550 19932 15506
rect 19892 14544 19944 14550
rect 19892 14486 19944 14492
rect 19996 13394 20024 17462
rect 20272 16590 20300 19722
rect 20352 18964 20404 18970
rect 20352 18906 20404 18912
rect 20260 16584 20312 16590
rect 20260 16526 20312 16532
rect 20364 16250 20392 18906
rect 20548 18358 20576 21898
rect 20732 21690 20760 22918
rect 20824 22234 20852 23054
rect 21100 22574 21128 23122
rect 21088 22568 21140 22574
rect 21088 22510 21140 22516
rect 20812 22228 20864 22234
rect 20812 22170 20864 22176
rect 21100 22030 21128 22510
rect 20812 22024 20864 22030
rect 20812 21966 20864 21972
rect 21088 22024 21140 22030
rect 21088 21966 21140 21972
rect 20720 21684 20772 21690
rect 20720 21626 20772 21632
rect 20824 21010 20852 21966
rect 21284 21894 21312 26794
rect 21376 25362 21404 30110
rect 21468 28218 21496 32846
rect 21546 32056 21602 32065
rect 21546 31991 21602 32000
rect 21560 31958 21588 31991
rect 21548 31952 21600 31958
rect 21548 31894 21600 31900
rect 21652 31414 21680 33254
rect 21730 33008 21786 33017
rect 21730 32943 21786 32952
rect 21744 32910 21772 32943
rect 21732 32904 21784 32910
rect 21732 32846 21784 32852
rect 21836 32502 21864 37062
rect 22100 36100 22152 36106
rect 22100 36042 22152 36048
rect 21916 35760 21968 35766
rect 21916 35702 21968 35708
rect 21928 34202 21956 35702
rect 22008 35216 22060 35222
rect 22006 35184 22008 35193
rect 22060 35184 22062 35193
rect 22006 35119 22062 35128
rect 22112 34542 22140 36042
rect 22204 35018 22232 37674
rect 22192 35012 22244 35018
rect 22192 34954 22244 34960
rect 22100 34536 22152 34542
rect 22100 34478 22152 34484
rect 22008 34400 22060 34406
rect 22008 34342 22060 34348
rect 21916 34196 21968 34202
rect 21916 34138 21968 34144
rect 21916 32904 21968 32910
rect 21916 32846 21968 32852
rect 21928 32774 21956 32846
rect 21916 32768 21968 32774
rect 21916 32710 21968 32716
rect 21824 32496 21876 32502
rect 21824 32438 21876 32444
rect 21824 32224 21876 32230
rect 21824 32166 21876 32172
rect 21836 31754 21864 32166
rect 21744 31726 21864 31754
rect 21640 31408 21692 31414
rect 21640 31350 21692 31356
rect 21456 28212 21508 28218
rect 21456 28154 21508 28160
rect 21640 28144 21692 28150
rect 21640 28086 21692 28092
rect 21548 26512 21600 26518
rect 21548 26454 21600 26460
rect 21364 25356 21416 25362
rect 21364 25298 21416 25304
rect 21364 21956 21416 21962
rect 21364 21898 21416 21904
rect 20904 21888 20956 21894
rect 20904 21830 20956 21836
rect 21272 21888 21324 21894
rect 21272 21830 21324 21836
rect 20812 21004 20864 21010
rect 20812 20946 20864 20952
rect 20628 19304 20680 19310
rect 20628 19246 20680 19252
rect 20720 19304 20772 19310
rect 20720 19246 20772 19252
rect 20536 18352 20588 18358
rect 20536 18294 20588 18300
rect 20548 17882 20576 18294
rect 20536 17876 20588 17882
rect 20536 17818 20588 17824
rect 20640 17338 20668 19246
rect 20732 18426 20760 19246
rect 20916 19174 20944 21830
rect 21376 20602 21404 21898
rect 21364 20596 21416 20602
rect 21364 20538 21416 20544
rect 21456 19848 21508 19854
rect 21456 19790 21508 19796
rect 21180 19440 21232 19446
rect 21180 19382 21232 19388
rect 21192 19310 21220 19382
rect 21180 19304 21232 19310
rect 21180 19246 21232 19252
rect 20904 19168 20956 19174
rect 20904 19110 20956 19116
rect 21364 18964 21416 18970
rect 21364 18906 21416 18912
rect 20996 18760 21048 18766
rect 20996 18702 21048 18708
rect 20720 18420 20772 18426
rect 20720 18362 20772 18368
rect 20732 17610 20760 18362
rect 21008 18154 21036 18702
rect 20996 18148 21048 18154
rect 20996 18090 21048 18096
rect 20720 17604 20772 17610
rect 20720 17546 20772 17552
rect 20628 17332 20680 17338
rect 20628 17274 20680 17280
rect 20732 17270 20760 17546
rect 20720 17264 20772 17270
rect 20720 17206 20772 17212
rect 20628 17196 20680 17202
rect 20628 17138 20680 17144
rect 20444 16992 20496 16998
rect 20444 16934 20496 16940
rect 20352 16244 20404 16250
rect 20352 16186 20404 16192
rect 20456 15978 20484 16934
rect 20536 16448 20588 16454
rect 20536 16390 20588 16396
rect 20444 15972 20496 15978
rect 20444 15914 20496 15920
rect 20548 15570 20576 16390
rect 20536 15564 20588 15570
rect 20536 15506 20588 15512
rect 20536 15428 20588 15434
rect 20536 15370 20588 15376
rect 20548 14006 20576 15370
rect 20640 15162 20668 17138
rect 20812 16652 20864 16658
rect 20812 16594 20864 16600
rect 20904 16652 20956 16658
rect 20904 16594 20956 16600
rect 20718 16552 20774 16561
rect 20718 16487 20774 16496
rect 20732 15502 20760 16487
rect 20720 15496 20772 15502
rect 20720 15438 20772 15444
rect 20628 15156 20680 15162
rect 20628 15098 20680 15104
rect 20536 14000 20588 14006
rect 20536 13942 20588 13948
rect 20640 13870 20668 15098
rect 20260 13864 20312 13870
rect 20260 13806 20312 13812
rect 20628 13864 20680 13870
rect 20628 13806 20680 13812
rect 19708 13388 19760 13394
rect 19708 13330 19760 13336
rect 19984 13388 20036 13394
rect 19984 13330 20036 13336
rect 19892 13320 19944 13326
rect 19892 13262 19944 13268
rect 19904 12986 19932 13262
rect 19984 13252 20036 13258
rect 19984 13194 20036 13200
rect 19892 12980 19944 12986
rect 19892 12922 19944 12928
rect 19800 12164 19852 12170
rect 19800 12106 19852 12112
rect 19708 11756 19760 11762
rect 19708 11698 19760 11704
rect 19720 11558 19748 11698
rect 19708 11552 19760 11558
rect 19708 11494 19760 11500
rect 19524 10804 19576 10810
rect 19524 10746 19576 10752
rect 19616 10804 19668 10810
rect 19616 10746 19668 10752
rect 19720 10606 19748 11494
rect 19708 10600 19760 10606
rect 19708 10542 19760 10548
rect 19812 7886 19840 12106
rect 19800 7880 19852 7886
rect 19800 7822 19852 7828
rect 19524 5296 19576 5302
rect 19524 5238 19576 5244
rect 19340 5160 19392 5166
rect 19340 5102 19392 5108
rect 19248 4140 19300 4146
rect 19248 4082 19300 4088
rect 19156 3664 19208 3670
rect 19156 3606 19208 3612
rect 18972 3460 19024 3466
rect 18972 3402 19024 3408
rect 17950 3292 18258 3301
rect 17950 3290 17956 3292
rect 18012 3290 18036 3292
rect 18092 3290 18116 3292
rect 18172 3290 18196 3292
rect 18252 3290 18258 3292
rect 18012 3238 18014 3290
rect 18194 3238 18196 3290
rect 17950 3236 17956 3238
rect 18012 3236 18036 3238
rect 18092 3236 18116 3238
rect 18172 3236 18196 3238
rect 18252 3236 18258 3238
rect 17950 3227 18258 3236
rect 17868 3052 17920 3058
rect 17868 2994 17920 3000
rect 18512 3052 18564 3058
rect 18512 2994 18564 3000
rect 18524 2514 18552 2994
rect 18604 2848 18656 2854
rect 18604 2790 18656 2796
rect 18512 2508 18564 2514
rect 18512 2450 18564 2456
rect 18328 2304 18380 2310
rect 18328 2246 18380 2252
rect 17950 2204 18258 2213
rect 17950 2202 17956 2204
rect 18012 2202 18036 2204
rect 18092 2202 18116 2204
rect 18172 2202 18196 2204
rect 18252 2202 18258 2204
rect 18012 2150 18014 2202
rect 18194 2150 18196 2202
rect 17950 2148 17956 2150
rect 18012 2148 18036 2150
rect 18092 2148 18116 2150
rect 18172 2148 18196 2150
rect 18252 2148 18258 2150
rect 17950 2139 18258 2148
rect 17788 1686 17908 1714
rect 17880 800 17908 1686
rect 18340 1170 18368 2246
rect 18248 1142 18368 1170
rect 18248 800 18276 1142
rect 18616 800 18644 2790
rect 18984 800 19012 3402
rect 19352 800 19380 5102
rect 19536 3942 19564 5238
rect 19892 4684 19944 4690
rect 19892 4626 19944 4632
rect 19524 3936 19576 3942
rect 19524 3878 19576 3884
rect 19708 2916 19760 2922
rect 19708 2858 19760 2864
rect 19720 800 19748 2858
rect 19904 2854 19932 4626
rect 19996 4146 20024 13194
rect 20272 11830 20300 13806
rect 20824 13462 20852 16594
rect 20916 14414 20944 16594
rect 21008 16046 21036 18090
rect 21086 16552 21142 16561
rect 21086 16487 21088 16496
rect 21140 16487 21142 16496
rect 21088 16458 21140 16464
rect 21376 16182 21404 18906
rect 21468 17882 21496 19790
rect 21560 18834 21588 26454
rect 21652 25226 21680 28086
rect 21744 25430 21772 31726
rect 22020 29306 22048 34342
rect 22100 33856 22152 33862
rect 22100 33798 22152 33804
rect 22112 31414 22140 33798
rect 22204 33454 22232 34954
rect 22296 33538 22324 38134
rect 22376 37664 22428 37670
rect 22376 37606 22428 37612
rect 22388 35057 22416 37606
rect 22572 37330 22600 43182
rect 22664 42362 22692 44270
rect 22756 42634 22784 46310
rect 22950 46268 23258 46277
rect 22950 46266 22956 46268
rect 23012 46266 23036 46268
rect 23092 46266 23116 46268
rect 23172 46266 23196 46268
rect 23252 46266 23258 46268
rect 23012 46214 23014 46266
rect 23194 46214 23196 46266
rect 22950 46212 22956 46214
rect 23012 46212 23036 46214
rect 23092 46212 23116 46214
rect 23172 46212 23196 46214
rect 23252 46212 23258 46214
rect 22950 46203 23258 46212
rect 22836 45824 22888 45830
rect 22836 45766 22888 45772
rect 22744 42628 22796 42634
rect 22744 42570 22796 42576
rect 22848 42514 22876 45766
rect 22950 45180 23258 45189
rect 22950 45178 22956 45180
rect 23012 45178 23036 45180
rect 23092 45178 23116 45180
rect 23172 45178 23196 45180
rect 23252 45178 23258 45180
rect 23012 45126 23014 45178
rect 23194 45126 23196 45178
rect 22950 45124 22956 45126
rect 23012 45124 23036 45126
rect 23092 45124 23116 45126
rect 23172 45124 23196 45126
rect 23252 45124 23258 45126
rect 22950 45115 23258 45124
rect 22950 44092 23258 44101
rect 22950 44090 22956 44092
rect 23012 44090 23036 44092
rect 23092 44090 23116 44092
rect 23172 44090 23196 44092
rect 23252 44090 23258 44092
rect 23012 44038 23014 44090
rect 23194 44038 23196 44090
rect 22950 44036 22956 44038
rect 23012 44036 23036 44038
rect 23092 44036 23116 44038
rect 23172 44036 23196 44038
rect 23252 44036 23258 44038
rect 22950 44027 23258 44036
rect 22950 43004 23258 43013
rect 22950 43002 22956 43004
rect 23012 43002 23036 43004
rect 23092 43002 23116 43004
rect 23172 43002 23196 43004
rect 23252 43002 23258 43004
rect 23012 42950 23014 43002
rect 23194 42950 23196 43002
rect 22950 42948 22956 42950
rect 23012 42948 23036 42950
rect 23092 42948 23116 42950
rect 23172 42948 23196 42950
rect 23252 42948 23258 42950
rect 22950 42939 23258 42948
rect 23020 42764 23072 42770
rect 23020 42706 23072 42712
rect 22756 42486 22876 42514
rect 22652 42356 22704 42362
rect 22652 42298 22704 42304
rect 22652 42220 22704 42226
rect 22652 42162 22704 42168
rect 22664 40526 22692 42162
rect 22756 41682 22784 42486
rect 23032 42129 23060 42706
rect 23204 42696 23256 42702
rect 23204 42638 23256 42644
rect 23216 42401 23244 42638
rect 23202 42392 23258 42401
rect 23202 42327 23258 42336
rect 23018 42120 23074 42129
rect 23018 42055 23074 42064
rect 23308 42022 23336 47534
rect 23388 44736 23440 44742
rect 23388 44678 23440 44684
rect 23296 42016 23348 42022
rect 23296 41958 23348 41964
rect 22950 41916 23258 41925
rect 22950 41914 22956 41916
rect 23012 41914 23036 41916
rect 23092 41914 23116 41916
rect 23172 41914 23196 41916
rect 23252 41914 23258 41916
rect 23012 41862 23014 41914
rect 23194 41862 23196 41914
rect 22950 41860 22956 41862
rect 23012 41860 23036 41862
rect 23092 41860 23116 41862
rect 23172 41860 23196 41862
rect 23252 41860 23258 41862
rect 22950 41851 23258 41860
rect 22928 41744 22980 41750
rect 22928 41686 22980 41692
rect 23204 41744 23256 41750
rect 23204 41686 23256 41692
rect 22744 41676 22796 41682
rect 22744 41618 22796 41624
rect 22744 41472 22796 41478
rect 22744 41414 22796 41420
rect 22940 41414 22968 41686
rect 22652 40520 22704 40526
rect 22652 40462 22704 40468
rect 22664 40186 22692 40462
rect 22652 40180 22704 40186
rect 22652 40122 22704 40128
rect 22756 39642 22784 41414
rect 22848 41386 22968 41414
rect 22848 40526 22876 41386
rect 23216 41206 23244 41686
rect 23204 41200 23256 41206
rect 23204 41142 23256 41148
rect 22950 40828 23258 40837
rect 22950 40826 22956 40828
rect 23012 40826 23036 40828
rect 23092 40826 23116 40828
rect 23172 40826 23196 40828
rect 23252 40826 23258 40828
rect 23012 40774 23014 40826
rect 23194 40774 23196 40826
rect 22950 40772 22956 40774
rect 23012 40772 23036 40774
rect 23092 40772 23116 40774
rect 23172 40772 23196 40774
rect 23252 40772 23258 40774
rect 22950 40763 23258 40772
rect 22836 40520 22888 40526
rect 22836 40462 22888 40468
rect 22928 40452 22980 40458
rect 22928 40394 22980 40400
rect 22940 40050 22968 40394
rect 22928 40044 22980 40050
rect 22928 39986 22980 39992
rect 22836 39840 22888 39846
rect 22836 39782 22888 39788
rect 22744 39636 22796 39642
rect 22744 39578 22796 39584
rect 22848 39098 22876 39782
rect 22950 39740 23258 39749
rect 22950 39738 22956 39740
rect 23012 39738 23036 39740
rect 23092 39738 23116 39740
rect 23172 39738 23196 39740
rect 23252 39738 23258 39740
rect 23012 39686 23014 39738
rect 23194 39686 23196 39738
rect 22950 39684 22956 39686
rect 23012 39684 23036 39686
rect 23092 39684 23116 39686
rect 23172 39684 23196 39686
rect 23252 39684 23258 39686
rect 22950 39675 23258 39684
rect 22836 39092 22888 39098
rect 22836 39034 22888 39040
rect 22950 38652 23258 38661
rect 22950 38650 22956 38652
rect 23012 38650 23036 38652
rect 23092 38650 23116 38652
rect 23172 38650 23196 38652
rect 23252 38650 23258 38652
rect 23012 38598 23014 38650
rect 23194 38598 23196 38650
rect 22950 38596 22956 38598
rect 23012 38596 23036 38598
rect 23092 38596 23116 38598
rect 23172 38596 23196 38598
rect 23252 38596 23258 38598
rect 22950 38587 23258 38596
rect 22836 38276 22888 38282
rect 22836 38218 22888 38224
rect 23204 38276 23256 38282
rect 23204 38218 23256 38224
rect 22744 38208 22796 38214
rect 22744 38150 22796 38156
rect 22650 38040 22706 38049
rect 22650 37975 22652 37984
rect 22704 37975 22706 37984
rect 22652 37946 22704 37952
rect 22560 37324 22612 37330
rect 22560 37266 22612 37272
rect 22664 37126 22692 37946
rect 22652 37120 22704 37126
rect 22652 37062 22704 37068
rect 22560 36916 22612 36922
rect 22560 36858 22612 36864
rect 22468 35624 22520 35630
rect 22468 35566 22520 35572
rect 22374 35048 22430 35057
rect 22374 34983 22430 34992
rect 22376 34944 22428 34950
rect 22376 34886 22428 34892
rect 22388 33658 22416 34886
rect 22376 33652 22428 33658
rect 22376 33594 22428 33600
rect 22296 33510 22416 33538
rect 22192 33448 22244 33454
rect 22192 33390 22244 33396
rect 22190 33144 22246 33153
rect 22190 33079 22246 33088
rect 22204 32434 22232 33079
rect 22284 32768 22336 32774
rect 22284 32710 22336 32716
rect 22192 32428 22244 32434
rect 22192 32370 22244 32376
rect 22296 31754 22324 32710
rect 22388 32434 22416 33510
rect 22480 33114 22508 35566
rect 22572 34746 22600 36858
rect 22652 36712 22704 36718
rect 22652 36654 22704 36660
rect 22664 36378 22692 36654
rect 22652 36372 22704 36378
rect 22652 36314 22704 36320
rect 22652 36032 22704 36038
rect 22652 35974 22704 35980
rect 22664 35834 22692 35974
rect 22652 35828 22704 35834
rect 22652 35770 22704 35776
rect 22650 35048 22706 35057
rect 22650 34983 22706 34992
rect 22560 34740 22612 34746
rect 22560 34682 22612 34688
rect 22560 34400 22612 34406
rect 22560 34342 22612 34348
rect 22468 33108 22520 33114
rect 22468 33050 22520 33056
rect 22468 32768 22520 32774
rect 22468 32710 22520 32716
rect 22376 32428 22428 32434
rect 22376 32370 22428 32376
rect 22480 32314 22508 32710
rect 22388 32286 22508 32314
rect 22284 31748 22336 31754
rect 22284 31690 22336 31696
rect 22192 31476 22244 31482
rect 22192 31418 22244 31424
rect 22100 31408 22152 31414
rect 22100 31350 22152 31356
rect 22204 31226 22232 31418
rect 22112 31198 22232 31226
rect 21824 29300 21876 29306
rect 21824 29242 21876 29248
rect 22008 29300 22060 29306
rect 22008 29242 22060 29248
rect 21836 28422 21864 29242
rect 21916 29028 21968 29034
rect 21916 28970 21968 28976
rect 21824 28416 21876 28422
rect 21824 28358 21876 28364
rect 21824 26444 21876 26450
rect 21824 26386 21876 26392
rect 21732 25424 21784 25430
rect 21732 25366 21784 25372
rect 21640 25220 21692 25226
rect 21640 25162 21692 25168
rect 21652 24954 21680 25162
rect 21640 24948 21692 24954
rect 21640 24890 21692 24896
rect 21652 23866 21680 24890
rect 21836 24154 21864 26386
rect 21928 24274 21956 28970
rect 22008 28008 22060 28014
rect 22008 27950 22060 27956
rect 22020 27470 22048 27950
rect 22112 27674 22140 31198
rect 22388 30954 22416 32286
rect 22468 32224 22520 32230
rect 22468 32166 22520 32172
rect 22296 30926 22416 30954
rect 22192 30864 22244 30870
rect 22192 30806 22244 30812
rect 22204 28150 22232 30806
rect 22192 28144 22244 28150
rect 22192 28086 22244 28092
rect 22100 27668 22152 27674
rect 22100 27610 22152 27616
rect 22192 27600 22244 27606
rect 22192 27542 22244 27548
rect 22008 27464 22060 27470
rect 22008 27406 22060 27412
rect 22020 26926 22048 27406
rect 22008 26920 22060 26926
rect 22008 26862 22060 26868
rect 22100 26580 22152 26586
rect 22100 26522 22152 26528
rect 22112 25242 22140 26522
rect 22204 26042 22232 27542
rect 22296 27010 22324 30926
rect 22480 29186 22508 32166
rect 22572 31482 22600 34342
rect 22664 34218 22692 34983
rect 22756 34377 22784 38150
rect 22848 37806 22876 38218
rect 22928 38208 22980 38214
rect 22928 38150 22980 38156
rect 22940 37942 22968 38150
rect 22928 37936 22980 37942
rect 22928 37878 22980 37884
rect 22836 37800 22888 37806
rect 22836 37742 22888 37748
rect 22848 36718 22876 37742
rect 23216 37738 23244 38218
rect 23204 37732 23256 37738
rect 23204 37674 23256 37680
rect 22950 37564 23258 37573
rect 22950 37562 22956 37564
rect 23012 37562 23036 37564
rect 23092 37562 23116 37564
rect 23172 37562 23196 37564
rect 23252 37562 23258 37564
rect 23012 37510 23014 37562
rect 23194 37510 23196 37562
rect 22950 37508 22956 37510
rect 23012 37508 23036 37510
rect 23092 37508 23116 37510
rect 23172 37508 23196 37510
rect 23252 37508 23258 37510
rect 22950 37499 23258 37508
rect 23308 37346 23336 41958
rect 23400 40594 23428 44678
rect 23480 43240 23532 43246
rect 23480 43182 23532 43188
rect 23492 42158 23520 43182
rect 23480 42152 23532 42158
rect 23480 42094 23532 42100
rect 23492 41750 23520 42094
rect 23480 41744 23532 41750
rect 23480 41686 23532 41692
rect 23584 40662 23612 53926
rect 23676 53106 23704 55186
rect 24504 54330 24532 56199
rect 24674 55448 24730 55457
rect 24674 55383 24730 55392
rect 24688 54330 24716 55383
rect 24766 54632 24822 54641
rect 24766 54567 24822 54576
rect 24492 54324 24544 54330
rect 24492 54266 24544 54272
rect 24676 54324 24728 54330
rect 24676 54266 24728 54272
rect 24504 53582 24532 54266
rect 24780 53582 24808 54567
rect 25044 54188 25096 54194
rect 25044 54130 25096 54136
rect 25056 53825 25084 54130
rect 25042 53816 25098 53825
rect 25042 53751 25098 53760
rect 25318 53816 25374 53825
rect 25318 53751 25374 53760
rect 24492 53576 24544 53582
rect 24492 53518 24544 53524
rect 24768 53576 24820 53582
rect 24768 53518 24820 53524
rect 23940 53440 23992 53446
rect 23940 53382 23992 53388
rect 23664 53100 23716 53106
rect 23664 53042 23716 53048
rect 23952 53009 23980 53382
rect 23938 53000 23994 53009
rect 23938 52935 23994 52944
rect 23940 52896 23992 52902
rect 23940 52838 23992 52844
rect 23756 47048 23808 47054
rect 23756 46990 23808 46996
rect 23768 42650 23796 46990
rect 23848 46912 23900 46918
rect 23848 46854 23900 46860
rect 23860 45830 23888 46854
rect 23952 45966 23980 52838
rect 24780 52698 24808 53518
rect 25044 53440 25096 53446
rect 25044 53382 25096 53388
rect 25056 53281 25084 53382
rect 25042 53272 25098 53281
rect 25042 53207 25098 53216
rect 25044 53100 25096 53106
rect 25044 53042 25096 53048
rect 25056 53009 25084 53042
rect 25042 53000 25098 53009
rect 25042 52935 25098 52944
rect 24860 52896 24912 52902
rect 24860 52838 24912 52844
rect 24768 52692 24820 52698
rect 24768 52634 24820 52640
rect 24768 52488 24820 52494
rect 24768 52430 24820 52436
rect 24780 52193 24808 52430
rect 24766 52184 24822 52193
rect 24766 52119 24822 52128
rect 24308 50720 24360 50726
rect 24308 50662 24360 50668
rect 23940 45960 23992 45966
rect 23940 45902 23992 45908
rect 24032 45960 24084 45966
rect 24032 45902 24084 45908
rect 23848 45824 23900 45830
rect 23848 45766 23900 45772
rect 23860 45558 23888 45766
rect 23848 45552 23900 45558
rect 23848 45494 23900 45500
rect 23860 45422 23888 45494
rect 23848 45416 23900 45422
rect 23848 45358 23900 45364
rect 23860 45082 23888 45358
rect 23848 45076 23900 45082
rect 23848 45018 23900 45024
rect 23860 44810 23888 45018
rect 23848 44804 23900 44810
rect 23848 44746 23900 44752
rect 23860 44470 23888 44746
rect 24044 44742 24072 45902
rect 24216 45824 24268 45830
rect 24216 45766 24268 45772
rect 24124 44872 24176 44878
rect 24124 44814 24176 44820
rect 24032 44736 24084 44742
rect 24032 44678 24084 44684
rect 23848 44464 23900 44470
rect 23848 44406 23900 44412
rect 23860 43722 23888 44406
rect 24032 44192 24084 44198
rect 24136 44180 24164 44814
rect 24084 44152 24164 44180
rect 24032 44134 24084 44140
rect 23848 43716 23900 43722
rect 23848 43658 23900 43664
rect 23940 43648 23992 43654
rect 23940 43590 23992 43596
rect 23848 43240 23900 43246
rect 23848 43182 23900 43188
rect 23676 42622 23796 42650
rect 23676 42106 23704 42622
rect 23756 42560 23808 42566
rect 23756 42502 23808 42508
rect 23768 42294 23796 42502
rect 23756 42288 23808 42294
rect 23756 42230 23808 42236
rect 23676 42078 23796 42106
rect 23664 41676 23716 41682
rect 23664 41618 23716 41624
rect 23572 40656 23624 40662
rect 23572 40598 23624 40604
rect 23388 40588 23440 40594
rect 23388 40530 23440 40536
rect 23388 40452 23440 40458
rect 23388 40394 23440 40400
rect 23400 37942 23428 40394
rect 23572 40384 23624 40390
rect 23572 40326 23624 40332
rect 23480 38344 23532 38350
rect 23480 38286 23532 38292
rect 23388 37936 23440 37942
rect 23388 37878 23440 37884
rect 23400 37670 23428 37878
rect 23388 37664 23440 37670
rect 23388 37606 23440 37612
rect 23386 37496 23442 37505
rect 23386 37431 23442 37440
rect 23112 37324 23164 37330
rect 23112 37266 23164 37272
rect 23216 37318 23336 37346
rect 23124 36718 23152 37266
rect 23216 36922 23244 37318
rect 23296 37256 23348 37262
rect 23296 37198 23348 37204
rect 23204 36916 23256 36922
rect 23204 36858 23256 36864
rect 22836 36712 22888 36718
rect 22836 36654 22888 36660
rect 23112 36712 23164 36718
rect 23112 36654 23164 36660
rect 22848 35766 22876 36654
rect 22950 36476 23258 36485
rect 22950 36474 22956 36476
rect 23012 36474 23036 36476
rect 23092 36474 23116 36476
rect 23172 36474 23196 36476
rect 23252 36474 23258 36476
rect 23012 36422 23014 36474
rect 23194 36422 23196 36474
rect 22950 36420 22956 36422
rect 23012 36420 23036 36422
rect 23092 36420 23116 36422
rect 23172 36420 23196 36422
rect 23252 36420 23258 36422
rect 22950 36411 23258 36420
rect 22928 35828 22980 35834
rect 22928 35770 22980 35776
rect 22836 35760 22888 35766
rect 22836 35702 22888 35708
rect 22940 35578 22968 35770
rect 23308 35714 23336 37198
rect 23400 36854 23428 37431
rect 23492 37126 23520 38286
rect 23480 37120 23532 37126
rect 23480 37062 23532 37068
rect 23388 36848 23440 36854
rect 23388 36790 23440 36796
rect 23480 36712 23532 36718
rect 23400 36672 23480 36700
rect 23400 35850 23428 36672
rect 23480 36654 23532 36660
rect 23400 35834 23520 35850
rect 23400 35828 23532 35834
rect 23400 35822 23480 35828
rect 23480 35770 23532 35776
rect 23124 35686 23336 35714
rect 23388 35760 23440 35766
rect 23388 35702 23440 35708
rect 23124 35630 23152 35686
rect 22848 35550 22968 35578
rect 23112 35624 23164 35630
rect 23112 35566 23164 35572
rect 22742 34368 22798 34377
rect 22742 34303 22798 34312
rect 22664 34190 22784 34218
rect 22652 34128 22704 34134
rect 22652 34070 22704 34076
rect 22664 33114 22692 34070
rect 22652 33108 22704 33114
rect 22652 33050 22704 33056
rect 22756 32994 22784 34190
rect 22848 33046 22876 35550
rect 22950 35388 23258 35397
rect 22950 35386 22956 35388
rect 23012 35386 23036 35388
rect 23092 35386 23116 35388
rect 23172 35386 23196 35388
rect 23252 35386 23258 35388
rect 23012 35334 23014 35386
rect 23194 35334 23196 35386
rect 22950 35332 22956 35334
rect 23012 35332 23036 35334
rect 23092 35332 23116 35334
rect 23172 35332 23196 35334
rect 23252 35332 23258 35334
rect 22950 35323 23258 35332
rect 23202 35184 23258 35193
rect 23400 35170 23428 35702
rect 23308 35154 23428 35170
rect 23202 35119 23258 35128
rect 23296 35148 23428 35154
rect 23216 34388 23244 35119
rect 23348 35142 23428 35148
rect 23296 35090 23348 35096
rect 23216 34360 23336 34388
rect 22950 34300 23258 34309
rect 22950 34298 22956 34300
rect 23012 34298 23036 34300
rect 23092 34298 23116 34300
rect 23172 34298 23196 34300
rect 23252 34298 23258 34300
rect 23012 34246 23014 34298
rect 23194 34246 23196 34298
rect 22950 34244 22956 34246
rect 23012 34244 23036 34246
rect 23092 34244 23116 34246
rect 23172 34244 23196 34246
rect 23252 34244 23258 34246
rect 22950 34235 23258 34244
rect 22926 34096 22982 34105
rect 22926 34031 22928 34040
rect 22980 34031 22982 34040
rect 22928 34002 22980 34008
rect 22950 33212 23258 33221
rect 22950 33210 22956 33212
rect 23012 33210 23036 33212
rect 23092 33210 23116 33212
rect 23172 33210 23196 33212
rect 23252 33210 23258 33212
rect 23012 33158 23014 33210
rect 23194 33158 23196 33210
rect 22950 33156 22956 33158
rect 23012 33156 23036 33158
rect 23092 33156 23116 33158
rect 23172 33156 23196 33158
rect 23252 33156 23258 33158
rect 22950 33147 23258 33156
rect 22664 32978 22784 32994
rect 22836 33040 22888 33046
rect 23020 33040 23072 33046
rect 22836 32982 22888 32988
rect 23018 33008 23020 33017
rect 23072 33008 23074 33017
rect 22652 32972 22784 32978
rect 22704 32966 22784 32972
rect 23018 32943 23074 32952
rect 22652 32914 22704 32920
rect 22664 32774 22692 32914
rect 23308 32892 23336 34360
rect 23400 33454 23428 35142
rect 23584 34610 23612 40326
rect 23676 39506 23704 41618
rect 23664 39500 23716 39506
rect 23664 39442 23716 39448
rect 23768 39114 23796 42078
rect 23860 41818 23888 43182
rect 23952 42906 23980 43590
rect 23940 42900 23992 42906
rect 23940 42842 23992 42848
rect 24044 42838 24072 44134
rect 24228 43790 24256 45766
rect 24320 44554 24348 50662
rect 24492 50176 24544 50182
rect 24492 50118 24544 50124
rect 24504 49774 24532 50118
rect 24492 49768 24544 49774
rect 24492 49710 24544 49716
rect 24504 48113 24532 49710
rect 24676 48680 24728 48686
rect 24676 48622 24728 48628
rect 24490 48104 24546 48113
rect 24490 48039 24546 48048
rect 24400 46980 24452 46986
rect 24400 46922 24452 46928
rect 24584 46980 24636 46986
rect 24584 46922 24636 46928
rect 24412 45801 24440 46922
rect 24596 46510 24624 46922
rect 24584 46504 24636 46510
rect 24584 46446 24636 46452
rect 24492 46368 24544 46374
rect 24492 46310 24544 46316
rect 24398 45792 24454 45801
rect 24398 45727 24454 45736
rect 24504 45422 24532 46310
rect 24492 45416 24544 45422
rect 24492 45358 24544 45364
rect 24320 44526 24440 44554
rect 24308 44396 24360 44402
rect 24308 44338 24360 44344
rect 24216 43784 24268 43790
rect 24216 43726 24268 43732
rect 24216 43648 24268 43654
rect 24216 43590 24268 43596
rect 24124 43376 24176 43382
rect 24228 43364 24256 43590
rect 24176 43336 24256 43364
rect 24124 43318 24176 43324
rect 24124 42900 24176 42906
rect 24124 42842 24176 42848
rect 24032 42832 24084 42838
rect 24032 42774 24084 42780
rect 23848 41812 23900 41818
rect 23848 41754 23900 41760
rect 24136 41698 24164 42842
rect 24228 42294 24256 43336
rect 24216 42288 24268 42294
rect 24216 42230 24268 42236
rect 24228 42022 24256 42230
rect 24216 42016 24268 42022
rect 24216 41958 24268 41964
rect 24044 41670 24164 41698
rect 24044 40662 24072 41670
rect 24124 41608 24176 41614
rect 24124 41550 24176 41556
rect 24136 40934 24164 41550
rect 24228 41138 24256 41958
rect 24216 41132 24268 41138
rect 24216 41074 24268 41080
rect 24124 40928 24176 40934
rect 24124 40870 24176 40876
rect 23940 40656 23992 40662
rect 23940 40598 23992 40604
rect 24032 40656 24084 40662
rect 24032 40598 24084 40604
rect 23676 39086 23796 39114
rect 23676 37398 23704 39086
rect 23952 38654 23980 40598
rect 24032 40520 24084 40526
rect 24032 40462 24084 40468
rect 24044 39137 24072 40462
rect 24136 40089 24164 40870
rect 24216 40520 24268 40526
rect 24216 40462 24268 40468
rect 24122 40080 24178 40089
rect 24122 40015 24178 40024
rect 24030 39128 24086 39137
rect 24030 39063 24086 39072
rect 24032 38752 24084 38758
rect 24032 38694 24084 38700
rect 23768 38626 23980 38654
rect 23664 37392 23716 37398
rect 23664 37334 23716 37340
rect 23664 36032 23716 36038
rect 23664 35974 23716 35980
rect 23676 35494 23704 35974
rect 23664 35488 23716 35494
rect 23664 35430 23716 35436
rect 23572 34604 23624 34610
rect 23572 34546 23624 34552
rect 23572 34400 23624 34406
rect 23572 34342 23624 34348
rect 23480 33584 23532 33590
rect 23584 33561 23612 34342
rect 23768 33946 23796 38626
rect 24044 38418 24072 38694
rect 24032 38412 24084 38418
rect 24032 38354 24084 38360
rect 24228 38010 24256 40462
rect 24320 38457 24348 44338
rect 24412 41449 24440 44526
rect 24504 44033 24532 45358
rect 24596 44849 24624 46446
rect 24582 44840 24638 44849
rect 24582 44775 24638 44784
rect 24584 44328 24636 44334
rect 24584 44270 24636 44276
rect 24490 44024 24546 44033
rect 24490 43959 24546 43968
rect 24492 43852 24544 43858
rect 24492 43794 24544 43800
rect 24504 42362 24532 43794
rect 24596 43450 24624 44270
rect 24584 43444 24636 43450
rect 24584 43386 24636 43392
rect 24596 43217 24624 43386
rect 24582 43208 24638 43217
rect 24582 43143 24638 43152
rect 24492 42356 24544 42362
rect 24492 42298 24544 42304
rect 24398 41440 24454 41449
rect 24398 41375 24454 41384
rect 24400 41132 24452 41138
rect 24400 41074 24452 41080
rect 24412 40118 24440 41074
rect 24504 40526 24532 42298
rect 24584 41608 24636 41614
rect 24584 41550 24636 41556
rect 24596 41274 24624 41550
rect 24584 41268 24636 41274
rect 24584 41210 24636 41216
rect 24492 40520 24544 40526
rect 24492 40462 24544 40468
rect 24400 40112 24452 40118
rect 24400 40054 24452 40060
rect 24412 39030 24440 40054
rect 24400 39024 24452 39030
rect 24400 38966 24452 38972
rect 24492 38956 24544 38962
rect 24492 38898 24544 38904
rect 24306 38448 24362 38457
rect 24306 38383 24362 38392
rect 24400 38412 24452 38418
rect 24400 38354 24452 38360
rect 24216 38004 24268 38010
rect 24216 37946 24268 37952
rect 23848 37800 23900 37806
rect 23848 37742 23900 37748
rect 23860 37466 23888 37742
rect 23940 37664 23992 37670
rect 23940 37606 23992 37612
rect 23848 37460 23900 37466
rect 23848 37402 23900 37408
rect 23848 37120 23900 37126
rect 23848 37062 23900 37068
rect 23860 36174 23888 37062
rect 23952 36242 23980 37606
rect 24412 37262 24440 38354
rect 24504 37670 24532 38898
rect 24688 38554 24716 48622
rect 24768 48544 24820 48550
rect 24768 48486 24820 48492
rect 24780 48006 24808 48486
rect 24768 48000 24820 48006
rect 24768 47942 24820 47948
rect 24780 46617 24808 47942
rect 24766 46608 24822 46617
rect 24766 46543 24822 46552
rect 24768 46504 24820 46510
rect 24768 46446 24820 46452
rect 24780 45665 24808 46446
rect 24766 45656 24822 45665
rect 24766 45591 24822 45600
rect 24768 45416 24820 45422
rect 24768 45358 24820 45364
rect 24780 44305 24808 45358
rect 24766 44296 24822 44305
rect 24766 44231 24822 44240
rect 24768 43784 24820 43790
rect 24768 43726 24820 43732
rect 24780 40769 24808 43726
rect 24872 42809 24900 52838
rect 25136 52624 25188 52630
rect 25136 52566 25188 52572
rect 24952 51264 25004 51270
rect 24952 51206 25004 51212
rect 24964 42906 24992 51206
rect 25044 50924 25096 50930
rect 25044 50866 25096 50872
rect 25056 50561 25084 50866
rect 25042 50552 25098 50561
rect 25042 50487 25098 50496
rect 25148 43926 25176 52566
rect 25332 52154 25360 53751
rect 25320 52148 25372 52154
rect 25320 52090 25372 52096
rect 25504 51808 25556 51814
rect 25504 51750 25556 51756
rect 25516 51406 25544 51750
rect 25504 51400 25556 51406
rect 25502 51368 25504 51377
rect 25556 51368 25558 51377
rect 25502 51303 25558 51312
rect 25320 50312 25372 50318
rect 25320 50254 25372 50260
rect 25332 49745 25360 50254
rect 25318 49736 25374 49745
rect 25318 49671 25374 49680
rect 25320 49224 25372 49230
rect 25320 49166 25372 49172
rect 25332 48929 25360 49166
rect 25318 48920 25374 48929
rect 25318 48855 25374 48864
rect 25504 48000 25556 48006
rect 25504 47942 25556 47948
rect 25516 47666 25544 47942
rect 25504 47660 25556 47666
rect 25504 47602 25556 47608
rect 25516 47297 25544 47602
rect 25502 47288 25558 47297
rect 25502 47223 25558 47232
rect 25228 45824 25280 45830
rect 25228 45766 25280 45772
rect 25240 45490 25268 45766
rect 25228 45484 25280 45490
rect 25228 45426 25280 45432
rect 25136 43920 25188 43926
rect 25136 43862 25188 43868
rect 25148 43314 25176 43862
rect 25228 43648 25280 43654
rect 25228 43590 25280 43596
rect 25136 43308 25188 43314
rect 25136 43250 25188 43256
rect 24952 42900 25004 42906
rect 24952 42842 25004 42848
rect 24858 42800 24914 42809
rect 24858 42735 24914 42744
rect 24766 40760 24822 40769
rect 24766 40695 24822 40704
rect 24872 40526 24900 42735
rect 25136 42696 25188 42702
rect 25136 42638 25188 42644
rect 25044 41744 25096 41750
rect 25044 41686 25096 41692
rect 24952 41064 25004 41070
rect 24952 41006 25004 41012
rect 24860 40520 24912 40526
rect 24860 40462 24912 40468
rect 24860 40384 24912 40390
rect 24860 40326 24912 40332
rect 24768 39296 24820 39302
rect 24768 39238 24820 39244
rect 24676 38548 24728 38554
rect 24676 38490 24728 38496
rect 24584 38480 24636 38486
rect 24584 38422 24636 38428
rect 24492 37664 24544 37670
rect 24492 37606 24544 37612
rect 24400 37256 24452 37262
rect 24400 37198 24452 37204
rect 24412 36922 24440 37198
rect 24596 37126 24624 38422
rect 24676 38276 24728 38282
rect 24676 38218 24728 38224
rect 24688 37194 24716 38218
rect 24676 37188 24728 37194
rect 24676 37130 24728 37136
rect 24584 37120 24636 37126
rect 24584 37062 24636 37068
rect 24400 36916 24452 36922
rect 24400 36858 24452 36864
rect 24400 36780 24452 36786
rect 24400 36722 24452 36728
rect 23940 36236 23992 36242
rect 23940 36178 23992 36184
rect 23848 36168 23900 36174
rect 23848 36110 23900 36116
rect 24412 36038 24440 36722
rect 24688 36689 24716 37130
rect 24674 36680 24730 36689
rect 24674 36615 24730 36624
rect 24492 36304 24544 36310
rect 24492 36246 24544 36252
rect 24400 36032 24452 36038
rect 24400 35974 24452 35980
rect 24412 35154 24440 35974
rect 24400 35148 24452 35154
rect 24400 35090 24452 35096
rect 24032 34944 24084 34950
rect 24032 34886 24084 34892
rect 23848 34196 23900 34202
rect 23848 34138 23900 34144
rect 23676 33918 23796 33946
rect 23480 33526 23532 33532
rect 23570 33552 23626 33561
rect 23388 33448 23440 33454
rect 23388 33390 23440 33396
rect 22756 32864 23336 32892
rect 22652 32768 22704 32774
rect 22652 32710 22704 32716
rect 22652 31816 22704 31822
rect 22652 31758 22704 31764
rect 22560 31476 22612 31482
rect 22560 31418 22612 31424
rect 22664 30054 22692 31758
rect 22756 30938 22784 32864
rect 23204 32768 23256 32774
rect 23204 32710 23256 32716
rect 23216 32502 23244 32710
rect 23204 32496 23256 32502
rect 23204 32438 23256 32444
rect 22836 32224 22888 32230
rect 22836 32166 22888 32172
rect 22744 30932 22796 30938
rect 22744 30874 22796 30880
rect 22744 30796 22796 30802
rect 22744 30738 22796 30744
rect 22652 30048 22704 30054
rect 22652 29990 22704 29996
rect 22560 29640 22612 29646
rect 22560 29582 22612 29588
rect 22388 29158 22508 29186
rect 22388 27334 22416 29158
rect 22468 29096 22520 29102
rect 22468 29038 22520 29044
rect 22376 27328 22428 27334
rect 22376 27270 22428 27276
rect 22296 26982 22416 27010
rect 22284 26920 22336 26926
rect 22284 26862 22336 26868
rect 22192 26036 22244 26042
rect 22192 25978 22244 25984
rect 22296 25498 22324 26862
rect 22388 26314 22416 26982
rect 22480 26450 22508 29038
rect 22572 28762 22600 29582
rect 22756 29170 22784 30738
rect 22744 29164 22796 29170
rect 22744 29106 22796 29112
rect 22848 29016 22876 32166
rect 22950 32124 23258 32133
rect 22950 32122 22956 32124
rect 23012 32122 23036 32124
rect 23092 32122 23116 32124
rect 23172 32122 23196 32124
rect 23252 32122 23258 32124
rect 23012 32070 23014 32122
rect 23194 32070 23196 32122
rect 22950 32068 22956 32070
rect 23012 32068 23036 32070
rect 23092 32068 23116 32070
rect 23172 32068 23196 32070
rect 23252 32068 23258 32070
rect 22950 32059 23258 32068
rect 23296 31952 23348 31958
rect 23296 31894 23348 31900
rect 22950 31036 23258 31045
rect 22950 31034 22956 31036
rect 23012 31034 23036 31036
rect 23092 31034 23116 31036
rect 23172 31034 23196 31036
rect 23252 31034 23258 31036
rect 23012 30982 23014 31034
rect 23194 30982 23196 31034
rect 22950 30980 22956 30982
rect 23012 30980 23036 30982
rect 23092 30980 23116 30982
rect 23172 30980 23196 30982
rect 23252 30980 23258 30982
rect 22950 30971 23258 30980
rect 22950 29948 23258 29957
rect 22950 29946 22956 29948
rect 23012 29946 23036 29948
rect 23092 29946 23116 29948
rect 23172 29946 23196 29948
rect 23252 29946 23258 29948
rect 23012 29894 23014 29946
rect 23194 29894 23196 29946
rect 22950 29892 22956 29894
rect 23012 29892 23036 29894
rect 23092 29892 23116 29894
rect 23172 29892 23196 29894
rect 23252 29892 23258 29894
rect 22950 29883 23258 29892
rect 23308 29714 23336 31894
rect 23400 31142 23428 33390
rect 23492 31958 23520 33526
rect 23570 33487 23626 33496
rect 23676 33046 23704 33918
rect 23756 33448 23808 33454
rect 23756 33390 23808 33396
rect 23664 33040 23716 33046
rect 23664 32982 23716 32988
rect 23768 32026 23796 33390
rect 23756 32020 23808 32026
rect 23756 31962 23808 31968
rect 23480 31952 23532 31958
rect 23480 31894 23532 31900
rect 23664 31884 23716 31890
rect 23664 31826 23716 31832
rect 23676 31142 23704 31826
rect 23860 31482 23888 34138
rect 24044 34066 24072 34886
rect 24412 34678 24440 35090
rect 24400 34672 24452 34678
rect 24400 34614 24452 34620
rect 24032 34060 24084 34066
rect 24032 34002 24084 34008
rect 23940 33856 23992 33862
rect 23940 33798 23992 33804
rect 23848 31476 23900 31482
rect 23848 31418 23900 31424
rect 23848 31340 23900 31346
rect 23848 31282 23900 31288
rect 23388 31136 23440 31142
rect 23388 31078 23440 31084
rect 23664 31136 23716 31142
rect 23664 31078 23716 31084
rect 23400 30258 23428 31078
rect 23676 30326 23704 31078
rect 23664 30320 23716 30326
rect 23664 30262 23716 30268
rect 23860 30274 23888 31282
rect 23952 30734 23980 33798
rect 24504 31346 24532 36246
rect 24676 36168 24728 36174
rect 24676 36110 24728 36116
rect 24688 36038 24716 36110
rect 24676 36032 24728 36038
rect 24676 35974 24728 35980
rect 24688 35057 24716 35974
rect 24674 35048 24730 35057
rect 24674 34983 24730 34992
rect 24676 34536 24728 34542
rect 24676 34478 24728 34484
rect 24584 33856 24636 33862
rect 24584 33798 24636 33804
rect 24492 31340 24544 31346
rect 24492 31282 24544 31288
rect 24308 31136 24360 31142
rect 24308 31078 24360 31084
rect 23940 30728 23992 30734
rect 23940 30670 23992 30676
rect 23940 30320 23992 30326
rect 23860 30268 23940 30274
rect 23860 30262 23992 30268
rect 23388 30252 23440 30258
rect 23388 30194 23440 30200
rect 23388 30048 23440 30054
rect 23388 29990 23440 29996
rect 23400 29714 23428 29990
rect 23296 29708 23348 29714
rect 23296 29650 23348 29656
rect 23388 29708 23440 29714
rect 23388 29650 23440 29656
rect 23296 29096 23348 29102
rect 23296 29038 23348 29044
rect 22756 28988 22876 29016
rect 22560 28756 22612 28762
rect 22560 28698 22612 28704
rect 22560 28144 22612 28150
rect 22560 28086 22612 28092
rect 22468 26444 22520 26450
rect 22468 26386 22520 26392
rect 22572 26314 22600 28086
rect 22652 27532 22704 27538
rect 22652 27474 22704 27480
rect 22664 27402 22692 27474
rect 22652 27396 22704 27402
rect 22652 27338 22704 27344
rect 22664 27130 22692 27338
rect 22652 27124 22704 27130
rect 22652 27066 22704 27072
rect 22756 26382 22784 28988
rect 22950 28860 23258 28869
rect 22950 28858 22956 28860
rect 23012 28858 23036 28860
rect 23092 28858 23116 28860
rect 23172 28858 23196 28860
rect 23252 28858 23258 28860
rect 23012 28806 23014 28858
rect 23194 28806 23196 28858
rect 22950 28804 22956 28806
rect 23012 28804 23036 28806
rect 23092 28804 23116 28806
rect 23172 28804 23196 28806
rect 23252 28804 23258 28806
rect 22950 28795 23258 28804
rect 22836 27872 22888 27878
rect 22836 27814 22888 27820
rect 22848 27402 22876 27814
rect 22950 27772 23258 27781
rect 22950 27770 22956 27772
rect 23012 27770 23036 27772
rect 23092 27770 23116 27772
rect 23172 27770 23196 27772
rect 23252 27770 23258 27772
rect 23012 27718 23014 27770
rect 23194 27718 23196 27770
rect 22950 27716 22956 27718
rect 23012 27716 23036 27718
rect 23092 27716 23116 27718
rect 23172 27716 23196 27718
rect 23252 27716 23258 27718
rect 22950 27707 23258 27716
rect 23308 27538 23336 29038
rect 23676 28626 23704 30262
rect 23860 30246 23980 30262
rect 23664 28620 23716 28626
rect 23664 28562 23716 28568
rect 23756 28416 23808 28422
rect 23756 28358 23808 28364
rect 23768 28218 23796 28358
rect 23756 28212 23808 28218
rect 23756 28154 23808 28160
rect 23860 27878 23888 30246
rect 23940 29844 23992 29850
rect 23940 29786 23992 29792
rect 23952 29306 23980 29786
rect 23940 29300 23992 29306
rect 23940 29242 23992 29248
rect 24124 29164 24176 29170
rect 24124 29106 24176 29112
rect 23848 27872 23900 27878
rect 23848 27814 23900 27820
rect 24136 27713 24164 29106
rect 24122 27704 24178 27713
rect 24122 27639 24178 27648
rect 23296 27532 23348 27538
rect 23296 27474 23348 27480
rect 22836 27396 22888 27402
rect 22836 27338 22888 27344
rect 22848 27062 22876 27338
rect 22836 27056 22888 27062
rect 22836 26998 22888 27004
rect 22848 26926 22876 26998
rect 22836 26920 22888 26926
rect 22836 26862 22888 26868
rect 22836 26784 22888 26790
rect 22836 26726 22888 26732
rect 22744 26376 22796 26382
rect 22744 26318 22796 26324
rect 22376 26308 22428 26314
rect 22376 26250 22428 26256
rect 22560 26308 22612 26314
rect 22560 26250 22612 26256
rect 22468 26240 22520 26246
rect 22468 26182 22520 26188
rect 22376 25696 22428 25702
rect 22376 25638 22428 25644
rect 22284 25492 22336 25498
rect 22284 25434 22336 25440
rect 22112 25214 22324 25242
rect 22100 25152 22152 25158
rect 22100 25094 22152 25100
rect 22112 24750 22140 25094
rect 22100 24744 22152 24750
rect 22100 24686 22152 24692
rect 21916 24268 21968 24274
rect 21916 24210 21968 24216
rect 21836 24126 21956 24154
rect 21732 24064 21784 24070
rect 21732 24006 21784 24012
rect 21640 23860 21692 23866
rect 21640 23802 21692 23808
rect 21652 23322 21680 23802
rect 21640 23316 21692 23322
rect 21640 23258 21692 23264
rect 21652 21962 21680 23258
rect 21640 21956 21692 21962
rect 21640 21898 21692 21904
rect 21652 21146 21680 21898
rect 21640 21140 21692 21146
rect 21640 21082 21692 21088
rect 21652 20942 21680 21082
rect 21640 20936 21692 20942
rect 21640 20878 21692 20884
rect 21640 20800 21692 20806
rect 21640 20742 21692 20748
rect 21652 20466 21680 20742
rect 21640 20460 21692 20466
rect 21640 20402 21692 20408
rect 21744 19666 21772 24006
rect 21824 21344 21876 21350
rect 21824 21286 21876 21292
rect 21652 19638 21772 19666
rect 21548 18828 21600 18834
rect 21548 18770 21600 18776
rect 21456 17876 21508 17882
rect 21456 17818 21508 17824
rect 21468 17134 21496 17818
rect 21456 17128 21508 17134
rect 21456 17070 21508 17076
rect 21364 16176 21416 16182
rect 21364 16118 21416 16124
rect 21272 16108 21324 16114
rect 21272 16050 21324 16056
rect 20996 16040 21048 16046
rect 20996 15982 21048 15988
rect 20996 15700 21048 15706
rect 20996 15642 21048 15648
rect 20904 14408 20956 14414
rect 20904 14350 20956 14356
rect 20812 13456 20864 13462
rect 20812 13398 20864 13404
rect 20536 13252 20588 13258
rect 20536 13194 20588 13200
rect 20352 12912 20404 12918
rect 20352 12854 20404 12860
rect 20364 12646 20392 12854
rect 20352 12640 20404 12646
rect 20352 12582 20404 12588
rect 20260 11824 20312 11830
rect 20260 11766 20312 11772
rect 20364 11762 20392 12582
rect 20352 11756 20404 11762
rect 20352 11698 20404 11704
rect 20444 8356 20496 8362
rect 20444 8298 20496 8304
rect 20260 7744 20312 7750
rect 20260 7686 20312 7692
rect 20272 6322 20300 7686
rect 20456 7478 20484 8298
rect 20444 7472 20496 7478
rect 20444 7414 20496 7420
rect 20260 6316 20312 6322
rect 20260 6258 20312 6264
rect 20444 5772 20496 5778
rect 20444 5714 20496 5720
rect 19984 4140 20036 4146
rect 19984 4082 20036 4088
rect 20076 4072 20128 4078
rect 20076 4014 20128 4020
rect 19892 2848 19944 2854
rect 19892 2790 19944 2796
rect 20088 800 20116 4014
rect 20456 800 20484 5714
rect 20548 5710 20576 13194
rect 20812 13184 20864 13190
rect 20812 13126 20864 13132
rect 20628 12776 20680 12782
rect 20628 12718 20680 12724
rect 20640 11898 20668 12718
rect 20720 12640 20772 12646
rect 20720 12582 20772 12588
rect 20628 11892 20680 11898
rect 20628 11834 20680 11840
rect 20732 10674 20760 12582
rect 20824 12102 20852 13126
rect 20916 12306 20944 14350
rect 21008 12434 21036 15642
rect 21180 15632 21232 15638
rect 21180 15574 21232 15580
rect 21088 15360 21140 15366
rect 21088 15302 21140 15308
rect 21100 15094 21128 15302
rect 21088 15088 21140 15094
rect 21088 15030 21140 15036
rect 21192 12986 21220 15574
rect 21284 15570 21312 16050
rect 21548 15904 21600 15910
rect 21548 15846 21600 15852
rect 21272 15564 21324 15570
rect 21272 15506 21324 15512
rect 21364 15360 21416 15366
rect 21364 15302 21416 15308
rect 21180 12980 21232 12986
rect 21180 12922 21232 12928
rect 21008 12406 21128 12434
rect 20904 12300 20956 12306
rect 20904 12242 20956 12248
rect 20812 12096 20864 12102
rect 20812 12038 20864 12044
rect 21100 11082 21128 12406
rect 21180 12164 21232 12170
rect 21180 12106 21232 12112
rect 21192 11898 21220 12106
rect 21180 11892 21232 11898
rect 21180 11834 21232 11840
rect 21192 11762 21220 11834
rect 21180 11756 21232 11762
rect 21180 11698 21232 11704
rect 21088 11076 21140 11082
rect 21088 11018 21140 11024
rect 21100 10810 21128 11018
rect 21088 10804 21140 10810
rect 21088 10746 21140 10752
rect 20720 10668 20772 10674
rect 20720 10610 20772 10616
rect 20628 10532 20680 10538
rect 20628 10474 20680 10480
rect 20640 9586 20668 10474
rect 21180 10464 21232 10470
rect 21180 10406 21232 10412
rect 20628 9580 20680 9586
rect 20628 9522 20680 9528
rect 21192 7886 21220 10406
rect 21376 8566 21404 15302
rect 21456 15156 21508 15162
rect 21456 15098 21508 15104
rect 21468 14822 21496 15098
rect 21456 14816 21508 14822
rect 21456 14758 21508 14764
rect 21560 12306 21588 15846
rect 21652 15502 21680 19638
rect 21732 19508 21784 19514
rect 21732 19450 21784 19456
rect 21744 19310 21772 19450
rect 21732 19304 21784 19310
rect 21732 19246 21784 19252
rect 21744 18766 21772 19246
rect 21732 18760 21784 18766
rect 21732 18702 21784 18708
rect 21744 18222 21772 18702
rect 21732 18216 21784 18222
rect 21732 18158 21784 18164
rect 21744 17678 21772 18158
rect 21732 17672 21784 17678
rect 21732 17614 21784 17620
rect 21744 16658 21772 17614
rect 21732 16652 21784 16658
rect 21732 16594 21784 16600
rect 21640 15496 21692 15502
rect 21640 15438 21692 15444
rect 21836 15026 21864 21286
rect 21928 19242 21956 24126
rect 22100 23724 22152 23730
rect 22100 23666 22152 23672
rect 22112 22574 22140 23666
rect 22100 22568 22152 22574
rect 22100 22510 22152 22516
rect 22112 22234 22140 22510
rect 22100 22228 22152 22234
rect 22100 22170 22152 22176
rect 22296 20466 22324 25214
rect 22388 24206 22416 25638
rect 22376 24200 22428 24206
rect 22376 24142 22428 24148
rect 22480 21690 22508 26182
rect 22558 26072 22614 26081
rect 22558 26007 22614 26016
rect 22572 24818 22600 26007
rect 22560 24812 22612 24818
rect 22560 24754 22612 24760
rect 22848 24750 22876 26726
rect 22950 26684 23258 26693
rect 22950 26682 22956 26684
rect 23012 26682 23036 26684
rect 23092 26682 23116 26684
rect 23172 26682 23196 26684
rect 23252 26682 23258 26684
rect 23012 26630 23014 26682
rect 23194 26630 23196 26682
rect 22950 26628 22956 26630
rect 23012 26628 23036 26630
rect 23092 26628 23116 26630
rect 23172 26628 23196 26630
rect 23252 26628 23258 26630
rect 22950 26619 23258 26628
rect 23308 25922 23336 27474
rect 24320 27062 24348 31078
rect 24492 30592 24544 30598
rect 24492 30534 24544 30540
rect 24308 27056 24360 27062
rect 24308 26998 24360 27004
rect 23386 26888 23442 26897
rect 23386 26823 23442 26832
rect 23400 25974 23428 26823
rect 24032 26444 24084 26450
rect 24032 26386 24084 26392
rect 23216 25894 23336 25922
rect 23388 25968 23440 25974
rect 23388 25910 23440 25916
rect 23216 25838 23244 25894
rect 23204 25832 23256 25838
rect 23204 25774 23256 25780
rect 22950 25596 23258 25605
rect 22950 25594 22956 25596
rect 23012 25594 23036 25596
rect 23092 25594 23116 25596
rect 23172 25594 23196 25596
rect 23252 25594 23258 25596
rect 23012 25542 23014 25594
rect 23194 25542 23196 25594
rect 22950 25540 22956 25542
rect 23012 25540 23036 25542
rect 23092 25540 23116 25542
rect 23172 25540 23196 25542
rect 23252 25540 23258 25542
rect 22950 25531 23258 25540
rect 23308 24886 23336 25894
rect 23572 25424 23624 25430
rect 23572 25366 23624 25372
rect 23296 24880 23348 24886
rect 23296 24822 23348 24828
rect 22836 24744 22888 24750
rect 22836 24686 22888 24692
rect 22652 24064 22704 24070
rect 22652 24006 22704 24012
rect 22468 21684 22520 21690
rect 22468 21626 22520 21632
rect 22560 21140 22612 21146
rect 22560 21082 22612 21088
rect 22284 20460 22336 20466
rect 22284 20402 22336 20408
rect 22192 19712 22244 19718
rect 22192 19654 22244 19660
rect 22008 19508 22060 19514
rect 22008 19450 22060 19456
rect 21916 19236 21968 19242
rect 21916 19178 21968 19184
rect 21928 18970 21956 19178
rect 21916 18964 21968 18970
rect 21916 18906 21968 18912
rect 22020 18834 22048 19450
rect 22008 18828 22060 18834
rect 22008 18770 22060 18776
rect 22020 17202 22048 18770
rect 22204 17746 22232 19654
rect 22572 19446 22600 21082
rect 22664 19718 22692 24006
rect 22744 23792 22796 23798
rect 22744 23734 22796 23740
rect 22756 23662 22784 23734
rect 22848 23730 22876 24686
rect 22950 24508 23258 24517
rect 22950 24506 22956 24508
rect 23012 24506 23036 24508
rect 23092 24506 23116 24508
rect 23172 24506 23196 24508
rect 23252 24506 23258 24508
rect 23012 24454 23014 24506
rect 23194 24454 23196 24506
rect 22950 24452 22956 24454
rect 23012 24452 23036 24454
rect 23092 24452 23116 24454
rect 23172 24452 23196 24454
rect 23252 24452 23258 24454
rect 22950 24443 23258 24452
rect 23480 24336 23532 24342
rect 23480 24278 23532 24284
rect 22836 23724 22888 23730
rect 22836 23666 22888 23672
rect 22744 23656 22796 23662
rect 22744 23598 22796 23604
rect 22756 22098 22784 23598
rect 22950 23420 23258 23429
rect 22950 23418 22956 23420
rect 23012 23418 23036 23420
rect 23092 23418 23116 23420
rect 23172 23418 23196 23420
rect 23252 23418 23258 23420
rect 23012 23366 23014 23418
rect 23194 23366 23196 23418
rect 22950 23364 22956 23366
rect 23012 23364 23036 23366
rect 23092 23364 23116 23366
rect 23172 23364 23196 23366
rect 23252 23364 23258 23366
rect 22950 23355 23258 23364
rect 23492 23254 23520 24278
rect 23584 24206 23612 25366
rect 23940 25152 23992 25158
rect 23940 25094 23992 25100
rect 23664 24948 23716 24954
rect 23664 24890 23716 24896
rect 23572 24200 23624 24206
rect 23572 24142 23624 24148
rect 23676 23798 23704 24890
rect 23756 24608 23808 24614
rect 23756 24550 23808 24556
rect 23768 24274 23796 24550
rect 23756 24268 23808 24274
rect 23756 24210 23808 24216
rect 23664 23792 23716 23798
rect 23664 23734 23716 23740
rect 23664 23656 23716 23662
rect 23664 23598 23716 23604
rect 23846 23624 23902 23633
rect 23480 23248 23532 23254
rect 23480 23190 23532 23196
rect 23572 22976 23624 22982
rect 23572 22918 23624 22924
rect 23294 22808 23350 22817
rect 23294 22743 23350 22752
rect 22950 22332 23258 22341
rect 22950 22330 22956 22332
rect 23012 22330 23036 22332
rect 23092 22330 23116 22332
rect 23172 22330 23196 22332
rect 23252 22330 23258 22332
rect 23012 22278 23014 22330
rect 23194 22278 23196 22330
rect 22950 22276 22956 22278
rect 23012 22276 23036 22278
rect 23092 22276 23116 22278
rect 23172 22276 23196 22278
rect 23252 22276 23258 22278
rect 22950 22267 23258 22276
rect 23204 22228 23256 22234
rect 23204 22170 23256 22176
rect 22744 22092 22796 22098
rect 22744 22034 22796 22040
rect 23216 21554 23244 22170
rect 23204 21548 23256 21554
rect 23204 21490 23256 21496
rect 22950 21244 23258 21253
rect 22950 21242 22956 21244
rect 23012 21242 23036 21244
rect 23092 21242 23116 21244
rect 23172 21242 23196 21244
rect 23252 21242 23258 21244
rect 23012 21190 23014 21242
rect 23194 21190 23196 21242
rect 22950 21188 22956 21190
rect 23012 21188 23036 21190
rect 23092 21188 23116 21190
rect 23172 21188 23196 21190
rect 23252 21188 23258 21190
rect 22950 21179 23258 21188
rect 23308 20398 23336 22743
rect 23388 22024 23440 22030
rect 23388 21966 23440 21972
rect 23400 21690 23428 21966
rect 23388 21684 23440 21690
rect 23388 21626 23440 21632
rect 23584 21350 23612 22918
rect 23572 21344 23624 21350
rect 23572 21286 23624 21292
rect 23386 21176 23442 21185
rect 23386 21111 23442 21120
rect 23400 20534 23428 21111
rect 23388 20528 23440 20534
rect 23388 20470 23440 20476
rect 23296 20392 23348 20398
rect 23296 20334 23348 20340
rect 22836 20324 22888 20330
rect 22836 20266 22888 20272
rect 22744 19780 22796 19786
rect 22744 19722 22796 19728
rect 22652 19712 22704 19718
rect 22652 19654 22704 19660
rect 22560 19440 22612 19446
rect 22560 19382 22612 19388
rect 22572 19334 22600 19382
rect 22572 19310 22692 19334
rect 22572 19306 22704 19310
rect 22652 19304 22704 19306
rect 22652 19246 22704 19252
rect 22284 18896 22336 18902
rect 22284 18838 22336 18844
rect 22192 17740 22244 17746
rect 22192 17682 22244 17688
rect 22296 17626 22324 18838
rect 22296 17598 22600 17626
rect 22192 17264 22244 17270
rect 22192 17206 22244 17212
rect 22008 17196 22060 17202
rect 22008 17138 22060 17144
rect 22008 16992 22060 16998
rect 22008 16934 22060 16940
rect 22020 16658 22048 16934
rect 22008 16652 22060 16658
rect 22008 16594 22060 16600
rect 22204 16250 22232 17206
rect 22468 16652 22520 16658
rect 22468 16594 22520 16600
rect 22480 16250 22508 16594
rect 22192 16244 22244 16250
rect 22192 16186 22244 16192
rect 22468 16244 22520 16250
rect 22468 16186 22520 16192
rect 22284 15360 22336 15366
rect 22284 15302 22336 15308
rect 21824 15020 21876 15026
rect 21824 14962 21876 14968
rect 21916 15020 21968 15026
rect 21916 14962 21968 14968
rect 21928 14618 21956 14962
rect 22192 14952 22244 14958
rect 22192 14894 22244 14900
rect 21916 14612 21968 14618
rect 21916 14554 21968 14560
rect 22100 14272 22152 14278
rect 22100 14214 22152 14220
rect 21916 14068 21968 14074
rect 21916 14010 21968 14016
rect 21548 12300 21600 12306
rect 21548 12242 21600 12248
rect 21824 12232 21876 12238
rect 21824 12174 21876 12180
rect 21836 11830 21864 12174
rect 21824 11824 21876 11830
rect 21824 11766 21876 11772
rect 21732 11348 21784 11354
rect 21732 11290 21784 11296
rect 21744 11150 21772 11290
rect 21732 11144 21784 11150
rect 21732 11086 21784 11092
rect 21928 10062 21956 14010
rect 22112 13326 22140 14214
rect 22100 13320 22152 13326
rect 22100 13262 22152 13268
rect 22008 12776 22060 12782
rect 22112 12730 22140 13262
rect 22204 12850 22232 14894
rect 22296 14482 22324 15302
rect 22284 14476 22336 14482
rect 22284 14418 22336 14424
rect 22572 13938 22600 17598
rect 22652 16516 22704 16522
rect 22652 16458 22704 16464
rect 22664 16250 22692 16458
rect 22652 16244 22704 16250
rect 22652 16186 22704 16192
rect 22664 14822 22692 16186
rect 22756 15502 22784 19722
rect 22848 17270 22876 20266
rect 22950 20156 23258 20165
rect 22950 20154 22956 20156
rect 23012 20154 23036 20156
rect 23092 20154 23116 20156
rect 23172 20154 23196 20156
rect 23252 20154 23258 20156
rect 23012 20102 23014 20154
rect 23194 20102 23196 20154
rect 22950 20100 22956 20102
rect 23012 20100 23036 20102
rect 23092 20100 23116 20102
rect 23172 20100 23196 20102
rect 23252 20100 23258 20102
rect 22950 20091 23258 20100
rect 23572 19304 23624 19310
rect 23572 19246 23624 19252
rect 22950 19068 23258 19077
rect 22950 19066 22956 19068
rect 23012 19066 23036 19068
rect 23092 19066 23116 19068
rect 23172 19066 23196 19068
rect 23252 19066 23258 19068
rect 23012 19014 23014 19066
rect 23194 19014 23196 19066
rect 22950 19012 22956 19014
rect 23012 19012 23036 19014
rect 23092 19012 23116 19014
rect 23172 19012 23196 19014
rect 23252 19012 23258 19014
rect 22950 19003 23258 19012
rect 23584 18698 23612 19246
rect 23572 18692 23624 18698
rect 23572 18634 23624 18640
rect 23388 18216 23440 18222
rect 23388 18158 23440 18164
rect 22950 17980 23258 17989
rect 22950 17978 22956 17980
rect 23012 17978 23036 17980
rect 23092 17978 23116 17980
rect 23172 17978 23196 17980
rect 23252 17978 23258 17980
rect 23012 17926 23014 17978
rect 23194 17926 23196 17978
rect 22950 17924 22956 17926
rect 23012 17924 23036 17926
rect 23092 17924 23116 17926
rect 23172 17924 23196 17926
rect 23252 17924 23258 17926
rect 22950 17915 23258 17924
rect 23400 17921 23428 18158
rect 23386 17912 23442 17921
rect 23386 17847 23442 17856
rect 23584 17814 23612 18634
rect 23676 18290 23704 23598
rect 23846 23559 23902 23568
rect 23860 23118 23888 23559
rect 23848 23112 23900 23118
rect 23848 23054 23900 23060
rect 23664 18284 23716 18290
rect 23664 18226 23716 18232
rect 23664 17876 23716 17882
rect 23664 17818 23716 17824
rect 23572 17808 23624 17814
rect 23572 17750 23624 17756
rect 22836 17264 22888 17270
rect 22836 17206 22888 17212
rect 23388 17060 23440 17066
rect 23388 17002 23440 17008
rect 22950 16892 23258 16901
rect 22950 16890 22956 16892
rect 23012 16890 23036 16892
rect 23092 16890 23116 16892
rect 23172 16890 23196 16892
rect 23252 16890 23258 16892
rect 23012 16838 23014 16890
rect 23194 16838 23196 16890
rect 22950 16836 22956 16838
rect 23012 16836 23036 16838
rect 23092 16836 23116 16838
rect 23172 16836 23196 16838
rect 23252 16836 23258 16838
rect 22950 16827 23258 16836
rect 22950 15804 23258 15813
rect 22950 15802 22956 15804
rect 23012 15802 23036 15804
rect 23092 15802 23116 15804
rect 23172 15802 23196 15804
rect 23252 15802 23258 15804
rect 23012 15750 23014 15802
rect 23194 15750 23196 15802
rect 22950 15748 22956 15750
rect 23012 15748 23036 15750
rect 23092 15748 23116 15750
rect 23172 15748 23196 15750
rect 23252 15748 23258 15750
rect 22950 15739 23258 15748
rect 22744 15496 22796 15502
rect 22744 15438 22796 15444
rect 22744 14884 22796 14890
rect 22744 14826 22796 14832
rect 22652 14816 22704 14822
rect 22652 14758 22704 14764
rect 22664 14346 22692 14758
rect 22652 14340 22704 14346
rect 22652 14282 22704 14288
rect 22560 13932 22612 13938
rect 22560 13874 22612 13880
rect 22192 12844 22244 12850
rect 22192 12786 22244 12792
rect 22060 12724 22140 12730
rect 22008 12718 22140 12724
rect 22020 12702 22140 12718
rect 22100 12640 22152 12646
rect 22100 12582 22152 12588
rect 22008 12096 22060 12102
rect 22008 12038 22060 12044
rect 21916 10056 21968 10062
rect 21916 9998 21968 10004
rect 21824 9920 21876 9926
rect 21824 9862 21876 9868
rect 21364 8560 21416 8566
rect 21364 8502 21416 8508
rect 21272 8356 21324 8362
rect 21272 8298 21324 8304
rect 21180 7880 21232 7886
rect 21180 7822 21232 7828
rect 20720 7404 20772 7410
rect 20720 7346 20772 7352
rect 20628 7200 20680 7206
rect 20628 7142 20680 7148
rect 20640 5710 20668 7142
rect 20732 5914 20760 7346
rect 20720 5908 20772 5914
rect 20720 5850 20772 5856
rect 20536 5704 20588 5710
rect 20536 5646 20588 5652
rect 20628 5704 20680 5710
rect 20628 5646 20680 5652
rect 20720 4684 20772 4690
rect 20720 4626 20772 4632
rect 20628 4548 20680 4554
rect 20628 4490 20680 4496
rect 20640 2990 20668 4490
rect 20628 2984 20680 2990
rect 20628 2926 20680 2932
rect 20732 2922 20760 4626
rect 21284 4622 21312 8298
rect 21640 7336 21692 7342
rect 21640 7278 21692 7284
rect 21548 5772 21600 5778
rect 21548 5714 21600 5720
rect 21272 4616 21324 4622
rect 21272 4558 21324 4564
rect 21180 4004 21232 4010
rect 21180 3946 21232 3952
rect 20720 2916 20772 2922
rect 20720 2858 20772 2864
rect 20812 2848 20864 2854
rect 20812 2790 20864 2796
rect 20824 800 20852 2790
rect 21192 800 21220 3946
rect 21560 800 21588 5714
rect 21652 2417 21680 7278
rect 21732 6248 21784 6254
rect 21732 6190 21784 6196
rect 21744 3058 21772 6190
rect 21836 5642 21864 9862
rect 22020 9654 22048 12038
rect 22008 9648 22060 9654
rect 22008 9590 22060 9596
rect 22008 6724 22060 6730
rect 22008 6666 22060 6672
rect 21916 6248 21968 6254
rect 21916 6190 21968 6196
rect 21824 5636 21876 5642
rect 21824 5578 21876 5584
rect 21732 3052 21784 3058
rect 21732 2994 21784 3000
rect 21638 2408 21694 2417
rect 21638 2343 21694 2352
rect 21928 800 21956 6190
rect 22020 3398 22048 6666
rect 22112 5234 22140 12582
rect 22664 12102 22692 14282
rect 22652 12096 22704 12102
rect 22652 12038 22704 12044
rect 22664 11642 22692 12038
rect 22756 11762 22784 14826
rect 22950 14716 23258 14725
rect 22950 14714 22956 14716
rect 23012 14714 23036 14716
rect 23092 14714 23116 14716
rect 23172 14714 23196 14716
rect 23252 14714 23258 14716
rect 23012 14662 23014 14714
rect 23194 14662 23196 14714
rect 22950 14660 22956 14662
rect 23012 14660 23036 14662
rect 23092 14660 23116 14662
rect 23172 14660 23196 14662
rect 23252 14660 23258 14662
rect 22950 14651 23258 14660
rect 22836 14068 22888 14074
rect 22836 14010 22888 14016
rect 22744 11756 22796 11762
rect 22744 11698 22796 11704
rect 22664 11614 22784 11642
rect 22192 11280 22244 11286
rect 22192 11222 22244 11228
rect 22204 6322 22232 11222
rect 22560 10464 22612 10470
rect 22560 10406 22612 10412
rect 22376 8492 22428 8498
rect 22376 8434 22428 8440
rect 22284 7336 22336 7342
rect 22284 7278 22336 7284
rect 22192 6316 22244 6322
rect 22192 6258 22244 6264
rect 22192 6180 22244 6186
rect 22192 6122 22244 6128
rect 22100 5228 22152 5234
rect 22100 5170 22152 5176
rect 22098 4040 22154 4049
rect 22098 3975 22154 3984
rect 22112 3942 22140 3975
rect 22100 3936 22152 3942
rect 22100 3878 22152 3884
rect 22204 3466 22232 6122
rect 22192 3460 22244 3466
rect 22192 3402 22244 3408
rect 22008 3392 22060 3398
rect 22008 3334 22060 3340
rect 22296 800 22324 7278
rect 22388 4826 22416 8434
rect 22468 5160 22520 5166
rect 22468 5102 22520 5108
rect 22376 4820 22428 4826
rect 22376 4762 22428 4768
rect 22480 2854 22508 5102
rect 22572 4690 22600 10406
rect 22652 10056 22704 10062
rect 22652 9998 22704 10004
rect 22664 9722 22692 9998
rect 22652 9716 22704 9722
rect 22652 9658 22704 9664
rect 22756 9602 22784 11614
rect 22848 10062 22876 14010
rect 22950 13628 23258 13637
rect 22950 13626 22956 13628
rect 23012 13626 23036 13628
rect 23092 13626 23116 13628
rect 23172 13626 23196 13628
rect 23252 13626 23258 13628
rect 23012 13574 23014 13626
rect 23194 13574 23196 13626
rect 22950 13572 22956 13574
rect 23012 13572 23036 13574
rect 23092 13572 23116 13574
rect 23172 13572 23196 13574
rect 23252 13572 23258 13574
rect 22950 13563 23258 13572
rect 23400 12850 23428 17002
rect 23676 16046 23704 17818
rect 23952 17202 23980 25094
rect 24044 23866 24072 26386
rect 24124 25900 24176 25906
rect 24124 25842 24176 25848
rect 24032 23860 24084 23866
rect 24032 23802 24084 23808
rect 24136 22778 24164 25842
rect 24504 25294 24532 30534
rect 24596 29238 24624 33798
rect 24584 29232 24636 29238
rect 24584 29174 24636 29180
rect 24688 28150 24716 34478
rect 24780 33998 24808 39238
rect 24872 38894 24900 40326
rect 24860 38888 24912 38894
rect 24860 38830 24912 38836
rect 24860 38752 24912 38758
rect 24860 38694 24912 38700
rect 24872 37942 24900 38694
rect 24964 37992 24992 41006
rect 25056 39506 25084 41686
rect 25148 39506 25176 42638
rect 25240 41206 25268 43590
rect 25596 43308 25648 43314
rect 25596 43250 25648 43256
rect 25412 43172 25464 43178
rect 25412 43114 25464 43120
rect 25320 43104 25372 43110
rect 25320 43046 25372 43052
rect 25332 42702 25360 43046
rect 25320 42696 25372 42702
rect 25320 42638 25372 42644
rect 25228 41200 25280 41206
rect 25228 41142 25280 41148
rect 25320 41132 25372 41138
rect 25320 41074 25372 41080
rect 25228 39976 25280 39982
rect 25228 39918 25280 39924
rect 25044 39500 25096 39506
rect 25044 39442 25096 39448
rect 25136 39500 25188 39506
rect 25136 39442 25188 39448
rect 25240 39098 25268 39918
rect 25332 39914 25360 41074
rect 25320 39908 25372 39914
rect 25320 39850 25372 39856
rect 25228 39092 25280 39098
rect 25228 39034 25280 39040
rect 25332 38321 25360 39850
rect 25424 38350 25452 43114
rect 25504 40928 25556 40934
rect 25504 40870 25556 40876
rect 25412 38344 25464 38350
rect 25318 38312 25374 38321
rect 25412 38286 25464 38292
rect 25318 38247 25374 38256
rect 24964 37964 25084 37992
rect 24860 37936 24912 37942
rect 24860 37878 24912 37884
rect 24872 36922 24900 37878
rect 25056 37262 25084 37964
rect 24952 37256 25004 37262
rect 24952 37198 25004 37204
rect 25044 37256 25096 37262
rect 25044 37198 25096 37204
rect 24964 37074 24992 37198
rect 24964 37046 25084 37074
rect 24860 36916 24912 36922
rect 24860 36858 24912 36864
rect 24860 36780 24912 36786
rect 24860 36722 24912 36728
rect 24872 36038 24900 36722
rect 25056 36378 25084 37046
rect 25044 36372 25096 36378
rect 25044 36314 25096 36320
rect 24860 36032 24912 36038
rect 24860 35974 24912 35980
rect 24872 35873 24900 35974
rect 24858 35864 24914 35873
rect 24858 35799 24914 35808
rect 24768 33992 24820 33998
rect 24768 33934 24820 33940
rect 25056 33658 25084 36314
rect 25516 36242 25544 40870
rect 25608 38214 25636 43250
rect 25596 38208 25648 38214
rect 25596 38150 25648 38156
rect 25504 36236 25556 36242
rect 25504 36178 25556 36184
rect 25136 36032 25188 36038
rect 25136 35974 25188 35980
rect 25044 33652 25096 33658
rect 25044 33594 25096 33600
rect 24860 33516 24912 33522
rect 24860 33458 24912 33464
rect 24872 31754 24900 33458
rect 24872 31726 24992 31754
rect 24964 31142 24992 31726
rect 24952 31136 25004 31142
rect 24952 31078 25004 31084
rect 24964 30394 24992 31078
rect 25148 30802 25176 35974
rect 25412 35760 25464 35766
rect 25412 35702 25464 35708
rect 25228 35624 25280 35630
rect 25228 35566 25280 35572
rect 25240 35290 25268 35566
rect 25424 35494 25452 35702
rect 25412 35488 25464 35494
rect 25412 35430 25464 35436
rect 25228 35284 25280 35290
rect 25228 35226 25280 35232
rect 25424 34678 25452 35430
rect 25412 34672 25464 34678
rect 25412 34614 25464 34620
rect 25320 34604 25372 34610
rect 25320 34546 25372 34552
rect 25332 34241 25360 34546
rect 25318 34232 25374 34241
rect 25424 34202 25452 34614
rect 25318 34167 25320 34176
rect 25372 34167 25374 34176
rect 25412 34196 25464 34202
rect 25320 34138 25372 34144
rect 25412 34138 25464 34144
rect 25410 33416 25466 33425
rect 25410 33351 25466 33360
rect 25320 32904 25372 32910
rect 25320 32846 25372 32852
rect 25332 32609 25360 32846
rect 25318 32600 25374 32609
rect 25318 32535 25374 32544
rect 25424 32434 25452 33351
rect 25412 32428 25464 32434
rect 25412 32370 25464 32376
rect 25320 31816 25372 31822
rect 25318 31784 25320 31793
rect 25372 31784 25374 31793
rect 25318 31719 25374 31728
rect 25320 31340 25372 31346
rect 25320 31282 25372 31288
rect 25332 30977 25360 31282
rect 25318 30968 25374 30977
rect 25318 30903 25320 30912
rect 25372 30903 25374 30912
rect 25320 30874 25372 30880
rect 25136 30796 25188 30802
rect 25136 30738 25188 30744
rect 25504 30728 25556 30734
rect 25504 30670 25556 30676
rect 25136 30592 25188 30598
rect 25134 30560 25136 30569
rect 25188 30560 25190 30569
rect 25134 30495 25190 30504
rect 24952 30388 25004 30394
rect 24952 30330 25004 30336
rect 25412 30184 25464 30190
rect 25318 30152 25374 30161
rect 25412 30126 25464 30132
rect 25318 30087 25374 30096
rect 25332 29646 25360 30087
rect 25320 29640 25372 29646
rect 25320 29582 25372 29588
rect 24768 29572 24820 29578
rect 24768 29514 24820 29520
rect 24780 28558 24808 29514
rect 25332 29306 25360 29582
rect 25320 29300 25372 29306
rect 25320 29242 25372 29248
rect 25044 29028 25096 29034
rect 25044 28970 25096 28976
rect 24768 28552 24820 28558
rect 24768 28494 24820 28500
rect 24768 28416 24820 28422
rect 24768 28358 24820 28364
rect 24676 28144 24728 28150
rect 24676 28086 24728 28092
rect 24584 26376 24636 26382
rect 24584 26318 24636 26324
rect 24492 25288 24544 25294
rect 24492 25230 24544 25236
rect 24596 24614 24624 26318
rect 24676 25152 24728 25158
rect 24676 25094 24728 25100
rect 24584 24608 24636 24614
rect 24584 24550 24636 24556
rect 24400 24064 24452 24070
rect 24400 24006 24452 24012
rect 24124 22772 24176 22778
rect 24124 22714 24176 22720
rect 24032 22568 24084 22574
rect 24032 22510 24084 22516
rect 24044 22098 24072 22510
rect 24032 22092 24084 22098
rect 24032 22034 24084 22040
rect 24124 21888 24176 21894
rect 24124 21830 24176 21836
rect 23940 17196 23992 17202
rect 23940 17138 23992 17144
rect 23848 16788 23900 16794
rect 23848 16730 23900 16736
rect 23664 16040 23716 16046
rect 23664 15982 23716 15988
rect 23480 15904 23532 15910
rect 23480 15846 23532 15852
rect 23388 12844 23440 12850
rect 23388 12786 23440 12792
rect 22950 12540 23258 12549
rect 22950 12538 22956 12540
rect 23012 12538 23036 12540
rect 23092 12538 23116 12540
rect 23172 12538 23196 12540
rect 23252 12538 23258 12540
rect 23012 12486 23014 12538
rect 23194 12486 23196 12538
rect 22950 12484 22956 12486
rect 23012 12484 23036 12486
rect 23092 12484 23116 12486
rect 23172 12484 23196 12486
rect 23252 12484 23258 12486
rect 22950 12475 23258 12484
rect 23492 12238 23520 15846
rect 23860 13938 23888 16730
rect 24136 16114 24164 21830
rect 24308 19712 24360 19718
rect 24308 19654 24360 19660
rect 24124 16108 24176 16114
rect 24124 16050 24176 16056
rect 24320 15026 24348 19654
rect 24412 18290 24440 24006
rect 24584 23860 24636 23866
rect 24584 23802 24636 23808
rect 24596 23322 24624 23802
rect 24584 23316 24636 23322
rect 24584 23258 24636 23264
rect 24596 22094 24624 23258
rect 24688 23050 24716 25094
rect 24676 23044 24728 23050
rect 24676 22986 24728 22992
rect 24780 22642 24808 28358
rect 24952 26852 25004 26858
rect 24952 26794 25004 26800
rect 24858 24440 24914 24449
rect 24858 24375 24914 24384
rect 24872 24274 24900 24375
rect 24860 24268 24912 24274
rect 24860 24210 24912 24216
rect 24768 22636 24820 22642
rect 24768 22578 24820 22584
rect 24504 22066 24624 22094
rect 24504 21486 24532 22066
rect 24858 21992 24914 22001
rect 24858 21927 24914 21936
rect 24492 21480 24544 21486
rect 24492 21422 24544 21428
rect 24872 21010 24900 21927
rect 24860 21004 24912 21010
rect 24860 20946 24912 20952
rect 24964 20466 24992 26794
rect 25056 24138 25084 28970
rect 25226 28520 25282 28529
rect 25226 28455 25228 28464
rect 25280 28455 25282 28464
rect 25228 28426 25280 28432
rect 25240 28218 25268 28426
rect 25228 28212 25280 28218
rect 25228 28154 25280 28160
rect 25136 28008 25188 28014
rect 25136 27950 25188 27956
rect 25148 26586 25176 27950
rect 25228 27940 25280 27946
rect 25228 27882 25280 27888
rect 25136 26580 25188 26586
rect 25136 26522 25188 26528
rect 25136 25832 25188 25838
rect 25136 25774 25188 25780
rect 25148 25265 25176 25774
rect 25134 25256 25190 25265
rect 25134 25191 25190 25200
rect 25136 24948 25188 24954
rect 25136 24890 25188 24896
rect 25148 24410 25176 24890
rect 25136 24404 25188 24410
rect 25136 24346 25188 24352
rect 25044 24132 25096 24138
rect 25044 24074 25096 24080
rect 25148 22778 25176 24346
rect 25136 22772 25188 22778
rect 25136 22714 25188 22720
rect 25148 22234 25176 22714
rect 25136 22228 25188 22234
rect 25136 22170 25188 22176
rect 25148 21622 25176 22170
rect 25136 21616 25188 21622
rect 25136 21558 25188 21564
rect 25240 20942 25268 27882
rect 25320 27396 25372 27402
rect 25320 27338 25372 27344
rect 25228 20936 25280 20942
rect 25228 20878 25280 20884
rect 24952 20460 25004 20466
rect 24952 20402 25004 20408
rect 24950 20360 25006 20369
rect 24950 20295 25006 20304
rect 24964 19922 24992 20295
rect 24952 19916 25004 19922
rect 24952 19858 25004 19864
rect 25332 19854 25360 27338
rect 25424 23798 25452 30126
rect 25516 29345 25544 30670
rect 25502 29336 25558 29345
rect 25502 29271 25504 29280
rect 25556 29271 25558 29280
rect 25504 29242 25556 29248
rect 25412 23792 25464 23798
rect 25412 23734 25464 23740
rect 25320 19848 25372 19854
rect 25320 19790 25372 19796
rect 24766 19544 24822 19553
rect 24766 19479 24822 19488
rect 24584 18760 24636 18766
rect 24584 18702 24636 18708
rect 24674 18728 24730 18737
rect 24400 18284 24452 18290
rect 24400 18226 24452 18232
rect 24596 17882 24624 18702
rect 24674 18663 24730 18672
rect 24584 17876 24636 17882
rect 24584 17818 24636 17824
rect 24688 17134 24716 18663
rect 24780 18222 24808 19479
rect 24768 18216 24820 18222
rect 24768 18158 24820 18164
rect 24676 17128 24728 17134
rect 24676 17070 24728 17076
rect 24766 17096 24822 17105
rect 24766 17031 24822 17040
rect 24584 16448 24636 16454
rect 24584 16390 24636 16396
rect 24596 15502 24624 16390
rect 24674 16280 24730 16289
rect 24674 16215 24730 16224
rect 24584 15496 24636 15502
rect 24584 15438 24636 15444
rect 24308 15020 24360 15026
rect 24308 14962 24360 14968
rect 24688 14958 24716 16215
rect 24780 16046 24808 17031
rect 24768 16040 24820 16046
rect 24768 15982 24820 15988
rect 24950 15464 25006 15473
rect 24950 15399 24952 15408
rect 25004 15399 25006 15408
rect 24952 15370 25004 15376
rect 24676 14952 24728 14958
rect 24676 14894 24728 14900
rect 23940 14884 23992 14890
rect 23940 14826 23992 14832
rect 23848 13932 23900 13938
rect 23848 13874 23900 13880
rect 23480 12232 23532 12238
rect 23480 12174 23532 12180
rect 23296 12096 23348 12102
rect 23296 12038 23348 12044
rect 22950 11452 23258 11461
rect 22950 11450 22956 11452
rect 23012 11450 23036 11452
rect 23092 11450 23116 11452
rect 23172 11450 23196 11452
rect 23252 11450 23258 11452
rect 23012 11398 23014 11450
rect 23194 11398 23196 11450
rect 22950 11396 22956 11398
rect 23012 11396 23036 11398
rect 23092 11396 23116 11398
rect 23172 11396 23196 11398
rect 23252 11396 23258 11398
rect 22950 11387 23258 11396
rect 22950 10364 23258 10373
rect 22950 10362 22956 10364
rect 23012 10362 23036 10364
rect 23092 10362 23116 10364
rect 23172 10362 23196 10364
rect 23252 10362 23258 10364
rect 23012 10310 23014 10362
rect 23194 10310 23196 10362
rect 22950 10308 22956 10310
rect 23012 10308 23036 10310
rect 23092 10308 23116 10310
rect 23172 10308 23196 10310
rect 23252 10308 23258 10310
rect 22950 10299 23258 10308
rect 22836 10056 22888 10062
rect 22836 9998 22888 10004
rect 22664 9574 22784 9602
rect 22560 4684 22612 4690
rect 22560 4626 22612 4632
rect 22664 3194 22692 9574
rect 22836 9444 22888 9450
rect 22836 9386 22888 9392
rect 22744 8424 22796 8430
rect 22744 8366 22796 8372
rect 22756 3233 22784 8366
rect 22848 4146 22876 9386
rect 22950 9276 23258 9285
rect 22950 9274 22956 9276
rect 23012 9274 23036 9276
rect 23092 9274 23116 9276
rect 23172 9274 23196 9276
rect 23252 9274 23258 9276
rect 23012 9222 23014 9274
rect 23194 9222 23196 9274
rect 22950 9220 22956 9222
rect 23012 9220 23036 9222
rect 23092 9220 23116 9222
rect 23172 9220 23196 9222
rect 23252 9220 23258 9222
rect 22950 9211 23258 9220
rect 23308 8974 23336 12038
rect 23388 11280 23440 11286
rect 23388 11222 23440 11228
rect 23296 8968 23348 8974
rect 23296 8910 23348 8916
rect 23296 8832 23348 8838
rect 23296 8774 23348 8780
rect 22950 8188 23258 8197
rect 22950 8186 22956 8188
rect 23012 8186 23036 8188
rect 23092 8186 23116 8188
rect 23172 8186 23196 8188
rect 23252 8186 23258 8188
rect 23012 8134 23014 8186
rect 23194 8134 23196 8186
rect 22950 8132 22956 8134
rect 23012 8132 23036 8134
rect 23092 8132 23116 8134
rect 23172 8132 23196 8134
rect 23252 8132 23258 8134
rect 22950 8123 23258 8132
rect 23308 8106 23336 8774
rect 23400 8498 23428 11222
rect 23848 11076 23900 11082
rect 23848 11018 23900 11024
rect 23572 9920 23624 9926
rect 23572 9862 23624 9868
rect 23480 9376 23532 9382
rect 23480 9318 23532 9324
rect 23388 8492 23440 8498
rect 23388 8434 23440 8440
rect 23308 8078 23428 8106
rect 23296 7948 23348 7954
rect 23296 7890 23348 7896
rect 22950 7100 23258 7109
rect 22950 7098 22956 7100
rect 23012 7098 23036 7100
rect 23092 7098 23116 7100
rect 23172 7098 23196 7100
rect 23252 7098 23258 7100
rect 23012 7046 23014 7098
rect 23194 7046 23196 7098
rect 22950 7044 22956 7046
rect 23012 7044 23036 7046
rect 23092 7044 23116 7046
rect 23172 7044 23196 7046
rect 23252 7044 23258 7046
rect 22950 7035 23258 7044
rect 22950 6012 23258 6021
rect 22950 6010 22956 6012
rect 23012 6010 23036 6012
rect 23092 6010 23116 6012
rect 23172 6010 23196 6012
rect 23252 6010 23258 6012
rect 23012 5958 23014 6010
rect 23194 5958 23196 6010
rect 22950 5956 22956 5958
rect 23012 5956 23036 5958
rect 23092 5956 23116 5958
rect 23172 5956 23196 5958
rect 23252 5956 23258 5958
rect 22950 5947 23258 5956
rect 22950 4924 23258 4933
rect 22950 4922 22956 4924
rect 23012 4922 23036 4924
rect 23092 4922 23116 4924
rect 23172 4922 23196 4924
rect 23252 4922 23258 4924
rect 23012 4870 23014 4922
rect 23194 4870 23196 4922
rect 22950 4868 22956 4870
rect 23012 4868 23036 4870
rect 23092 4868 23116 4870
rect 23172 4868 23196 4870
rect 23252 4868 23258 4870
rect 22950 4859 23258 4868
rect 23308 4842 23336 7890
rect 23400 6798 23428 8078
rect 23388 6792 23440 6798
rect 23388 6734 23440 6740
rect 23492 6322 23520 9318
rect 23584 7886 23612 9862
rect 23860 9586 23888 11018
rect 23952 10674 23980 14826
rect 25134 14648 25190 14657
rect 25134 14583 25190 14592
rect 25148 14006 25176 14583
rect 25136 14000 25188 14006
rect 25136 13942 25188 13948
rect 24766 13832 24822 13841
rect 24766 13767 24822 13776
rect 24780 12782 24808 13767
rect 24952 13252 25004 13258
rect 24952 13194 25004 13200
rect 24964 13025 24992 13194
rect 24950 13016 25006 13025
rect 24950 12951 25006 12960
rect 24768 12776 24820 12782
rect 24768 12718 24820 12724
rect 24860 12368 24912 12374
rect 24860 12310 24912 12316
rect 24766 11384 24822 11393
rect 24766 11319 24822 11328
rect 23940 10668 23992 10674
rect 23940 10610 23992 10616
rect 24780 10606 24808 11319
rect 24768 10600 24820 10606
rect 24674 10568 24730 10577
rect 24768 10542 24820 10548
rect 24674 10503 24730 10512
rect 23848 9580 23900 9586
rect 23848 9522 23900 9528
rect 24688 9518 24716 10503
rect 24676 9512 24728 9518
rect 24676 9454 24728 9460
rect 24872 8974 24900 12310
rect 25134 12200 25190 12209
rect 25134 12135 25190 12144
rect 25148 11830 25176 12135
rect 25136 11824 25188 11830
rect 25136 11766 25188 11772
rect 24952 9988 25004 9994
rect 24952 9930 25004 9936
rect 24964 9761 24992 9930
rect 24950 9752 25006 9761
rect 24950 9687 25006 9696
rect 24860 8968 24912 8974
rect 24860 8910 24912 8916
rect 25134 8936 25190 8945
rect 25134 8871 25190 8880
rect 23940 8832 23992 8838
rect 23940 8774 23992 8780
rect 23572 7880 23624 7886
rect 23572 7822 23624 7828
rect 23480 6316 23532 6322
rect 23480 6258 23532 6264
rect 23952 5234 23980 8774
rect 25148 8566 25176 8871
rect 25136 8560 25188 8566
rect 25136 8502 25188 8508
rect 25134 8120 25190 8129
rect 25134 8055 25190 8064
rect 24676 7744 24728 7750
rect 24676 7686 24728 7692
rect 23940 5228 23992 5234
rect 23940 5170 23992 5176
rect 23386 4856 23442 4865
rect 23308 4814 23386 4842
rect 23386 4791 23442 4800
rect 24688 4622 24716 7686
rect 25148 7478 25176 8055
rect 25136 7472 25188 7478
rect 25136 7414 25188 7420
rect 24766 7304 24822 7313
rect 24766 7239 24822 7248
rect 24780 6254 24808 7239
rect 25780 6724 25832 6730
rect 25780 6666 25832 6672
rect 25792 6497 25820 6666
rect 25778 6488 25834 6497
rect 25778 6423 25834 6432
rect 24768 6248 24820 6254
rect 24768 6190 24820 6196
rect 24766 5672 24822 5681
rect 24766 5607 24822 5616
rect 24780 5166 24808 5607
rect 24768 5160 24820 5166
rect 24768 5102 24820 5108
rect 24676 4616 24728 4622
rect 24676 4558 24728 4564
rect 22836 4140 22888 4146
rect 22836 4082 22888 4088
rect 22950 3836 23258 3845
rect 22950 3834 22956 3836
rect 23012 3834 23036 3836
rect 23092 3834 23116 3836
rect 23172 3834 23196 3836
rect 23252 3834 23258 3836
rect 23012 3782 23014 3834
rect 23194 3782 23196 3834
rect 22950 3780 22956 3782
rect 23012 3780 23036 3782
rect 23092 3780 23116 3782
rect 23172 3780 23196 3782
rect 23252 3780 23258 3782
rect 22950 3771 23258 3780
rect 23754 3496 23810 3505
rect 23754 3431 23810 3440
rect 24952 3460 25004 3466
rect 22836 3392 22888 3398
rect 22836 3334 22888 3340
rect 23572 3392 23624 3398
rect 23572 3334 23624 3340
rect 22742 3224 22798 3233
rect 22652 3188 22704 3194
rect 22742 3159 22798 3168
rect 22652 3130 22704 3136
rect 22652 3052 22704 3058
rect 22652 2994 22704 3000
rect 22468 2848 22520 2854
rect 22468 2790 22520 2796
rect 22664 800 22692 2994
rect 22848 2530 22876 3334
rect 23584 3126 23612 3334
rect 23572 3120 23624 3126
rect 23572 3062 23624 3068
rect 23388 2984 23440 2990
rect 23388 2926 23440 2932
rect 22950 2748 23258 2757
rect 22950 2746 22956 2748
rect 23012 2746 23036 2748
rect 23092 2746 23116 2748
rect 23172 2746 23196 2748
rect 23252 2746 23258 2748
rect 23012 2694 23014 2746
rect 23194 2694 23196 2746
rect 22950 2692 22956 2694
rect 23012 2692 23036 2694
rect 23092 2692 23116 2694
rect 23172 2692 23196 2694
rect 23252 2692 23258 2694
rect 22950 2683 23258 2692
rect 22848 2502 23060 2530
rect 23032 800 23060 2502
rect 23400 800 23428 2926
rect 23768 800 23796 3431
rect 24952 3402 25004 3408
rect 24124 3392 24176 3398
rect 24124 3334 24176 3340
rect 24136 800 24164 3334
rect 13188 734 13400 762
rect 13450 0 13506 800
rect 13818 0 13874 800
rect 14186 0 14242 800
rect 14554 0 14610 800
rect 14922 0 14978 800
rect 15290 0 15346 800
rect 15658 0 15714 800
rect 16026 0 16082 800
rect 16394 0 16450 800
rect 16762 0 16818 800
rect 17130 0 17186 800
rect 17498 0 17554 800
rect 17866 0 17922 800
rect 18234 0 18290 800
rect 18602 0 18658 800
rect 18970 0 19026 800
rect 19338 0 19394 800
rect 19706 0 19762 800
rect 20074 0 20130 800
rect 20442 0 20498 800
rect 20810 0 20866 800
rect 21178 0 21234 800
rect 21546 0 21602 800
rect 21914 0 21970 800
rect 22282 0 22338 800
rect 22650 0 22706 800
rect 23018 0 23074 800
rect 23386 0 23442 800
rect 23754 0 23810 800
rect 24122 0 24178 800
rect 24490 0 24546 800
rect 24858 0 24914 800
rect 24964 785 24992 3402
rect 25320 2440 25372 2446
rect 25320 2382 25372 2388
rect 25332 1601 25360 2382
rect 25318 1592 25374 1601
rect 25318 1527 25374 1536
rect 24950 776 25006 785
rect 24950 711 25006 720
<< via2 >>
rect 2778 55392 2834 55448
rect 2956 53882 3012 53884
rect 3036 53882 3092 53884
rect 3116 53882 3172 53884
rect 3196 53882 3252 53884
rect 2956 53830 3002 53882
rect 3002 53830 3012 53882
rect 3036 53830 3066 53882
rect 3066 53830 3078 53882
rect 3078 53830 3092 53882
rect 3116 53830 3130 53882
rect 3130 53830 3142 53882
rect 3142 53830 3172 53882
rect 3196 53830 3206 53882
rect 3206 53830 3252 53882
rect 2956 53828 3012 53830
rect 3036 53828 3092 53830
rect 3116 53828 3172 53830
rect 3196 53828 3252 53830
rect 2956 52794 3012 52796
rect 3036 52794 3092 52796
rect 3116 52794 3172 52796
rect 3196 52794 3252 52796
rect 2956 52742 3002 52794
rect 3002 52742 3012 52794
rect 3036 52742 3066 52794
rect 3066 52742 3078 52794
rect 3078 52742 3092 52794
rect 3116 52742 3130 52794
rect 3130 52742 3142 52794
rect 3142 52742 3172 52794
rect 3196 52742 3206 52794
rect 3206 52742 3252 52794
rect 2956 52740 3012 52742
rect 3036 52740 3092 52742
rect 3116 52740 3172 52742
rect 3196 52740 3252 52742
rect 3422 52964 3478 53000
rect 3422 52944 3424 52964
rect 3424 52944 3476 52964
rect 3476 52944 3478 52964
rect 2956 51706 3012 51708
rect 3036 51706 3092 51708
rect 3116 51706 3172 51708
rect 3196 51706 3252 51708
rect 2956 51654 3002 51706
rect 3002 51654 3012 51706
rect 3036 51654 3066 51706
rect 3066 51654 3078 51706
rect 3078 51654 3092 51706
rect 3116 51654 3130 51706
rect 3130 51654 3142 51706
rect 3142 51654 3172 51706
rect 3196 51654 3206 51706
rect 3206 51654 3252 51706
rect 2956 51652 3012 51654
rect 3036 51652 3092 51654
rect 3116 51652 3172 51654
rect 3196 51652 3252 51654
rect 2956 50618 3012 50620
rect 3036 50618 3092 50620
rect 3116 50618 3172 50620
rect 3196 50618 3252 50620
rect 2956 50566 3002 50618
rect 3002 50566 3012 50618
rect 3036 50566 3066 50618
rect 3066 50566 3078 50618
rect 3078 50566 3092 50618
rect 3116 50566 3130 50618
rect 3130 50566 3142 50618
rect 3142 50566 3172 50618
rect 3196 50566 3206 50618
rect 3206 50566 3252 50618
rect 2956 50564 3012 50566
rect 3036 50564 3092 50566
rect 3116 50564 3172 50566
rect 3196 50564 3252 50566
rect 3974 50360 4030 50416
rect 2956 49530 3012 49532
rect 3036 49530 3092 49532
rect 3116 49530 3172 49532
rect 3196 49530 3252 49532
rect 2956 49478 3002 49530
rect 3002 49478 3012 49530
rect 3036 49478 3066 49530
rect 3066 49478 3078 49530
rect 3078 49478 3092 49530
rect 3116 49478 3130 49530
rect 3130 49478 3142 49530
rect 3142 49478 3172 49530
rect 3196 49478 3206 49530
rect 3206 49478 3252 49530
rect 2956 49476 3012 49478
rect 3036 49476 3092 49478
rect 3116 49476 3172 49478
rect 3196 49476 3252 49478
rect 2956 48442 3012 48444
rect 3036 48442 3092 48444
rect 3116 48442 3172 48444
rect 3196 48442 3252 48444
rect 2956 48390 3002 48442
rect 3002 48390 3012 48442
rect 3036 48390 3066 48442
rect 3066 48390 3078 48442
rect 3078 48390 3092 48442
rect 3116 48390 3130 48442
rect 3130 48390 3142 48442
rect 3142 48390 3172 48442
rect 3196 48390 3206 48442
rect 3206 48390 3252 48442
rect 2956 48388 3012 48390
rect 3036 48388 3092 48390
rect 3116 48388 3172 48390
rect 3196 48388 3252 48390
rect 2956 47354 3012 47356
rect 3036 47354 3092 47356
rect 3116 47354 3172 47356
rect 3196 47354 3252 47356
rect 2956 47302 3002 47354
rect 3002 47302 3012 47354
rect 3036 47302 3066 47354
rect 3066 47302 3078 47354
rect 3078 47302 3092 47354
rect 3116 47302 3130 47354
rect 3130 47302 3142 47354
rect 3142 47302 3172 47354
rect 3196 47302 3206 47354
rect 3206 47302 3252 47354
rect 2956 47300 3012 47302
rect 3036 47300 3092 47302
rect 3116 47300 3172 47302
rect 3196 47300 3252 47302
rect 2956 46266 3012 46268
rect 3036 46266 3092 46268
rect 3116 46266 3172 46268
rect 3196 46266 3252 46268
rect 2956 46214 3002 46266
rect 3002 46214 3012 46266
rect 3036 46214 3066 46266
rect 3066 46214 3078 46266
rect 3078 46214 3092 46266
rect 3116 46214 3130 46266
rect 3130 46214 3142 46266
rect 3142 46214 3172 46266
rect 3196 46214 3206 46266
rect 3206 46214 3252 46266
rect 2956 46212 3012 46214
rect 3036 46212 3092 46214
rect 3116 46212 3172 46214
rect 3196 46212 3252 46214
rect 2956 45178 3012 45180
rect 3036 45178 3092 45180
rect 3116 45178 3172 45180
rect 3196 45178 3252 45180
rect 2956 45126 3002 45178
rect 3002 45126 3012 45178
rect 3036 45126 3066 45178
rect 3066 45126 3078 45178
rect 3078 45126 3092 45178
rect 3116 45126 3130 45178
rect 3130 45126 3142 45178
rect 3142 45126 3172 45178
rect 3196 45126 3206 45178
rect 3206 45126 3252 45178
rect 2956 45124 3012 45126
rect 3036 45124 3092 45126
rect 3116 45124 3172 45126
rect 3196 45124 3252 45126
rect 2956 44090 3012 44092
rect 3036 44090 3092 44092
rect 3116 44090 3172 44092
rect 3196 44090 3252 44092
rect 2956 44038 3002 44090
rect 3002 44038 3012 44090
rect 3036 44038 3066 44090
rect 3066 44038 3078 44090
rect 3078 44038 3092 44090
rect 3116 44038 3130 44090
rect 3130 44038 3142 44090
rect 3142 44038 3172 44090
rect 3196 44038 3206 44090
rect 3206 44038 3252 44090
rect 2956 44036 3012 44038
rect 3036 44036 3092 44038
rect 3116 44036 3172 44038
rect 3196 44036 3252 44038
rect 1306 43152 1362 43208
rect 2956 43002 3012 43004
rect 3036 43002 3092 43004
rect 3116 43002 3172 43004
rect 3196 43002 3252 43004
rect 2956 42950 3002 43002
rect 3002 42950 3012 43002
rect 3036 42950 3066 43002
rect 3066 42950 3078 43002
rect 3078 42950 3092 43002
rect 3116 42950 3130 43002
rect 3130 42950 3142 43002
rect 3142 42950 3172 43002
rect 3196 42950 3206 43002
rect 3206 42950 3252 43002
rect 2956 42948 3012 42950
rect 3036 42948 3092 42950
rect 3116 42948 3172 42950
rect 3196 42948 3252 42950
rect 2956 41914 3012 41916
rect 3036 41914 3092 41916
rect 3116 41914 3172 41916
rect 3196 41914 3252 41916
rect 2956 41862 3002 41914
rect 3002 41862 3012 41914
rect 3036 41862 3066 41914
rect 3066 41862 3078 41914
rect 3078 41862 3092 41914
rect 3116 41862 3130 41914
rect 3130 41862 3142 41914
rect 3142 41862 3172 41914
rect 3196 41862 3206 41914
rect 3206 41862 3252 41914
rect 2956 41860 3012 41862
rect 3036 41860 3092 41862
rect 3116 41860 3172 41862
rect 3196 41860 3252 41862
rect 2956 40826 3012 40828
rect 3036 40826 3092 40828
rect 3116 40826 3172 40828
rect 3196 40826 3252 40828
rect 2956 40774 3002 40826
rect 3002 40774 3012 40826
rect 3036 40774 3066 40826
rect 3066 40774 3078 40826
rect 3078 40774 3092 40826
rect 3116 40774 3130 40826
rect 3130 40774 3142 40826
rect 3142 40774 3172 40826
rect 3196 40774 3206 40826
rect 3206 40774 3252 40826
rect 2956 40772 3012 40774
rect 3036 40772 3092 40774
rect 3116 40772 3172 40774
rect 3196 40772 3252 40774
rect 1306 40704 1362 40760
rect 2956 39738 3012 39740
rect 3036 39738 3092 39740
rect 3116 39738 3172 39740
rect 3196 39738 3252 39740
rect 2956 39686 3002 39738
rect 3002 39686 3012 39738
rect 3036 39686 3066 39738
rect 3066 39686 3078 39738
rect 3078 39686 3092 39738
rect 3116 39686 3130 39738
rect 3130 39686 3142 39738
rect 3142 39686 3172 39738
rect 3196 39686 3206 39738
rect 3206 39686 3252 39738
rect 2956 39684 3012 39686
rect 3036 39684 3092 39686
rect 3116 39684 3172 39686
rect 3196 39684 3252 39686
rect 2956 38650 3012 38652
rect 3036 38650 3092 38652
rect 3116 38650 3172 38652
rect 3196 38650 3252 38652
rect 2956 38598 3002 38650
rect 3002 38598 3012 38650
rect 3036 38598 3066 38650
rect 3066 38598 3078 38650
rect 3078 38598 3092 38650
rect 3116 38598 3130 38650
rect 3130 38598 3142 38650
rect 3142 38598 3172 38650
rect 3196 38598 3206 38650
rect 3206 38598 3252 38650
rect 2956 38596 3012 38598
rect 3036 38596 3092 38598
rect 3116 38596 3172 38598
rect 3196 38596 3252 38598
rect 1306 38292 1308 38312
rect 1308 38292 1360 38312
rect 1360 38292 1362 38312
rect 1306 38256 1362 38292
rect 2956 37562 3012 37564
rect 3036 37562 3092 37564
rect 3116 37562 3172 37564
rect 3196 37562 3252 37564
rect 2956 37510 3002 37562
rect 3002 37510 3012 37562
rect 3036 37510 3066 37562
rect 3066 37510 3078 37562
rect 3078 37510 3092 37562
rect 3116 37510 3130 37562
rect 3130 37510 3142 37562
rect 3142 37510 3172 37562
rect 3196 37510 3206 37562
rect 3206 37510 3252 37562
rect 2956 37508 3012 37510
rect 3036 37508 3092 37510
rect 3116 37508 3172 37510
rect 3196 37508 3252 37510
rect 2956 36474 3012 36476
rect 3036 36474 3092 36476
rect 3116 36474 3172 36476
rect 3196 36474 3252 36476
rect 2956 36422 3002 36474
rect 3002 36422 3012 36474
rect 3036 36422 3066 36474
rect 3066 36422 3078 36474
rect 3078 36422 3092 36474
rect 3116 36422 3130 36474
rect 3130 36422 3142 36474
rect 3142 36422 3172 36474
rect 3196 36422 3206 36474
rect 3206 36422 3252 36474
rect 2956 36420 3012 36422
rect 3036 36420 3092 36422
rect 3116 36420 3172 36422
rect 3196 36420 3252 36422
rect 1306 33360 1362 33416
rect 1766 35808 1822 35864
rect 2956 35386 3012 35388
rect 3036 35386 3092 35388
rect 3116 35386 3172 35388
rect 3196 35386 3252 35388
rect 2956 35334 3002 35386
rect 3002 35334 3012 35386
rect 3036 35334 3066 35386
rect 3066 35334 3078 35386
rect 3078 35334 3092 35386
rect 3116 35334 3130 35386
rect 3130 35334 3142 35386
rect 3142 35334 3172 35386
rect 3196 35334 3206 35386
rect 3206 35334 3252 35386
rect 2956 35332 3012 35334
rect 3036 35332 3092 35334
rect 3116 35332 3172 35334
rect 3196 35332 3252 35334
rect 2956 34298 3012 34300
rect 3036 34298 3092 34300
rect 3116 34298 3172 34300
rect 3196 34298 3252 34300
rect 2956 34246 3002 34298
rect 3002 34246 3012 34298
rect 3036 34246 3066 34298
rect 3066 34246 3078 34298
rect 3078 34246 3092 34298
rect 3116 34246 3130 34298
rect 3130 34246 3142 34298
rect 3142 34246 3172 34298
rect 3196 34246 3206 34298
rect 3206 34246 3252 34298
rect 2956 34244 3012 34246
rect 3036 34244 3092 34246
rect 3116 34244 3172 34246
rect 3196 34244 3252 34246
rect 2956 33210 3012 33212
rect 3036 33210 3092 33212
rect 3116 33210 3172 33212
rect 3196 33210 3252 33212
rect 2956 33158 3002 33210
rect 3002 33158 3012 33210
rect 3036 33158 3066 33210
rect 3066 33158 3078 33210
rect 3078 33158 3092 33210
rect 3116 33158 3130 33210
rect 3130 33158 3142 33210
rect 3142 33158 3172 33210
rect 3196 33158 3206 33210
rect 3206 33158 3252 33210
rect 2956 33156 3012 33158
rect 3036 33156 3092 33158
rect 3116 33156 3172 33158
rect 3196 33156 3252 33158
rect 2956 32122 3012 32124
rect 3036 32122 3092 32124
rect 3116 32122 3172 32124
rect 3196 32122 3252 32124
rect 2956 32070 3002 32122
rect 3002 32070 3012 32122
rect 3036 32070 3066 32122
rect 3066 32070 3078 32122
rect 3078 32070 3092 32122
rect 3116 32070 3130 32122
rect 3130 32070 3142 32122
rect 3142 32070 3172 32122
rect 3196 32070 3206 32122
rect 3206 32070 3252 32122
rect 2956 32068 3012 32070
rect 3036 32068 3092 32070
rect 3116 32068 3172 32070
rect 3196 32068 3252 32070
rect 2956 31034 3012 31036
rect 3036 31034 3092 31036
rect 3116 31034 3172 31036
rect 3196 31034 3252 31036
rect 2956 30982 3002 31034
rect 3002 30982 3012 31034
rect 3036 30982 3066 31034
rect 3066 30982 3078 31034
rect 3078 30982 3092 31034
rect 3116 30982 3130 31034
rect 3130 30982 3142 31034
rect 3142 30982 3172 31034
rect 3196 30982 3206 31034
rect 3206 30982 3252 31034
rect 2956 30980 3012 30982
rect 3036 30980 3092 30982
rect 3116 30980 3172 30982
rect 3196 30980 3252 30982
rect 2778 30912 2834 30968
rect 2956 29946 3012 29948
rect 3036 29946 3092 29948
rect 3116 29946 3172 29948
rect 3196 29946 3252 29948
rect 2956 29894 3002 29946
rect 3002 29894 3012 29946
rect 3036 29894 3066 29946
rect 3066 29894 3078 29946
rect 3078 29894 3092 29946
rect 3116 29894 3130 29946
rect 3130 29894 3142 29946
rect 3142 29894 3172 29946
rect 3196 29894 3206 29946
rect 3206 29894 3252 29946
rect 2956 29892 3012 29894
rect 3036 29892 3092 29894
rect 3116 29892 3172 29894
rect 3196 29892 3252 29894
rect 2956 28858 3012 28860
rect 3036 28858 3092 28860
rect 3116 28858 3172 28860
rect 3196 28858 3252 28860
rect 2956 28806 3002 28858
rect 3002 28806 3012 28858
rect 3036 28806 3066 28858
rect 3066 28806 3078 28858
rect 3078 28806 3092 28858
rect 3116 28806 3130 28858
rect 3130 28806 3142 28858
rect 3142 28806 3172 28858
rect 3196 28806 3206 28858
rect 3206 28806 3252 28858
rect 2956 28804 3012 28806
rect 3036 28804 3092 28806
rect 3116 28804 3172 28806
rect 3196 28804 3252 28806
rect 2870 28464 2926 28520
rect 1306 21120 1362 21176
rect 2778 26016 2834 26072
rect 2956 27770 3012 27772
rect 3036 27770 3092 27772
rect 3116 27770 3172 27772
rect 3196 27770 3252 27772
rect 2956 27718 3002 27770
rect 3002 27718 3012 27770
rect 3036 27718 3066 27770
rect 3066 27718 3078 27770
rect 3078 27718 3092 27770
rect 3116 27718 3130 27770
rect 3130 27718 3142 27770
rect 3142 27718 3172 27770
rect 3196 27718 3206 27770
rect 3206 27718 3252 27770
rect 2956 27716 3012 27718
rect 3036 27716 3092 27718
rect 3116 27716 3172 27718
rect 3196 27716 3252 27718
rect 4066 48048 4122 48104
rect 4066 45620 4122 45656
rect 4066 45600 4068 45620
rect 4068 45600 4120 45620
rect 4120 45600 4122 45620
rect 2956 26682 3012 26684
rect 3036 26682 3092 26684
rect 3116 26682 3172 26684
rect 3196 26682 3252 26684
rect 2956 26630 3002 26682
rect 3002 26630 3012 26682
rect 3036 26630 3066 26682
rect 3066 26630 3078 26682
rect 3078 26630 3092 26682
rect 3116 26630 3130 26682
rect 3130 26630 3142 26682
rect 3142 26630 3172 26682
rect 3196 26630 3206 26682
rect 3206 26630 3252 26682
rect 2956 26628 3012 26630
rect 3036 26628 3092 26630
rect 3116 26628 3172 26630
rect 3196 26628 3252 26630
rect 2956 25594 3012 25596
rect 3036 25594 3092 25596
rect 3116 25594 3172 25596
rect 3196 25594 3252 25596
rect 2956 25542 3002 25594
rect 3002 25542 3012 25594
rect 3036 25542 3066 25594
rect 3066 25542 3078 25594
rect 3078 25542 3092 25594
rect 3116 25542 3130 25594
rect 3130 25542 3142 25594
rect 3142 25542 3172 25594
rect 3196 25542 3206 25594
rect 3206 25542 3252 25594
rect 2956 25540 3012 25542
rect 3036 25540 3092 25542
rect 3116 25540 3172 25542
rect 3196 25540 3252 25542
rect 2956 24506 3012 24508
rect 3036 24506 3092 24508
rect 3116 24506 3172 24508
rect 3196 24506 3252 24508
rect 2956 24454 3002 24506
rect 3002 24454 3012 24506
rect 3036 24454 3066 24506
rect 3066 24454 3078 24506
rect 3078 24454 3092 24506
rect 3116 24454 3130 24506
rect 3130 24454 3142 24506
rect 3142 24454 3172 24506
rect 3196 24454 3206 24506
rect 3206 24454 3252 24506
rect 2956 24452 3012 24454
rect 3036 24452 3092 24454
rect 3116 24452 3172 24454
rect 3196 24452 3252 24454
rect 2870 23568 2926 23624
rect 1306 18672 1362 18728
rect 1306 16224 1362 16280
rect 2956 23418 3012 23420
rect 3036 23418 3092 23420
rect 3116 23418 3172 23420
rect 3196 23418 3252 23420
rect 2956 23366 3002 23418
rect 3002 23366 3012 23418
rect 3036 23366 3066 23418
rect 3066 23366 3078 23418
rect 3078 23366 3092 23418
rect 3116 23366 3130 23418
rect 3130 23366 3142 23418
rect 3142 23366 3172 23418
rect 3196 23366 3206 23418
rect 3206 23366 3252 23418
rect 2956 23364 3012 23366
rect 3036 23364 3092 23366
rect 3116 23364 3172 23366
rect 3196 23364 3252 23366
rect 2956 22330 3012 22332
rect 3036 22330 3092 22332
rect 3116 22330 3172 22332
rect 3196 22330 3252 22332
rect 2956 22278 3002 22330
rect 3002 22278 3012 22330
rect 3036 22278 3066 22330
rect 3066 22278 3078 22330
rect 3078 22278 3092 22330
rect 3116 22278 3130 22330
rect 3130 22278 3142 22330
rect 3142 22278 3172 22330
rect 3196 22278 3206 22330
rect 3206 22278 3252 22330
rect 2956 22276 3012 22278
rect 3036 22276 3092 22278
rect 3116 22276 3172 22278
rect 3196 22276 3252 22278
rect 2956 21242 3012 21244
rect 3036 21242 3092 21244
rect 3116 21242 3172 21244
rect 3196 21242 3252 21244
rect 2956 21190 3002 21242
rect 3002 21190 3012 21242
rect 3036 21190 3066 21242
rect 3066 21190 3078 21242
rect 3078 21190 3092 21242
rect 3116 21190 3130 21242
rect 3130 21190 3142 21242
rect 3142 21190 3172 21242
rect 3196 21190 3206 21242
rect 3206 21190 3252 21242
rect 2956 21188 3012 21190
rect 3036 21188 3092 21190
rect 3116 21188 3172 21190
rect 3196 21188 3252 21190
rect 2956 20154 3012 20156
rect 3036 20154 3092 20156
rect 3116 20154 3172 20156
rect 3196 20154 3252 20156
rect 2956 20102 3002 20154
rect 3002 20102 3012 20154
rect 3036 20102 3066 20154
rect 3066 20102 3078 20154
rect 3078 20102 3092 20154
rect 3116 20102 3130 20154
rect 3130 20102 3142 20154
rect 3142 20102 3172 20154
rect 3196 20102 3206 20154
rect 3206 20102 3252 20154
rect 2956 20100 3012 20102
rect 3036 20100 3092 20102
rect 3116 20100 3172 20102
rect 3196 20100 3252 20102
rect 2956 19066 3012 19068
rect 3036 19066 3092 19068
rect 3116 19066 3172 19068
rect 3196 19066 3252 19068
rect 2956 19014 3002 19066
rect 3002 19014 3012 19066
rect 3036 19014 3066 19066
rect 3066 19014 3078 19066
rect 3078 19014 3092 19066
rect 3116 19014 3130 19066
rect 3130 19014 3142 19066
rect 3142 19014 3172 19066
rect 3196 19014 3206 19066
rect 3206 19014 3252 19066
rect 2956 19012 3012 19014
rect 3036 19012 3092 19014
rect 3116 19012 3172 19014
rect 3196 19012 3252 19014
rect 2956 17978 3012 17980
rect 3036 17978 3092 17980
rect 3116 17978 3172 17980
rect 3196 17978 3252 17980
rect 2956 17926 3002 17978
rect 3002 17926 3012 17978
rect 3036 17926 3066 17978
rect 3066 17926 3078 17978
rect 3078 17926 3092 17978
rect 3116 17926 3130 17978
rect 3130 17926 3142 17978
rect 3142 17926 3172 17978
rect 3196 17926 3206 17978
rect 3206 17926 3252 17978
rect 2956 17924 3012 17926
rect 3036 17924 3092 17926
rect 3116 17924 3172 17926
rect 3196 17924 3252 17926
rect 2956 16890 3012 16892
rect 3036 16890 3092 16892
rect 3116 16890 3172 16892
rect 3196 16890 3252 16892
rect 2956 16838 3002 16890
rect 3002 16838 3012 16890
rect 3036 16838 3066 16890
rect 3066 16838 3078 16890
rect 3078 16838 3092 16890
rect 3116 16838 3130 16890
rect 3130 16838 3142 16890
rect 3142 16838 3172 16890
rect 3196 16838 3206 16890
rect 3206 16838 3252 16890
rect 2956 16836 3012 16838
rect 3036 16836 3092 16838
rect 3116 16836 3172 16838
rect 3196 16836 3252 16838
rect 2956 15802 3012 15804
rect 3036 15802 3092 15804
rect 3116 15802 3172 15804
rect 3196 15802 3252 15804
rect 2956 15750 3002 15802
rect 3002 15750 3012 15802
rect 3036 15750 3066 15802
rect 3066 15750 3078 15802
rect 3078 15750 3092 15802
rect 3116 15750 3130 15802
rect 3130 15750 3142 15802
rect 3142 15750 3172 15802
rect 3196 15750 3206 15802
rect 3206 15750 3252 15802
rect 2956 15748 3012 15750
rect 3036 15748 3092 15750
rect 3116 15748 3172 15750
rect 3196 15748 3252 15750
rect 2956 14714 3012 14716
rect 3036 14714 3092 14716
rect 3116 14714 3172 14716
rect 3196 14714 3252 14716
rect 2956 14662 3002 14714
rect 3002 14662 3012 14714
rect 3036 14662 3066 14714
rect 3066 14662 3078 14714
rect 3078 14662 3092 14714
rect 3116 14662 3130 14714
rect 3130 14662 3142 14714
rect 3142 14662 3172 14714
rect 3196 14662 3206 14714
rect 3206 14662 3252 14714
rect 2956 14660 3012 14662
rect 3036 14660 3092 14662
rect 3116 14660 3172 14662
rect 3196 14660 3252 14662
rect 1306 13812 1308 13832
rect 1308 13812 1360 13832
rect 1360 13812 1362 13832
rect 1306 13776 1362 13812
rect 2956 13626 3012 13628
rect 3036 13626 3092 13628
rect 3116 13626 3172 13628
rect 3196 13626 3252 13628
rect 2956 13574 3002 13626
rect 3002 13574 3012 13626
rect 3036 13574 3066 13626
rect 3066 13574 3078 13626
rect 3078 13574 3092 13626
rect 3116 13574 3130 13626
rect 3130 13574 3142 13626
rect 3142 13574 3172 13626
rect 3196 13574 3206 13626
rect 3206 13574 3252 13626
rect 2956 13572 3012 13574
rect 3036 13572 3092 13574
rect 3116 13572 3172 13574
rect 3196 13572 3252 13574
rect 2956 12538 3012 12540
rect 3036 12538 3092 12540
rect 3116 12538 3172 12540
rect 3196 12538 3252 12540
rect 2956 12486 3002 12538
rect 3002 12486 3012 12538
rect 3036 12486 3066 12538
rect 3066 12486 3078 12538
rect 3078 12486 3092 12538
rect 3116 12486 3130 12538
rect 3130 12486 3142 12538
rect 3142 12486 3172 12538
rect 3196 12486 3206 12538
rect 3206 12486 3252 12538
rect 2956 12484 3012 12486
rect 3036 12484 3092 12486
rect 3116 12484 3172 12486
rect 3196 12484 3252 12486
rect 2956 11450 3012 11452
rect 3036 11450 3092 11452
rect 3116 11450 3172 11452
rect 3196 11450 3252 11452
rect 2956 11398 3002 11450
rect 3002 11398 3012 11450
rect 3036 11398 3066 11450
rect 3066 11398 3078 11450
rect 3078 11398 3092 11450
rect 3116 11398 3130 11450
rect 3130 11398 3142 11450
rect 3142 11398 3172 11450
rect 3196 11398 3206 11450
rect 3206 11398 3252 11450
rect 2956 11396 3012 11398
rect 3036 11396 3092 11398
rect 3116 11396 3172 11398
rect 3196 11396 3252 11398
rect 2778 11328 2834 11384
rect 2956 10362 3012 10364
rect 3036 10362 3092 10364
rect 3116 10362 3172 10364
rect 3196 10362 3252 10364
rect 2956 10310 3002 10362
rect 3002 10310 3012 10362
rect 3036 10310 3066 10362
rect 3066 10310 3078 10362
rect 3078 10310 3092 10362
rect 3116 10310 3130 10362
rect 3130 10310 3142 10362
rect 3142 10310 3172 10362
rect 3196 10310 3206 10362
rect 3206 10310 3252 10362
rect 2956 10308 3012 10310
rect 3036 10308 3092 10310
rect 3116 10308 3172 10310
rect 3196 10308 3252 10310
rect 2956 9274 3012 9276
rect 3036 9274 3092 9276
rect 3116 9274 3172 9276
rect 3196 9274 3252 9276
rect 2956 9222 3002 9274
rect 3002 9222 3012 9274
rect 3036 9222 3066 9274
rect 3066 9222 3078 9274
rect 3078 9222 3092 9274
rect 3116 9222 3130 9274
rect 3130 9222 3142 9274
rect 3142 9222 3172 9274
rect 3196 9222 3206 9274
rect 3206 9222 3252 9274
rect 2956 9220 3012 9222
rect 3036 9220 3092 9222
rect 3116 9220 3172 9222
rect 3196 9220 3252 9222
rect 2870 8880 2926 8936
rect 2956 8186 3012 8188
rect 3036 8186 3092 8188
rect 3116 8186 3172 8188
rect 3196 8186 3252 8188
rect 2956 8134 3002 8186
rect 3002 8134 3012 8186
rect 3036 8134 3066 8186
rect 3066 8134 3078 8186
rect 3078 8134 3092 8186
rect 3116 8134 3130 8186
rect 3130 8134 3142 8186
rect 3142 8134 3172 8186
rect 3196 8134 3206 8186
rect 3206 8134 3252 8186
rect 2956 8132 3012 8134
rect 3036 8132 3092 8134
rect 3116 8132 3172 8134
rect 3196 8132 3252 8134
rect 2956 7098 3012 7100
rect 3036 7098 3092 7100
rect 3116 7098 3172 7100
rect 3196 7098 3252 7100
rect 2956 7046 3002 7098
rect 3002 7046 3012 7098
rect 3036 7046 3066 7098
rect 3066 7046 3078 7098
rect 3078 7046 3092 7098
rect 3116 7046 3130 7098
rect 3130 7046 3142 7098
rect 3142 7046 3172 7098
rect 3196 7046 3206 7098
rect 3206 7046 3252 7098
rect 2956 7044 3012 7046
rect 3036 7044 3092 7046
rect 3116 7044 3172 7046
rect 3196 7044 3252 7046
rect 3054 6432 3110 6488
rect 2956 6010 3012 6012
rect 3036 6010 3092 6012
rect 3116 6010 3172 6012
rect 3196 6010 3252 6012
rect 2956 5958 3002 6010
rect 3002 5958 3012 6010
rect 3036 5958 3066 6010
rect 3066 5958 3078 6010
rect 3078 5958 3092 6010
rect 3116 5958 3130 6010
rect 3130 5958 3142 6010
rect 3142 5958 3172 6010
rect 3196 5958 3206 6010
rect 3206 5958 3252 6010
rect 2956 5956 3012 5958
rect 3036 5956 3092 5958
rect 3116 5956 3172 5958
rect 3196 5956 3252 5958
rect 2956 4922 3012 4924
rect 3036 4922 3092 4924
rect 3116 4922 3172 4924
rect 3196 4922 3252 4924
rect 2956 4870 3002 4922
rect 3002 4870 3012 4922
rect 3036 4870 3066 4922
rect 3066 4870 3078 4922
rect 3078 4870 3092 4922
rect 3116 4870 3130 4922
rect 3130 4870 3142 4922
rect 3142 4870 3172 4922
rect 3196 4870 3206 4922
rect 3206 4870 3252 4922
rect 2956 4868 3012 4870
rect 3036 4868 3092 4870
rect 3116 4868 3172 4870
rect 3196 4868 3252 4870
rect 2870 4020 2872 4040
rect 2872 4020 2924 4040
rect 2924 4020 2926 4040
rect 2870 3984 2926 4020
rect 2956 3834 3012 3836
rect 3036 3834 3092 3836
rect 3116 3834 3172 3836
rect 3196 3834 3252 3836
rect 2956 3782 3002 3834
rect 3002 3782 3012 3834
rect 3036 3782 3066 3834
rect 3066 3782 3078 3834
rect 3078 3782 3092 3834
rect 3116 3782 3130 3834
rect 3130 3782 3142 3834
rect 3142 3782 3172 3834
rect 3196 3782 3206 3834
rect 3206 3782 3252 3834
rect 2956 3780 3012 3782
rect 3036 3780 3092 3782
rect 3116 3780 3172 3782
rect 3196 3780 3252 3782
rect 2956 2746 3012 2748
rect 3036 2746 3092 2748
rect 3116 2746 3172 2748
rect 3196 2746 3252 2748
rect 2956 2694 3002 2746
rect 3002 2694 3012 2746
rect 3036 2694 3066 2746
rect 3066 2694 3078 2746
rect 3078 2694 3092 2746
rect 3116 2694 3130 2746
rect 3130 2694 3142 2746
rect 3142 2694 3172 2746
rect 3196 2694 3206 2746
rect 3206 2694 3252 2746
rect 2956 2692 3012 2694
rect 3036 2692 3092 2694
rect 3116 2692 3172 2694
rect 3196 2692 3252 2694
rect 2870 1536 2926 1592
rect 7956 54426 8012 54428
rect 8036 54426 8092 54428
rect 8116 54426 8172 54428
rect 8196 54426 8252 54428
rect 7956 54374 8002 54426
rect 8002 54374 8012 54426
rect 8036 54374 8066 54426
rect 8066 54374 8078 54426
rect 8078 54374 8092 54426
rect 8116 54374 8130 54426
rect 8130 54374 8142 54426
rect 8142 54374 8172 54426
rect 8196 54374 8206 54426
rect 8206 54374 8252 54426
rect 7956 54372 8012 54374
rect 8036 54372 8092 54374
rect 8116 54372 8172 54374
rect 8196 54372 8252 54374
rect 7956 53338 8012 53340
rect 8036 53338 8092 53340
rect 8116 53338 8172 53340
rect 8196 53338 8252 53340
rect 7956 53286 8002 53338
rect 8002 53286 8012 53338
rect 8036 53286 8066 53338
rect 8066 53286 8078 53338
rect 8078 53286 8092 53338
rect 8116 53286 8130 53338
rect 8130 53286 8142 53338
rect 8142 53286 8172 53338
rect 8196 53286 8206 53338
rect 8206 53286 8252 53338
rect 7956 53284 8012 53286
rect 8036 53284 8092 53286
rect 8116 53284 8172 53286
rect 8196 53284 8252 53286
rect 7956 52250 8012 52252
rect 8036 52250 8092 52252
rect 8116 52250 8172 52252
rect 8196 52250 8252 52252
rect 7956 52198 8002 52250
rect 8002 52198 8012 52250
rect 8036 52198 8066 52250
rect 8066 52198 8078 52250
rect 8078 52198 8092 52250
rect 8116 52198 8130 52250
rect 8130 52198 8142 52250
rect 8142 52198 8172 52250
rect 8196 52198 8206 52250
rect 8206 52198 8252 52250
rect 7956 52196 8012 52198
rect 8036 52196 8092 52198
rect 8116 52196 8172 52198
rect 8196 52196 8252 52198
rect 7956 51162 8012 51164
rect 8036 51162 8092 51164
rect 8116 51162 8172 51164
rect 8196 51162 8252 51164
rect 7956 51110 8002 51162
rect 8002 51110 8012 51162
rect 8036 51110 8066 51162
rect 8066 51110 8078 51162
rect 8078 51110 8092 51162
rect 8116 51110 8130 51162
rect 8130 51110 8142 51162
rect 8142 51110 8172 51162
rect 8196 51110 8206 51162
rect 8206 51110 8252 51162
rect 7956 51108 8012 51110
rect 8036 51108 8092 51110
rect 8116 51108 8172 51110
rect 8196 51108 8252 51110
rect 7956 50074 8012 50076
rect 8036 50074 8092 50076
rect 8116 50074 8172 50076
rect 8196 50074 8252 50076
rect 7956 50022 8002 50074
rect 8002 50022 8012 50074
rect 8036 50022 8066 50074
rect 8066 50022 8078 50074
rect 8078 50022 8092 50074
rect 8116 50022 8130 50074
rect 8130 50022 8142 50074
rect 8142 50022 8172 50074
rect 8196 50022 8206 50074
rect 8206 50022 8252 50074
rect 7956 50020 8012 50022
rect 8036 50020 8092 50022
rect 8116 50020 8172 50022
rect 8196 50020 8252 50022
rect 7956 48986 8012 48988
rect 8036 48986 8092 48988
rect 8116 48986 8172 48988
rect 8196 48986 8252 48988
rect 7956 48934 8002 48986
rect 8002 48934 8012 48986
rect 8036 48934 8066 48986
rect 8066 48934 8078 48986
rect 8078 48934 8092 48986
rect 8116 48934 8130 48986
rect 8130 48934 8142 48986
rect 8142 48934 8172 48986
rect 8196 48934 8206 48986
rect 8206 48934 8252 48986
rect 7956 48932 8012 48934
rect 8036 48932 8092 48934
rect 8116 48932 8172 48934
rect 8196 48932 8252 48934
rect 7956 47898 8012 47900
rect 8036 47898 8092 47900
rect 8116 47898 8172 47900
rect 8196 47898 8252 47900
rect 7956 47846 8002 47898
rect 8002 47846 8012 47898
rect 8036 47846 8066 47898
rect 8066 47846 8078 47898
rect 8078 47846 8092 47898
rect 8116 47846 8130 47898
rect 8130 47846 8142 47898
rect 8142 47846 8172 47898
rect 8196 47846 8206 47898
rect 8206 47846 8252 47898
rect 7956 47844 8012 47846
rect 8036 47844 8092 47846
rect 8116 47844 8172 47846
rect 8196 47844 8252 47846
rect 7956 46810 8012 46812
rect 8036 46810 8092 46812
rect 8116 46810 8172 46812
rect 8196 46810 8252 46812
rect 7956 46758 8002 46810
rect 8002 46758 8012 46810
rect 8036 46758 8066 46810
rect 8066 46758 8078 46810
rect 8078 46758 8092 46810
rect 8116 46758 8130 46810
rect 8130 46758 8142 46810
rect 8142 46758 8172 46810
rect 8196 46758 8206 46810
rect 8206 46758 8252 46810
rect 7956 46756 8012 46758
rect 8036 46756 8092 46758
rect 8116 46756 8172 46758
rect 8196 46756 8252 46758
rect 7956 45722 8012 45724
rect 8036 45722 8092 45724
rect 8116 45722 8172 45724
rect 8196 45722 8252 45724
rect 7956 45670 8002 45722
rect 8002 45670 8012 45722
rect 8036 45670 8066 45722
rect 8066 45670 8078 45722
rect 8078 45670 8092 45722
rect 8116 45670 8130 45722
rect 8130 45670 8142 45722
rect 8142 45670 8172 45722
rect 8196 45670 8206 45722
rect 8206 45670 8252 45722
rect 7956 45668 8012 45670
rect 8036 45668 8092 45670
rect 8116 45668 8172 45670
rect 8196 45668 8252 45670
rect 7956 44634 8012 44636
rect 8036 44634 8092 44636
rect 8116 44634 8172 44636
rect 8196 44634 8252 44636
rect 7956 44582 8002 44634
rect 8002 44582 8012 44634
rect 8036 44582 8066 44634
rect 8066 44582 8078 44634
rect 8078 44582 8092 44634
rect 8116 44582 8130 44634
rect 8130 44582 8142 44634
rect 8142 44582 8172 44634
rect 8196 44582 8206 44634
rect 8206 44582 8252 44634
rect 7956 44580 8012 44582
rect 8036 44580 8092 44582
rect 8116 44580 8172 44582
rect 8196 44580 8252 44582
rect 7956 43546 8012 43548
rect 8036 43546 8092 43548
rect 8116 43546 8172 43548
rect 8196 43546 8252 43548
rect 7956 43494 8002 43546
rect 8002 43494 8012 43546
rect 8036 43494 8066 43546
rect 8066 43494 8078 43546
rect 8078 43494 8092 43546
rect 8116 43494 8130 43546
rect 8130 43494 8142 43546
rect 8142 43494 8172 43546
rect 8196 43494 8206 43546
rect 8206 43494 8252 43546
rect 7956 43492 8012 43494
rect 8036 43492 8092 43494
rect 8116 43492 8172 43494
rect 8196 43492 8252 43494
rect 7956 42458 8012 42460
rect 8036 42458 8092 42460
rect 8116 42458 8172 42460
rect 8196 42458 8252 42460
rect 7956 42406 8002 42458
rect 8002 42406 8012 42458
rect 8036 42406 8066 42458
rect 8066 42406 8078 42458
rect 8078 42406 8092 42458
rect 8116 42406 8130 42458
rect 8130 42406 8142 42458
rect 8142 42406 8172 42458
rect 8196 42406 8206 42458
rect 8206 42406 8252 42458
rect 7956 42404 8012 42406
rect 8036 42404 8092 42406
rect 8116 42404 8172 42406
rect 8196 42404 8252 42406
rect 7956 41370 8012 41372
rect 8036 41370 8092 41372
rect 8116 41370 8172 41372
rect 8196 41370 8252 41372
rect 7956 41318 8002 41370
rect 8002 41318 8012 41370
rect 8036 41318 8066 41370
rect 8066 41318 8078 41370
rect 8078 41318 8092 41370
rect 8116 41318 8130 41370
rect 8130 41318 8142 41370
rect 8142 41318 8172 41370
rect 8196 41318 8206 41370
rect 8206 41318 8252 41370
rect 7956 41316 8012 41318
rect 8036 41316 8092 41318
rect 8116 41316 8172 41318
rect 8196 41316 8252 41318
rect 7956 40282 8012 40284
rect 8036 40282 8092 40284
rect 8116 40282 8172 40284
rect 8196 40282 8252 40284
rect 7956 40230 8002 40282
rect 8002 40230 8012 40282
rect 8036 40230 8066 40282
rect 8066 40230 8078 40282
rect 8078 40230 8092 40282
rect 8116 40230 8130 40282
rect 8130 40230 8142 40282
rect 8142 40230 8172 40282
rect 8196 40230 8206 40282
rect 8206 40230 8252 40282
rect 7956 40228 8012 40230
rect 8036 40228 8092 40230
rect 8116 40228 8172 40230
rect 8196 40228 8252 40230
rect 7956 39194 8012 39196
rect 8036 39194 8092 39196
rect 8116 39194 8172 39196
rect 8196 39194 8252 39196
rect 7956 39142 8002 39194
rect 8002 39142 8012 39194
rect 8036 39142 8066 39194
rect 8066 39142 8078 39194
rect 8078 39142 8092 39194
rect 8116 39142 8130 39194
rect 8130 39142 8142 39194
rect 8142 39142 8172 39194
rect 8196 39142 8206 39194
rect 8206 39142 8252 39194
rect 7956 39140 8012 39142
rect 8036 39140 8092 39142
rect 8116 39140 8172 39142
rect 8196 39140 8252 39142
rect 7956 38106 8012 38108
rect 8036 38106 8092 38108
rect 8116 38106 8172 38108
rect 8196 38106 8252 38108
rect 7956 38054 8002 38106
rect 8002 38054 8012 38106
rect 8036 38054 8066 38106
rect 8066 38054 8078 38106
rect 8078 38054 8092 38106
rect 8116 38054 8130 38106
rect 8130 38054 8142 38106
rect 8142 38054 8172 38106
rect 8196 38054 8206 38106
rect 8206 38054 8252 38106
rect 7956 38052 8012 38054
rect 8036 38052 8092 38054
rect 8116 38052 8172 38054
rect 8196 38052 8252 38054
rect 7956 37018 8012 37020
rect 8036 37018 8092 37020
rect 8116 37018 8172 37020
rect 8196 37018 8252 37020
rect 7956 36966 8002 37018
rect 8002 36966 8012 37018
rect 8036 36966 8066 37018
rect 8066 36966 8078 37018
rect 8078 36966 8092 37018
rect 8116 36966 8130 37018
rect 8130 36966 8142 37018
rect 8142 36966 8172 37018
rect 8196 36966 8206 37018
rect 8206 36966 8252 37018
rect 7956 36964 8012 36966
rect 8036 36964 8092 36966
rect 8116 36964 8172 36966
rect 8196 36964 8252 36966
rect 7956 35930 8012 35932
rect 8036 35930 8092 35932
rect 8116 35930 8172 35932
rect 8196 35930 8252 35932
rect 7956 35878 8002 35930
rect 8002 35878 8012 35930
rect 8036 35878 8066 35930
rect 8066 35878 8078 35930
rect 8078 35878 8092 35930
rect 8116 35878 8130 35930
rect 8130 35878 8142 35930
rect 8142 35878 8172 35930
rect 8196 35878 8206 35930
rect 8206 35878 8252 35930
rect 7956 35876 8012 35878
rect 8036 35876 8092 35878
rect 8116 35876 8172 35878
rect 8196 35876 8252 35878
rect 7956 34842 8012 34844
rect 8036 34842 8092 34844
rect 8116 34842 8172 34844
rect 8196 34842 8252 34844
rect 7956 34790 8002 34842
rect 8002 34790 8012 34842
rect 8036 34790 8066 34842
rect 8066 34790 8078 34842
rect 8078 34790 8092 34842
rect 8116 34790 8130 34842
rect 8130 34790 8142 34842
rect 8142 34790 8172 34842
rect 8196 34790 8206 34842
rect 8206 34790 8252 34842
rect 7956 34788 8012 34790
rect 8036 34788 8092 34790
rect 8116 34788 8172 34790
rect 8196 34788 8252 34790
rect 9770 44684 9772 44704
rect 9772 44684 9824 44704
rect 9824 44684 9826 44704
rect 9770 44648 9826 44684
rect 10230 44240 10286 44296
rect 7956 33754 8012 33756
rect 8036 33754 8092 33756
rect 8116 33754 8172 33756
rect 8196 33754 8252 33756
rect 7956 33702 8002 33754
rect 8002 33702 8012 33754
rect 8036 33702 8066 33754
rect 8066 33702 8078 33754
rect 8078 33702 8092 33754
rect 8116 33702 8130 33754
rect 8130 33702 8142 33754
rect 8142 33702 8172 33754
rect 8196 33702 8206 33754
rect 8206 33702 8252 33754
rect 7956 33700 8012 33702
rect 8036 33700 8092 33702
rect 8116 33700 8172 33702
rect 8196 33700 8252 33702
rect 7010 19216 7066 19272
rect 7956 32666 8012 32668
rect 8036 32666 8092 32668
rect 8116 32666 8172 32668
rect 8196 32666 8252 32668
rect 7956 32614 8002 32666
rect 8002 32614 8012 32666
rect 8036 32614 8066 32666
rect 8066 32614 8078 32666
rect 8078 32614 8092 32666
rect 8116 32614 8130 32666
rect 8130 32614 8142 32666
rect 8142 32614 8172 32666
rect 8196 32614 8206 32666
rect 8206 32614 8252 32666
rect 7956 32612 8012 32614
rect 8036 32612 8092 32614
rect 8116 32612 8172 32614
rect 8196 32612 8252 32614
rect 7956 31578 8012 31580
rect 8036 31578 8092 31580
rect 8116 31578 8172 31580
rect 8196 31578 8252 31580
rect 7956 31526 8002 31578
rect 8002 31526 8012 31578
rect 8036 31526 8066 31578
rect 8066 31526 8078 31578
rect 8078 31526 8092 31578
rect 8116 31526 8130 31578
rect 8130 31526 8142 31578
rect 8142 31526 8172 31578
rect 8196 31526 8206 31578
rect 8206 31526 8252 31578
rect 7956 31524 8012 31526
rect 8036 31524 8092 31526
rect 8116 31524 8172 31526
rect 8196 31524 8252 31526
rect 7956 30490 8012 30492
rect 8036 30490 8092 30492
rect 8116 30490 8172 30492
rect 8196 30490 8252 30492
rect 7956 30438 8002 30490
rect 8002 30438 8012 30490
rect 8036 30438 8066 30490
rect 8066 30438 8078 30490
rect 8078 30438 8092 30490
rect 8116 30438 8130 30490
rect 8130 30438 8142 30490
rect 8142 30438 8172 30490
rect 8196 30438 8206 30490
rect 8206 30438 8252 30490
rect 7956 30436 8012 30438
rect 8036 30436 8092 30438
rect 8116 30436 8172 30438
rect 8196 30436 8252 30438
rect 7956 29402 8012 29404
rect 8036 29402 8092 29404
rect 8116 29402 8172 29404
rect 8196 29402 8252 29404
rect 7956 29350 8002 29402
rect 8002 29350 8012 29402
rect 8036 29350 8066 29402
rect 8066 29350 8078 29402
rect 8078 29350 8092 29402
rect 8116 29350 8130 29402
rect 8130 29350 8142 29402
rect 8142 29350 8172 29402
rect 8196 29350 8206 29402
rect 8206 29350 8252 29402
rect 7956 29348 8012 29350
rect 8036 29348 8092 29350
rect 8116 29348 8172 29350
rect 8196 29348 8252 29350
rect 7956 28314 8012 28316
rect 8036 28314 8092 28316
rect 8116 28314 8172 28316
rect 8196 28314 8252 28316
rect 7956 28262 8002 28314
rect 8002 28262 8012 28314
rect 8036 28262 8066 28314
rect 8066 28262 8078 28314
rect 8078 28262 8092 28314
rect 8116 28262 8130 28314
rect 8130 28262 8142 28314
rect 8142 28262 8172 28314
rect 8196 28262 8206 28314
rect 8206 28262 8252 28314
rect 7956 28260 8012 28262
rect 8036 28260 8092 28262
rect 8116 28260 8172 28262
rect 8196 28260 8252 28262
rect 7956 27226 8012 27228
rect 8036 27226 8092 27228
rect 8116 27226 8172 27228
rect 8196 27226 8252 27228
rect 7956 27174 8002 27226
rect 8002 27174 8012 27226
rect 8036 27174 8066 27226
rect 8066 27174 8078 27226
rect 8078 27174 8092 27226
rect 8116 27174 8130 27226
rect 8130 27174 8142 27226
rect 8142 27174 8172 27226
rect 8196 27174 8206 27226
rect 8206 27174 8252 27226
rect 7956 27172 8012 27174
rect 8036 27172 8092 27174
rect 8116 27172 8172 27174
rect 8196 27172 8252 27174
rect 7956 26138 8012 26140
rect 8036 26138 8092 26140
rect 8116 26138 8172 26140
rect 8196 26138 8252 26140
rect 7956 26086 8002 26138
rect 8002 26086 8012 26138
rect 8036 26086 8066 26138
rect 8066 26086 8078 26138
rect 8078 26086 8092 26138
rect 8116 26086 8130 26138
rect 8130 26086 8142 26138
rect 8142 26086 8172 26138
rect 8196 26086 8206 26138
rect 8206 26086 8252 26138
rect 7956 26084 8012 26086
rect 8036 26084 8092 26086
rect 8116 26084 8172 26086
rect 8196 26084 8252 26086
rect 7956 25050 8012 25052
rect 8036 25050 8092 25052
rect 8116 25050 8172 25052
rect 8196 25050 8252 25052
rect 7956 24998 8002 25050
rect 8002 24998 8012 25050
rect 8036 24998 8066 25050
rect 8066 24998 8078 25050
rect 8078 24998 8092 25050
rect 8116 24998 8130 25050
rect 8130 24998 8142 25050
rect 8142 24998 8172 25050
rect 8196 24998 8206 25050
rect 8206 24998 8252 25050
rect 7956 24996 8012 24998
rect 8036 24996 8092 24998
rect 8116 24996 8172 24998
rect 8196 24996 8252 24998
rect 12956 53882 13012 53884
rect 13036 53882 13092 53884
rect 13116 53882 13172 53884
rect 13196 53882 13252 53884
rect 12956 53830 13002 53882
rect 13002 53830 13012 53882
rect 13036 53830 13066 53882
rect 13066 53830 13078 53882
rect 13078 53830 13092 53882
rect 13116 53830 13130 53882
rect 13130 53830 13142 53882
rect 13142 53830 13172 53882
rect 13196 53830 13206 53882
rect 13206 53830 13252 53882
rect 12956 53828 13012 53830
rect 13036 53828 13092 53830
rect 13116 53828 13172 53830
rect 13196 53828 13252 53830
rect 12956 52794 13012 52796
rect 13036 52794 13092 52796
rect 13116 52794 13172 52796
rect 13196 52794 13252 52796
rect 12956 52742 13002 52794
rect 13002 52742 13012 52794
rect 13036 52742 13066 52794
rect 13066 52742 13078 52794
rect 13078 52742 13092 52794
rect 13116 52742 13130 52794
rect 13130 52742 13142 52794
rect 13142 52742 13172 52794
rect 13196 52742 13206 52794
rect 13206 52742 13252 52794
rect 12956 52740 13012 52742
rect 13036 52740 13092 52742
rect 13116 52740 13172 52742
rect 13196 52740 13252 52742
rect 11610 44684 11612 44704
rect 11612 44684 11664 44704
rect 11664 44684 11666 44704
rect 11610 44648 11666 44684
rect 11610 44260 11666 44296
rect 11610 44240 11612 44260
rect 11612 44240 11664 44260
rect 11664 44240 11666 44260
rect 15750 53932 15752 53952
rect 15752 53932 15804 53952
rect 15804 53932 15806 53952
rect 15750 53896 15806 53932
rect 13634 52556 13690 52592
rect 13634 52536 13636 52556
rect 13636 52536 13688 52556
rect 13688 52536 13690 52556
rect 14002 52536 14058 52592
rect 12956 51706 13012 51708
rect 13036 51706 13092 51708
rect 13116 51706 13172 51708
rect 13196 51706 13252 51708
rect 12956 51654 13002 51706
rect 13002 51654 13012 51706
rect 13036 51654 13066 51706
rect 13066 51654 13078 51706
rect 13078 51654 13092 51706
rect 13116 51654 13130 51706
rect 13130 51654 13142 51706
rect 13142 51654 13172 51706
rect 13196 51654 13206 51706
rect 13206 51654 13252 51706
rect 12956 51652 13012 51654
rect 13036 51652 13092 51654
rect 13116 51652 13172 51654
rect 13196 51652 13252 51654
rect 12956 50618 13012 50620
rect 13036 50618 13092 50620
rect 13116 50618 13172 50620
rect 13196 50618 13252 50620
rect 12956 50566 13002 50618
rect 13002 50566 13012 50618
rect 13036 50566 13066 50618
rect 13066 50566 13078 50618
rect 13078 50566 13092 50618
rect 13116 50566 13130 50618
rect 13130 50566 13142 50618
rect 13142 50566 13172 50618
rect 13196 50566 13206 50618
rect 13206 50566 13252 50618
rect 12956 50564 13012 50566
rect 13036 50564 13092 50566
rect 13116 50564 13172 50566
rect 13196 50564 13252 50566
rect 12956 49530 13012 49532
rect 13036 49530 13092 49532
rect 13116 49530 13172 49532
rect 13196 49530 13252 49532
rect 12956 49478 13002 49530
rect 13002 49478 13012 49530
rect 13036 49478 13066 49530
rect 13066 49478 13078 49530
rect 13078 49478 13092 49530
rect 13116 49478 13130 49530
rect 13130 49478 13142 49530
rect 13142 49478 13172 49530
rect 13196 49478 13206 49530
rect 13206 49478 13252 49530
rect 12956 49476 13012 49478
rect 13036 49476 13092 49478
rect 13116 49476 13172 49478
rect 13196 49476 13252 49478
rect 12956 48442 13012 48444
rect 13036 48442 13092 48444
rect 13116 48442 13172 48444
rect 13196 48442 13252 48444
rect 12956 48390 13002 48442
rect 13002 48390 13012 48442
rect 13036 48390 13066 48442
rect 13066 48390 13078 48442
rect 13078 48390 13092 48442
rect 13116 48390 13130 48442
rect 13130 48390 13142 48442
rect 13142 48390 13172 48442
rect 13196 48390 13206 48442
rect 13206 48390 13252 48442
rect 12956 48388 13012 48390
rect 13036 48388 13092 48390
rect 13116 48388 13172 48390
rect 13196 48388 13252 48390
rect 11794 45328 11850 45384
rect 10598 37324 10654 37360
rect 10598 37304 10600 37324
rect 10600 37304 10652 37324
rect 10652 37304 10654 37324
rect 10138 36760 10194 36816
rect 7956 23962 8012 23964
rect 8036 23962 8092 23964
rect 8116 23962 8172 23964
rect 8196 23962 8252 23964
rect 7956 23910 8002 23962
rect 8002 23910 8012 23962
rect 8036 23910 8066 23962
rect 8066 23910 8078 23962
rect 8078 23910 8092 23962
rect 8116 23910 8130 23962
rect 8130 23910 8142 23962
rect 8142 23910 8172 23962
rect 8196 23910 8206 23962
rect 8206 23910 8252 23962
rect 7956 23908 8012 23910
rect 8036 23908 8092 23910
rect 8116 23908 8172 23910
rect 8196 23908 8252 23910
rect 7956 22874 8012 22876
rect 8036 22874 8092 22876
rect 8116 22874 8172 22876
rect 8196 22874 8252 22876
rect 7956 22822 8002 22874
rect 8002 22822 8012 22874
rect 8036 22822 8066 22874
rect 8066 22822 8078 22874
rect 8078 22822 8092 22874
rect 8116 22822 8130 22874
rect 8130 22822 8142 22874
rect 8142 22822 8172 22874
rect 8196 22822 8206 22874
rect 8206 22822 8252 22874
rect 7956 22820 8012 22822
rect 8036 22820 8092 22822
rect 8116 22820 8172 22822
rect 8196 22820 8252 22822
rect 7956 21786 8012 21788
rect 8036 21786 8092 21788
rect 8116 21786 8172 21788
rect 8196 21786 8252 21788
rect 7956 21734 8002 21786
rect 8002 21734 8012 21786
rect 8036 21734 8066 21786
rect 8066 21734 8078 21786
rect 8078 21734 8092 21786
rect 8116 21734 8130 21786
rect 8130 21734 8142 21786
rect 8142 21734 8172 21786
rect 8196 21734 8206 21786
rect 8206 21734 8252 21786
rect 7956 21732 8012 21734
rect 8036 21732 8092 21734
rect 8116 21732 8172 21734
rect 8196 21732 8252 21734
rect 7956 20698 8012 20700
rect 8036 20698 8092 20700
rect 8116 20698 8172 20700
rect 8196 20698 8252 20700
rect 7956 20646 8002 20698
rect 8002 20646 8012 20698
rect 8036 20646 8066 20698
rect 8066 20646 8078 20698
rect 8078 20646 8092 20698
rect 8116 20646 8130 20698
rect 8130 20646 8142 20698
rect 8142 20646 8172 20698
rect 8196 20646 8206 20698
rect 8206 20646 8252 20698
rect 7956 20644 8012 20646
rect 8036 20644 8092 20646
rect 8116 20644 8172 20646
rect 8196 20644 8252 20646
rect 7956 19610 8012 19612
rect 8036 19610 8092 19612
rect 8116 19610 8172 19612
rect 8196 19610 8252 19612
rect 7956 19558 8002 19610
rect 8002 19558 8012 19610
rect 8036 19558 8066 19610
rect 8066 19558 8078 19610
rect 8078 19558 8092 19610
rect 8116 19558 8130 19610
rect 8130 19558 8142 19610
rect 8142 19558 8172 19610
rect 8196 19558 8206 19610
rect 8206 19558 8252 19610
rect 7956 19556 8012 19558
rect 8036 19556 8092 19558
rect 8116 19556 8172 19558
rect 8196 19556 8252 19558
rect 7956 18522 8012 18524
rect 8036 18522 8092 18524
rect 8116 18522 8172 18524
rect 8196 18522 8252 18524
rect 7956 18470 8002 18522
rect 8002 18470 8012 18522
rect 8036 18470 8066 18522
rect 8066 18470 8078 18522
rect 8078 18470 8092 18522
rect 8116 18470 8130 18522
rect 8130 18470 8142 18522
rect 8142 18470 8172 18522
rect 8196 18470 8206 18522
rect 8206 18470 8252 18522
rect 7956 18468 8012 18470
rect 8036 18468 8092 18470
rect 8116 18468 8172 18470
rect 8196 18468 8252 18470
rect 7956 17434 8012 17436
rect 8036 17434 8092 17436
rect 8116 17434 8172 17436
rect 8196 17434 8252 17436
rect 7956 17382 8002 17434
rect 8002 17382 8012 17434
rect 8036 17382 8066 17434
rect 8066 17382 8078 17434
rect 8078 17382 8092 17434
rect 8116 17382 8130 17434
rect 8130 17382 8142 17434
rect 8142 17382 8172 17434
rect 8196 17382 8206 17434
rect 8206 17382 8252 17434
rect 7956 17380 8012 17382
rect 8036 17380 8092 17382
rect 8116 17380 8172 17382
rect 8196 17380 8252 17382
rect 7956 16346 8012 16348
rect 8036 16346 8092 16348
rect 8116 16346 8172 16348
rect 8196 16346 8252 16348
rect 7956 16294 8002 16346
rect 8002 16294 8012 16346
rect 8036 16294 8066 16346
rect 8066 16294 8078 16346
rect 8078 16294 8092 16346
rect 8116 16294 8130 16346
rect 8130 16294 8142 16346
rect 8142 16294 8172 16346
rect 8196 16294 8206 16346
rect 8206 16294 8252 16346
rect 7956 16292 8012 16294
rect 8036 16292 8092 16294
rect 8116 16292 8172 16294
rect 8196 16292 8252 16294
rect 7956 15258 8012 15260
rect 8036 15258 8092 15260
rect 8116 15258 8172 15260
rect 8196 15258 8252 15260
rect 7956 15206 8002 15258
rect 8002 15206 8012 15258
rect 8036 15206 8066 15258
rect 8066 15206 8078 15258
rect 8078 15206 8092 15258
rect 8116 15206 8130 15258
rect 8130 15206 8142 15258
rect 8142 15206 8172 15258
rect 8196 15206 8206 15258
rect 8206 15206 8252 15258
rect 7956 15204 8012 15206
rect 8036 15204 8092 15206
rect 8116 15204 8172 15206
rect 8196 15204 8252 15206
rect 7956 14170 8012 14172
rect 8036 14170 8092 14172
rect 8116 14170 8172 14172
rect 8196 14170 8252 14172
rect 7956 14118 8002 14170
rect 8002 14118 8012 14170
rect 8036 14118 8066 14170
rect 8066 14118 8078 14170
rect 8078 14118 8092 14170
rect 8116 14118 8130 14170
rect 8130 14118 8142 14170
rect 8142 14118 8172 14170
rect 8196 14118 8206 14170
rect 8206 14118 8252 14170
rect 7956 14116 8012 14118
rect 8036 14116 8092 14118
rect 8116 14116 8172 14118
rect 8196 14116 8252 14118
rect 7956 13082 8012 13084
rect 8036 13082 8092 13084
rect 8116 13082 8172 13084
rect 8196 13082 8252 13084
rect 7956 13030 8002 13082
rect 8002 13030 8012 13082
rect 8036 13030 8066 13082
rect 8066 13030 8078 13082
rect 8078 13030 8092 13082
rect 8116 13030 8130 13082
rect 8130 13030 8142 13082
rect 8142 13030 8172 13082
rect 8196 13030 8206 13082
rect 8206 13030 8252 13082
rect 7956 13028 8012 13030
rect 8036 13028 8092 13030
rect 8116 13028 8172 13030
rect 8196 13028 8252 13030
rect 7956 11994 8012 11996
rect 8036 11994 8092 11996
rect 8116 11994 8172 11996
rect 8196 11994 8252 11996
rect 7956 11942 8002 11994
rect 8002 11942 8012 11994
rect 8036 11942 8066 11994
rect 8066 11942 8078 11994
rect 8078 11942 8092 11994
rect 8116 11942 8130 11994
rect 8130 11942 8142 11994
rect 8142 11942 8172 11994
rect 8196 11942 8206 11994
rect 8206 11942 8252 11994
rect 7956 11940 8012 11942
rect 8036 11940 8092 11942
rect 8116 11940 8172 11942
rect 8196 11940 8252 11942
rect 7956 10906 8012 10908
rect 8036 10906 8092 10908
rect 8116 10906 8172 10908
rect 8196 10906 8252 10908
rect 7956 10854 8002 10906
rect 8002 10854 8012 10906
rect 8036 10854 8066 10906
rect 8066 10854 8078 10906
rect 8078 10854 8092 10906
rect 8116 10854 8130 10906
rect 8130 10854 8142 10906
rect 8142 10854 8172 10906
rect 8196 10854 8206 10906
rect 8206 10854 8252 10906
rect 7956 10852 8012 10854
rect 8036 10852 8092 10854
rect 8116 10852 8172 10854
rect 8196 10852 8252 10854
rect 7956 9818 8012 9820
rect 8036 9818 8092 9820
rect 8116 9818 8172 9820
rect 8196 9818 8252 9820
rect 7956 9766 8002 9818
rect 8002 9766 8012 9818
rect 8036 9766 8066 9818
rect 8066 9766 8078 9818
rect 8078 9766 8092 9818
rect 8116 9766 8130 9818
rect 8130 9766 8142 9818
rect 8142 9766 8172 9818
rect 8196 9766 8206 9818
rect 8206 9766 8252 9818
rect 7956 9764 8012 9766
rect 8036 9764 8092 9766
rect 8116 9764 8172 9766
rect 8196 9764 8252 9766
rect 7956 8730 8012 8732
rect 8036 8730 8092 8732
rect 8116 8730 8172 8732
rect 8196 8730 8252 8732
rect 7956 8678 8002 8730
rect 8002 8678 8012 8730
rect 8036 8678 8066 8730
rect 8066 8678 8078 8730
rect 8078 8678 8092 8730
rect 8116 8678 8130 8730
rect 8130 8678 8142 8730
rect 8142 8678 8172 8730
rect 8196 8678 8206 8730
rect 8206 8678 8252 8730
rect 7956 8676 8012 8678
rect 8036 8676 8092 8678
rect 8116 8676 8172 8678
rect 8196 8676 8252 8678
rect 7956 7642 8012 7644
rect 8036 7642 8092 7644
rect 8116 7642 8172 7644
rect 8196 7642 8252 7644
rect 7956 7590 8002 7642
rect 8002 7590 8012 7642
rect 8036 7590 8066 7642
rect 8066 7590 8078 7642
rect 8078 7590 8092 7642
rect 8116 7590 8130 7642
rect 8130 7590 8142 7642
rect 8142 7590 8172 7642
rect 8196 7590 8206 7642
rect 8206 7590 8252 7642
rect 7956 7588 8012 7590
rect 8036 7588 8092 7590
rect 8116 7588 8172 7590
rect 8196 7588 8252 7590
rect 7956 6554 8012 6556
rect 8036 6554 8092 6556
rect 8116 6554 8172 6556
rect 8196 6554 8252 6556
rect 7956 6502 8002 6554
rect 8002 6502 8012 6554
rect 8036 6502 8066 6554
rect 8066 6502 8078 6554
rect 8078 6502 8092 6554
rect 8116 6502 8130 6554
rect 8130 6502 8142 6554
rect 8142 6502 8172 6554
rect 8196 6502 8206 6554
rect 8206 6502 8252 6554
rect 7956 6500 8012 6502
rect 8036 6500 8092 6502
rect 8116 6500 8172 6502
rect 8196 6500 8252 6502
rect 7956 5466 8012 5468
rect 8036 5466 8092 5468
rect 8116 5466 8172 5468
rect 8196 5466 8252 5468
rect 7956 5414 8002 5466
rect 8002 5414 8012 5466
rect 8036 5414 8066 5466
rect 8066 5414 8078 5466
rect 8078 5414 8092 5466
rect 8116 5414 8130 5466
rect 8130 5414 8142 5466
rect 8142 5414 8172 5466
rect 8196 5414 8206 5466
rect 8206 5414 8252 5466
rect 7956 5412 8012 5414
rect 8036 5412 8092 5414
rect 8116 5412 8172 5414
rect 8196 5412 8252 5414
rect 7956 4378 8012 4380
rect 8036 4378 8092 4380
rect 8116 4378 8172 4380
rect 8196 4378 8252 4380
rect 7956 4326 8002 4378
rect 8002 4326 8012 4378
rect 8036 4326 8066 4378
rect 8066 4326 8078 4378
rect 8078 4326 8092 4378
rect 8116 4326 8130 4378
rect 8130 4326 8142 4378
rect 8142 4326 8172 4378
rect 8196 4326 8206 4378
rect 8206 4326 8252 4378
rect 7956 4324 8012 4326
rect 8036 4324 8092 4326
rect 8116 4324 8172 4326
rect 8196 4324 8252 4326
rect 8482 4120 8538 4176
rect 7956 3290 8012 3292
rect 8036 3290 8092 3292
rect 8116 3290 8172 3292
rect 8196 3290 8252 3292
rect 7956 3238 8002 3290
rect 8002 3238 8012 3290
rect 8036 3238 8066 3290
rect 8066 3238 8078 3290
rect 8078 3238 8092 3290
rect 8116 3238 8130 3290
rect 8130 3238 8142 3290
rect 8142 3238 8172 3290
rect 8196 3238 8206 3290
rect 8206 3238 8252 3290
rect 7956 3236 8012 3238
rect 8036 3236 8092 3238
rect 8116 3236 8172 3238
rect 8196 3236 8252 3238
rect 7956 2202 8012 2204
rect 8036 2202 8092 2204
rect 8116 2202 8172 2204
rect 8196 2202 8252 2204
rect 7956 2150 8002 2202
rect 8002 2150 8012 2202
rect 8036 2150 8066 2202
rect 8066 2150 8078 2202
rect 8078 2150 8092 2202
rect 8116 2150 8130 2202
rect 8130 2150 8142 2202
rect 8142 2150 8172 2202
rect 8196 2150 8206 2202
rect 8206 2150 8252 2202
rect 7956 2148 8012 2150
rect 8036 2148 8092 2150
rect 8116 2148 8172 2150
rect 8196 2148 8252 2150
rect 11242 36372 11298 36408
rect 11242 36352 11244 36372
rect 11244 36352 11296 36372
rect 11296 36352 11298 36372
rect 11334 32972 11390 33008
rect 11334 32952 11336 32972
rect 11336 32952 11388 32972
rect 11388 32952 11390 32972
rect 11978 30796 12034 30832
rect 11978 30776 11980 30796
rect 11980 30776 12032 30796
rect 12032 30776 12034 30796
rect 12956 47354 13012 47356
rect 13036 47354 13092 47356
rect 13116 47354 13172 47356
rect 13196 47354 13252 47356
rect 12956 47302 13002 47354
rect 13002 47302 13012 47354
rect 13036 47302 13066 47354
rect 13066 47302 13078 47354
rect 13078 47302 13092 47354
rect 13116 47302 13130 47354
rect 13130 47302 13142 47354
rect 13142 47302 13172 47354
rect 13196 47302 13206 47354
rect 13206 47302 13252 47354
rect 12956 47300 13012 47302
rect 13036 47300 13092 47302
rect 13116 47300 13172 47302
rect 13196 47300 13252 47302
rect 12956 46266 13012 46268
rect 13036 46266 13092 46268
rect 13116 46266 13172 46268
rect 13196 46266 13252 46268
rect 12956 46214 13002 46266
rect 13002 46214 13012 46266
rect 13036 46214 13066 46266
rect 13066 46214 13078 46266
rect 13078 46214 13092 46266
rect 13116 46214 13130 46266
rect 13130 46214 13142 46266
rect 13142 46214 13172 46266
rect 13196 46214 13206 46266
rect 13206 46214 13252 46266
rect 12956 46212 13012 46214
rect 13036 46212 13092 46214
rect 13116 46212 13172 46214
rect 13196 46212 13252 46214
rect 12956 45178 13012 45180
rect 13036 45178 13092 45180
rect 13116 45178 13172 45180
rect 13196 45178 13252 45180
rect 12956 45126 13002 45178
rect 13002 45126 13012 45178
rect 13036 45126 13066 45178
rect 13066 45126 13078 45178
rect 13078 45126 13092 45178
rect 13116 45126 13130 45178
rect 13130 45126 13142 45178
rect 13142 45126 13172 45178
rect 13196 45126 13206 45178
rect 13206 45126 13252 45178
rect 12956 45124 13012 45126
rect 13036 45124 13092 45126
rect 13116 45124 13172 45126
rect 13196 45124 13252 45126
rect 12956 44090 13012 44092
rect 13036 44090 13092 44092
rect 13116 44090 13172 44092
rect 13196 44090 13252 44092
rect 12956 44038 13002 44090
rect 13002 44038 13012 44090
rect 13036 44038 13066 44090
rect 13066 44038 13078 44090
rect 13078 44038 13092 44090
rect 13116 44038 13130 44090
rect 13130 44038 13142 44090
rect 13142 44038 13172 44090
rect 13196 44038 13206 44090
rect 13206 44038 13252 44090
rect 12956 44036 13012 44038
rect 13036 44036 13092 44038
rect 13116 44036 13172 44038
rect 13196 44036 13252 44038
rect 12956 43002 13012 43004
rect 13036 43002 13092 43004
rect 13116 43002 13172 43004
rect 13196 43002 13252 43004
rect 12956 42950 13002 43002
rect 13002 42950 13012 43002
rect 13036 42950 13066 43002
rect 13066 42950 13078 43002
rect 13078 42950 13092 43002
rect 13116 42950 13130 43002
rect 13130 42950 13142 43002
rect 13142 42950 13172 43002
rect 13196 42950 13206 43002
rect 13206 42950 13252 43002
rect 12956 42948 13012 42950
rect 13036 42948 13092 42950
rect 13116 42948 13172 42950
rect 13196 42948 13252 42950
rect 12956 41914 13012 41916
rect 13036 41914 13092 41916
rect 13116 41914 13172 41916
rect 13196 41914 13252 41916
rect 12956 41862 13002 41914
rect 13002 41862 13012 41914
rect 13036 41862 13066 41914
rect 13066 41862 13078 41914
rect 13078 41862 13092 41914
rect 13116 41862 13130 41914
rect 13130 41862 13142 41914
rect 13142 41862 13172 41914
rect 13196 41862 13206 41914
rect 13206 41862 13252 41914
rect 12956 41860 13012 41862
rect 13036 41860 13092 41862
rect 13116 41860 13172 41862
rect 13196 41860 13252 41862
rect 12622 38256 12678 38312
rect 12956 40826 13012 40828
rect 13036 40826 13092 40828
rect 13116 40826 13172 40828
rect 13196 40826 13252 40828
rect 12956 40774 13002 40826
rect 13002 40774 13012 40826
rect 13036 40774 13066 40826
rect 13066 40774 13078 40826
rect 13078 40774 13092 40826
rect 13116 40774 13130 40826
rect 13130 40774 13142 40826
rect 13142 40774 13172 40826
rect 13196 40774 13206 40826
rect 13206 40774 13252 40826
rect 12956 40772 13012 40774
rect 13036 40772 13092 40774
rect 13116 40772 13172 40774
rect 13196 40772 13252 40774
rect 12956 39738 13012 39740
rect 13036 39738 13092 39740
rect 13116 39738 13172 39740
rect 13196 39738 13252 39740
rect 12956 39686 13002 39738
rect 13002 39686 13012 39738
rect 13036 39686 13066 39738
rect 13066 39686 13078 39738
rect 13078 39686 13092 39738
rect 13116 39686 13130 39738
rect 13130 39686 13142 39738
rect 13142 39686 13172 39738
rect 13196 39686 13206 39738
rect 13206 39686 13252 39738
rect 12956 39684 13012 39686
rect 13036 39684 13092 39686
rect 13116 39684 13172 39686
rect 13196 39684 13252 39686
rect 12956 38650 13012 38652
rect 13036 38650 13092 38652
rect 13116 38650 13172 38652
rect 13196 38650 13252 38652
rect 12956 38598 13002 38650
rect 13002 38598 13012 38650
rect 13036 38598 13066 38650
rect 13066 38598 13078 38650
rect 13078 38598 13092 38650
rect 13116 38598 13130 38650
rect 13130 38598 13142 38650
rect 13142 38598 13172 38650
rect 13196 38598 13206 38650
rect 13206 38598 13252 38650
rect 12956 38596 13012 38598
rect 13036 38596 13092 38598
rect 13116 38596 13172 38598
rect 13196 38596 13252 38598
rect 12956 37562 13012 37564
rect 13036 37562 13092 37564
rect 13116 37562 13172 37564
rect 13196 37562 13252 37564
rect 12956 37510 13002 37562
rect 13002 37510 13012 37562
rect 13036 37510 13066 37562
rect 13066 37510 13078 37562
rect 13078 37510 13092 37562
rect 13116 37510 13130 37562
rect 13130 37510 13142 37562
rect 13142 37510 13172 37562
rect 13196 37510 13206 37562
rect 13206 37510 13252 37562
rect 12956 37508 13012 37510
rect 13036 37508 13092 37510
rect 13116 37508 13172 37510
rect 13196 37508 13252 37510
rect 12530 35536 12586 35592
rect 13358 37324 13414 37360
rect 13358 37304 13360 37324
rect 13360 37304 13412 37324
rect 13412 37304 13414 37324
rect 12530 33260 12532 33280
rect 12532 33260 12584 33280
rect 12584 33260 12586 33280
rect 12530 33224 12586 33260
rect 12956 36474 13012 36476
rect 13036 36474 13092 36476
rect 13116 36474 13172 36476
rect 13196 36474 13252 36476
rect 12956 36422 13002 36474
rect 13002 36422 13012 36474
rect 13036 36422 13066 36474
rect 13066 36422 13078 36474
rect 13078 36422 13092 36474
rect 13116 36422 13130 36474
rect 13130 36422 13142 36474
rect 13142 36422 13172 36474
rect 13196 36422 13206 36474
rect 13206 36422 13252 36474
rect 12956 36420 13012 36422
rect 13036 36420 13092 36422
rect 13116 36420 13172 36422
rect 13196 36420 13252 36422
rect 12956 35386 13012 35388
rect 13036 35386 13092 35388
rect 13116 35386 13172 35388
rect 13196 35386 13252 35388
rect 12956 35334 13002 35386
rect 13002 35334 13012 35386
rect 13036 35334 13066 35386
rect 13066 35334 13078 35386
rect 13078 35334 13092 35386
rect 13116 35334 13130 35386
rect 13130 35334 13142 35386
rect 13142 35334 13172 35386
rect 13196 35334 13206 35386
rect 13206 35334 13252 35386
rect 12956 35332 13012 35334
rect 13036 35332 13092 35334
rect 13116 35332 13172 35334
rect 13196 35332 13252 35334
rect 12956 34298 13012 34300
rect 13036 34298 13092 34300
rect 13116 34298 13172 34300
rect 13196 34298 13252 34300
rect 12956 34246 13002 34298
rect 13002 34246 13012 34298
rect 13036 34246 13066 34298
rect 13066 34246 13078 34298
rect 13078 34246 13092 34298
rect 13116 34246 13130 34298
rect 13130 34246 13142 34298
rect 13142 34246 13172 34298
rect 13196 34246 13206 34298
rect 13206 34246 13252 34298
rect 12956 34244 13012 34246
rect 13036 34244 13092 34246
rect 13116 34244 13172 34246
rect 13196 34244 13252 34246
rect 13818 35980 13820 36000
rect 13820 35980 13872 36000
rect 13872 35980 13874 36000
rect 13818 35944 13874 35980
rect 13634 35400 13690 35456
rect 12956 33210 13012 33212
rect 13036 33210 13092 33212
rect 13116 33210 13172 33212
rect 13196 33210 13252 33212
rect 12956 33158 13002 33210
rect 13002 33158 13012 33210
rect 13036 33158 13066 33210
rect 13066 33158 13078 33210
rect 13078 33158 13092 33210
rect 13116 33158 13130 33210
rect 13130 33158 13142 33210
rect 13142 33158 13172 33210
rect 13196 33158 13206 33210
rect 13206 33158 13252 33210
rect 12956 33156 13012 33158
rect 13036 33156 13092 33158
rect 13116 33156 13172 33158
rect 13196 33156 13252 33158
rect 13266 32544 13322 32600
rect 12956 32122 13012 32124
rect 13036 32122 13092 32124
rect 13116 32122 13172 32124
rect 13196 32122 13252 32124
rect 12956 32070 13002 32122
rect 13002 32070 13012 32122
rect 13036 32070 13066 32122
rect 13066 32070 13078 32122
rect 13078 32070 13092 32122
rect 13116 32070 13130 32122
rect 13130 32070 13142 32122
rect 13142 32070 13172 32122
rect 13196 32070 13206 32122
rect 13206 32070 13252 32122
rect 12956 32068 13012 32070
rect 13036 32068 13092 32070
rect 13116 32068 13172 32070
rect 13196 32068 13252 32070
rect 11426 24792 11482 24848
rect 11794 23196 11796 23216
rect 11796 23196 11848 23216
rect 11848 23196 11850 23216
rect 11794 23160 11850 23196
rect 12956 31034 13012 31036
rect 13036 31034 13092 31036
rect 13116 31034 13172 31036
rect 13196 31034 13252 31036
rect 12956 30982 13002 31034
rect 13002 30982 13012 31034
rect 13036 30982 13066 31034
rect 13066 30982 13078 31034
rect 13078 30982 13092 31034
rect 13116 30982 13130 31034
rect 13130 30982 13142 31034
rect 13142 30982 13172 31034
rect 13196 30982 13206 31034
rect 13206 30982 13252 31034
rect 12956 30980 13012 30982
rect 13036 30980 13092 30982
rect 13116 30980 13172 30982
rect 13196 30980 13252 30982
rect 12956 29946 13012 29948
rect 13036 29946 13092 29948
rect 13116 29946 13172 29948
rect 13196 29946 13252 29948
rect 12956 29894 13002 29946
rect 13002 29894 13012 29946
rect 13036 29894 13066 29946
rect 13066 29894 13078 29946
rect 13078 29894 13092 29946
rect 13116 29894 13130 29946
rect 13130 29894 13142 29946
rect 13142 29894 13172 29946
rect 13196 29894 13206 29946
rect 13206 29894 13252 29946
rect 12956 29892 13012 29894
rect 13036 29892 13092 29894
rect 13116 29892 13172 29894
rect 13196 29892 13252 29894
rect 12956 28858 13012 28860
rect 13036 28858 13092 28860
rect 13116 28858 13172 28860
rect 13196 28858 13252 28860
rect 12956 28806 13002 28858
rect 13002 28806 13012 28858
rect 13036 28806 13066 28858
rect 13066 28806 13078 28858
rect 13078 28806 13092 28858
rect 13116 28806 13130 28858
rect 13130 28806 13142 28858
rect 13142 28806 13172 28858
rect 13196 28806 13206 28858
rect 13206 28806 13252 28858
rect 12956 28804 13012 28806
rect 13036 28804 13092 28806
rect 13116 28804 13172 28806
rect 13196 28804 13252 28806
rect 12956 27770 13012 27772
rect 13036 27770 13092 27772
rect 13116 27770 13172 27772
rect 13196 27770 13252 27772
rect 12956 27718 13002 27770
rect 13002 27718 13012 27770
rect 13036 27718 13066 27770
rect 13066 27718 13078 27770
rect 13078 27718 13092 27770
rect 13116 27718 13130 27770
rect 13130 27718 13142 27770
rect 13142 27718 13172 27770
rect 13196 27718 13206 27770
rect 13206 27718 13252 27770
rect 12956 27716 13012 27718
rect 13036 27716 13092 27718
rect 13116 27716 13172 27718
rect 13196 27716 13252 27718
rect 12956 26682 13012 26684
rect 13036 26682 13092 26684
rect 13116 26682 13172 26684
rect 13196 26682 13252 26684
rect 12956 26630 13002 26682
rect 13002 26630 13012 26682
rect 13036 26630 13066 26682
rect 13066 26630 13078 26682
rect 13078 26630 13092 26682
rect 13116 26630 13130 26682
rect 13130 26630 13142 26682
rect 13142 26630 13172 26682
rect 13196 26630 13206 26682
rect 13206 26630 13252 26682
rect 12956 26628 13012 26630
rect 13036 26628 13092 26630
rect 13116 26628 13172 26630
rect 13196 26628 13252 26630
rect 12956 25594 13012 25596
rect 13036 25594 13092 25596
rect 13116 25594 13172 25596
rect 13196 25594 13252 25596
rect 12956 25542 13002 25594
rect 13002 25542 13012 25594
rect 13036 25542 13066 25594
rect 13066 25542 13078 25594
rect 13078 25542 13092 25594
rect 13116 25542 13130 25594
rect 13130 25542 13142 25594
rect 13142 25542 13172 25594
rect 13196 25542 13206 25594
rect 13206 25542 13252 25594
rect 12956 25540 13012 25542
rect 13036 25540 13092 25542
rect 13116 25540 13172 25542
rect 13196 25540 13252 25542
rect 12956 24506 13012 24508
rect 13036 24506 13092 24508
rect 13116 24506 13172 24508
rect 13196 24506 13252 24508
rect 12956 24454 13002 24506
rect 13002 24454 13012 24506
rect 13036 24454 13066 24506
rect 13066 24454 13078 24506
rect 13078 24454 13092 24506
rect 13116 24454 13130 24506
rect 13130 24454 13142 24506
rect 13142 24454 13172 24506
rect 13196 24454 13206 24506
rect 13206 24454 13252 24506
rect 12956 24452 13012 24454
rect 13036 24452 13092 24454
rect 13116 24452 13172 24454
rect 13196 24452 13252 24454
rect 12956 23418 13012 23420
rect 13036 23418 13092 23420
rect 13116 23418 13172 23420
rect 13196 23418 13252 23420
rect 12956 23366 13002 23418
rect 13002 23366 13012 23418
rect 13036 23366 13066 23418
rect 13066 23366 13078 23418
rect 13078 23366 13092 23418
rect 13116 23366 13130 23418
rect 13130 23366 13142 23418
rect 13142 23366 13172 23418
rect 13196 23366 13206 23418
rect 13206 23366 13252 23418
rect 12956 23364 13012 23366
rect 13036 23364 13092 23366
rect 13116 23364 13172 23366
rect 13196 23364 13252 23366
rect 12438 21528 12494 21584
rect 12346 18300 12348 18320
rect 12348 18300 12400 18320
rect 12400 18300 12402 18320
rect 12346 18264 12402 18300
rect 12956 22330 13012 22332
rect 13036 22330 13092 22332
rect 13116 22330 13172 22332
rect 13196 22330 13252 22332
rect 12956 22278 13002 22330
rect 13002 22278 13012 22330
rect 13036 22278 13066 22330
rect 13066 22278 13078 22330
rect 13078 22278 13092 22330
rect 13116 22278 13130 22330
rect 13130 22278 13142 22330
rect 13142 22278 13172 22330
rect 13196 22278 13206 22330
rect 13206 22278 13252 22330
rect 12956 22276 13012 22278
rect 13036 22276 13092 22278
rect 13116 22276 13172 22278
rect 13196 22276 13252 22278
rect 12956 21242 13012 21244
rect 13036 21242 13092 21244
rect 13116 21242 13172 21244
rect 13196 21242 13252 21244
rect 12956 21190 13002 21242
rect 13002 21190 13012 21242
rect 13036 21190 13066 21242
rect 13066 21190 13078 21242
rect 13078 21190 13092 21242
rect 13116 21190 13130 21242
rect 13130 21190 13142 21242
rect 13142 21190 13172 21242
rect 13196 21190 13206 21242
rect 13206 21190 13252 21242
rect 12956 21188 13012 21190
rect 13036 21188 13092 21190
rect 13116 21188 13172 21190
rect 13196 21188 13252 21190
rect 12956 20154 13012 20156
rect 13036 20154 13092 20156
rect 13116 20154 13172 20156
rect 13196 20154 13252 20156
rect 12956 20102 13002 20154
rect 13002 20102 13012 20154
rect 13036 20102 13066 20154
rect 13066 20102 13078 20154
rect 13078 20102 13092 20154
rect 13116 20102 13130 20154
rect 13130 20102 13142 20154
rect 13142 20102 13172 20154
rect 13196 20102 13206 20154
rect 13206 20102 13252 20154
rect 12956 20100 13012 20102
rect 13036 20100 13092 20102
rect 13116 20100 13172 20102
rect 13196 20100 13252 20102
rect 12438 16768 12494 16824
rect 11058 7928 11114 7984
rect 11886 3188 11942 3224
rect 11886 3168 11888 3188
rect 11888 3168 11940 3188
rect 11940 3168 11942 3188
rect 12956 19066 13012 19068
rect 13036 19066 13092 19068
rect 13116 19066 13172 19068
rect 13196 19066 13252 19068
rect 12956 19014 13002 19066
rect 13002 19014 13012 19066
rect 13036 19014 13066 19066
rect 13066 19014 13078 19066
rect 13078 19014 13092 19066
rect 13116 19014 13130 19066
rect 13130 19014 13142 19066
rect 13142 19014 13172 19066
rect 13196 19014 13206 19066
rect 13206 19014 13252 19066
rect 12956 19012 13012 19014
rect 13036 19012 13092 19014
rect 13116 19012 13172 19014
rect 13196 19012 13252 19014
rect 12956 17978 13012 17980
rect 13036 17978 13092 17980
rect 13116 17978 13172 17980
rect 13196 17978 13252 17980
rect 12956 17926 13002 17978
rect 13002 17926 13012 17978
rect 13036 17926 13066 17978
rect 13066 17926 13078 17978
rect 13078 17926 13092 17978
rect 13116 17926 13130 17978
rect 13130 17926 13142 17978
rect 13142 17926 13172 17978
rect 13196 17926 13206 17978
rect 13206 17926 13252 17978
rect 12956 17924 13012 17926
rect 13036 17924 13092 17926
rect 13116 17924 13172 17926
rect 13196 17924 13252 17926
rect 12956 16890 13012 16892
rect 13036 16890 13092 16892
rect 13116 16890 13172 16892
rect 13196 16890 13252 16892
rect 12956 16838 13002 16890
rect 13002 16838 13012 16890
rect 13036 16838 13066 16890
rect 13066 16838 13078 16890
rect 13078 16838 13092 16890
rect 13116 16838 13130 16890
rect 13130 16838 13142 16890
rect 13142 16838 13172 16890
rect 13196 16838 13206 16890
rect 13206 16838 13252 16890
rect 12956 16836 13012 16838
rect 13036 16836 13092 16838
rect 13116 16836 13172 16838
rect 13196 16836 13252 16838
rect 12806 16788 12862 16824
rect 12806 16768 12808 16788
rect 12808 16768 12860 16788
rect 12860 16768 12862 16788
rect 12956 15802 13012 15804
rect 13036 15802 13092 15804
rect 13116 15802 13172 15804
rect 13196 15802 13252 15804
rect 12956 15750 13002 15802
rect 13002 15750 13012 15802
rect 13036 15750 13066 15802
rect 13066 15750 13078 15802
rect 13078 15750 13092 15802
rect 13116 15750 13130 15802
rect 13130 15750 13142 15802
rect 13142 15750 13172 15802
rect 13196 15750 13206 15802
rect 13206 15750 13252 15802
rect 12956 15748 13012 15750
rect 13036 15748 13092 15750
rect 13116 15748 13172 15750
rect 13196 15748 13252 15750
rect 12956 14714 13012 14716
rect 13036 14714 13092 14716
rect 13116 14714 13172 14716
rect 13196 14714 13252 14716
rect 12956 14662 13002 14714
rect 13002 14662 13012 14714
rect 13036 14662 13066 14714
rect 13066 14662 13078 14714
rect 13078 14662 13092 14714
rect 13116 14662 13130 14714
rect 13130 14662 13142 14714
rect 13142 14662 13172 14714
rect 13196 14662 13206 14714
rect 13206 14662 13252 14714
rect 12956 14660 13012 14662
rect 13036 14660 13092 14662
rect 13116 14660 13172 14662
rect 13196 14660 13252 14662
rect 13726 23704 13782 23760
rect 13634 21528 13690 21584
rect 13542 18828 13598 18864
rect 13542 18808 13544 18828
rect 13544 18808 13596 18828
rect 13596 18808 13598 18828
rect 13726 19252 13728 19272
rect 13728 19252 13780 19272
rect 13780 19252 13782 19272
rect 13726 19216 13782 19252
rect 12956 13626 13012 13628
rect 13036 13626 13092 13628
rect 13116 13626 13172 13628
rect 13196 13626 13252 13628
rect 12956 13574 13002 13626
rect 13002 13574 13012 13626
rect 13036 13574 13066 13626
rect 13066 13574 13078 13626
rect 13078 13574 13092 13626
rect 13116 13574 13130 13626
rect 13130 13574 13142 13626
rect 13142 13574 13172 13626
rect 13196 13574 13206 13626
rect 13206 13574 13252 13626
rect 12956 13572 13012 13574
rect 13036 13572 13092 13574
rect 13116 13572 13172 13574
rect 13196 13572 13252 13574
rect 13358 13096 13414 13152
rect 12956 12538 13012 12540
rect 13036 12538 13092 12540
rect 13116 12538 13172 12540
rect 13196 12538 13252 12540
rect 12956 12486 13002 12538
rect 13002 12486 13012 12538
rect 13036 12486 13066 12538
rect 13066 12486 13078 12538
rect 13078 12486 13092 12538
rect 13116 12486 13130 12538
rect 13130 12486 13142 12538
rect 13142 12486 13172 12538
rect 13196 12486 13206 12538
rect 13206 12486 13252 12538
rect 12956 12484 13012 12486
rect 13036 12484 13092 12486
rect 13116 12484 13172 12486
rect 13196 12484 13252 12486
rect 12956 11450 13012 11452
rect 13036 11450 13092 11452
rect 13116 11450 13172 11452
rect 13196 11450 13252 11452
rect 12956 11398 13002 11450
rect 13002 11398 13012 11450
rect 13036 11398 13066 11450
rect 13066 11398 13078 11450
rect 13078 11398 13092 11450
rect 13116 11398 13130 11450
rect 13130 11398 13142 11450
rect 13142 11398 13172 11450
rect 13196 11398 13206 11450
rect 13206 11398 13252 11450
rect 12956 11396 13012 11398
rect 13036 11396 13092 11398
rect 13116 11396 13172 11398
rect 13196 11396 13252 11398
rect 12956 10362 13012 10364
rect 13036 10362 13092 10364
rect 13116 10362 13172 10364
rect 13196 10362 13252 10364
rect 12956 10310 13002 10362
rect 13002 10310 13012 10362
rect 13036 10310 13066 10362
rect 13066 10310 13078 10362
rect 13078 10310 13092 10362
rect 13116 10310 13130 10362
rect 13130 10310 13142 10362
rect 13142 10310 13172 10362
rect 13196 10310 13206 10362
rect 13206 10310 13252 10362
rect 12956 10308 13012 10310
rect 13036 10308 13092 10310
rect 13116 10308 13172 10310
rect 13196 10308 13252 10310
rect 12956 9274 13012 9276
rect 13036 9274 13092 9276
rect 13116 9274 13172 9276
rect 13196 9274 13252 9276
rect 12956 9222 13002 9274
rect 13002 9222 13012 9274
rect 13036 9222 13066 9274
rect 13066 9222 13078 9274
rect 13078 9222 13092 9274
rect 13116 9222 13130 9274
rect 13130 9222 13142 9274
rect 13142 9222 13172 9274
rect 13196 9222 13206 9274
rect 13206 9222 13252 9274
rect 12956 9220 13012 9222
rect 13036 9220 13092 9222
rect 13116 9220 13172 9222
rect 13196 9220 13252 9222
rect 12956 8186 13012 8188
rect 13036 8186 13092 8188
rect 13116 8186 13172 8188
rect 13196 8186 13252 8188
rect 12956 8134 13002 8186
rect 13002 8134 13012 8186
rect 13036 8134 13066 8186
rect 13066 8134 13078 8186
rect 13078 8134 13092 8186
rect 13116 8134 13130 8186
rect 13130 8134 13142 8186
rect 13142 8134 13172 8186
rect 13196 8134 13206 8186
rect 13206 8134 13252 8186
rect 12956 8132 13012 8134
rect 13036 8132 13092 8134
rect 13116 8132 13172 8134
rect 13196 8132 13252 8134
rect 12956 7098 13012 7100
rect 13036 7098 13092 7100
rect 13116 7098 13172 7100
rect 13196 7098 13252 7100
rect 12956 7046 13002 7098
rect 13002 7046 13012 7098
rect 13036 7046 13066 7098
rect 13066 7046 13078 7098
rect 13078 7046 13092 7098
rect 13116 7046 13130 7098
rect 13130 7046 13142 7098
rect 13142 7046 13172 7098
rect 13196 7046 13206 7098
rect 13206 7046 13252 7098
rect 12956 7044 13012 7046
rect 13036 7044 13092 7046
rect 13116 7044 13172 7046
rect 13196 7044 13252 7046
rect 12956 6010 13012 6012
rect 13036 6010 13092 6012
rect 13116 6010 13172 6012
rect 13196 6010 13252 6012
rect 12956 5958 13002 6010
rect 13002 5958 13012 6010
rect 13036 5958 13066 6010
rect 13066 5958 13078 6010
rect 13078 5958 13092 6010
rect 13116 5958 13130 6010
rect 13130 5958 13142 6010
rect 13142 5958 13172 6010
rect 13196 5958 13206 6010
rect 13206 5958 13252 6010
rect 12956 5956 13012 5958
rect 13036 5956 13092 5958
rect 13116 5956 13172 5958
rect 13196 5956 13252 5958
rect 12956 4922 13012 4924
rect 13036 4922 13092 4924
rect 13116 4922 13172 4924
rect 13196 4922 13252 4924
rect 12956 4870 13002 4922
rect 13002 4870 13012 4922
rect 13036 4870 13066 4922
rect 13066 4870 13078 4922
rect 13078 4870 13092 4922
rect 13116 4870 13130 4922
rect 13130 4870 13142 4922
rect 13142 4870 13172 4922
rect 13196 4870 13206 4922
rect 13206 4870 13252 4922
rect 12956 4868 13012 4870
rect 13036 4868 13092 4870
rect 13116 4868 13172 4870
rect 13196 4868 13252 4870
rect 12956 3834 13012 3836
rect 13036 3834 13092 3836
rect 13116 3834 13172 3836
rect 13196 3834 13252 3836
rect 12956 3782 13002 3834
rect 13002 3782 13012 3834
rect 13036 3782 13066 3834
rect 13066 3782 13078 3834
rect 13078 3782 13092 3834
rect 13116 3782 13130 3834
rect 13130 3782 13142 3834
rect 13142 3782 13172 3834
rect 13196 3782 13206 3834
rect 13206 3782 13252 3834
rect 12956 3780 13012 3782
rect 13036 3780 13092 3782
rect 13116 3780 13172 3782
rect 13196 3780 13252 3782
rect 12956 2746 13012 2748
rect 13036 2746 13092 2748
rect 13116 2746 13172 2748
rect 13196 2746 13252 2748
rect 12956 2694 13002 2746
rect 13002 2694 13012 2746
rect 13036 2694 13066 2746
rect 13066 2694 13078 2746
rect 13078 2694 13092 2746
rect 13116 2694 13130 2746
rect 13130 2694 13142 2746
rect 13142 2694 13172 2746
rect 13196 2694 13206 2746
rect 13206 2694 13252 2746
rect 12956 2692 13012 2694
rect 13036 2692 13092 2694
rect 13116 2692 13172 2694
rect 13196 2692 13252 2694
rect 15750 52536 15806 52592
rect 15106 38392 15162 38448
rect 16854 52536 16910 52592
rect 14830 32816 14886 32872
rect 15934 38700 15936 38720
rect 15936 38700 15988 38720
rect 15988 38700 15990 38720
rect 15934 38664 15990 38700
rect 15382 30540 15384 30560
rect 15384 30540 15436 30560
rect 15436 30540 15438 30560
rect 15382 30504 15438 30540
rect 15290 29280 15346 29336
rect 15750 31728 15806 31784
rect 16578 40604 16580 40624
rect 16580 40604 16632 40624
rect 16632 40604 16634 40624
rect 16578 40568 16634 40604
rect 16670 36780 16726 36816
rect 16670 36760 16672 36780
rect 16672 36760 16724 36780
rect 16724 36760 16726 36780
rect 16946 40432 17002 40488
rect 16854 37712 16910 37768
rect 17956 54426 18012 54428
rect 18036 54426 18092 54428
rect 18116 54426 18172 54428
rect 18196 54426 18252 54428
rect 17956 54374 18002 54426
rect 18002 54374 18012 54426
rect 18036 54374 18066 54426
rect 18066 54374 18078 54426
rect 18078 54374 18092 54426
rect 18116 54374 18130 54426
rect 18130 54374 18142 54426
rect 18142 54374 18172 54426
rect 18196 54374 18206 54426
rect 18206 54374 18252 54426
rect 17956 54372 18012 54374
rect 18036 54372 18092 54374
rect 18116 54372 18172 54374
rect 18196 54372 18252 54374
rect 24490 56208 24546 56264
rect 17956 53338 18012 53340
rect 18036 53338 18092 53340
rect 18116 53338 18172 53340
rect 18196 53338 18252 53340
rect 17956 53286 18002 53338
rect 18002 53286 18012 53338
rect 18036 53286 18066 53338
rect 18066 53286 18078 53338
rect 18078 53286 18092 53338
rect 18116 53286 18130 53338
rect 18130 53286 18142 53338
rect 18142 53286 18172 53338
rect 18196 53286 18206 53338
rect 18206 53286 18252 53338
rect 17956 53284 18012 53286
rect 18036 53284 18092 53286
rect 18116 53284 18172 53286
rect 18196 53284 18252 53286
rect 17956 52250 18012 52252
rect 18036 52250 18092 52252
rect 18116 52250 18172 52252
rect 18196 52250 18252 52252
rect 17956 52198 18002 52250
rect 18002 52198 18012 52250
rect 18036 52198 18066 52250
rect 18066 52198 18078 52250
rect 18078 52198 18092 52250
rect 18116 52198 18130 52250
rect 18130 52198 18142 52250
rect 18142 52198 18172 52250
rect 18196 52198 18206 52250
rect 18206 52198 18252 52250
rect 17956 52196 18012 52198
rect 18036 52196 18092 52198
rect 18116 52196 18172 52198
rect 18196 52196 18252 52198
rect 17956 51162 18012 51164
rect 18036 51162 18092 51164
rect 18116 51162 18172 51164
rect 18196 51162 18252 51164
rect 17956 51110 18002 51162
rect 18002 51110 18012 51162
rect 18036 51110 18066 51162
rect 18066 51110 18078 51162
rect 18078 51110 18092 51162
rect 18116 51110 18130 51162
rect 18130 51110 18142 51162
rect 18142 51110 18172 51162
rect 18196 51110 18206 51162
rect 18206 51110 18252 51162
rect 17956 51108 18012 51110
rect 18036 51108 18092 51110
rect 18116 51108 18172 51110
rect 18196 51108 18252 51110
rect 17956 50074 18012 50076
rect 18036 50074 18092 50076
rect 18116 50074 18172 50076
rect 18196 50074 18252 50076
rect 17956 50022 18002 50074
rect 18002 50022 18012 50074
rect 18036 50022 18066 50074
rect 18066 50022 18078 50074
rect 18078 50022 18092 50074
rect 18116 50022 18130 50074
rect 18130 50022 18142 50074
rect 18142 50022 18172 50074
rect 18196 50022 18206 50074
rect 18206 50022 18252 50074
rect 17956 50020 18012 50022
rect 18036 50020 18092 50022
rect 18116 50020 18172 50022
rect 18196 50020 18252 50022
rect 17956 48986 18012 48988
rect 18036 48986 18092 48988
rect 18116 48986 18172 48988
rect 18196 48986 18252 48988
rect 17956 48934 18002 48986
rect 18002 48934 18012 48986
rect 18036 48934 18066 48986
rect 18066 48934 18078 48986
rect 18078 48934 18092 48986
rect 18116 48934 18130 48986
rect 18130 48934 18142 48986
rect 18142 48934 18172 48986
rect 18196 48934 18206 48986
rect 18206 48934 18252 48986
rect 17956 48932 18012 48934
rect 18036 48932 18092 48934
rect 18116 48932 18172 48934
rect 18196 48932 18252 48934
rect 17956 47898 18012 47900
rect 18036 47898 18092 47900
rect 18116 47898 18172 47900
rect 18196 47898 18252 47900
rect 17956 47846 18002 47898
rect 18002 47846 18012 47898
rect 18036 47846 18066 47898
rect 18066 47846 18078 47898
rect 18078 47846 18092 47898
rect 18116 47846 18130 47898
rect 18130 47846 18142 47898
rect 18142 47846 18172 47898
rect 18196 47846 18206 47898
rect 18206 47846 18252 47898
rect 17956 47844 18012 47846
rect 18036 47844 18092 47846
rect 18116 47844 18172 47846
rect 18196 47844 18252 47846
rect 17956 46810 18012 46812
rect 18036 46810 18092 46812
rect 18116 46810 18172 46812
rect 18196 46810 18252 46812
rect 17956 46758 18002 46810
rect 18002 46758 18012 46810
rect 18036 46758 18066 46810
rect 18066 46758 18078 46810
rect 18078 46758 18092 46810
rect 18116 46758 18130 46810
rect 18130 46758 18142 46810
rect 18142 46758 18172 46810
rect 18196 46758 18206 46810
rect 18206 46758 18252 46810
rect 17956 46756 18012 46758
rect 18036 46756 18092 46758
rect 18116 46756 18172 46758
rect 18196 46756 18252 46758
rect 17956 45722 18012 45724
rect 18036 45722 18092 45724
rect 18116 45722 18172 45724
rect 18196 45722 18252 45724
rect 17956 45670 18002 45722
rect 18002 45670 18012 45722
rect 18036 45670 18066 45722
rect 18066 45670 18078 45722
rect 18078 45670 18092 45722
rect 18116 45670 18130 45722
rect 18130 45670 18142 45722
rect 18142 45670 18172 45722
rect 18196 45670 18206 45722
rect 18206 45670 18252 45722
rect 17956 45668 18012 45670
rect 18036 45668 18092 45670
rect 18116 45668 18172 45670
rect 18196 45668 18252 45670
rect 17956 44634 18012 44636
rect 18036 44634 18092 44636
rect 18116 44634 18172 44636
rect 18196 44634 18252 44636
rect 17956 44582 18002 44634
rect 18002 44582 18012 44634
rect 18036 44582 18066 44634
rect 18066 44582 18078 44634
rect 18078 44582 18092 44634
rect 18116 44582 18130 44634
rect 18130 44582 18142 44634
rect 18142 44582 18172 44634
rect 18196 44582 18206 44634
rect 18206 44582 18252 44634
rect 17956 44580 18012 44582
rect 18036 44580 18092 44582
rect 18116 44580 18172 44582
rect 18196 44580 18252 44582
rect 17130 37576 17186 37632
rect 17956 43546 18012 43548
rect 18036 43546 18092 43548
rect 18116 43546 18172 43548
rect 18196 43546 18252 43548
rect 17956 43494 18002 43546
rect 18002 43494 18012 43546
rect 18036 43494 18066 43546
rect 18066 43494 18078 43546
rect 18078 43494 18092 43546
rect 18116 43494 18130 43546
rect 18130 43494 18142 43546
rect 18142 43494 18172 43546
rect 18196 43494 18206 43546
rect 18206 43494 18252 43546
rect 17956 43492 18012 43494
rect 18036 43492 18092 43494
rect 18116 43492 18172 43494
rect 18196 43492 18252 43494
rect 17956 42458 18012 42460
rect 18036 42458 18092 42460
rect 18116 42458 18172 42460
rect 18196 42458 18252 42460
rect 17956 42406 18002 42458
rect 18002 42406 18012 42458
rect 18036 42406 18066 42458
rect 18066 42406 18078 42458
rect 18078 42406 18092 42458
rect 18116 42406 18130 42458
rect 18130 42406 18142 42458
rect 18142 42406 18172 42458
rect 18196 42406 18206 42458
rect 18206 42406 18252 42458
rect 17956 42404 18012 42406
rect 18036 42404 18092 42406
rect 18116 42404 18172 42406
rect 18196 42404 18252 42406
rect 18510 46996 18512 47016
rect 18512 46996 18564 47016
rect 18564 46996 18566 47016
rect 18510 46960 18566 46996
rect 17956 41370 18012 41372
rect 18036 41370 18092 41372
rect 18116 41370 18172 41372
rect 18196 41370 18252 41372
rect 17956 41318 18002 41370
rect 18002 41318 18012 41370
rect 18036 41318 18066 41370
rect 18066 41318 18078 41370
rect 18078 41318 18092 41370
rect 18116 41318 18130 41370
rect 18130 41318 18142 41370
rect 18142 41318 18172 41370
rect 18196 41318 18206 41370
rect 18206 41318 18252 41370
rect 17956 41316 18012 41318
rect 18036 41316 18092 41318
rect 18116 41316 18172 41318
rect 18196 41316 18252 41318
rect 17956 40282 18012 40284
rect 18036 40282 18092 40284
rect 18116 40282 18172 40284
rect 18196 40282 18252 40284
rect 17956 40230 18002 40282
rect 18002 40230 18012 40282
rect 18036 40230 18066 40282
rect 18066 40230 18078 40282
rect 18078 40230 18092 40282
rect 18116 40230 18130 40282
rect 18130 40230 18142 40282
rect 18142 40230 18172 40282
rect 18196 40230 18206 40282
rect 18206 40230 18252 40282
rect 17956 40228 18012 40230
rect 18036 40228 18092 40230
rect 18116 40228 18172 40230
rect 18196 40228 18252 40230
rect 18234 40024 18290 40080
rect 17956 39194 18012 39196
rect 18036 39194 18092 39196
rect 18116 39194 18172 39196
rect 18196 39194 18252 39196
rect 17956 39142 18002 39194
rect 18002 39142 18012 39194
rect 18036 39142 18066 39194
rect 18066 39142 18078 39194
rect 18078 39142 18092 39194
rect 18116 39142 18130 39194
rect 18130 39142 18142 39194
rect 18142 39142 18172 39194
rect 18196 39142 18206 39194
rect 18206 39142 18252 39194
rect 17956 39140 18012 39142
rect 18036 39140 18092 39142
rect 18116 39140 18172 39142
rect 18196 39140 18252 39142
rect 17956 38106 18012 38108
rect 18036 38106 18092 38108
rect 18116 38106 18172 38108
rect 18196 38106 18252 38108
rect 17956 38054 18002 38106
rect 18002 38054 18012 38106
rect 18036 38054 18066 38106
rect 18066 38054 18078 38106
rect 18078 38054 18092 38106
rect 18116 38054 18130 38106
rect 18130 38054 18142 38106
rect 18142 38054 18172 38106
rect 18196 38054 18206 38106
rect 18206 38054 18252 38106
rect 17956 38052 18012 38054
rect 18036 38052 18092 38054
rect 18116 38052 18172 38054
rect 18196 38052 18252 38054
rect 14278 15136 14334 15192
rect 14738 18572 14740 18592
rect 14740 18572 14792 18592
rect 14792 18572 14794 18592
rect 14738 18536 14794 18572
rect 15382 28192 15438 28248
rect 15750 23160 15806 23216
rect 15014 15700 15070 15736
rect 15014 15680 15016 15700
rect 15016 15680 15068 15700
rect 15068 15680 15070 15700
rect 14922 14068 14978 14104
rect 14922 14048 14924 14068
rect 14924 14048 14976 14068
rect 14976 14048 14978 14068
rect 16118 26732 16120 26752
rect 16120 26732 16172 26752
rect 16172 26732 16174 26752
rect 16118 26696 16174 26732
rect 16118 22208 16174 22264
rect 15842 21140 15898 21176
rect 15842 21120 15844 21140
rect 15844 21120 15896 21140
rect 15896 21120 15898 21140
rect 15934 20440 15990 20496
rect 16762 29452 16764 29472
rect 16764 29452 16816 29472
rect 16816 29452 16818 29472
rect 16762 29416 16818 29452
rect 17682 33108 17738 33144
rect 17682 33088 17684 33108
rect 17684 33088 17736 33108
rect 17736 33088 17738 33108
rect 17956 37018 18012 37020
rect 18036 37018 18092 37020
rect 18116 37018 18172 37020
rect 18196 37018 18252 37020
rect 17956 36966 18002 37018
rect 18002 36966 18012 37018
rect 18036 36966 18066 37018
rect 18066 36966 18078 37018
rect 18078 36966 18092 37018
rect 18116 36966 18130 37018
rect 18130 36966 18142 37018
rect 18142 36966 18172 37018
rect 18196 36966 18206 37018
rect 18206 36966 18252 37018
rect 17956 36964 18012 36966
rect 18036 36964 18092 36966
rect 18116 36964 18172 36966
rect 18196 36964 18252 36966
rect 18326 36624 18382 36680
rect 17956 35930 18012 35932
rect 18036 35930 18092 35932
rect 18116 35930 18172 35932
rect 18196 35930 18252 35932
rect 17956 35878 18002 35930
rect 18002 35878 18012 35930
rect 18036 35878 18066 35930
rect 18066 35878 18078 35930
rect 18078 35878 18092 35930
rect 18116 35878 18130 35930
rect 18130 35878 18142 35930
rect 18142 35878 18172 35930
rect 18196 35878 18206 35930
rect 18206 35878 18252 35930
rect 17956 35876 18012 35878
rect 18036 35876 18092 35878
rect 18116 35876 18172 35878
rect 18196 35876 18252 35878
rect 19614 46552 19670 46608
rect 19338 44684 19340 44704
rect 19340 44684 19392 44704
rect 19392 44684 19394 44704
rect 19338 44648 19394 44684
rect 17956 34842 18012 34844
rect 18036 34842 18092 34844
rect 18116 34842 18172 34844
rect 18196 34842 18252 34844
rect 17956 34790 18002 34842
rect 18002 34790 18012 34842
rect 18036 34790 18066 34842
rect 18066 34790 18078 34842
rect 18078 34790 18092 34842
rect 18116 34790 18130 34842
rect 18130 34790 18142 34842
rect 18142 34790 18172 34842
rect 18196 34790 18206 34842
rect 18206 34790 18252 34842
rect 17956 34788 18012 34790
rect 18036 34788 18092 34790
rect 18116 34788 18172 34790
rect 18196 34788 18252 34790
rect 17314 29300 17370 29336
rect 17314 29280 17316 29300
rect 17316 29280 17368 29300
rect 17368 29280 17370 29300
rect 17956 33754 18012 33756
rect 18036 33754 18092 33756
rect 18116 33754 18172 33756
rect 18196 33754 18252 33756
rect 17956 33702 18002 33754
rect 18002 33702 18012 33754
rect 18036 33702 18066 33754
rect 18066 33702 18078 33754
rect 18078 33702 18092 33754
rect 18116 33702 18130 33754
rect 18130 33702 18142 33754
rect 18142 33702 18172 33754
rect 18196 33702 18206 33754
rect 18206 33702 18252 33754
rect 17956 33700 18012 33702
rect 18036 33700 18092 33702
rect 18116 33700 18172 33702
rect 18196 33700 18252 33702
rect 17956 32666 18012 32668
rect 18036 32666 18092 32668
rect 18116 32666 18172 32668
rect 18196 32666 18252 32668
rect 17956 32614 18002 32666
rect 18002 32614 18012 32666
rect 18036 32614 18066 32666
rect 18066 32614 18078 32666
rect 18078 32614 18092 32666
rect 18116 32614 18130 32666
rect 18130 32614 18142 32666
rect 18142 32614 18172 32666
rect 18196 32614 18206 32666
rect 18206 32614 18252 32666
rect 17956 32612 18012 32614
rect 18036 32612 18092 32614
rect 18116 32612 18172 32614
rect 18196 32612 18252 32614
rect 17314 28364 17316 28384
rect 17316 28364 17368 28384
rect 17368 28364 17370 28384
rect 17314 28328 17370 28364
rect 17314 26868 17316 26888
rect 17316 26868 17368 26888
rect 17368 26868 17370 26888
rect 17314 26832 17370 26868
rect 16670 21120 16726 21176
rect 16210 16244 16266 16280
rect 16210 16224 16212 16244
rect 16212 16224 16264 16244
rect 16264 16224 16266 16244
rect 16026 11228 16028 11248
rect 16028 11228 16080 11248
rect 16080 11228 16082 11248
rect 16026 11192 16082 11228
rect 17682 28364 17684 28384
rect 17684 28364 17736 28384
rect 17736 28364 17738 28384
rect 17682 28328 17738 28364
rect 17682 28212 17738 28248
rect 17682 28192 17684 28212
rect 17684 28192 17736 28212
rect 17736 28192 17738 28212
rect 17956 31578 18012 31580
rect 18036 31578 18092 31580
rect 18116 31578 18172 31580
rect 18196 31578 18252 31580
rect 17956 31526 18002 31578
rect 18002 31526 18012 31578
rect 18036 31526 18066 31578
rect 18066 31526 18078 31578
rect 18078 31526 18092 31578
rect 18116 31526 18130 31578
rect 18130 31526 18142 31578
rect 18142 31526 18172 31578
rect 18196 31526 18206 31578
rect 18206 31526 18252 31578
rect 17956 31524 18012 31526
rect 18036 31524 18092 31526
rect 18116 31524 18172 31526
rect 18196 31524 18252 31526
rect 17956 30490 18012 30492
rect 18036 30490 18092 30492
rect 18116 30490 18172 30492
rect 18196 30490 18252 30492
rect 17956 30438 18002 30490
rect 18002 30438 18012 30490
rect 18036 30438 18066 30490
rect 18066 30438 18078 30490
rect 18078 30438 18092 30490
rect 18116 30438 18130 30490
rect 18130 30438 18142 30490
rect 18142 30438 18172 30490
rect 18196 30438 18206 30490
rect 18206 30438 18252 30490
rect 17956 30436 18012 30438
rect 18036 30436 18092 30438
rect 18116 30436 18172 30438
rect 18196 30436 18252 30438
rect 17956 29402 18012 29404
rect 18036 29402 18092 29404
rect 18116 29402 18172 29404
rect 18196 29402 18252 29404
rect 17956 29350 18002 29402
rect 18002 29350 18012 29402
rect 18036 29350 18066 29402
rect 18066 29350 18078 29402
rect 18078 29350 18092 29402
rect 18116 29350 18130 29402
rect 18130 29350 18142 29402
rect 18142 29350 18172 29402
rect 18196 29350 18206 29402
rect 18206 29350 18252 29402
rect 17956 29348 18012 29350
rect 18036 29348 18092 29350
rect 18116 29348 18172 29350
rect 18196 29348 18252 29350
rect 17956 28314 18012 28316
rect 18036 28314 18092 28316
rect 18116 28314 18172 28316
rect 18196 28314 18252 28316
rect 17956 28262 18002 28314
rect 18002 28262 18012 28314
rect 18036 28262 18066 28314
rect 18066 28262 18078 28314
rect 18078 28262 18092 28314
rect 18116 28262 18130 28314
rect 18130 28262 18142 28314
rect 18142 28262 18172 28314
rect 18196 28262 18206 28314
rect 18206 28262 18252 28314
rect 17956 28260 18012 28262
rect 18036 28260 18092 28262
rect 18116 28260 18172 28262
rect 18196 28260 18252 28262
rect 17956 27226 18012 27228
rect 18036 27226 18092 27228
rect 18116 27226 18172 27228
rect 18196 27226 18252 27228
rect 17956 27174 18002 27226
rect 18002 27174 18012 27226
rect 18036 27174 18066 27226
rect 18066 27174 18078 27226
rect 18078 27174 18092 27226
rect 18116 27174 18130 27226
rect 18130 27174 18142 27226
rect 18142 27174 18172 27226
rect 18196 27174 18206 27226
rect 18206 27174 18252 27226
rect 17956 27172 18012 27174
rect 18036 27172 18092 27174
rect 18116 27172 18172 27174
rect 18196 27172 18252 27174
rect 17956 26138 18012 26140
rect 18036 26138 18092 26140
rect 18116 26138 18172 26140
rect 18196 26138 18252 26140
rect 17956 26086 18002 26138
rect 18002 26086 18012 26138
rect 18036 26086 18066 26138
rect 18066 26086 18078 26138
rect 18078 26086 18092 26138
rect 18116 26086 18130 26138
rect 18130 26086 18142 26138
rect 18142 26086 18172 26138
rect 18196 26086 18206 26138
rect 18206 26086 18252 26138
rect 17956 26084 18012 26086
rect 18036 26084 18092 26086
rect 18116 26084 18172 26086
rect 18196 26084 18252 26086
rect 18602 31884 18658 31920
rect 18602 31864 18604 31884
rect 18604 31864 18656 31884
rect 18656 31864 18658 31884
rect 20626 46688 20682 46744
rect 18970 37440 19026 37496
rect 19246 37576 19302 37632
rect 19062 37304 19118 37360
rect 18694 29996 18696 30016
rect 18696 29996 18748 30016
rect 18748 29996 18750 30016
rect 18694 29960 18750 29996
rect 17956 25050 18012 25052
rect 18036 25050 18092 25052
rect 18116 25050 18172 25052
rect 18196 25050 18252 25052
rect 17956 24998 18002 25050
rect 18002 24998 18012 25050
rect 18036 24998 18066 25050
rect 18066 24998 18078 25050
rect 18078 24998 18092 25050
rect 18116 24998 18130 25050
rect 18130 24998 18142 25050
rect 18142 24998 18172 25050
rect 18196 24998 18206 25050
rect 18206 24998 18252 25050
rect 17956 24996 18012 24998
rect 18036 24996 18092 24998
rect 18116 24996 18172 24998
rect 18196 24996 18252 24998
rect 17956 23962 18012 23964
rect 18036 23962 18092 23964
rect 18116 23962 18172 23964
rect 18196 23962 18252 23964
rect 17956 23910 18002 23962
rect 18002 23910 18012 23962
rect 18036 23910 18066 23962
rect 18066 23910 18078 23962
rect 18078 23910 18092 23962
rect 18116 23910 18130 23962
rect 18130 23910 18142 23962
rect 18142 23910 18172 23962
rect 18196 23910 18206 23962
rect 18206 23910 18252 23962
rect 17956 23908 18012 23910
rect 18036 23908 18092 23910
rect 18116 23908 18172 23910
rect 18196 23908 18252 23910
rect 17956 22874 18012 22876
rect 18036 22874 18092 22876
rect 18116 22874 18172 22876
rect 18196 22874 18252 22876
rect 17956 22822 18002 22874
rect 18002 22822 18012 22874
rect 18036 22822 18066 22874
rect 18066 22822 18078 22874
rect 18078 22822 18092 22874
rect 18116 22822 18130 22874
rect 18130 22822 18142 22874
rect 18142 22822 18172 22874
rect 18196 22822 18206 22874
rect 18206 22822 18252 22874
rect 17956 22820 18012 22822
rect 18036 22820 18092 22822
rect 18116 22820 18172 22822
rect 18196 22820 18252 22822
rect 17956 21786 18012 21788
rect 18036 21786 18092 21788
rect 18116 21786 18172 21788
rect 18196 21786 18252 21788
rect 17956 21734 18002 21786
rect 18002 21734 18012 21786
rect 18036 21734 18066 21786
rect 18066 21734 18078 21786
rect 18078 21734 18092 21786
rect 18116 21734 18130 21786
rect 18130 21734 18142 21786
rect 18142 21734 18172 21786
rect 18196 21734 18206 21786
rect 18206 21734 18252 21786
rect 17956 21732 18012 21734
rect 18036 21732 18092 21734
rect 18116 21732 18172 21734
rect 18196 21732 18252 21734
rect 17956 20698 18012 20700
rect 18036 20698 18092 20700
rect 18116 20698 18172 20700
rect 18196 20698 18252 20700
rect 17956 20646 18002 20698
rect 18002 20646 18012 20698
rect 18036 20646 18066 20698
rect 18066 20646 18078 20698
rect 18078 20646 18092 20698
rect 18116 20646 18130 20698
rect 18130 20646 18142 20698
rect 18142 20646 18172 20698
rect 18196 20646 18206 20698
rect 18206 20646 18252 20698
rect 17956 20644 18012 20646
rect 18036 20644 18092 20646
rect 18116 20644 18172 20646
rect 18196 20644 18252 20646
rect 17590 18672 17646 18728
rect 17956 19610 18012 19612
rect 18036 19610 18092 19612
rect 18116 19610 18172 19612
rect 18196 19610 18252 19612
rect 17956 19558 18002 19610
rect 18002 19558 18012 19610
rect 18036 19558 18066 19610
rect 18066 19558 18078 19610
rect 18078 19558 18092 19610
rect 18116 19558 18130 19610
rect 18130 19558 18142 19610
rect 18142 19558 18172 19610
rect 18196 19558 18206 19610
rect 18206 19558 18252 19610
rect 17956 19556 18012 19558
rect 18036 19556 18092 19558
rect 18116 19556 18172 19558
rect 18196 19556 18252 19558
rect 18326 18672 18382 18728
rect 17956 18522 18012 18524
rect 18036 18522 18092 18524
rect 18116 18522 18172 18524
rect 18196 18522 18252 18524
rect 17956 18470 18002 18522
rect 18002 18470 18012 18522
rect 18036 18470 18066 18522
rect 18066 18470 18078 18522
rect 18078 18470 18092 18522
rect 18116 18470 18130 18522
rect 18130 18470 18142 18522
rect 18142 18470 18172 18522
rect 18196 18470 18206 18522
rect 18206 18470 18252 18522
rect 17956 18468 18012 18470
rect 18036 18468 18092 18470
rect 18116 18468 18172 18470
rect 18196 18468 18252 18470
rect 17956 17434 18012 17436
rect 18036 17434 18092 17436
rect 18116 17434 18172 17436
rect 18196 17434 18252 17436
rect 17956 17382 18002 17434
rect 18002 17382 18012 17434
rect 18036 17382 18066 17434
rect 18066 17382 18078 17434
rect 18078 17382 18092 17434
rect 18116 17382 18130 17434
rect 18130 17382 18142 17434
rect 18142 17382 18172 17434
rect 18196 17382 18206 17434
rect 18206 17382 18252 17434
rect 17956 17380 18012 17382
rect 18036 17380 18092 17382
rect 18116 17380 18172 17382
rect 18196 17380 18252 17382
rect 17956 16346 18012 16348
rect 18036 16346 18092 16348
rect 18116 16346 18172 16348
rect 18196 16346 18252 16348
rect 17956 16294 18002 16346
rect 18002 16294 18012 16346
rect 18036 16294 18066 16346
rect 18066 16294 18078 16346
rect 18078 16294 18092 16346
rect 18116 16294 18130 16346
rect 18130 16294 18142 16346
rect 18142 16294 18172 16346
rect 18196 16294 18206 16346
rect 18206 16294 18252 16346
rect 17956 16292 18012 16294
rect 18036 16292 18092 16294
rect 18116 16292 18172 16294
rect 18196 16292 18252 16294
rect 17956 15258 18012 15260
rect 18036 15258 18092 15260
rect 18116 15258 18172 15260
rect 18196 15258 18252 15260
rect 17956 15206 18002 15258
rect 18002 15206 18012 15258
rect 18036 15206 18066 15258
rect 18066 15206 18078 15258
rect 18078 15206 18092 15258
rect 18116 15206 18130 15258
rect 18130 15206 18142 15258
rect 18142 15206 18172 15258
rect 18196 15206 18206 15258
rect 18206 15206 18252 15258
rect 17956 15204 18012 15206
rect 18036 15204 18092 15206
rect 18116 15204 18172 15206
rect 18196 15204 18252 15206
rect 17956 14170 18012 14172
rect 18036 14170 18092 14172
rect 18116 14170 18172 14172
rect 18196 14170 18252 14172
rect 17956 14118 18002 14170
rect 18002 14118 18012 14170
rect 18036 14118 18066 14170
rect 18066 14118 18078 14170
rect 18078 14118 18092 14170
rect 18116 14118 18130 14170
rect 18130 14118 18142 14170
rect 18142 14118 18172 14170
rect 18196 14118 18206 14170
rect 18206 14118 18252 14170
rect 17956 14116 18012 14118
rect 18036 14116 18092 14118
rect 18116 14116 18172 14118
rect 18196 14116 18252 14118
rect 17956 13082 18012 13084
rect 18036 13082 18092 13084
rect 18116 13082 18172 13084
rect 18196 13082 18252 13084
rect 17956 13030 18002 13082
rect 18002 13030 18012 13082
rect 18036 13030 18066 13082
rect 18066 13030 18078 13082
rect 18078 13030 18092 13082
rect 18116 13030 18130 13082
rect 18130 13030 18142 13082
rect 18142 13030 18172 13082
rect 18196 13030 18206 13082
rect 18206 13030 18252 13082
rect 17956 13028 18012 13030
rect 18036 13028 18092 13030
rect 18116 13028 18172 13030
rect 18196 13028 18252 13030
rect 18418 14456 18474 14512
rect 17956 11994 18012 11996
rect 18036 11994 18092 11996
rect 18116 11994 18172 11996
rect 18196 11994 18252 11996
rect 17956 11942 18002 11994
rect 18002 11942 18012 11994
rect 18036 11942 18066 11994
rect 18066 11942 18078 11994
rect 18078 11942 18092 11994
rect 18116 11942 18130 11994
rect 18130 11942 18142 11994
rect 18142 11942 18172 11994
rect 18196 11942 18206 11994
rect 18206 11942 18252 11994
rect 17956 11940 18012 11942
rect 18036 11940 18092 11942
rect 18116 11940 18172 11942
rect 18196 11940 18252 11942
rect 17956 10906 18012 10908
rect 18036 10906 18092 10908
rect 18116 10906 18172 10908
rect 18196 10906 18252 10908
rect 17956 10854 18002 10906
rect 18002 10854 18012 10906
rect 18036 10854 18066 10906
rect 18066 10854 18078 10906
rect 18078 10854 18092 10906
rect 18116 10854 18130 10906
rect 18130 10854 18142 10906
rect 18142 10854 18172 10906
rect 18196 10854 18206 10906
rect 18206 10854 18252 10906
rect 17956 10852 18012 10854
rect 18036 10852 18092 10854
rect 18116 10852 18172 10854
rect 18196 10852 18252 10854
rect 19338 37304 19394 37360
rect 19154 36624 19210 36680
rect 19614 36080 19670 36136
rect 20534 42064 20590 42120
rect 20166 40432 20222 40488
rect 19798 33496 19854 33552
rect 18878 18672 18934 18728
rect 17956 9818 18012 9820
rect 18036 9818 18092 9820
rect 18116 9818 18172 9820
rect 18196 9818 18252 9820
rect 17956 9766 18002 9818
rect 18002 9766 18012 9818
rect 18036 9766 18066 9818
rect 18066 9766 18078 9818
rect 18078 9766 18092 9818
rect 18116 9766 18130 9818
rect 18130 9766 18142 9818
rect 18142 9766 18172 9818
rect 18196 9766 18206 9818
rect 18206 9766 18252 9818
rect 17956 9764 18012 9766
rect 18036 9764 18092 9766
rect 18116 9764 18172 9766
rect 18196 9764 18252 9766
rect 17956 8730 18012 8732
rect 18036 8730 18092 8732
rect 18116 8730 18172 8732
rect 18196 8730 18252 8732
rect 17956 8678 18002 8730
rect 18002 8678 18012 8730
rect 18036 8678 18066 8730
rect 18066 8678 18078 8730
rect 18078 8678 18092 8730
rect 18116 8678 18130 8730
rect 18130 8678 18142 8730
rect 18142 8678 18172 8730
rect 18196 8678 18206 8730
rect 18206 8678 18252 8730
rect 17956 8676 18012 8678
rect 18036 8676 18092 8678
rect 18116 8676 18172 8678
rect 18196 8676 18252 8678
rect 17956 7642 18012 7644
rect 18036 7642 18092 7644
rect 18116 7642 18172 7644
rect 18196 7642 18252 7644
rect 17956 7590 18002 7642
rect 18002 7590 18012 7642
rect 18036 7590 18066 7642
rect 18066 7590 18078 7642
rect 18078 7590 18092 7642
rect 18116 7590 18130 7642
rect 18130 7590 18142 7642
rect 18142 7590 18172 7642
rect 18196 7590 18206 7642
rect 18206 7590 18252 7642
rect 17956 7588 18012 7590
rect 18036 7588 18092 7590
rect 18116 7588 18172 7590
rect 18196 7588 18252 7590
rect 17956 6554 18012 6556
rect 18036 6554 18092 6556
rect 18116 6554 18172 6556
rect 18196 6554 18252 6556
rect 17956 6502 18002 6554
rect 18002 6502 18012 6554
rect 18036 6502 18066 6554
rect 18066 6502 18078 6554
rect 18078 6502 18092 6554
rect 18116 6502 18130 6554
rect 18130 6502 18142 6554
rect 18142 6502 18172 6554
rect 18196 6502 18206 6554
rect 18206 6502 18252 6554
rect 17956 6500 18012 6502
rect 18036 6500 18092 6502
rect 18116 6500 18172 6502
rect 18196 6500 18252 6502
rect 17956 5466 18012 5468
rect 18036 5466 18092 5468
rect 18116 5466 18172 5468
rect 18196 5466 18252 5468
rect 17956 5414 18002 5466
rect 18002 5414 18012 5466
rect 18036 5414 18066 5466
rect 18066 5414 18078 5466
rect 18078 5414 18092 5466
rect 18116 5414 18130 5466
rect 18130 5414 18142 5466
rect 18142 5414 18172 5466
rect 18196 5414 18206 5466
rect 18206 5414 18252 5466
rect 17956 5412 18012 5414
rect 18036 5412 18092 5414
rect 18116 5412 18172 5414
rect 18196 5412 18252 5414
rect 20074 36352 20130 36408
rect 19890 30540 19892 30560
rect 19892 30540 19944 30560
rect 19944 30540 19946 30560
rect 19890 30504 19946 30540
rect 19798 29960 19854 30016
rect 19798 29008 19854 29064
rect 21086 43152 21142 43208
rect 22006 45872 22062 45928
rect 22374 53932 22376 53952
rect 22376 53932 22428 53952
rect 22428 53932 22430 53952
rect 22374 53896 22430 53932
rect 21914 43152 21970 43208
rect 22006 42764 22062 42800
rect 22006 42744 22008 42764
rect 22008 42744 22060 42764
rect 22060 42744 22062 42764
rect 21086 36524 21088 36544
rect 21088 36524 21140 36544
rect 21140 36524 21142 36544
rect 21086 36488 21142 36524
rect 21454 36352 21510 36408
rect 22956 53882 23012 53884
rect 23036 53882 23092 53884
rect 23116 53882 23172 53884
rect 23196 53882 23252 53884
rect 22956 53830 23002 53882
rect 23002 53830 23012 53882
rect 23036 53830 23066 53882
rect 23066 53830 23078 53882
rect 23078 53830 23092 53882
rect 23116 53830 23130 53882
rect 23130 53830 23142 53882
rect 23142 53830 23172 53882
rect 23196 53830 23206 53882
rect 23206 53830 23252 53882
rect 22956 53828 23012 53830
rect 23036 53828 23092 53830
rect 23116 53828 23172 53830
rect 23196 53828 23252 53830
rect 22190 42608 22246 42664
rect 22282 42336 22338 42392
rect 22098 41520 22154 41576
rect 22098 41248 22154 41304
rect 22098 40180 22154 40216
rect 22098 40160 22100 40180
rect 22100 40160 22152 40180
rect 22152 40160 22154 40180
rect 22956 52794 23012 52796
rect 23036 52794 23092 52796
rect 23116 52794 23172 52796
rect 23196 52794 23252 52796
rect 22956 52742 23002 52794
rect 23002 52742 23012 52794
rect 23036 52742 23066 52794
rect 23066 52742 23078 52794
rect 23078 52742 23092 52794
rect 23116 52742 23130 52794
rect 23130 52742 23142 52794
rect 23142 52742 23172 52794
rect 23196 52742 23206 52794
rect 23206 52742 23252 52794
rect 22956 52740 23012 52742
rect 23036 52740 23092 52742
rect 23116 52740 23172 52742
rect 23196 52740 23252 52742
rect 22956 51706 23012 51708
rect 23036 51706 23092 51708
rect 23116 51706 23172 51708
rect 23196 51706 23252 51708
rect 22956 51654 23002 51706
rect 23002 51654 23012 51706
rect 23036 51654 23066 51706
rect 23066 51654 23078 51706
rect 23078 51654 23092 51706
rect 23116 51654 23130 51706
rect 23130 51654 23142 51706
rect 23142 51654 23172 51706
rect 23196 51654 23206 51706
rect 23206 51654 23252 51706
rect 22956 51652 23012 51654
rect 23036 51652 23092 51654
rect 23116 51652 23172 51654
rect 23196 51652 23252 51654
rect 22956 50618 23012 50620
rect 23036 50618 23092 50620
rect 23116 50618 23172 50620
rect 23196 50618 23252 50620
rect 22956 50566 23002 50618
rect 23002 50566 23012 50618
rect 23036 50566 23066 50618
rect 23066 50566 23078 50618
rect 23078 50566 23092 50618
rect 23116 50566 23130 50618
rect 23130 50566 23142 50618
rect 23142 50566 23172 50618
rect 23196 50566 23206 50618
rect 23206 50566 23252 50618
rect 22956 50564 23012 50566
rect 23036 50564 23092 50566
rect 23116 50564 23172 50566
rect 23196 50564 23252 50566
rect 22956 49530 23012 49532
rect 23036 49530 23092 49532
rect 23116 49530 23172 49532
rect 23196 49530 23252 49532
rect 22956 49478 23002 49530
rect 23002 49478 23012 49530
rect 23036 49478 23066 49530
rect 23066 49478 23078 49530
rect 23078 49478 23092 49530
rect 23116 49478 23130 49530
rect 23130 49478 23142 49530
rect 23142 49478 23172 49530
rect 23196 49478 23206 49530
rect 23206 49478 23252 49530
rect 22956 49476 23012 49478
rect 23036 49476 23092 49478
rect 23116 49476 23172 49478
rect 23196 49476 23252 49478
rect 22956 48442 23012 48444
rect 23036 48442 23092 48444
rect 23116 48442 23172 48444
rect 23196 48442 23252 48444
rect 22956 48390 23002 48442
rect 23002 48390 23012 48442
rect 23036 48390 23066 48442
rect 23066 48390 23078 48442
rect 23078 48390 23092 48442
rect 23116 48390 23130 48442
rect 23130 48390 23142 48442
rect 23142 48390 23172 48442
rect 23196 48390 23206 48442
rect 23206 48390 23252 48442
rect 22956 48388 23012 48390
rect 23036 48388 23092 48390
rect 23116 48388 23172 48390
rect 23196 48388 23252 48390
rect 22956 47354 23012 47356
rect 23036 47354 23092 47356
rect 23116 47354 23172 47356
rect 23196 47354 23252 47356
rect 22956 47302 23002 47354
rect 23002 47302 23012 47354
rect 23036 47302 23066 47354
rect 23066 47302 23078 47354
rect 23078 47302 23092 47354
rect 23116 47302 23130 47354
rect 23130 47302 23142 47354
rect 23142 47302 23172 47354
rect 23196 47302 23206 47354
rect 23206 47302 23252 47354
rect 22956 47300 23012 47302
rect 23036 47300 23092 47302
rect 23116 47300 23172 47302
rect 23196 47300 23252 47302
rect 22098 37712 22154 37768
rect 21270 33360 21326 33416
rect 21178 30504 21234 30560
rect 20442 27124 20498 27160
rect 20442 27104 20444 27124
rect 20444 27104 20496 27124
rect 20496 27104 20498 27124
rect 20718 28056 20774 28112
rect 17956 4378 18012 4380
rect 18036 4378 18092 4380
rect 18116 4378 18172 4380
rect 18196 4378 18252 4380
rect 17956 4326 18002 4378
rect 18002 4326 18012 4378
rect 18036 4326 18066 4378
rect 18066 4326 18078 4378
rect 18078 4326 18092 4378
rect 18116 4326 18130 4378
rect 18130 4326 18142 4378
rect 18142 4326 18172 4378
rect 18196 4326 18206 4378
rect 18206 4326 18252 4378
rect 17956 4324 18012 4326
rect 18036 4324 18092 4326
rect 18116 4324 18172 4326
rect 18196 4324 18252 4326
rect 20810 26580 20866 26616
rect 20810 26560 20812 26580
rect 20812 26560 20864 26580
rect 20864 26560 20866 26580
rect 21546 32000 21602 32056
rect 21730 32952 21786 33008
rect 22006 35164 22008 35184
rect 22008 35164 22060 35184
rect 22060 35164 22062 35184
rect 22006 35128 22062 35164
rect 20718 16496 20774 16552
rect 17956 3290 18012 3292
rect 18036 3290 18092 3292
rect 18116 3290 18172 3292
rect 18196 3290 18252 3292
rect 17956 3238 18002 3290
rect 18002 3238 18012 3290
rect 18036 3238 18066 3290
rect 18066 3238 18078 3290
rect 18078 3238 18092 3290
rect 18116 3238 18130 3290
rect 18130 3238 18142 3290
rect 18142 3238 18172 3290
rect 18196 3238 18206 3290
rect 18206 3238 18252 3290
rect 17956 3236 18012 3238
rect 18036 3236 18092 3238
rect 18116 3236 18172 3238
rect 18196 3236 18252 3238
rect 17956 2202 18012 2204
rect 18036 2202 18092 2204
rect 18116 2202 18172 2204
rect 18196 2202 18252 2204
rect 17956 2150 18002 2202
rect 18002 2150 18012 2202
rect 18036 2150 18066 2202
rect 18066 2150 18078 2202
rect 18078 2150 18092 2202
rect 18116 2150 18130 2202
rect 18130 2150 18142 2202
rect 18142 2150 18172 2202
rect 18196 2150 18206 2202
rect 18206 2150 18252 2202
rect 17956 2148 18012 2150
rect 18036 2148 18092 2150
rect 18116 2148 18172 2150
rect 18196 2148 18252 2150
rect 21086 16516 21142 16552
rect 21086 16496 21088 16516
rect 21088 16496 21140 16516
rect 21140 16496 21142 16516
rect 22956 46266 23012 46268
rect 23036 46266 23092 46268
rect 23116 46266 23172 46268
rect 23196 46266 23252 46268
rect 22956 46214 23002 46266
rect 23002 46214 23012 46266
rect 23036 46214 23066 46266
rect 23066 46214 23078 46266
rect 23078 46214 23092 46266
rect 23116 46214 23130 46266
rect 23130 46214 23142 46266
rect 23142 46214 23172 46266
rect 23196 46214 23206 46266
rect 23206 46214 23252 46266
rect 22956 46212 23012 46214
rect 23036 46212 23092 46214
rect 23116 46212 23172 46214
rect 23196 46212 23252 46214
rect 22956 45178 23012 45180
rect 23036 45178 23092 45180
rect 23116 45178 23172 45180
rect 23196 45178 23252 45180
rect 22956 45126 23002 45178
rect 23002 45126 23012 45178
rect 23036 45126 23066 45178
rect 23066 45126 23078 45178
rect 23078 45126 23092 45178
rect 23116 45126 23130 45178
rect 23130 45126 23142 45178
rect 23142 45126 23172 45178
rect 23196 45126 23206 45178
rect 23206 45126 23252 45178
rect 22956 45124 23012 45126
rect 23036 45124 23092 45126
rect 23116 45124 23172 45126
rect 23196 45124 23252 45126
rect 22956 44090 23012 44092
rect 23036 44090 23092 44092
rect 23116 44090 23172 44092
rect 23196 44090 23252 44092
rect 22956 44038 23002 44090
rect 23002 44038 23012 44090
rect 23036 44038 23066 44090
rect 23066 44038 23078 44090
rect 23078 44038 23092 44090
rect 23116 44038 23130 44090
rect 23130 44038 23142 44090
rect 23142 44038 23172 44090
rect 23196 44038 23206 44090
rect 23206 44038 23252 44090
rect 22956 44036 23012 44038
rect 23036 44036 23092 44038
rect 23116 44036 23172 44038
rect 23196 44036 23252 44038
rect 22956 43002 23012 43004
rect 23036 43002 23092 43004
rect 23116 43002 23172 43004
rect 23196 43002 23252 43004
rect 22956 42950 23002 43002
rect 23002 42950 23012 43002
rect 23036 42950 23066 43002
rect 23066 42950 23078 43002
rect 23078 42950 23092 43002
rect 23116 42950 23130 43002
rect 23130 42950 23142 43002
rect 23142 42950 23172 43002
rect 23196 42950 23206 43002
rect 23206 42950 23252 43002
rect 22956 42948 23012 42950
rect 23036 42948 23092 42950
rect 23116 42948 23172 42950
rect 23196 42948 23252 42950
rect 23202 42336 23258 42392
rect 23018 42064 23074 42120
rect 22956 41914 23012 41916
rect 23036 41914 23092 41916
rect 23116 41914 23172 41916
rect 23196 41914 23252 41916
rect 22956 41862 23002 41914
rect 23002 41862 23012 41914
rect 23036 41862 23066 41914
rect 23066 41862 23078 41914
rect 23078 41862 23092 41914
rect 23116 41862 23130 41914
rect 23130 41862 23142 41914
rect 23142 41862 23172 41914
rect 23196 41862 23206 41914
rect 23206 41862 23252 41914
rect 22956 41860 23012 41862
rect 23036 41860 23092 41862
rect 23116 41860 23172 41862
rect 23196 41860 23252 41862
rect 22956 40826 23012 40828
rect 23036 40826 23092 40828
rect 23116 40826 23172 40828
rect 23196 40826 23252 40828
rect 22956 40774 23002 40826
rect 23002 40774 23012 40826
rect 23036 40774 23066 40826
rect 23066 40774 23078 40826
rect 23078 40774 23092 40826
rect 23116 40774 23130 40826
rect 23130 40774 23142 40826
rect 23142 40774 23172 40826
rect 23196 40774 23206 40826
rect 23206 40774 23252 40826
rect 22956 40772 23012 40774
rect 23036 40772 23092 40774
rect 23116 40772 23172 40774
rect 23196 40772 23252 40774
rect 22956 39738 23012 39740
rect 23036 39738 23092 39740
rect 23116 39738 23172 39740
rect 23196 39738 23252 39740
rect 22956 39686 23002 39738
rect 23002 39686 23012 39738
rect 23036 39686 23066 39738
rect 23066 39686 23078 39738
rect 23078 39686 23092 39738
rect 23116 39686 23130 39738
rect 23130 39686 23142 39738
rect 23142 39686 23172 39738
rect 23196 39686 23206 39738
rect 23206 39686 23252 39738
rect 22956 39684 23012 39686
rect 23036 39684 23092 39686
rect 23116 39684 23172 39686
rect 23196 39684 23252 39686
rect 22956 38650 23012 38652
rect 23036 38650 23092 38652
rect 23116 38650 23172 38652
rect 23196 38650 23252 38652
rect 22956 38598 23002 38650
rect 23002 38598 23012 38650
rect 23036 38598 23066 38650
rect 23066 38598 23078 38650
rect 23078 38598 23092 38650
rect 23116 38598 23130 38650
rect 23130 38598 23142 38650
rect 23142 38598 23172 38650
rect 23196 38598 23206 38650
rect 23206 38598 23252 38650
rect 22956 38596 23012 38598
rect 23036 38596 23092 38598
rect 23116 38596 23172 38598
rect 23196 38596 23252 38598
rect 22650 38004 22706 38040
rect 22650 37984 22652 38004
rect 22652 37984 22704 38004
rect 22704 37984 22706 38004
rect 22374 34992 22430 35048
rect 22190 33088 22246 33144
rect 22650 34992 22706 35048
rect 22956 37562 23012 37564
rect 23036 37562 23092 37564
rect 23116 37562 23172 37564
rect 23196 37562 23252 37564
rect 22956 37510 23002 37562
rect 23002 37510 23012 37562
rect 23036 37510 23066 37562
rect 23066 37510 23078 37562
rect 23078 37510 23092 37562
rect 23116 37510 23130 37562
rect 23130 37510 23142 37562
rect 23142 37510 23172 37562
rect 23196 37510 23206 37562
rect 23206 37510 23252 37562
rect 22956 37508 23012 37510
rect 23036 37508 23092 37510
rect 23116 37508 23172 37510
rect 23196 37508 23252 37510
rect 24674 55392 24730 55448
rect 24766 54576 24822 54632
rect 25042 53760 25098 53816
rect 25318 53760 25374 53816
rect 23938 52944 23994 53000
rect 25042 53216 25098 53272
rect 25042 52944 25098 53000
rect 24766 52128 24822 52184
rect 23386 37440 23442 37496
rect 22956 36474 23012 36476
rect 23036 36474 23092 36476
rect 23116 36474 23172 36476
rect 23196 36474 23252 36476
rect 22956 36422 23002 36474
rect 23002 36422 23012 36474
rect 23036 36422 23066 36474
rect 23066 36422 23078 36474
rect 23078 36422 23092 36474
rect 23116 36422 23130 36474
rect 23130 36422 23142 36474
rect 23142 36422 23172 36474
rect 23196 36422 23206 36474
rect 23206 36422 23252 36474
rect 22956 36420 23012 36422
rect 23036 36420 23092 36422
rect 23116 36420 23172 36422
rect 23196 36420 23252 36422
rect 22742 34312 22798 34368
rect 22956 35386 23012 35388
rect 23036 35386 23092 35388
rect 23116 35386 23172 35388
rect 23196 35386 23252 35388
rect 22956 35334 23002 35386
rect 23002 35334 23012 35386
rect 23036 35334 23066 35386
rect 23066 35334 23078 35386
rect 23078 35334 23092 35386
rect 23116 35334 23130 35386
rect 23130 35334 23142 35386
rect 23142 35334 23172 35386
rect 23196 35334 23206 35386
rect 23206 35334 23252 35386
rect 22956 35332 23012 35334
rect 23036 35332 23092 35334
rect 23116 35332 23172 35334
rect 23196 35332 23252 35334
rect 23202 35128 23258 35184
rect 22956 34298 23012 34300
rect 23036 34298 23092 34300
rect 23116 34298 23172 34300
rect 23196 34298 23252 34300
rect 22956 34246 23002 34298
rect 23002 34246 23012 34298
rect 23036 34246 23066 34298
rect 23066 34246 23078 34298
rect 23078 34246 23092 34298
rect 23116 34246 23130 34298
rect 23130 34246 23142 34298
rect 23142 34246 23172 34298
rect 23196 34246 23206 34298
rect 23206 34246 23252 34298
rect 22956 34244 23012 34246
rect 23036 34244 23092 34246
rect 23116 34244 23172 34246
rect 23196 34244 23252 34246
rect 22926 34060 22982 34096
rect 22926 34040 22928 34060
rect 22928 34040 22980 34060
rect 22980 34040 22982 34060
rect 22956 33210 23012 33212
rect 23036 33210 23092 33212
rect 23116 33210 23172 33212
rect 23196 33210 23252 33212
rect 22956 33158 23002 33210
rect 23002 33158 23012 33210
rect 23036 33158 23066 33210
rect 23066 33158 23078 33210
rect 23078 33158 23092 33210
rect 23116 33158 23130 33210
rect 23130 33158 23142 33210
rect 23142 33158 23172 33210
rect 23196 33158 23206 33210
rect 23206 33158 23252 33210
rect 22956 33156 23012 33158
rect 23036 33156 23092 33158
rect 23116 33156 23172 33158
rect 23196 33156 23252 33158
rect 23018 32988 23020 33008
rect 23020 32988 23072 33008
rect 23072 32988 23074 33008
rect 23018 32952 23074 32988
rect 24490 48048 24546 48104
rect 24398 45736 24454 45792
rect 24122 40024 24178 40080
rect 24030 39072 24086 39128
rect 24582 44784 24638 44840
rect 24490 43968 24546 44024
rect 24582 43152 24638 43208
rect 24398 41384 24454 41440
rect 24306 38392 24362 38448
rect 24766 46552 24822 46608
rect 24766 45600 24822 45656
rect 24766 44240 24822 44296
rect 25042 50496 25098 50552
rect 25502 51348 25504 51368
rect 25504 51348 25556 51368
rect 25556 51348 25558 51368
rect 25502 51312 25558 51348
rect 25318 49680 25374 49736
rect 25318 48864 25374 48920
rect 25502 47232 25558 47288
rect 24858 42744 24914 42800
rect 24766 40704 24822 40760
rect 24674 36624 24730 36680
rect 22956 32122 23012 32124
rect 23036 32122 23092 32124
rect 23116 32122 23172 32124
rect 23196 32122 23252 32124
rect 22956 32070 23002 32122
rect 23002 32070 23012 32122
rect 23036 32070 23066 32122
rect 23066 32070 23078 32122
rect 23078 32070 23092 32122
rect 23116 32070 23130 32122
rect 23130 32070 23142 32122
rect 23142 32070 23172 32122
rect 23196 32070 23206 32122
rect 23206 32070 23252 32122
rect 22956 32068 23012 32070
rect 23036 32068 23092 32070
rect 23116 32068 23172 32070
rect 23196 32068 23252 32070
rect 22956 31034 23012 31036
rect 23036 31034 23092 31036
rect 23116 31034 23172 31036
rect 23196 31034 23252 31036
rect 22956 30982 23002 31034
rect 23002 30982 23012 31034
rect 23036 30982 23066 31034
rect 23066 30982 23078 31034
rect 23078 30982 23092 31034
rect 23116 30982 23130 31034
rect 23130 30982 23142 31034
rect 23142 30982 23172 31034
rect 23196 30982 23206 31034
rect 23206 30982 23252 31034
rect 22956 30980 23012 30982
rect 23036 30980 23092 30982
rect 23116 30980 23172 30982
rect 23196 30980 23252 30982
rect 22956 29946 23012 29948
rect 23036 29946 23092 29948
rect 23116 29946 23172 29948
rect 23196 29946 23252 29948
rect 22956 29894 23002 29946
rect 23002 29894 23012 29946
rect 23036 29894 23066 29946
rect 23066 29894 23078 29946
rect 23078 29894 23092 29946
rect 23116 29894 23130 29946
rect 23130 29894 23142 29946
rect 23142 29894 23172 29946
rect 23196 29894 23206 29946
rect 23206 29894 23252 29946
rect 22956 29892 23012 29894
rect 23036 29892 23092 29894
rect 23116 29892 23172 29894
rect 23196 29892 23252 29894
rect 23570 33496 23626 33552
rect 24674 34992 24730 35048
rect 22956 28858 23012 28860
rect 23036 28858 23092 28860
rect 23116 28858 23172 28860
rect 23196 28858 23252 28860
rect 22956 28806 23002 28858
rect 23002 28806 23012 28858
rect 23036 28806 23066 28858
rect 23066 28806 23078 28858
rect 23078 28806 23092 28858
rect 23116 28806 23130 28858
rect 23130 28806 23142 28858
rect 23142 28806 23172 28858
rect 23196 28806 23206 28858
rect 23206 28806 23252 28858
rect 22956 28804 23012 28806
rect 23036 28804 23092 28806
rect 23116 28804 23172 28806
rect 23196 28804 23252 28806
rect 22956 27770 23012 27772
rect 23036 27770 23092 27772
rect 23116 27770 23172 27772
rect 23196 27770 23252 27772
rect 22956 27718 23002 27770
rect 23002 27718 23012 27770
rect 23036 27718 23066 27770
rect 23066 27718 23078 27770
rect 23078 27718 23092 27770
rect 23116 27718 23130 27770
rect 23130 27718 23142 27770
rect 23142 27718 23172 27770
rect 23196 27718 23206 27770
rect 23206 27718 23252 27770
rect 22956 27716 23012 27718
rect 23036 27716 23092 27718
rect 23116 27716 23172 27718
rect 23196 27716 23252 27718
rect 24122 27648 24178 27704
rect 22558 26016 22614 26072
rect 22956 26682 23012 26684
rect 23036 26682 23092 26684
rect 23116 26682 23172 26684
rect 23196 26682 23252 26684
rect 22956 26630 23002 26682
rect 23002 26630 23012 26682
rect 23036 26630 23066 26682
rect 23066 26630 23078 26682
rect 23078 26630 23092 26682
rect 23116 26630 23130 26682
rect 23130 26630 23142 26682
rect 23142 26630 23172 26682
rect 23196 26630 23206 26682
rect 23206 26630 23252 26682
rect 22956 26628 23012 26630
rect 23036 26628 23092 26630
rect 23116 26628 23172 26630
rect 23196 26628 23252 26630
rect 23386 26832 23442 26888
rect 22956 25594 23012 25596
rect 23036 25594 23092 25596
rect 23116 25594 23172 25596
rect 23196 25594 23252 25596
rect 22956 25542 23002 25594
rect 23002 25542 23012 25594
rect 23036 25542 23066 25594
rect 23066 25542 23078 25594
rect 23078 25542 23092 25594
rect 23116 25542 23130 25594
rect 23130 25542 23142 25594
rect 23142 25542 23172 25594
rect 23196 25542 23206 25594
rect 23206 25542 23252 25594
rect 22956 25540 23012 25542
rect 23036 25540 23092 25542
rect 23116 25540 23172 25542
rect 23196 25540 23252 25542
rect 22956 24506 23012 24508
rect 23036 24506 23092 24508
rect 23116 24506 23172 24508
rect 23196 24506 23252 24508
rect 22956 24454 23002 24506
rect 23002 24454 23012 24506
rect 23036 24454 23066 24506
rect 23066 24454 23078 24506
rect 23078 24454 23092 24506
rect 23116 24454 23130 24506
rect 23130 24454 23142 24506
rect 23142 24454 23172 24506
rect 23196 24454 23206 24506
rect 23206 24454 23252 24506
rect 22956 24452 23012 24454
rect 23036 24452 23092 24454
rect 23116 24452 23172 24454
rect 23196 24452 23252 24454
rect 22956 23418 23012 23420
rect 23036 23418 23092 23420
rect 23116 23418 23172 23420
rect 23196 23418 23252 23420
rect 22956 23366 23002 23418
rect 23002 23366 23012 23418
rect 23036 23366 23066 23418
rect 23066 23366 23078 23418
rect 23078 23366 23092 23418
rect 23116 23366 23130 23418
rect 23130 23366 23142 23418
rect 23142 23366 23172 23418
rect 23196 23366 23206 23418
rect 23206 23366 23252 23418
rect 22956 23364 23012 23366
rect 23036 23364 23092 23366
rect 23116 23364 23172 23366
rect 23196 23364 23252 23366
rect 23294 22752 23350 22808
rect 22956 22330 23012 22332
rect 23036 22330 23092 22332
rect 23116 22330 23172 22332
rect 23196 22330 23252 22332
rect 22956 22278 23002 22330
rect 23002 22278 23012 22330
rect 23036 22278 23066 22330
rect 23066 22278 23078 22330
rect 23078 22278 23092 22330
rect 23116 22278 23130 22330
rect 23130 22278 23142 22330
rect 23142 22278 23172 22330
rect 23196 22278 23206 22330
rect 23206 22278 23252 22330
rect 22956 22276 23012 22278
rect 23036 22276 23092 22278
rect 23116 22276 23172 22278
rect 23196 22276 23252 22278
rect 22956 21242 23012 21244
rect 23036 21242 23092 21244
rect 23116 21242 23172 21244
rect 23196 21242 23252 21244
rect 22956 21190 23002 21242
rect 23002 21190 23012 21242
rect 23036 21190 23066 21242
rect 23066 21190 23078 21242
rect 23078 21190 23092 21242
rect 23116 21190 23130 21242
rect 23130 21190 23142 21242
rect 23142 21190 23172 21242
rect 23196 21190 23206 21242
rect 23206 21190 23252 21242
rect 22956 21188 23012 21190
rect 23036 21188 23092 21190
rect 23116 21188 23172 21190
rect 23196 21188 23252 21190
rect 23386 21120 23442 21176
rect 22956 20154 23012 20156
rect 23036 20154 23092 20156
rect 23116 20154 23172 20156
rect 23196 20154 23252 20156
rect 22956 20102 23002 20154
rect 23002 20102 23012 20154
rect 23036 20102 23066 20154
rect 23066 20102 23078 20154
rect 23078 20102 23092 20154
rect 23116 20102 23130 20154
rect 23130 20102 23142 20154
rect 23142 20102 23172 20154
rect 23196 20102 23206 20154
rect 23206 20102 23252 20154
rect 22956 20100 23012 20102
rect 23036 20100 23092 20102
rect 23116 20100 23172 20102
rect 23196 20100 23252 20102
rect 22956 19066 23012 19068
rect 23036 19066 23092 19068
rect 23116 19066 23172 19068
rect 23196 19066 23252 19068
rect 22956 19014 23002 19066
rect 23002 19014 23012 19066
rect 23036 19014 23066 19066
rect 23066 19014 23078 19066
rect 23078 19014 23092 19066
rect 23116 19014 23130 19066
rect 23130 19014 23142 19066
rect 23142 19014 23172 19066
rect 23196 19014 23206 19066
rect 23206 19014 23252 19066
rect 22956 19012 23012 19014
rect 23036 19012 23092 19014
rect 23116 19012 23172 19014
rect 23196 19012 23252 19014
rect 22956 17978 23012 17980
rect 23036 17978 23092 17980
rect 23116 17978 23172 17980
rect 23196 17978 23252 17980
rect 22956 17926 23002 17978
rect 23002 17926 23012 17978
rect 23036 17926 23066 17978
rect 23066 17926 23078 17978
rect 23078 17926 23092 17978
rect 23116 17926 23130 17978
rect 23130 17926 23142 17978
rect 23142 17926 23172 17978
rect 23196 17926 23206 17978
rect 23206 17926 23252 17978
rect 22956 17924 23012 17926
rect 23036 17924 23092 17926
rect 23116 17924 23172 17926
rect 23196 17924 23252 17926
rect 23386 17856 23442 17912
rect 23846 23568 23902 23624
rect 22956 16890 23012 16892
rect 23036 16890 23092 16892
rect 23116 16890 23172 16892
rect 23196 16890 23252 16892
rect 22956 16838 23002 16890
rect 23002 16838 23012 16890
rect 23036 16838 23066 16890
rect 23066 16838 23078 16890
rect 23078 16838 23092 16890
rect 23116 16838 23130 16890
rect 23130 16838 23142 16890
rect 23142 16838 23172 16890
rect 23196 16838 23206 16890
rect 23206 16838 23252 16890
rect 22956 16836 23012 16838
rect 23036 16836 23092 16838
rect 23116 16836 23172 16838
rect 23196 16836 23252 16838
rect 22956 15802 23012 15804
rect 23036 15802 23092 15804
rect 23116 15802 23172 15804
rect 23196 15802 23252 15804
rect 22956 15750 23002 15802
rect 23002 15750 23012 15802
rect 23036 15750 23066 15802
rect 23066 15750 23078 15802
rect 23078 15750 23092 15802
rect 23116 15750 23130 15802
rect 23130 15750 23142 15802
rect 23142 15750 23172 15802
rect 23196 15750 23206 15802
rect 23206 15750 23252 15802
rect 22956 15748 23012 15750
rect 23036 15748 23092 15750
rect 23116 15748 23172 15750
rect 23196 15748 23252 15750
rect 21638 2352 21694 2408
rect 22956 14714 23012 14716
rect 23036 14714 23092 14716
rect 23116 14714 23172 14716
rect 23196 14714 23252 14716
rect 22956 14662 23002 14714
rect 23002 14662 23012 14714
rect 23036 14662 23066 14714
rect 23066 14662 23078 14714
rect 23078 14662 23092 14714
rect 23116 14662 23130 14714
rect 23130 14662 23142 14714
rect 23142 14662 23172 14714
rect 23196 14662 23206 14714
rect 23206 14662 23252 14714
rect 22956 14660 23012 14662
rect 23036 14660 23092 14662
rect 23116 14660 23172 14662
rect 23196 14660 23252 14662
rect 22098 3984 22154 4040
rect 22956 13626 23012 13628
rect 23036 13626 23092 13628
rect 23116 13626 23172 13628
rect 23196 13626 23252 13628
rect 22956 13574 23002 13626
rect 23002 13574 23012 13626
rect 23036 13574 23066 13626
rect 23066 13574 23078 13626
rect 23078 13574 23092 13626
rect 23116 13574 23130 13626
rect 23130 13574 23142 13626
rect 23142 13574 23172 13626
rect 23196 13574 23206 13626
rect 23206 13574 23252 13626
rect 22956 13572 23012 13574
rect 23036 13572 23092 13574
rect 23116 13572 23172 13574
rect 23196 13572 23252 13574
rect 25318 38256 25374 38312
rect 24858 35808 24914 35864
rect 25318 34196 25374 34232
rect 25318 34176 25320 34196
rect 25320 34176 25372 34196
rect 25372 34176 25374 34196
rect 25410 33360 25466 33416
rect 25318 32544 25374 32600
rect 25318 31764 25320 31784
rect 25320 31764 25372 31784
rect 25372 31764 25374 31784
rect 25318 31728 25374 31764
rect 25318 30932 25374 30968
rect 25318 30912 25320 30932
rect 25320 30912 25372 30932
rect 25372 30912 25374 30932
rect 25134 30540 25136 30560
rect 25136 30540 25188 30560
rect 25188 30540 25190 30560
rect 25134 30504 25190 30540
rect 25318 30096 25374 30152
rect 22956 12538 23012 12540
rect 23036 12538 23092 12540
rect 23116 12538 23172 12540
rect 23196 12538 23252 12540
rect 22956 12486 23002 12538
rect 23002 12486 23012 12538
rect 23036 12486 23066 12538
rect 23066 12486 23078 12538
rect 23078 12486 23092 12538
rect 23116 12486 23130 12538
rect 23130 12486 23142 12538
rect 23142 12486 23172 12538
rect 23196 12486 23206 12538
rect 23206 12486 23252 12538
rect 22956 12484 23012 12486
rect 23036 12484 23092 12486
rect 23116 12484 23172 12486
rect 23196 12484 23252 12486
rect 24858 24384 24914 24440
rect 24858 21936 24914 21992
rect 25226 28484 25282 28520
rect 25226 28464 25228 28484
rect 25228 28464 25280 28484
rect 25280 28464 25282 28484
rect 25134 25200 25190 25256
rect 24950 20304 25006 20360
rect 25502 29300 25558 29336
rect 25502 29280 25504 29300
rect 25504 29280 25556 29300
rect 25556 29280 25558 29300
rect 24766 19488 24822 19544
rect 24674 18672 24730 18728
rect 24766 17040 24822 17096
rect 24674 16224 24730 16280
rect 24950 15428 25006 15464
rect 24950 15408 24952 15428
rect 24952 15408 25004 15428
rect 25004 15408 25006 15428
rect 22956 11450 23012 11452
rect 23036 11450 23092 11452
rect 23116 11450 23172 11452
rect 23196 11450 23252 11452
rect 22956 11398 23002 11450
rect 23002 11398 23012 11450
rect 23036 11398 23066 11450
rect 23066 11398 23078 11450
rect 23078 11398 23092 11450
rect 23116 11398 23130 11450
rect 23130 11398 23142 11450
rect 23142 11398 23172 11450
rect 23196 11398 23206 11450
rect 23206 11398 23252 11450
rect 22956 11396 23012 11398
rect 23036 11396 23092 11398
rect 23116 11396 23172 11398
rect 23196 11396 23252 11398
rect 22956 10362 23012 10364
rect 23036 10362 23092 10364
rect 23116 10362 23172 10364
rect 23196 10362 23252 10364
rect 22956 10310 23002 10362
rect 23002 10310 23012 10362
rect 23036 10310 23066 10362
rect 23066 10310 23078 10362
rect 23078 10310 23092 10362
rect 23116 10310 23130 10362
rect 23130 10310 23142 10362
rect 23142 10310 23172 10362
rect 23196 10310 23206 10362
rect 23206 10310 23252 10362
rect 22956 10308 23012 10310
rect 23036 10308 23092 10310
rect 23116 10308 23172 10310
rect 23196 10308 23252 10310
rect 22956 9274 23012 9276
rect 23036 9274 23092 9276
rect 23116 9274 23172 9276
rect 23196 9274 23252 9276
rect 22956 9222 23002 9274
rect 23002 9222 23012 9274
rect 23036 9222 23066 9274
rect 23066 9222 23078 9274
rect 23078 9222 23092 9274
rect 23116 9222 23130 9274
rect 23130 9222 23142 9274
rect 23142 9222 23172 9274
rect 23196 9222 23206 9274
rect 23206 9222 23252 9274
rect 22956 9220 23012 9222
rect 23036 9220 23092 9222
rect 23116 9220 23172 9222
rect 23196 9220 23252 9222
rect 22956 8186 23012 8188
rect 23036 8186 23092 8188
rect 23116 8186 23172 8188
rect 23196 8186 23252 8188
rect 22956 8134 23002 8186
rect 23002 8134 23012 8186
rect 23036 8134 23066 8186
rect 23066 8134 23078 8186
rect 23078 8134 23092 8186
rect 23116 8134 23130 8186
rect 23130 8134 23142 8186
rect 23142 8134 23172 8186
rect 23196 8134 23206 8186
rect 23206 8134 23252 8186
rect 22956 8132 23012 8134
rect 23036 8132 23092 8134
rect 23116 8132 23172 8134
rect 23196 8132 23252 8134
rect 22956 7098 23012 7100
rect 23036 7098 23092 7100
rect 23116 7098 23172 7100
rect 23196 7098 23252 7100
rect 22956 7046 23002 7098
rect 23002 7046 23012 7098
rect 23036 7046 23066 7098
rect 23066 7046 23078 7098
rect 23078 7046 23092 7098
rect 23116 7046 23130 7098
rect 23130 7046 23142 7098
rect 23142 7046 23172 7098
rect 23196 7046 23206 7098
rect 23206 7046 23252 7098
rect 22956 7044 23012 7046
rect 23036 7044 23092 7046
rect 23116 7044 23172 7046
rect 23196 7044 23252 7046
rect 22956 6010 23012 6012
rect 23036 6010 23092 6012
rect 23116 6010 23172 6012
rect 23196 6010 23252 6012
rect 22956 5958 23002 6010
rect 23002 5958 23012 6010
rect 23036 5958 23066 6010
rect 23066 5958 23078 6010
rect 23078 5958 23092 6010
rect 23116 5958 23130 6010
rect 23130 5958 23142 6010
rect 23142 5958 23172 6010
rect 23196 5958 23206 6010
rect 23206 5958 23252 6010
rect 22956 5956 23012 5958
rect 23036 5956 23092 5958
rect 23116 5956 23172 5958
rect 23196 5956 23252 5958
rect 22956 4922 23012 4924
rect 23036 4922 23092 4924
rect 23116 4922 23172 4924
rect 23196 4922 23252 4924
rect 22956 4870 23002 4922
rect 23002 4870 23012 4922
rect 23036 4870 23066 4922
rect 23066 4870 23078 4922
rect 23078 4870 23092 4922
rect 23116 4870 23130 4922
rect 23130 4870 23142 4922
rect 23142 4870 23172 4922
rect 23196 4870 23206 4922
rect 23206 4870 23252 4922
rect 22956 4868 23012 4870
rect 23036 4868 23092 4870
rect 23116 4868 23172 4870
rect 23196 4868 23252 4870
rect 25134 14592 25190 14648
rect 24766 13776 24822 13832
rect 24950 12960 25006 13016
rect 24766 11328 24822 11384
rect 24674 10512 24730 10568
rect 25134 12144 25190 12200
rect 24950 9696 25006 9752
rect 25134 8880 25190 8936
rect 25134 8064 25190 8120
rect 23386 4800 23442 4856
rect 24766 7248 24822 7304
rect 25778 6432 25834 6488
rect 24766 5616 24822 5672
rect 22956 3834 23012 3836
rect 23036 3834 23092 3836
rect 23116 3834 23172 3836
rect 23196 3834 23252 3836
rect 22956 3782 23002 3834
rect 23002 3782 23012 3834
rect 23036 3782 23066 3834
rect 23066 3782 23078 3834
rect 23078 3782 23092 3834
rect 23116 3782 23130 3834
rect 23130 3782 23142 3834
rect 23142 3782 23172 3834
rect 23196 3782 23206 3834
rect 23206 3782 23252 3834
rect 22956 3780 23012 3782
rect 23036 3780 23092 3782
rect 23116 3780 23172 3782
rect 23196 3780 23252 3782
rect 23754 3440 23810 3496
rect 22742 3168 22798 3224
rect 22956 2746 23012 2748
rect 23036 2746 23092 2748
rect 23116 2746 23172 2748
rect 23196 2746 23252 2748
rect 22956 2694 23002 2746
rect 23002 2694 23012 2746
rect 23036 2694 23066 2746
rect 23066 2694 23078 2746
rect 23078 2694 23092 2746
rect 23116 2694 23130 2746
rect 23130 2694 23142 2746
rect 23142 2694 23172 2746
rect 23196 2694 23206 2746
rect 23206 2694 23252 2746
rect 22956 2692 23012 2694
rect 23036 2692 23092 2694
rect 23116 2692 23172 2694
rect 23196 2692 23252 2694
rect 25318 1536 25374 1592
rect 24950 720 25006 776
<< metal3 >>
rect 24485 56266 24551 56269
rect 26200 56266 27000 56296
rect 24485 56264 27000 56266
rect 24485 56208 24490 56264
rect 24546 56208 27000 56264
rect 24485 56206 27000 56208
rect 24485 56203 24551 56206
rect 26200 56176 27000 56206
rect 0 55450 800 55480
rect 2773 55450 2839 55453
rect 0 55448 2839 55450
rect 0 55392 2778 55448
rect 2834 55392 2839 55448
rect 0 55390 2839 55392
rect 0 55360 800 55390
rect 2773 55387 2839 55390
rect 24669 55450 24735 55453
rect 26200 55450 27000 55480
rect 24669 55448 27000 55450
rect 24669 55392 24674 55448
rect 24730 55392 27000 55448
rect 24669 55390 27000 55392
rect 24669 55387 24735 55390
rect 26200 55360 27000 55390
rect 24761 54634 24827 54637
rect 26200 54634 27000 54664
rect 24761 54632 27000 54634
rect 24761 54576 24766 54632
rect 24822 54576 27000 54632
rect 24761 54574 27000 54576
rect 24761 54571 24827 54574
rect 26200 54544 27000 54574
rect 7946 54432 8262 54433
rect 7946 54368 7952 54432
rect 8016 54368 8032 54432
rect 8096 54368 8112 54432
rect 8176 54368 8192 54432
rect 8256 54368 8262 54432
rect 7946 54367 8262 54368
rect 17946 54432 18262 54433
rect 17946 54368 17952 54432
rect 18016 54368 18032 54432
rect 18096 54368 18112 54432
rect 18176 54368 18192 54432
rect 18256 54368 18262 54432
rect 17946 54367 18262 54368
rect 15745 53954 15811 53957
rect 22369 53956 22435 53957
rect 15878 53954 15884 53956
rect 15745 53952 15884 53954
rect 15745 53896 15750 53952
rect 15806 53896 15884 53952
rect 15745 53894 15884 53896
rect 15745 53891 15811 53894
rect 15878 53892 15884 53894
rect 15948 53892 15954 53956
rect 22318 53954 22324 53956
rect 22278 53894 22324 53954
rect 22388 53952 22435 53956
rect 22430 53896 22435 53952
rect 22318 53892 22324 53894
rect 22388 53892 22435 53896
rect 22369 53891 22435 53892
rect 2946 53888 3262 53889
rect 2946 53824 2952 53888
rect 3016 53824 3032 53888
rect 3096 53824 3112 53888
rect 3176 53824 3192 53888
rect 3256 53824 3262 53888
rect 2946 53823 3262 53824
rect 12946 53888 13262 53889
rect 12946 53824 12952 53888
rect 13016 53824 13032 53888
rect 13096 53824 13112 53888
rect 13176 53824 13192 53888
rect 13256 53824 13262 53888
rect 12946 53823 13262 53824
rect 22946 53888 23262 53889
rect 22946 53824 22952 53888
rect 23016 53824 23032 53888
rect 23096 53824 23112 53888
rect 23176 53824 23192 53888
rect 23256 53824 23262 53888
rect 22946 53823 23262 53824
rect 25037 53818 25103 53821
rect 25313 53818 25379 53821
rect 26200 53818 27000 53848
rect 25037 53816 27000 53818
rect 25037 53760 25042 53816
rect 25098 53760 25318 53816
rect 25374 53760 27000 53816
rect 25037 53758 27000 53760
rect 25037 53755 25103 53758
rect 25313 53755 25379 53758
rect 26200 53728 27000 53758
rect 7946 53344 8262 53345
rect 7946 53280 7952 53344
rect 8016 53280 8032 53344
rect 8096 53280 8112 53344
rect 8176 53280 8192 53344
rect 8256 53280 8262 53344
rect 7946 53279 8262 53280
rect 17946 53344 18262 53345
rect 17946 53280 17952 53344
rect 18016 53280 18032 53344
rect 18096 53280 18112 53344
rect 18176 53280 18192 53344
rect 18256 53280 18262 53344
rect 17946 53279 18262 53280
rect 22502 53212 22508 53276
rect 22572 53274 22578 53276
rect 25037 53274 25103 53277
rect 22572 53272 25103 53274
rect 22572 53216 25042 53272
rect 25098 53216 25103 53272
rect 22572 53214 25103 53216
rect 22572 53212 22578 53214
rect 25037 53211 25103 53214
rect 0 53002 800 53032
rect 3417 53002 3483 53005
rect 0 53000 3483 53002
rect 0 52944 3422 53000
rect 3478 52944 3483 53000
rect 0 52942 3483 52944
rect 0 52912 800 52942
rect 3417 52939 3483 52942
rect 21030 52940 21036 53004
rect 21100 53002 21106 53004
rect 23933 53002 23999 53005
rect 21100 53000 23999 53002
rect 21100 52944 23938 53000
rect 23994 52944 23999 53000
rect 21100 52942 23999 52944
rect 21100 52940 21106 52942
rect 23933 52939 23999 52942
rect 25037 53002 25103 53005
rect 26200 53002 27000 53032
rect 25037 53000 27000 53002
rect 25037 52944 25042 53000
rect 25098 52944 27000 53000
rect 25037 52942 27000 52944
rect 25037 52939 25103 52942
rect 26200 52912 27000 52942
rect 2946 52800 3262 52801
rect 2946 52736 2952 52800
rect 3016 52736 3032 52800
rect 3096 52736 3112 52800
rect 3176 52736 3192 52800
rect 3256 52736 3262 52800
rect 2946 52735 3262 52736
rect 12946 52800 13262 52801
rect 12946 52736 12952 52800
rect 13016 52736 13032 52800
rect 13096 52736 13112 52800
rect 13176 52736 13192 52800
rect 13256 52736 13262 52800
rect 12946 52735 13262 52736
rect 22946 52800 23262 52801
rect 22946 52736 22952 52800
rect 23016 52736 23032 52800
rect 23096 52736 23112 52800
rect 23176 52736 23192 52800
rect 23256 52736 23262 52800
rect 22946 52735 23262 52736
rect 13629 52594 13695 52597
rect 13997 52596 14063 52597
rect 13854 52594 13860 52596
rect 13629 52592 13860 52594
rect 13629 52536 13634 52592
rect 13690 52536 13860 52592
rect 13629 52534 13860 52536
rect 13629 52531 13695 52534
rect 13854 52532 13860 52534
rect 13924 52532 13930 52596
rect 13997 52592 14044 52596
rect 14108 52594 14114 52596
rect 13997 52536 14002 52592
rect 13997 52532 14044 52536
rect 14108 52534 14154 52594
rect 14108 52532 14114 52534
rect 15326 52532 15332 52596
rect 15396 52594 15402 52596
rect 15745 52594 15811 52597
rect 15396 52592 15811 52594
rect 15396 52536 15750 52592
rect 15806 52536 15811 52592
rect 15396 52534 15811 52536
rect 15396 52532 15402 52534
rect 13997 52531 14063 52532
rect 15745 52531 15811 52534
rect 16849 52594 16915 52597
rect 17718 52594 17724 52596
rect 16849 52592 17724 52594
rect 16849 52536 16854 52592
rect 16910 52536 17724 52592
rect 16849 52534 17724 52536
rect 16849 52531 16915 52534
rect 17718 52532 17724 52534
rect 17788 52532 17794 52596
rect 7946 52256 8262 52257
rect 7946 52192 7952 52256
rect 8016 52192 8032 52256
rect 8096 52192 8112 52256
rect 8176 52192 8192 52256
rect 8256 52192 8262 52256
rect 7946 52191 8262 52192
rect 17946 52256 18262 52257
rect 17946 52192 17952 52256
rect 18016 52192 18032 52256
rect 18096 52192 18112 52256
rect 18176 52192 18192 52256
rect 18256 52192 18262 52256
rect 17946 52191 18262 52192
rect 24761 52186 24827 52189
rect 26200 52186 27000 52216
rect 24761 52184 27000 52186
rect 24761 52128 24766 52184
rect 24822 52128 27000 52184
rect 24761 52126 27000 52128
rect 24761 52123 24827 52126
rect 26200 52096 27000 52126
rect 2946 51712 3262 51713
rect 2946 51648 2952 51712
rect 3016 51648 3032 51712
rect 3096 51648 3112 51712
rect 3176 51648 3192 51712
rect 3256 51648 3262 51712
rect 2946 51647 3262 51648
rect 12946 51712 13262 51713
rect 12946 51648 12952 51712
rect 13016 51648 13032 51712
rect 13096 51648 13112 51712
rect 13176 51648 13192 51712
rect 13256 51648 13262 51712
rect 12946 51647 13262 51648
rect 22946 51712 23262 51713
rect 22946 51648 22952 51712
rect 23016 51648 23032 51712
rect 23096 51648 23112 51712
rect 23176 51648 23192 51712
rect 23256 51648 23262 51712
rect 22946 51647 23262 51648
rect 25497 51370 25563 51373
rect 26200 51370 27000 51400
rect 25497 51368 27000 51370
rect 25497 51312 25502 51368
rect 25558 51312 27000 51368
rect 25497 51310 27000 51312
rect 25497 51307 25563 51310
rect 26200 51280 27000 51310
rect 7946 51168 8262 51169
rect 7946 51104 7952 51168
rect 8016 51104 8032 51168
rect 8096 51104 8112 51168
rect 8176 51104 8192 51168
rect 8256 51104 8262 51168
rect 7946 51103 8262 51104
rect 17946 51168 18262 51169
rect 17946 51104 17952 51168
rect 18016 51104 18032 51168
rect 18096 51104 18112 51168
rect 18176 51104 18192 51168
rect 18256 51104 18262 51168
rect 17946 51103 18262 51104
rect 2946 50624 3262 50625
rect 0 50554 800 50584
rect 2946 50560 2952 50624
rect 3016 50560 3032 50624
rect 3096 50560 3112 50624
rect 3176 50560 3192 50624
rect 3256 50560 3262 50624
rect 2946 50559 3262 50560
rect 12946 50624 13262 50625
rect 12946 50560 12952 50624
rect 13016 50560 13032 50624
rect 13096 50560 13112 50624
rect 13176 50560 13192 50624
rect 13256 50560 13262 50624
rect 12946 50559 13262 50560
rect 22946 50624 23262 50625
rect 22946 50560 22952 50624
rect 23016 50560 23032 50624
rect 23096 50560 23112 50624
rect 23176 50560 23192 50624
rect 23256 50560 23262 50624
rect 22946 50559 23262 50560
rect 25037 50554 25103 50557
rect 26200 50554 27000 50584
rect 0 50494 1778 50554
rect 0 50464 800 50494
rect 1718 50418 1778 50494
rect 25037 50552 27000 50554
rect 25037 50496 25042 50552
rect 25098 50496 27000 50552
rect 25037 50494 27000 50496
rect 25037 50491 25103 50494
rect 26200 50464 27000 50494
rect 3969 50418 4035 50421
rect 1718 50416 4035 50418
rect 1718 50360 3974 50416
rect 4030 50360 4035 50416
rect 1718 50358 4035 50360
rect 3969 50355 4035 50358
rect 7946 50080 8262 50081
rect 7946 50016 7952 50080
rect 8016 50016 8032 50080
rect 8096 50016 8112 50080
rect 8176 50016 8192 50080
rect 8256 50016 8262 50080
rect 7946 50015 8262 50016
rect 17946 50080 18262 50081
rect 17946 50016 17952 50080
rect 18016 50016 18032 50080
rect 18096 50016 18112 50080
rect 18176 50016 18192 50080
rect 18256 50016 18262 50080
rect 17946 50015 18262 50016
rect 25313 49738 25379 49741
rect 26200 49738 27000 49768
rect 25313 49736 27000 49738
rect 25313 49680 25318 49736
rect 25374 49680 27000 49736
rect 25313 49678 27000 49680
rect 25313 49675 25379 49678
rect 26200 49648 27000 49678
rect 2946 49536 3262 49537
rect 2946 49472 2952 49536
rect 3016 49472 3032 49536
rect 3096 49472 3112 49536
rect 3176 49472 3192 49536
rect 3256 49472 3262 49536
rect 2946 49471 3262 49472
rect 12946 49536 13262 49537
rect 12946 49472 12952 49536
rect 13016 49472 13032 49536
rect 13096 49472 13112 49536
rect 13176 49472 13192 49536
rect 13256 49472 13262 49536
rect 12946 49471 13262 49472
rect 22946 49536 23262 49537
rect 22946 49472 22952 49536
rect 23016 49472 23032 49536
rect 23096 49472 23112 49536
rect 23176 49472 23192 49536
rect 23256 49472 23262 49536
rect 22946 49471 23262 49472
rect 7946 48992 8262 48993
rect 7946 48928 7952 48992
rect 8016 48928 8032 48992
rect 8096 48928 8112 48992
rect 8176 48928 8192 48992
rect 8256 48928 8262 48992
rect 7946 48927 8262 48928
rect 17946 48992 18262 48993
rect 17946 48928 17952 48992
rect 18016 48928 18032 48992
rect 18096 48928 18112 48992
rect 18176 48928 18192 48992
rect 18256 48928 18262 48992
rect 17946 48927 18262 48928
rect 25313 48922 25379 48925
rect 26200 48922 27000 48952
rect 25313 48920 27000 48922
rect 25313 48864 25318 48920
rect 25374 48864 27000 48920
rect 25313 48862 27000 48864
rect 25313 48859 25379 48862
rect 26200 48832 27000 48862
rect 2946 48448 3262 48449
rect 2946 48384 2952 48448
rect 3016 48384 3032 48448
rect 3096 48384 3112 48448
rect 3176 48384 3192 48448
rect 3256 48384 3262 48448
rect 2946 48383 3262 48384
rect 12946 48448 13262 48449
rect 12946 48384 12952 48448
rect 13016 48384 13032 48448
rect 13096 48384 13112 48448
rect 13176 48384 13192 48448
rect 13256 48384 13262 48448
rect 12946 48383 13262 48384
rect 22946 48448 23262 48449
rect 22946 48384 22952 48448
rect 23016 48384 23032 48448
rect 23096 48384 23112 48448
rect 23176 48384 23192 48448
rect 23256 48384 23262 48448
rect 22946 48383 23262 48384
rect 0 48106 800 48136
rect 4061 48106 4127 48109
rect 0 48104 4127 48106
rect 0 48048 4066 48104
rect 4122 48048 4127 48104
rect 0 48046 4127 48048
rect 0 48016 800 48046
rect 4061 48043 4127 48046
rect 24485 48106 24551 48109
rect 26200 48106 27000 48136
rect 24485 48104 27000 48106
rect 24485 48048 24490 48104
rect 24546 48048 27000 48104
rect 24485 48046 27000 48048
rect 24485 48043 24551 48046
rect 26200 48016 27000 48046
rect 7946 47904 8262 47905
rect 7946 47840 7952 47904
rect 8016 47840 8032 47904
rect 8096 47840 8112 47904
rect 8176 47840 8192 47904
rect 8256 47840 8262 47904
rect 7946 47839 8262 47840
rect 17946 47904 18262 47905
rect 17946 47840 17952 47904
rect 18016 47840 18032 47904
rect 18096 47840 18112 47904
rect 18176 47840 18192 47904
rect 18256 47840 18262 47904
rect 17946 47839 18262 47840
rect 2946 47360 3262 47361
rect 2946 47296 2952 47360
rect 3016 47296 3032 47360
rect 3096 47296 3112 47360
rect 3176 47296 3192 47360
rect 3256 47296 3262 47360
rect 2946 47295 3262 47296
rect 12946 47360 13262 47361
rect 12946 47296 12952 47360
rect 13016 47296 13032 47360
rect 13096 47296 13112 47360
rect 13176 47296 13192 47360
rect 13256 47296 13262 47360
rect 12946 47295 13262 47296
rect 22946 47360 23262 47361
rect 22946 47296 22952 47360
rect 23016 47296 23032 47360
rect 23096 47296 23112 47360
rect 23176 47296 23192 47360
rect 23256 47296 23262 47360
rect 22946 47295 23262 47296
rect 25497 47290 25563 47293
rect 26200 47290 27000 47320
rect 25497 47288 27000 47290
rect 25497 47232 25502 47288
rect 25558 47232 27000 47288
rect 25497 47230 27000 47232
rect 25497 47227 25563 47230
rect 26200 47200 27000 47230
rect 18505 47018 18571 47021
rect 19190 47018 19196 47020
rect 18505 47016 19196 47018
rect 18505 46960 18510 47016
rect 18566 46960 19196 47016
rect 18505 46958 19196 46960
rect 18505 46955 18571 46958
rect 19190 46956 19196 46958
rect 19260 46956 19266 47020
rect 7946 46816 8262 46817
rect 7946 46752 7952 46816
rect 8016 46752 8032 46816
rect 8096 46752 8112 46816
rect 8176 46752 8192 46816
rect 8256 46752 8262 46816
rect 7946 46751 8262 46752
rect 17946 46816 18262 46817
rect 17946 46752 17952 46816
rect 18016 46752 18032 46816
rect 18096 46752 18112 46816
rect 18176 46752 18192 46816
rect 18256 46752 18262 46816
rect 17946 46751 18262 46752
rect 20110 46684 20116 46748
rect 20180 46746 20186 46748
rect 20621 46746 20687 46749
rect 20180 46744 20687 46746
rect 20180 46688 20626 46744
rect 20682 46688 20687 46744
rect 20180 46686 20687 46688
rect 20180 46684 20186 46686
rect 20621 46683 20687 46686
rect 19609 46610 19675 46613
rect 19926 46610 19932 46612
rect 19609 46608 19932 46610
rect 19609 46552 19614 46608
rect 19670 46552 19932 46608
rect 19609 46550 19932 46552
rect 19609 46547 19675 46550
rect 19926 46548 19932 46550
rect 19996 46548 20002 46612
rect 24761 46610 24827 46613
rect 24761 46608 24962 46610
rect 24761 46552 24766 46608
rect 24822 46552 24962 46608
rect 24761 46550 24962 46552
rect 24761 46547 24827 46550
rect 24902 46474 24962 46550
rect 26200 46474 27000 46504
rect 24902 46414 27000 46474
rect 26200 46384 27000 46414
rect 2946 46272 3262 46273
rect 2946 46208 2952 46272
rect 3016 46208 3032 46272
rect 3096 46208 3112 46272
rect 3176 46208 3192 46272
rect 3256 46208 3262 46272
rect 2946 46207 3262 46208
rect 12946 46272 13262 46273
rect 12946 46208 12952 46272
rect 13016 46208 13032 46272
rect 13096 46208 13112 46272
rect 13176 46208 13192 46272
rect 13256 46208 13262 46272
rect 12946 46207 13262 46208
rect 22946 46272 23262 46273
rect 22946 46208 22952 46272
rect 23016 46208 23032 46272
rect 23096 46208 23112 46272
rect 23176 46208 23192 46272
rect 23256 46208 23262 46272
rect 22946 46207 23262 46208
rect 22001 45932 22067 45933
rect 21950 45930 21956 45932
rect 21910 45870 21956 45930
rect 22020 45928 22067 45932
rect 22062 45872 22067 45928
rect 21950 45868 21956 45870
rect 22020 45868 22067 45872
rect 22001 45867 22067 45868
rect 24393 45794 24459 45797
rect 24393 45792 24962 45794
rect 24393 45736 24398 45792
rect 24454 45736 24962 45792
rect 24393 45734 24962 45736
rect 24393 45731 24459 45734
rect 7946 45728 8262 45729
rect 0 45658 800 45688
rect 7946 45664 7952 45728
rect 8016 45664 8032 45728
rect 8096 45664 8112 45728
rect 8176 45664 8192 45728
rect 8256 45664 8262 45728
rect 7946 45663 8262 45664
rect 17946 45728 18262 45729
rect 17946 45664 17952 45728
rect 18016 45664 18032 45728
rect 18096 45664 18112 45728
rect 18176 45664 18192 45728
rect 18256 45664 18262 45728
rect 17946 45663 18262 45664
rect 4061 45658 4127 45661
rect 24761 45660 24827 45661
rect 24710 45658 24716 45660
rect 0 45656 4127 45658
rect 0 45600 4066 45656
rect 4122 45600 4127 45656
rect 0 45598 4127 45600
rect 24670 45598 24716 45658
rect 24780 45656 24827 45660
rect 24822 45600 24827 45656
rect 0 45568 800 45598
rect 4061 45595 4127 45598
rect 24710 45596 24716 45598
rect 24780 45596 24827 45600
rect 24902 45658 24962 45734
rect 26200 45658 27000 45688
rect 24902 45598 27000 45658
rect 24761 45595 24827 45596
rect 26200 45568 27000 45598
rect 11278 45324 11284 45388
rect 11348 45386 11354 45388
rect 11789 45386 11855 45389
rect 11348 45384 11855 45386
rect 11348 45328 11794 45384
rect 11850 45328 11855 45384
rect 11348 45326 11855 45328
rect 11348 45324 11354 45326
rect 11789 45323 11855 45326
rect 2946 45184 3262 45185
rect 2946 45120 2952 45184
rect 3016 45120 3032 45184
rect 3096 45120 3112 45184
rect 3176 45120 3192 45184
rect 3256 45120 3262 45184
rect 2946 45119 3262 45120
rect 12946 45184 13262 45185
rect 12946 45120 12952 45184
rect 13016 45120 13032 45184
rect 13096 45120 13112 45184
rect 13176 45120 13192 45184
rect 13256 45120 13262 45184
rect 12946 45119 13262 45120
rect 22946 45184 23262 45185
rect 22946 45120 22952 45184
rect 23016 45120 23032 45184
rect 23096 45120 23112 45184
rect 23176 45120 23192 45184
rect 23256 45120 23262 45184
rect 22946 45119 23262 45120
rect 24577 44842 24643 44845
rect 26200 44842 27000 44872
rect 24577 44840 27000 44842
rect 24577 44784 24582 44840
rect 24638 44784 27000 44840
rect 24577 44782 27000 44784
rect 24577 44779 24643 44782
rect 26200 44752 27000 44782
rect 9765 44708 9831 44709
rect 9765 44706 9812 44708
rect 9720 44704 9812 44706
rect 9720 44648 9770 44704
rect 9720 44646 9812 44648
rect 9765 44644 9812 44646
rect 9876 44644 9882 44708
rect 11462 44644 11468 44708
rect 11532 44706 11538 44708
rect 11605 44706 11671 44709
rect 11532 44704 11671 44706
rect 11532 44648 11610 44704
rect 11666 44648 11671 44704
rect 11532 44646 11671 44648
rect 11532 44644 11538 44646
rect 9765 44643 9831 44644
rect 11605 44643 11671 44646
rect 18454 44644 18460 44708
rect 18524 44706 18530 44708
rect 19333 44706 19399 44709
rect 18524 44704 19399 44706
rect 18524 44648 19338 44704
rect 19394 44648 19399 44704
rect 18524 44646 19399 44648
rect 18524 44644 18530 44646
rect 19333 44643 19399 44646
rect 7946 44640 8262 44641
rect 7946 44576 7952 44640
rect 8016 44576 8032 44640
rect 8096 44576 8112 44640
rect 8176 44576 8192 44640
rect 8256 44576 8262 44640
rect 7946 44575 8262 44576
rect 17946 44640 18262 44641
rect 17946 44576 17952 44640
rect 18016 44576 18032 44640
rect 18096 44576 18112 44640
rect 18176 44576 18192 44640
rect 18256 44576 18262 44640
rect 17946 44575 18262 44576
rect 10225 44298 10291 44301
rect 11605 44300 11671 44301
rect 10358 44298 10364 44300
rect 10225 44296 10364 44298
rect 10225 44240 10230 44296
rect 10286 44240 10364 44296
rect 10225 44238 10364 44240
rect 10225 44235 10291 44238
rect 10358 44236 10364 44238
rect 10428 44236 10434 44300
rect 11605 44298 11652 44300
rect 11560 44296 11652 44298
rect 11560 44240 11610 44296
rect 11560 44238 11652 44240
rect 11605 44236 11652 44238
rect 11716 44236 11722 44300
rect 24526 44236 24532 44300
rect 24596 44298 24602 44300
rect 24761 44298 24827 44301
rect 24596 44296 24827 44298
rect 24596 44240 24766 44296
rect 24822 44240 24827 44296
rect 24596 44238 24827 44240
rect 24596 44236 24602 44238
rect 11605 44235 11671 44236
rect 24761 44235 24827 44238
rect 2946 44096 3262 44097
rect 2946 44032 2952 44096
rect 3016 44032 3032 44096
rect 3096 44032 3112 44096
rect 3176 44032 3192 44096
rect 3256 44032 3262 44096
rect 2946 44031 3262 44032
rect 12946 44096 13262 44097
rect 12946 44032 12952 44096
rect 13016 44032 13032 44096
rect 13096 44032 13112 44096
rect 13176 44032 13192 44096
rect 13256 44032 13262 44096
rect 12946 44031 13262 44032
rect 22946 44096 23262 44097
rect 22946 44032 22952 44096
rect 23016 44032 23032 44096
rect 23096 44032 23112 44096
rect 23176 44032 23192 44096
rect 23256 44032 23262 44096
rect 22946 44031 23262 44032
rect 24485 44026 24551 44029
rect 26200 44026 27000 44056
rect 24485 44024 27000 44026
rect 24485 43968 24490 44024
rect 24546 43968 27000 44024
rect 24485 43966 27000 43968
rect 24485 43963 24551 43966
rect 26200 43936 27000 43966
rect 7946 43552 8262 43553
rect 7946 43488 7952 43552
rect 8016 43488 8032 43552
rect 8096 43488 8112 43552
rect 8176 43488 8192 43552
rect 8256 43488 8262 43552
rect 7946 43487 8262 43488
rect 17946 43552 18262 43553
rect 17946 43488 17952 43552
rect 18016 43488 18032 43552
rect 18096 43488 18112 43552
rect 18176 43488 18192 43552
rect 18256 43488 18262 43552
rect 17946 43487 18262 43488
rect 0 43210 800 43240
rect 1301 43210 1367 43213
rect 0 43208 1367 43210
rect 0 43152 1306 43208
rect 1362 43152 1367 43208
rect 0 43150 1367 43152
rect 0 43120 800 43150
rect 1301 43147 1367 43150
rect 17350 43148 17356 43212
rect 17420 43210 17426 43212
rect 21081 43210 21147 43213
rect 21909 43210 21975 43213
rect 17420 43208 21975 43210
rect 17420 43152 21086 43208
rect 21142 43152 21914 43208
rect 21970 43152 21975 43208
rect 17420 43150 21975 43152
rect 17420 43148 17426 43150
rect 21081 43147 21147 43150
rect 21909 43147 21975 43150
rect 24577 43210 24643 43213
rect 26200 43210 27000 43240
rect 24577 43208 27000 43210
rect 24577 43152 24582 43208
rect 24638 43152 27000 43208
rect 24577 43150 27000 43152
rect 24577 43147 24643 43150
rect 26200 43120 27000 43150
rect 2946 43008 3262 43009
rect 2946 42944 2952 43008
rect 3016 42944 3032 43008
rect 3096 42944 3112 43008
rect 3176 42944 3192 43008
rect 3256 42944 3262 43008
rect 2946 42943 3262 42944
rect 12946 43008 13262 43009
rect 12946 42944 12952 43008
rect 13016 42944 13032 43008
rect 13096 42944 13112 43008
rect 13176 42944 13192 43008
rect 13256 42944 13262 43008
rect 12946 42943 13262 42944
rect 22946 43008 23262 43009
rect 22946 42944 22952 43008
rect 23016 42944 23032 43008
rect 23096 42944 23112 43008
rect 23176 42944 23192 43008
rect 23256 42944 23262 43008
rect 22946 42943 23262 42944
rect 22001 42802 22067 42805
rect 24853 42802 24919 42805
rect 22001 42800 24919 42802
rect 22001 42744 22006 42800
rect 22062 42744 24858 42800
rect 24914 42744 24919 42800
rect 22001 42742 24919 42744
rect 22001 42739 22067 42742
rect 24853 42739 24919 42742
rect 22185 42666 22251 42669
rect 22142 42664 22251 42666
rect 22142 42608 22190 42664
rect 22246 42608 22251 42664
rect 22142 42603 22251 42608
rect 7946 42464 8262 42465
rect 7946 42400 7952 42464
rect 8016 42400 8032 42464
rect 8096 42400 8112 42464
rect 8176 42400 8192 42464
rect 8256 42400 8262 42464
rect 7946 42399 8262 42400
rect 17946 42464 18262 42465
rect 17946 42400 17952 42464
rect 18016 42400 18032 42464
rect 18096 42400 18112 42464
rect 18176 42400 18192 42464
rect 18256 42400 18262 42464
rect 17946 42399 18262 42400
rect 22142 42394 22202 42603
rect 22277 42394 22343 42397
rect 22142 42392 22343 42394
rect 22142 42336 22282 42392
rect 22338 42336 22343 42392
rect 22142 42334 22343 42336
rect 22277 42331 22343 42334
rect 23197 42394 23263 42397
rect 26200 42394 27000 42424
rect 23197 42392 27000 42394
rect 23197 42336 23202 42392
rect 23258 42336 27000 42392
rect 23197 42334 27000 42336
rect 23197 42331 23263 42334
rect 26200 42304 27000 42334
rect 20529 42122 20595 42125
rect 23013 42122 23079 42125
rect 20529 42120 23079 42122
rect 20529 42064 20534 42120
rect 20590 42064 23018 42120
rect 23074 42064 23079 42120
rect 20529 42062 23079 42064
rect 20529 42059 20595 42062
rect 23013 42059 23079 42062
rect 2946 41920 3262 41921
rect 2946 41856 2952 41920
rect 3016 41856 3032 41920
rect 3096 41856 3112 41920
rect 3176 41856 3192 41920
rect 3256 41856 3262 41920
rect 2946 41855 3262 41856
rect 12946 41920 13262 41921
rect 12946 41856 12952 41920
rect 13016 41856 13032 41920
rect 13096 41856 13112 41920
rect 13176 41856 13192 41920
rect 13256 41856 13262 41920
rect 12946 41855 13262 41856
rect 22946 41920 23262 41921
rect 22946 41856 22952 41920
rect 23016 41856 23032 41920
rect 23096 41856 23112 41920
rect 23176 41856 23192 41920
rect 23256 41856 23262 41920
rect 22946 41855 23262 41856
rect 22093 41578 22159 41581
rect 26200 41578 27000 41608
rect 22093 41576 27000 41578
rect 22093 41520 22098 41576
rect 22154 41520 27000 41576
rect 22093 41518 27000 41520
rect 22093 41515 22159 41518
rect 26200 41488 27000 41518
rect 22686 41442 22692 41444
rect 22142 41382 22692 41442
rect 7946 41376 8262 41377
rect 7946 41312 7952 41376
rect 8016 41312 8032 41376
rect 8096 41312 8112 41376
rect 8176 41312 8192 41376
rect 8256 41312 8262 41376
rect 7946 41311 8262 41312
rect 17946 41376 18262 41377
rect 17946 41312 17952 41376
rect 18016 41312 18032 41376
rect 18096 41312 18112 41376
rect 18176 41312 18192 41376
rect 18256 41312 18262 41376
rect 17946 41311 18262 41312
rect 22142 41309 22202 41382
rect 22686 41380 22692 41382
rect 22756 41442 22762 41444
rect 24393 41442 24459 41445
rect 22756 41440 24459 41442
rect 22756 41384 24398 41440
rect 24454 41384 24459 41440
rect 22756 41382 24459 41384
rect 22756 41380 22762 41382
rect 24393 41379 24459 41382
rect 22093 41304 22202 41309
rect 22093 41248 22098 41304
rect 22154 41248 22202 41304
rect 22093 41246 22202 41248
rect 22093 41243 22159 41246
rect 2946 40832 3262 40833
rect 0 40762 800 40792
rect 2946 40768 2952 40832
rect 3016 40768 3032 40832
rect 3096 40768 3112 40832
rect 3176 40768 3192 40832
rect 3256 40768 3262 40832
rect 2946 40767 3262 40768
rect 12946 40832 13262 40833
rect 12946 40768 12952 40832
rect 13016 40768 13032 40832
rect 13096 40768 13112 40832
rect 13176 40768 13192 40832
rect 13256 40768 13262 40832
rect 12946 40767 13262 40768
rect 22946 40832 23262 40833
rect 22946 40768 22952 40832
rect 23016 40768 23032 40832
rect 23096 40768 23112 40832
rect 23176 40768 23192 40832
rect 23256 40768 23262 40832
rect 22946 40767 23262 40768
rect 1301 40762 1367 40765
rect 0 40760 1367 40762
rect 0 40704 1306 40760
rect 1362 40704 1367 40760
rect 0 40702 1367 40704
rect 0 40672 800 40702
rect 1301 40699 1367 40702
rect 24761 40762 24827 40765
rect 26200 40762 27000 40792
rect 24761 40760 27000 40762
rect 24761 40704 24766 40760
rect 24822 40704 27000 40760
rect 24761 40702 27000 40704
rect 24761 40699 24827 40702
rect 26200 40672 27000 40702
rect 16573 40626 16639 40629
rect 17718 40626 17724 40628
rect 16573 40624 17724 40626
rect 16573 40568 16578 40624
rect 16634 40568 17724 40624
rect 16573 40566 17724 40568
rect 16573 40563 16639 40566
rect 17718 40564 17724 40566
rect 17788 40564 17794 40628
rect 16941 40490 17007 40493
rect 20161 40490 20227 40493
rect 16941 40488 20227 40490
rect 16941 40432 16946 40488
rect 17002 40432 20166 40488
rect 20222 40432 20227 40488
rect 16941 40430 20227 40432
rect 16941 40427 17007 40430
rect 20161 40427 20227 40430
rect 7946 40288 8262 40289
rect 7946 40224 7952 40288
rect 8016 40224 8032 40288
rect 8096 40224 8112 40288
rect 8176 40224 8192 40288
rect 8256 40224 8262 40288
rect 7946 40223 8262 40224
rect 17946 40288 18262 40289
rect 17946 40224 17952 40288
rect 18016 40224 18032 40288
rect 18096 40224 18112 40288
rect 18176 40224 18192 40288
rect 18256 40224 18262 40288
rect 17946 40223 18262 40224
rect 22093 40218 22159 40221
rect 22502 40218 22508 40220
rect 22093 40216 22508 40218
rect 22093 40160 22098 40216
rect 22154 40160 22508 40216
rect 22093 40158 22508 40160
rect 22093 40155 22159 40158
rect 22502 40156 22508 40158
rect 22572 40156 22578 40220
rect 18229 40082 18295 40085
rect 22134 40082 22140 40084
rect 18229 40080 22140 40082
rect 18229 40024 18234 40080
rect 18290 40024 22140 40080
rect 18229 40022 22140 40024
rect 18229 40019 18295 40022
rect 22134 40020 22140 40022
rect 22204 40020 22210 40084
rect 22318 40020 22324 40084
rect 22388 40082 22394 40084
rect 23422 40082 23428 40084
rect 22388 40022 23428 40082
rect 22388 40020 22394 40022
rect 23422 40020 23428 40022
rect 23492 40020 23498 40084
rect 24117 40082 24183 40085
rect 24117 40080 24226 40082
rect 24117 40024 24122 40080
rect 24178 40024 24226 40080
rect 24117 40019 24226 40024
rect 24166 39946 24226 40019
rect 26200 39946 27000 39976
rect 24166 39886 27000 39946
rect 26200 39856 27000 39886
rect 2946 39744 3262 39745
rect 2946 39680 2952 39744
rect 3016 39680 3032 39744
rect 3096 39680 3112 39744
rect 3176 39680 3192 39744
rect 3256 39680 3262 39744
rect 2946 39679 3262 39680
rect 12946 39744 13262 39745
rect 12946 39680 12952 39744
rect 13016 39680 13032 39744
rect 13096 39680 13112 39744
rect 13176 39680 13192 39744
rect 13256 39680 13262 39744
rect 12946 39679 13262 39680
rect 22946 39744 23262 39745
rect 22946 39680 22952 39744
rect 23016 39680 23032 39744
rect 23096 39680 23112 39744
rect 23176 39680 23192 39744
rect 23256 39680 23262 39744
rect 22946 39679 23262 39680
rect 7946 39200 8262 39201
rect 7946 39136 7952 39200
rect 8016 39136 8032 39200
rect 8096 39136 8112 39200
rect 8176 39136 8192 39200
rect 8256 39136 8262 39200
rect 7946 39135 8262 39136
rect 17946 39200 18262 39201
rect 17946 39136 17952 39200
rect 18016 39136 18032 39200
rect 18096 39136 18112 39200
rect 18176 39136 18192 39200
rect 18256 39136 18262 39200
rect 17946 39135 18262 39136
rect 24025 39130 24091 39133
rect 26200 39130 27000 39160
rect 24025 39128 27000 39130
rect 24025 39072 24030 39128
rect 24086 39072 27000 39128
rect 24025 39070 27000 39072
rect 24025 39067 24091 39070
rect 26200 39040 27000 39070
rect 15929 38722 15995 38725
rect 16062 38722 16068 38724
rect 15929 38720 16068 38722
rect 15929 38664 15934 38720
rect 15990 38664 16068 38720
rect 15929 38662 16068 38664
rect 15929 38659 15995 38662
rect 16062 38660 16068 38662
rect 16132 38660 16138 38724
rect 2946 38656 3262 38657
rect 2946 38592 2952 38656
rect 3016 38592 3032 38656
rect 3096 38592 3112 38656
rect 3176 38592 3192 38656
rect 3256 38592 3262 38656
rect 2946 38591 3262 38592
rect 12946 38656 13262 38657
rect 12946 38592 12952 38656
rect 13016 38592 13032 38656
rect 13096 38592 13112 38656
rect 13176 38592 13192 38656
rect 13256 38592 13262 38656
rect 12946 38591 13262 38592
rect 22946 38656 23262 38657
rect 22946 38592 22952 38656
rect 23016 38592 23032 38656
rect 23096 38592 23112 38656
rect 23176 38592 23192 38656
rect 23256 38592 23262 38656
rect 22946 38591 23262 38592
rect 15101 38450 15167 38453
rect 21582 38450 21588 38452
rect 15101 38448 21588 38450
rect 15101 38392 15106 38448
rect 15162 38392 21588 38448
rect 15101 38390 21588 38392
rect 15101 38387 15167 38390
rect 21582 38388 21588 38390
rect 21652 38450 21658 38452
rect 24301 38450 24367 38453
rect 21652 38448 24367 38450
rect 21652 38392 24306 38448
rect 24362 38392 24367 38448
rect 21652 38390 24367 38392
rect 21652 38388 21658 38390
rect 24301 38387 24367 38390
rect 0 38314 800 38344
rect 1301 38314 1367 38317
rect 12617 38316 12683 38317
rect 0 38312 1367 38314
rect 0 38256 1306 38312
rect 1362 38256 1367 38312
rect 0 38254 1367 38256
rect 0 38224 800 38254
rect 1301 38251 1367 38254
rect 12566 38252 12572 38316
rect 12636 38314 12683 38316
rect 25313 38314 25379 38317
rect 26200 38314 27000 38344
rect 12636 38312 12728 38314
rect 12678 38256 12728 38312
rect 12636 38254 12728 38256
rect 25313 38312 27000 38314
rect 25313 38256 25318 38312
rect 25374 38256 27000 38312
rect 25313 38254 27000 38256
rect 12636 38252 12683 38254
rect 12617 38251 12683 38252
rect 25313 38251 25379 38254
rect 26200 38224 27000 38254
rect 7946 38112 8262 38113
rect 7946 38048 7952 38112
rect 8016 38048 8032 38112
rect 8096 38048 8112 38112
rect 8176 38048 8192 38112
rect 8256 38048 8262 38112
rect 7946 38047 8262 38048
rect 17946 38112 18262 38113
rect 17946 38048 17952 38112
rect 18016 38048 18032 38112
rect 18096 38048 18112 38112
rect 18176 38048 18192 38112
rect 18256 38048 18262 38112
rect 17946 38047 18262 38048
rect 22645 38044 22711 38045
rect 22645 38040 22692 38044
rect 22756 38042 22762 38044
rect 22645 37984 22650 38040
rect 22645 37980 22692 37984
rect 22756 37982 22802 38042
rect 22756 37980 22762 37982
rect 22645 37979 22711 37980
rect 16849 37770 16915 37773
rect 22093 37770 22159 37773
rect 16849 37768 22159 37770
rect 16849 37712 16854 37768
rect 16910 37712 22098 37768
rect 22154 37712 22159 37768
rect 16849 37710 22159 37712
rect 16849 37707 16915 37710
rect 22093 37707 22159 37710
rect 17125 37634 17191 37637
rect 19241 37634 19307 37637
rect 17125 37632 19307 37634
rect 17125 37576 17130 37632
rect 17186 37576 19246 37632
rect 19302 37576 19307 37632
rect 17125 37574 19307 37576
rect 17125 37571 17191 37574
rect 19241 37571 19307 37574
rect 2946 37568 3262 37569
rect 2946 37504 2952 37568
rect 3016 37504 3032 37568
rect 3096 37504 3112 37568
rect 3176 37504 3192 37568
rect 3256 37504 3262 37568
rect 2946 37503 3262 37504
rect 12946 37568 13262 37569
rect 12946 37504 12952 37568
rect 13016 37504 13032 37568
rect 13096 37504 13112 37568
rect 13176 37504 13192 37568
rect 13256 37504 13262 37568
rect 12946 37503 13262 37504
rect 22946 37568 23262 37569
rect 22946 37504 22952 37568
rect 23016 37504 23032 37568
rect 23096 37504 23112 37568
rect 23176 37504 23192 37568
rect 23256 37504 23262 37568
rect 22946 37503 23262 37504
rect 18965 37498 19031 37501
rect 23381 37498 23447 37501
rect 26200 37498 27000 37528
rect 18965 37496 19074 37498
rect 18965 37440 18970 37496
rect 19026 37440 19074 37496
rect 18965 37435 19074 37440
rect 23381 37496 27000 37498
rect 23381 37440 23386 37496
rect 23442 37440 27000 37496
rect 23381 37438 27000 37440
rect 23381 37435 23447 37438
rect 19014 37365 19074 37435
rect 26200 37408 27000 37438
rect 10593 37362 10659 37365
rect 13353 37362 13419 37365
rect 10593 37360 13419 37362
rect 10593 37304 10598 37360
rect 10654 37304 13358 37360
rect 13414 37304 13419 37360
rect 10593 37302 13419 37304
rect 19014 37360 19123 37365
rect 19333 37364 19399 37365
rect 19333 37362 19380 37364
rect 19014 37304 19062 37360
rect 19118 37304 19123 37360
rect 19014 37302 19123 37304
rect 19288 37360 19380 37362
rect 19288 37304 19338 37360
rect 19288 37302 19380 37304
rect 10593 37299 10659 37302
rect 13353 37299 13419 37302
rect 19057 37299 19123 37302
rect 19333 37300 19380 37302
rect 19444 37300 19450 37364
rect 19333 37299 19399 37300
rect 7946 37024 8262 37025
rect 7946 36960 7952 37024
rect 8016 36960 8032 37024
rect 8096 36960 8112 37024
rect 8176 36960 8192 37024
rect 8256 36960 8262 37024
rect 7946 36959 8262 36960
rect 17946 37024 18262 37025
rect 17946 36960 17952 37024
rect 18016 36960 18032 37024
rect 18096 36960 18112 37024
rect 18176 36960 18192 37024
rect 18256 36960 18262 37024
rect 17946 36959 18262 36960
rect 9806 36756 9812 36820
rect 9876 36818 9882 36820
rect 10133 36818 10199 36821
rect 16665 36818 16731 36821
rect 9876 36816 16731 36818
rect 9876 36760 10138 36816
rect 10194 36760 16670 36816
rect 16726 36760 16731 36816
rect 9876 36758 16731 36760
rect 9876 36756 9882 36758
rect 10133 36755 10199 36758
rect 16665 36755 16731 36758
rect 18321 36682 18387 36685
rect 19149 36682 19215 36685
rect 18321 36680 19215 36682
rect 18321 36624 18326 36680
rect 18382 36624 19154 36680
rect 19210 36624 19215 36680
rect 18321 36622 19215 36624
rect 18321 36619 18387 36622
rect 19149 36619 19215 36622
rect 24669 36682 24735 36685
rect 26200 36682 27000 36712
rect 24669 36680 27000 36682
rect 24669 36624 24674 36680
rect 24730 36624 27000 36680
rect 24669 36622 27000 36624
rect 24669 36619 24735 36622
rect 26200 36592 27000 36622
rect 21081 36548 21147 36549
rect 21030 36484 21036 36548
rect 21100 36546 21147 36548
rect 21100 36544 21192 36546
rect 21142 36488 21192 36544
rect 21100 36486 21192 36488
rect 21100 36484 21147 36486
rect 21081 36483 21147 36484
rect 2946 36480 3262 36481
rect 2946 36416 2952 36480
rect 3016 36416 3032 36480
rect 3096 36416 3112 36480
rect 3176 36416 3192 36480
rect 3256 36416 3262 36480
rect 2946 36415 3262 36416
rect 12946 36480 13262 36481
rect 12946 36416 12952 36480
rect 13016 36416 13032 36480
rect 13096 36416 13112 36480
rect 13176 36416 13192 36480
rect 13256 36416 13262 36480
rect 12946 36415 13262 36416
rect 22946 36480 23262 36481
rect 22946 36416 22952 36480
rect 23016 36416 23032 36480
rect 23096 36416 23112 36480
rect 23176 36416 23192 36480
rect 23256 36416 23262 36480
rect 22946 36415 23262 36416
rect 11237 36412 11303 36413
rect 11237 36410 11284 36412
rect 11192 36408 11284 36410
rect 11192 36352 11242 36408
rect 11192 36350 11284 36352
rect 11237 36348 11284 36350
rect 11348 36348 11354 36412
rect 20069 36410 20135 36413
rect 21449 36410 21515 36413
rect 20069 36408 21515 36410
rect 20069 36352 20074 36408
rect 20130 36352 21454 36408
rect 21510 36352 21515 36408
rect 20069 36350 21515 36352
rect 11237 36347 11303 36348
rect 20069 36347 20135 36350
rect 21449 36347 21515 36350
rect 19609 36138 19675 36141
rect 14782 36136 19675 36138
rect 14782 36080 19614 36136
rect 19670 36080 19675 36136
rect 14782 36078 19675 36080
rect 13813 36002 13879 36005
rect 14782 36004 14842 36078
rect 19609 36075 19675 36078
rect 14774 36002 14780 36004
rect 13813 36000 14780 36002
rect 13813 35944 13818 36000
rect 13874 35944 14780 36000
rect 13813 35942 14780 35944
rect 13813 35939 13879 35942
rect 14774 35940 14780 35942
rect 14844 35940 14850 36004
rect 7946 35936 8262 35937
rect 0 35866 800 35896
rect 7946 35872 7952 35936
rect 8016 35872 8032 35936
rect 8096 35872 8112 35936
rect 8176 35872 8192 35936
rect 8256 35872 8262 35936
rect 7946 35871 8262 35872
rect 17946 35936 18262 35937
rect 17946 35872 17952 35936
rect 18016 35872 18032 35936
rect 18096 35872 18112 35936
rect 18176 35872 18192 35936
rect 18256 35872 18262 35936
rect 17946 35871 18262 35872
rect 1761 35866 1827 35869
rect 0 35864 1827 35866
rect 0 35808 1766 35864
rect 1822 35808 1827 35864
rect 0 35806 1827 35808
rect 0 35776 800 35806
rect 1761 35803 1827 35806
rect 24853 35866 24919 35869
rect 26200 35866 27000 35896
rect 24853 35864 27000 35866
rect 24853 35808 24858 35864
rect 24914 35808 27000 35864
rect 24853 35806 27000 35808
rect 24853 35803 24919 35806
rect 26200 35776 27000 35806
rect 12525 35594 12591 35597
rect 12525 35592 13554 35594
rect 12525 35536 12530 35592
rect 12586 35536 13554 35592
rect 12525 35534 13554 35536
rect 12525 35531 12591 35534
rect 13494 35458 13554 35534
rect 13629 35458 13695 35461
rect 13494 35456 13695 35458
rect 13494 35400 13634 35456
rect 13690 35400 13695 35456
rect 13494 35398 13695 35400
rect 13629 35395 13695 35398
rect 2946 35392 3262 35393
rect 2946 35328 2952 35392
rect 3016 35328 3032 35392
rect 3096 35328 3112 35392
rect 3176 35328 3192 35392
rect 3256 35328 3262 35392
rect 2946 35327 3262 35328
rect 12946 35392 13262 35393
rect 12946 35328 12952 35392
rect 13016 35328 13032 35392
rect 13096 35328 13112 35392
rect 13176 35328 13192 35392
rect 13256 35328 13262 35392
rect 12946 35327 13262 35328
rect 22946 35392 23262 35393
rect 22946 35328 22952 35392
rect 23016 35328 23032 35392
rect 23096 35328 23112 35392
rect 23176 35328 23192 35392
rect 23256 35328 23262 35392
rect 22946 35327 23262 35328
rect 22001 35186 22067 35189
rect 23197 35186 23263 35189
rect 24526 35186 24532 35188
rect 22001 35184 24532 35186
rect 22001 35128 22006 35184
rect 22062 35128 23202 35184
rect 23258 35128 24532 35184
rect 22001 35126 24532 35128
rect 22001 35123 22067 35126
rect 23197 35123 23263 35126
rect 24526 35124 24532 35126
rect 24596 35124 24602 35188
rect 22369 35050 22435 35053
rect 22645 35050 22711 35053
rect 22369 35048 22711 35050
rect 22369 34992 22374 35048
rect 22430 34992 22650 35048
rect 22706 34992 22711 35048
rect 22369 34990 22711 34992
rect 22369 34987 22435 34990
rect 22645 34987 22711 34990
rect 24669 35050 24735 35053
rect 26200 35050 27000 35080
rect 24669 35048 27000 35050
rect 24669 34992 24674 35048
rect 24730 34992 27000 35048
rect 24669 34990 27000 34992
rect 24669 34987 24735 34990
rect 26200 34960 27000 34990
rect 7946 34848 8262 34849
rect 7946 34784 7952 34848
rect 8016 34784 8032 34848
rect 8096 34784 8112 34848
rect 8176 34784 8192 34848
rect 8256 34784 8262 34848
rect 7946 34783 8262 34784
rect 17946 34848 18262 34849
rect 17946 34784 17952 34848
rect 18016 34784 18032 34848
rect 18096 34784 18112 34848
rect 18176 34784 18192 34848
rect 18256 34784 18262 34848
rect 17946 34783 18262 34784
rect 22737 34370 22803 34373
rect 22694 34368 22803 34370
rect 22694 34312 22742 34368
rect 22798 34312 22803 34368
rect 22694 34307 22803 34312
rect 2946 34304 3262 34305
rect 2946 34240 2952 34304
rect 3016 34240 3032 34304
rect 3096 34240 3112 34304
rect 3176 34240 3192 34304
rect 3256 34240 3262 34304
rect 2946 34239 3262 34240
rect 12946 34304 13262 34305
rect 12946 34240 12952 34304
rect 13016 34240 13032 34304
rect 13096 34240 13112 34304
rect 13176 34240 13192 34304
rect 13256 34240 13262 34304
rect 12946 34239 13262 34240
rect 22694 34098 22754 34307
rect 22946 34304 23262 34305
rect 22946 34240 22952 34304
rect 23016 34240 23032 34304
rect 23096 34240 23112 34304
rect 23176 34240 23192 34304
rect 23256 34240 23262 34304
rect 22946 34239 23262 34240
rect 25313 34234 25379 34237
rect 26200 34234 27000 34264
rect 25313 34232 27000 34234
rect 25313 34176 25318 34232
rect 25374 34176 27000 34232
rect 25313 34174 27000 34176
rect 25313 34171 25379 34174
rect 26200 34144 27000 34174
rect 22921 34098 22987 34101
rect 22694 34096 22987 34098
rect 22694 34040 22926 34096
rect 22982 34040 22987 34096
rect 22694 34038 22987 34040
rect 22921 34035 22987 34038
rect 7946 33760 8262 33761
rect 7946 33696 7952 33760
rect 8016 33696 8032 33760
rect 8096 33696 8112 33760
rect 8176 33696 8192 33760
rect 8256 33696 8262 33760
rect 7946 33695 8262 33696
rect 17946 33760 18262 33761
rect 17946 33696 17952 33760
rect 18016 33696 18032 33760
rect 18096 33696 18112 33760
rect 18176 33696 18192 33760
rect 18256 33696 18262 33760
rect 17946 33695 18262 33696
rect 19793 33554 19859 33557
rect 23565 33554 23631 33557
rect 19793 33552 23631 33554
rect 19793 33496 19798 33552
rect 19854 33496 23570 33552
rect 23626 33496 23631 33552
rect 19793 33494 23631 33496
rect 19793 33491 19859 33494
rect 23565 33491 23631 33494
rect 0 33418 800 33448
rect 1301 33418 1367 33421
rect 0 33416 1367 33418
rect 0 33360 1306 33416
rect 1362 33360 1367 33416
rect 0 33358 1367 33360
rect 0 33328 800 33358
rect 1301 33355 1367 33358
rect 21265 33418 21331 33421
rect 24710 33418 24716 33420
rect 21265 33416 24716 33418
rect 21265 33360 21270 33416
rect 21326 33360 24716 33416
rect 21265 33358 24716 33360
rect 21265 33355 21331 33358
rect 24710 33356 24716 33358
rect 24780 33356 24786 33420
rect 25405 33418 25471 33421
rect 26200 33418 27000 33448
rect 25405 33416 27000 33418
rect 25405 33360 25410 33416
rect 25466 33360 27000 33416
rect 25405 33358 27000 33360
rect 25405 33355 25471 33358
rect 26200 33328 27000 33358
rect 12525 33284 12591 33285
rect 12525 33282 12572 33284
rect 12480 33280 12572 33282
rect 12480 33224 12530 33280
rect 12480 33222 12572 33224
rect 12525 33220 12572 33222
rect 12636 33220 12642 33284
rect 12525 33219 12591 33220
rect 2946 33216 3262 33217
rect 2946 33152 2952 33216
rect 3016 33152 3032 33216
rect 3096 33152 3112 33216
rect 3176 33152 3192 33216
rect 3256 33152 3262 33216
rect 2946 33151 3262 33152
rect 12946 33216 13262 33217
rect 12946 33152 12952 33216
rect 13016 33152 13032 33216
rect 13096 33152 13112 33216
rect 13176 33152 13192 33216
rect 13256 33152 13262 33216
rect 12946 33151 13262 33152
rect 22946 33216 23262 33217
rect 22946 33152 22952 33216
rect 23016 33152 23032 33216
rect 23096 33152 23112 33216
rect 23176 33152 23192 33216
rect 23256 33152 23262 33216
rect 22946 33151 23262 33152
rect 17677 33146 17743 33149
rect 22185 33148 22251 33149
rect 19190 33146 19196 33148
rect 17677 33144 19196 33146
rect 17677 33088 17682 33144
rect 17738 33088 19196 33144
rect 17677 33086 19196 33088
rect 17677 33083 17743 33086
rect 19190 33084 19196 33086
rect 19260 33084 19266 33148
rect 22134 33146 22140 33148
rect 22094 33086 22140 33146
rect 22204 33144 22251 33148
rect 22246 33088 22251 33144
rect 22134 33084 22140 33086
rect 22204 33084 22251 33088
rect 22185 33083 22251 33084
rect 11329 33010 11395 33013
rect 11462 33010 11468 33012
rect 11329 33008 11468 33010
rect 11329 32952 11334 33008
rect 11390 32952 11468 33008
rect 11329 32950 11468 32952
rect 11329 32947 11395 32950
rect 11462 32948 11468 32950
rect 11532 32948 11538 33012
rect 21725 33010 21791 33013
rect 23013 33010 23079 33013
rect 23422 33010 23428 33012
rect 21725 33008 23428 33010
rect 21725 32952 21730 33008
rect 21786 32952 23018 33008
rect 23074 32952 23428 33008
rect 21725 32950 23428 32952
rect 21725 32947 21791 32950
rect 23013 32947 23079 32950
rect 23422 32948 23428 32950
rect 23492 32948 23498 33012
rect 13854 32812 13860 32876
rect 13924 32874 13930 32876
rect 14825 32874 14891 32877
rect 13924 32872 14891 32874
rect 13924 32816 14830 32872
rect 14886 32816 14891 32872
rect 13924 32814 14891 32816
rect 13924 32812 13930 32814
rect 14825 32811 14891 32814
rect 7946 32672 8262 32673
rect 7946 32608 7952 32672
rect 8016 32608 8032 32672
rect 8096 32608 8112 32672
rect 8176 32608 8192 32672
rect 8256 32608 8262 32672
rect 7946 32607 8262 32608
rect 17946 32672 18262 32673
rect 17946 32608 17952 32672
rect 18016 32608 18032 32672
rect 18096 32608 18112 32672
rect 18176 32608 18192 32672
rect 18256 32608 18262 32672
rect 17946 32607 18262 32608
rect 11646 32540 11652 32604
rect 11716 32602 11722 32604
rect 13261 32602 13327 32605
rect 11716 32600 13327 32602
rect 11716 32544 13266 32600
rect 13322 32544 13327 32600
rect 11716 32542 13327 32544
rect 11716 32540 11722 32542
rect 13261 32539 13327 32542
rect 25313 32602 25379 32605
rect 26200 32602 27000 32632
rect 25313 32600 27000 32602
rect 25313 32544 25318 32600
rect 25374 32544 27000 32600
rect 25313 32542 27000 32544
rect 25313 32539 25379 32542
rect 26200 32512 27000 32542
rect 2946 32128 3262 32129
rect 2946 32064 2952 32128
rect 3016 32064 3032 32128
rect 3096 32064 3112 32128
rect 3176 32064 3192 32128
rect 3256 32064 3262 32128
rect 2946 32063 3262 32064
rect 12946 32128 13262 32129
rect 12946 32064 12952 32128
rect 13016 32064 13032 32128
rect 13096 32064 13112 32128
rect 13176 32064 13192 32128
rect 13256 32064 13262 32128
rect 12946 32063 13262 32064
rect 22946 32128 23262 32129
rect 22946 32064 22952 32128
rect 23016 32064 23032 32128
rect 23096 32064 23112 32128
rect 23176 32064 23192 32128
rect 23256 32064 23262 32128
rect 22946 32063 23262 32064
rect 21541 32060 21607 32061
rect 21541 32058 21588 32060
rect 21496 32056 21588 32058
rect 21496 32000 21546 32056
rect 21496 31998 21588 32000
rect 21541 31996 21588 31998
rect 21652 31996 21658 32060
rect 21541 31995 21607 31996
rect 18597 31922 18663 31925
rect 20110 31922 20116 31924
rect 18597 31920 20116 31922
rect 18597 31864 18602 31920
rect 18658 31864 20116 31920
rect 18597 31862 20116 31864
rect 18597 31859 18663 31862
rect 20110 31860 20116 31862
rect 20180 31860 20186 31924
rect 15745 31786 15811 31789
rect 21030 31786 21036 31788
rect 15745 31784 21036 31786
rect 15745 31728 15750 31784
rect 15806 31728 21036 31784
rect 15745 31726 21036 31728
rect 15745 31723 15811 31726
rect 21030 31724 21036 31726
rect 21100 31724 21106 31788
rect 25313 31786 25379 31789
rect 26200 31786 27000 31816
rect 25313 31784 27000 31786
rect 25313 31728 25318 31784
rect 25374 31728 27000 31784
rect 25313 31726 27000 31728
rect 25313 31723 25379 31726
rect 26200 31696 27000 31726
rect 7946 31584 8262 31585
rect 7946 31520 7952 31584
rect 8016 31520 8032 31584
rect 8096 31520 8112 31584
rect 8176 31520 8192 31584
rect 8256 31520 8262 31584
rect 7946 31519 8262 31520
rect 17946 31584 18262 31585
rect 17946 31520 17952 31584
rect 18016 31520 18032 31584
rect 18096 31520 18112 31584
rect 18176 31520 18192 31584
rect 18256 31520 18262 31584
rect 17946 31519 18262 31520
rect 2946 31040 3262 31041
rect 0 30970 800 31000
rect 2946 30976 2952 31040
rect 3016 30976 3032 31040
rect 3096 30976 3112 31040
rect 3176 30976 3192 31040
rect 3256 30976 3262 31040
rect 2946 30975 3262 30976
rect 12946 31040 13262 31041
rect 12946 30976 12952 31040
rect 13016 30976 13032 31040
rect 13096 30976 13112 31040
rect 13176 30976 13192 31040
rect 13256 30976 13262 31040
rect 12946 30975 13262 30976
rect 22946 31040 23262 31041
rect 22946 30976 22952 31040
rect 23016 30976 23032 31040
rect 23096 30976 23112 31040
rect 23176 30976 23192 31040
rect 23256 30976 23262 31040
rect 22946 30975 23262 30976
rect 2773 30970 2839 30973
rect 0 30968 2839 30970
rect 0 30912 2778 30968
rect 2834 30912 2839 30968
rect 0 30910 2839 30912
rect 0 30880 800 30910
rect 2773 30907 2839 30910
rect 25313 30970 25379 30973
rect 26200 30970 27000 31000
rect 25313 30968 27000 30970
rect 25313 30912 25318 30968
rect 25374 30912 27000 30968
rect 25313 30910 27000 30912
rect 25313 30907 25379 30910
rect 26200 30880 27000 30910
rect 10358 30772 10364 30836
rect 10428 30834 10434 30836
rect 11973 30834 12039 30837
rect 19374 30834 19380 30836
rect 10428 30832 19380 30834
rect 10428 30776 11978 30832
rect 12034 30776 19380 30832
rect 10428 30774 19380 30776
rect 10428 30772 10434 30774
rect 11973 30771 12039 30774
rect 19374 30772 19380 30774
rect 19444 30772 19450 30836
rect 15377 30564 15443 30565
rect 15326 30500 15332 30564
rect 15396 30562 15443 30564
rect 19885 30564 19951 30565
rect 19885 30562 19932 30564
rect 15396 30560 15488 30562
rect 15438 30504 15488 30560
rect 15396 30502 15488 30504
rect 19840 30560 19932 30562
rect 19840 30504 19890 30560
rect 19840 30502 19932 30504
rect 15396 30500 15443 30502
rect 15377 30499 15443 30500
rect 19885 30500 19932 30502
rect 19996 30500 20002 30564
rect 21173 30562 21239 30565
rect 25129 30562 25195 30565
rect 21173 30560 25195 30562
rect 21173 30504 21178 30560
rect 21234 30504 25134 30560
rect 25190 30504 25195 30560
rect 21173 30502 25195 30504
rect 19885 30499 19951 30500
rect 21173 30499 21239 30502
rect 25129 30499 25195 30502
rect 7946 30496 8262 30497
rect 7946 30432 7952 30496
rect 8016 30432 8032 30496
rect 8096 30432 8112 30496
rect 8176 30432 8192 30496
rect 8256 30432 8262 30496
rect 7946 30431 8262 30432
rect 17946 30496 18262 30497
rect 17946 30432 17952 30496
rect 18016 30432 18032 30496
rect 18096 30432 18112 30496
rect 18176 30432 18192 30496
rect 18256 30432 18262 30496
rect 17946 30431 18262 30432
rect 25313 30154 25379 30157
rect 26200 30154 27000 30184
rect 25313 30152 27000 30154
rect 25313 30096 25318 30152
rect 25374 30096 27000 30152
rect 25313 30094 27000 30096
rect 25313 30091 25379 30094
rect 26200 30064 27000 30094
rect 18454 29956 18460 30020
rect 18524 30018 18530 30020
rect 18689 30018 18755 30021
rect 19793 30020 19859 30021
rect 18524 30016 18755 30018
rect 18524 29960 18694 30016
rect 18750 29960 18755 30016
rect 18524 29958 18755 29960
rect 18524 29956 18530 29958
rect 18689 29955 18755 29958
rect 19742 29956 19748 30020
rect 19812 30018 19859 30020
rect 19812 30016 19904 30018
rect 19854 29960 19904 30016
rect 19812 29958 19904 29960
rect 19812 29956 19859 29958
rect 19793 29955 19859 29956
rect 2946 29952 3262 29953
rect 2946 29888 2952 29952
rect 3016 29888 3032 29952
rect 3096 29888 3112 29952
rect 3176 29888 3192 29952
rect 3256 29888 3262 29952
rect 2946 29887 3262 29888
rect 12946 29952 13262 29953
rect 12946 29888 12952 29952
rect 13016 29888 13032 29952
rect 13096 29888 13112 29952
rect 13176 29888 13192 29952
rect 13256 29888 13262 29952
rect 12946 29887 13262 29888
rect 22946 29952 23262 29953
rect 22946 29888 22952 29952
rect 23016 29888 23032 29952
rect 23096 29888 23112 29952
rect 23176 29888 23192 29952
rect 23256 29888 23262 29952
rect 22946 29887 23262 29888
rect 16757 29476 16823 29477
rect 16757 29474 16804 29476
rect 16712 29472 16804 29474
rect 16712 29416 16762 29472
rect 16712 29414 16804 29416
rect 16757 29412 16804 29414
rect 16868 29412 16874 29476
rect 16757 29411 16823 29412
rect 7946 29408 8262 29409
rect 7946 29344 7952 29408
rect 8016 29344 8032 29408
rect 8096 29344 8112 29408
rect 8176 29344 8192 29408
rect 8256 29344 8262 29408
rect 7946 29343 8262 29344
rect 17946 29408 18262 29409
rect 17946 29344 17952 29408
rect 18016 29344 18032 29408
rect 18096 29344 18112 29408
rect 18176 29344 18192 29408
rect 18256 29344 18262 29408
rect 17946 29343 18262 29344
rect 15285 29338 15351 29341
rect 15878 29338 15884 29340
rect 15285 29336 15884 29338
rect 15285 29280 15290 29336
rect 15346 29280 15884 29336
rect 15285 29278 15884 29280
rect 15285 29275 15351 29278
rect 15878 29276 15884 29278
rect 15948 29338 15954 29340
rect 17309 29338 17375 29341
rect 15948 29336 17375 29338
rect 15948 29280 17314 29336
rect 17370 29280 17375 29336
rect 15948 29278 17375 29280
rect 15948 29276 15954 29278
rect 17309 29275 17375 29278
rect 25497 29338 25563 29341
rect 26200 29338 27000 29368
rect 25497 29336 27000 29338
rect 25497 29280 25502 29336
rect 25558 29280 27000 29336
rect 25497 29278 27000 29280
rect 25497 29275 25563 29278
rect 26200 29248 27000 29278
rect 15326 29004 15332 29068
rect 15396 29066 15402 29068
rect 16246 29066 16252 29068
rect 15396 29006 16252 29066
rect 15396 29004 15402 29006
rect 16246 29004 16252 29006
rect 16316 29066 16322 29068
rect 19793 29066 19859 29069
rect 16316 29064 19859 29066
rect 16316 29008 19798 29064
rect 19854 29008 19859 29064
rect 16316 29006 19859 29008
rect 16316 29004 16322 29006
rect 19793 29003 19859 29006
rect 2946 28864 3262 28865
rect 2946 28800 2952 28864
rect 3016 28800 3032 28864
rect 3096 28800 3112 28864
rect 3176 28800 3192 28864
rect 3256 28800 3262 28864
rect 2946 28799 3262 28800
rect 12946 28864 13262 28865
rect 12946 28800 12952 28864
rect 13016 28800 13032 28864
rect 13096 28800 13112 28864
rect 13176 28800 13192 28864
rect 13256 28800 13262 28864
rect 12946 28799 13262 28800
rect 22946 28864 23262 28865
rect 22946 28800 22952 28864
rect 23016 28800 23032 28864
rect 23096 28800 23112 28864
rect 23176 28800 23192 28864
rect 23256 28800 23262 28864
rect 22946 28799 23262 28800
rect 0 28522 800 28552
rect 2865 28522 2931 28525
rect 0 28520 2931 28522
rect 0 28464 2870 28520
rect 2926 28464 2931 28520
rect 0 28462 2931 28464
rect 0 28432 800 28462
rect 2865 28459 2931 28462
rect 25221 28522 25287 28525
rect 26200 28522 27000 28552
rect 25221 28520 27000 28522
rect 25221 28464 25226 28520
rect 25282 28464 27000 28520
rect 25221 28462 27000 28464
rect 25221 28459 25287 28462
rect 26200 28432 27000 28462
rect 17309 28388 17375 28389
rect 17309 28386 17356 28388
rect 17264 28384 17356 28386
rect 17264 28328 17314 28384
rect 17264 28326 17356 28328
rect 17309 28324 17356 28326
rect 17420 28324 17426 28388
rect 17534 28324 17540 28388
rect 17604 28386 17610 28388
rect 17677 28386 17743 28389
rect 17604 28384 17743 28386
rect 17604 28328 17682 28384
rect 17738 28328 17743 28384
rect 17604 28326 17743 28328
rect 17604 28324 17610 28326
rect 17309 28323 17375 28324
rect 17677 28323 17743 28326
rect 7946 28320 8262 28321
rect 7946 28256 7952 28320
rect 8016 28256 8032 28320
rect 8096 28256 8112 28320
rect 8176 28256 8192 28320
rect 8256 28256 8262 28320
rect 7946 28255 8262 28256
rect 17946 28320 18262 28321
rect 17946 28256 17952 28320
rect 18016 28256 18032 28320
rect 18096 28256 18112 28320
rect 18176 28256 18192 28320
rect 18256 28256 18262 28320
rect 17946 28255 18262 28256
rect 15377 28250 15443 28253
rect 17677 28252 17743 28253
rect 15694 28250 15700 28252
rect 15377 28248 15700 28250
rect 15377 28192 15382 28248
rect 15438 28192 15700 28248
rect 15377 28190 15700 28192
rect 15377 28187 15443 28190
rect 15694 28188 15700 28190
rect 15764 28188 15770 28252
rect 17677 28250 17724 28252
rect 17632 28248 17724 28250
rect 17632 28192 17682 28248
rect 17632 28190 17724 28192
rect 17677 28188 17724 28190
rect 17788 28188 17794 28252
rect 15702 28114 15762 28188
rect 17677 28187 17743 28188
rect 20713 28114 20779 28117
rect 15702 28112 20779 28114
rect 15702 28056 20718 28112
rect 20774 28056 20779 28112
rect 15702 28054 20779 28056
rect 20713 28051 20779 28054
rect 2946 27776 3262 27777
rect 2946 27712 2952 27776
rect 3016 27712 3032 27776
rect 3096 27712 3112 27776
rect 3176 27712 3192 27776
rect 3256 27712 3262 27776
rect 2946 27711 3262 27712
rect 12946 27776 13262 27777
rect 12946 27712 12952 27776
rect 13016 27712 13032 27776
rect 13096 27712 13112 27776
rect 13176 27712 13192 27776
rect 13256 27712 13262 27776
rect 12946 27711 13262 27712
rect 22946 27776 23262 27777
rect 22946 27712 22952 27776
rect 23016 27712 23032 27776
rect 23096 27712 23112 27776
rect 23176 27712 23192 27776
rect 23256 27712 23262 27776
rect 22946 27711 23262 27712
rect 24117 27706 24183 27709
rect 26200 27706 27000 27736
rect 24117 27704 27000 27706
rect 24117 27648 24122 27704
rect 24178 27648 27000 27704
rect 24117 27646 27000 27648
rect 24117 27643 24183 27646
rect 26200 27616 27000 27646
rect 7946 27232 8262 27233
rect 7946 27168 7952 27232
rect 8016 27168 8032 27232
rect 8096 27168 8112 27232
rect 8176 27168 8192 27232
rect 8256 27168 8262 27232
rect 7946 27167 8262 27168
rect 17946 27232 18262 27233
rect 17946 27168 17952 27232
rect 18016 27168 18032 27232
rect 18096 27168 18112 27232
rect 18176 27168 18192 27232
rect 18256 27168 18262 27232
rect 17946 27167 18262 27168
rect 20437 27162 20503 27165
rect 21950 27162 21956 27164
rect 20437 27160 21956 27162
rect 20437 27104 20442 27160
rect 20498 27104 21956 27160
rect 20437 27102 21956 27104
rect 20437 27099 20503 27102
rect 21950 27100 21956 27102
rect 22020 27100 22026 27164
rect 17309 26890 17375 26893
rect 19742 26890 19748 26892
rect 17309 26888 19748 26890
rect 17309 26832 17314 26888
rect 17370 26832 19748 26888
rect 17309 26830 19748 26832
rect 17309 26827 17375 26830
rect 19742 26828 19748 26830
rect 19812 26828 19818 26892
rect 23381 26890 23447 26893
rect 26200 26890 27000 26920
rect 23381 26888 27000 26890
rect 23381 26832 23386 26888
rect 23442 26832 27000 26888
rect 23381 26830 27000 26832
rect 23381 26827 23447 26830
rect 26200 26800 27000 26830
rect 14038 26692 14044 26756
rect 14108 26754 14114 26756
rect 14958 26754 14964 26756
rect 14108 26694 14964 26754
rect 14108 26692 14114 26694
rect 14958 26692 14964 26694
rect 15028 26754 15034 26756
rect 16113 26754 16179 26757
rect 15028 26752 16179 26754
rect 15028 26696 16118 26752
rect 16174 26696 16179 26752
rect 15028 26694 16179 26696
rect 15028 26692 15034 26694
rect 16113 26691 16179 26694
rect 2946 26688 3262 26689
rect 2946 26624 2952 26688
rect 3016 26624 3032 26688
rect 3096 26624 3112 26688
rect 3176 26624 3192 26688
rect 3256 26624 3262 26688
rect 2946 26623 3262 26624
rect 12946 26688 13262 26689
rect 12946 26624 12952 26688
rect 13016 26624 13032 26688
rect 13096 26624 13112 26688
rect 13176 26624 13192 26688
rect 13256 26624 13262 26688
rect 12946 26623 13262 26624
rect 22946 26688 23262 26689
rect 22946 26624 22952 26688
rect 23016 26624 23032 26688
rect 23096 26624 23112 26688
rect 23176 26624 23192 26688
rect 23256 26624 23262 26688
rect 22946 26623 23262 26624
rect 20805 26618 20871 26621
rect 21030 26618 21036 26620
rect 20805 26616 21036 26618
rect 20805 26560 20810 26616
rect 20866 26560 21036 26616
rect 20805 26558 21036 26560
rect 20805 26555 20871 26558
rect 21030 26556 21036 26558
rect 21100 26556 21106 26620
rect 7946 26144 8262 26145
rect 0 26074 800 26104
rect 7946 26080 7952 26144
rect 8016 26080 8032 26144
rect 8096 26080 8112 26144
rect 8176 26080 8192 26144
rect 8256 26080 8262 26144
rect 7946 26079 8262 26080
rect 17946 26144 18262 26145
rect 17946 26080 17952 26144
rect 18016 26080 18032 26144
rect 18096 26080 18112 26144
rect 18176 26080 18192 26144
rect 18256 26080 18262 26144
rect 17946 26079 18262 26080
rect 2773 26074 2839 26077
rect 0 26072 2839 26074
rect 0 26016 2778 26072
rect 2834 26016 2839 26072
rect 0 26014 2839 26016
rect 0 25984 800 26014
rect 2773 26011 2839 26014
rect 22553 26074 22619 26077
rect 26200 26074 27000 26104
rect 22553 26072 27000 26074
rect 22553 26016 22558 26072
rect 22614 26016 27000 26072
rect 22553 26014 27000 26016
rect 22553 26011 22619 26014
rect 26200 25984 27000 26014
rect 2946 25600 3262 25601
rect 2946 25536 2952 25600
rect 3016 25536 3032 25600
rect 3096 25536 3112 25600
rect 3176 25536 3192 25600
rect 3256 25536 3262 25600
rect 2946 25535 3262 25536
rect 12946 25600 13262 25601
rect 12946 25536 12952 25600
rect 13016 25536 13032 25600
rect 13096 25536 13112 25600
rect 13176 25536 13192 25600
rect 13256 25536 13262 25600
rect 12946 25535 13262 25536
rect 22946 25600 23262 25601
rect 22946 25536 22952 25600
rect 23016 25536 23032 25600
rect 23096 25536 23112 25600
rect 23176 25536 23192 25600
rect 23256 25536 23262 25600
rect 22946 25535 23262 25536
rect 25129 25258 25195 25261
rect 26200 25258 27000 25288
rect 25129 25256 27000 25258
rect 25129 25200 25134 25256
rect 25190 25200 27000 25256
rect 25129 25198 27000 25200
rect 25129 25195 25195 25198
rect 26200 25168 27000 25198
rect 7946 25056 8262 25057
rect 7946 24992 7952 25056
rect 8016 24992 8032 25056
rect 8096 24992 8112 25056
rect 8176 24992 8192 25056
rect 8256 24992 8262 25056
rect 7946 24991 8262 24992
rect 17946 25056 18262 25057
rect 17946 24992 17952 25056
rect 18016 24992 18032 25056
rect 18096 24992 18112 25056
rect 18176 24992 18192 25056
rect 18256 24992 18262 25056
rect 17946 24991 18262 24992
rect 9622 24788 9628 24852
rect 9692 24850 9698 24852
rect 11421 24850 11487 24853
rect 9692 24848 11487 24850
rect 9692 24792 11426 24848
rect 11482 24792 11487 24848
rect 9692 24790 11487 24792
rect 9692 24788 9698 24790
rect 11421 24787 11487 24790
rect 2946 24512 3262 24513
rect 2946 24448 2952 24512
rect 3016 24448 3032 24512
rect 3096 24448 3112 24512
rect 3176 24448 3192 24512
rect 3256 24448 3262 24512
rect 2946 24447 3262 24448
rect 12946 24512 13262 24513
rect 12946 24448 12952 24512
rect 13016 24448 13032 24512
rect 13096 24448 13112 24512
rect 13176 24448 13192 24512
rect 13256 24448 13262 24512
rect 12946 24447 13262 24448
rect 22946 24512 23262 24513
rect 22946 24448 22952 24512
rect 23016 24448 23032 24512
rect 23096 24448 23112 24512
rect 23176 24448 23192 24512
rect 23256 24448 23262 24512
rect 22946 24447 23262 24448
rect 24853 24442 24919 24445
rect 26200 24442 27000 24472
rect 24853 24440 27000 24442
rect 24853 24384 24858 24440
rect 24914 24384 27000 24440
rect 24853 24382 27000 24384
rect 24853 24379 24919 24382
rect 26200 24352 27000 24382
rect 7946 23968 8262 23969
rect 7946 23904 7952 23968
rect 8016 23904 8032 23968
rect 8096 23904 8112 23968
rect 8176 23904 8192 23968
rect 8256 23904 8262 23968
rect 7946 23903 8262 23904
rect 17946 23968 18262 23969
rect 17946 23904 17952 23968
rect 18016 23904 18032 23968
rect 18096 23904 18112 23968
rect 18176 23904 18192 23968
rect 18256 23904 18262 23968
rect 17946 23903 18262 23904
rect 13721 23762 13787 23765
rect 18454 23762 18460 23764
rect 13721 23760 18460 23762
rect 13721 23704 13726 23760
rect 13782 23704 18460 23760
rect 13721 23702 18460 23704
rect 13721 23699 13787 23702
rect 18454 23700 18460 23702
rect 18524 23700 18530 23764
rect 0 23626 800 23656
rect 2865 23626 2931 23629
rect 0 23624 2931 23626
rect 0 23568 2870 23624
rect 2926 23568 2931 23624
rect 0 23566 2931 23568
rect 0 23536 800 23566
rect 2865 23563 2931 23566
rect 23841 23626 23907 23629
rect 26200 23626 27000 23656
rect 23841 23624 27000 23626
rect 23841 23568 23846 23624
rect 23902 23568 27000 23624
rect 23841 23566 27000 23568
rect 23841 23563 23907 23566
rect 26200 23536 27000 23566
rect 2946 23424 3262 23425
rect 2946 23360 2952 23424
rect 3016 23360 3032 23424
rect 3096 23360 3112 23424
rect 3176 23360 3192 23424
rect 3256 23360 3262 23424
rect 2946 23359 3262 23360
rect 12946 23424 13262 23425
rect 12946 23360 12952 23424
rect 13016 23360 13032 23424
rect 13096 23360 13112 23424
rect 13176 23360 13192 23424
rect 13256 23360 13262 23424
rect 12946 23359 13262 23360
rect 22946 23424 23262 23425
rect 22946 23360 22952 23424
rect 23016 23360 23032 23424
rect 23096 23360 23112 23424
rect 23176 23360 23192 23424
rect 23256 23360 23262 23424
rect 22946 23359 23262 23360
rect 11789 23218 11855 23221
rect 15745 23218 15811 23221
rect 11789 23216 15811 23218
rect 11789 23160 11794 23216
rect 11850 23160 15750 23216
rect 15806 23160 15811 23216
rect 11789 23158 15811 23160
rect 11789 23155 11855 23158
rect 15745 23155 15811 23158
rect 7946 22880 8262 22881
rect 7946 22816 7952 22880
rect 8016 22816 8032 22880
rect 8096 22816 8112 22880
rect 8176 22816 8192 22880
rect 8256 22816 8262 22880
rect 7946 22815 8262 22816
rect 17946 22880 18262 22881
rect 17946 22816 17952 22880
rect 18016 22816 18032 22880
rect 18096 22816 18112 22880
rect 18176 22816 18192 22880
rect 18256 22816 18262 22880
rect 17946 22815 18262 22816
rect 23289 22810 23355 22813
rect 26200 22810 27000 22840
rect 23289 22808 27000 22810
rect 23289 22752 23294 22808
rect 23350 22752 27000 22808
rect 23289 22750 27000 22752
rect 23289 22747 23355 22750
rect 26200 22720 27000 22750
rect 2946 22336 3262 22337
rect 2946 22272 2952 22336
rect 3016 22272 3032 22336
rect 3096 22272 3112 22336
rect 3176 22272 3192 22336
rect 3256 22272 3262 22336
rect 2946 22271 3262 22272
rect 12946 22336 13262 22337
rect 12946 22272 12952 22336
rect 13016 22272 13032 22336
rect 13096 22272 13112 22336
rect 13176 22272 13192 22336
rect 13256 22272 13262 22336
rect 12946 22271 13262 22272
rect 22946 22336 23262 22337
rect 22946 22272 22952 22336
rect 23016 22272 23032 22336
rect 23096 22272 23112 22336
rect 23176 22272 23192 22336
rect 23256 22272 23262 22336
rect 22946 22271 23262 22272
rect 16113 22266 16179 22269
rect 21214 22266 21220 22268
rect 16113 22264 21220 22266
rect 16113 22208 16118 22264
rect 16174 22208 21220 22264
rect 16113 22206 21220 22208
rect 16113 22203 16179 22206
rect 21214 22204 21220 22206
rect 21284 22204 21290 22268
rect 24853 21994 24919 21997
rect 26200 21994 27000 22024
rect 24853 21992 27000 21994
rect 24853 21936 24858 21992
rect 24914 21936 27000 21992
rect 24853 21934 27000 21936
rect 24853 21931 24919 21934
rect 26200 21904 27000 21934
rect 7946 21792 8262 21793
rect 7946 21728 7952 21792
rect 8016 21728 8032 21792
rect 8096 21728 8112 21792
rect 8176 21728 8192 21792
rect 8256 21728 8262 21792
rect 7946 21727 8262 21728
rect 17946 21792 18262 21793
rect 17946 21728 17952 21792
rect 18016 21728 18032 21792
rect 18096 21728 18112 21792
rect 18176 21728 18192 21792
rect 18256 21728 18262 21792
rect 17946 21727 18262 21728
rect 12433 21586 12499 21589
rect 13629 21586 13695 21589
rect 12433 21584 13695 21586
rect 12433 21528 12438 21584
rect 12494 21528 13634 21584
rect 13690 21528 13695 21584
rect 12433 21526 13695 21528
rect 12433 21523 12499 21526
rect 13629 21523 13695 21526
rect 2946 21248 3262 21249
rect 0 21178 800 21208
rect 2946 21184 2952 21248
rect 3016 21184 3032 21248
rect 3096 21184 3112 21248
rect 3176 21184 3192 21248
rect 3256 21184 3262 21248
rect 2946 21183 3262 21184
rect 12946 21248 13262 21249
rect 12946 21184 12952 21248
rect 13016 21184 13032 21248
rect 13096 21184 13112 21248
rect 13176 21184 13192 21248
rect 13256 21184 13262 21248
rect 12946 21183 13262 21184
rect 22946 21248 23262 21249
rect 22946 21184 22952 21248
rect 23016 21184 23032 21248
rect 23096 21184 23112 21248
rect 23176 21184 23192 21248
rect 23256 21184 23262 21248
rect 22946 21183 23262 21184
rect 1301 21178 1367 21181
rect 0 21176 1367 21178
rect 0 21120 1306 21176
rect 1362 21120 1367 21176
rect 0 21118 1367 21120
rect 0 21088 800 21118
rect 1301 21115 1367 21118
rect 15837 21178 15903 21181
rect 16062 21178 16068 21180
rect 15837 21176 16068 21178
rect 15837 21120 15842 21176
rect 15898 21120 16068 21176
rect 15837 21118 16068 21120
rect 15837 21115 15903 21118
rect 16062 21116 16068 21118
rect 16132 21178 16138 21180
rect 16665 21178 16731 21181
rect 16132 21176 16731 21178
rect 16132 21120 16670 21176
rect 16726 21120 16731 21176
rect 16132 21118 16731 21120
rect 16132 21116 16138 21118
rect 16665 21115 16731 21118
rect 23381 21178 23447 21181
rect 26200 21178 27000 21208
rect 23381 21176 27000 21178
rect 23381 21120 23386 21176
rect 23442 21120 27000 21176
rect 23381 21118 27000 21120
rect 23381 21115 23447 21118
rect 26200 21088 27000 21118
rect 7946 20704 8262 20705
rect 7946 20640 7952 20704
rect 8016 20640 8032 20704
rect 8096 20640 8112 20704
rect 8176 20640 8192 20704
rect 8256 20640 8262 20704
rect 7946 20639 8262 20640
rect 17946 20704 18262 20705
rect 17946 20640 17952 20704
rect 18016 20640 18032 20704
rect 18096 20640 18112 20704
rect 18176 20640 18192 20704
rect 18256 20640 18262 20704
rect 17946 20639 18262 20640
rect 15929 20498 15995 20501
rect 20662 20498 20668 20500
rect 15929 20496 20668 20498
rect 15929 20440 15934 20496
rect 15990 20440 20668 20496
rect 15929 20438 20668 20440
rect 15929 20435 15995 20438
rect 20662 20436 20668 20438
rect 20732 20436 20738 20500
rect 24945 20362 25011 20365
rect 26200 20362 27000 20392
rect 24945 20360 27000 20362
rect 24945 20304 24950 20360
rect 25006 20304 27000 20360
rect 24945 20302 27000 20304
rect 24945 20299 25011 20302
rect 26200 20272 27000 20302
rect 2946 20160 3262 20161
rect 2946 20096 2952 20160
rect 3016 20096 3032 20160
rect 3096 20096 3112 20160
rect 3176 20096 3192 20160
rect 3256 20096 3262 20160
rect 2946 20095 3262 20096
rect 12946 20160 13262 20161
rect 12946 20096 12952 20160
rect 13016 20096 13032 20160
rect 13096 20096 13112 20160
rect 13176 20096 13192 20160
rect 13256 20096 13262 20160
rect 12946 20095 13262 20096
rect 22946 20160 23262 20161
rect 22946 20096 22952 20160
rect 23016 20096 23032 20160
rect 23096 20096 23112 20160
rect 23176 20096 23192 20160
rect 23256 20096 23262 20160
rect 22946 20095 23262 20096
rect 7946 19616 8262 19617
rect 7946 19552 7952 19616
rect 8016 19552 8032 19616
rect 8096 19552 8112 19616
rect 8176 19552 8192 19616
rect 8256 19552 8262 19616
rect 7946 19551 8262 19552
rect 17946 19616 18262 19617
rect 17946 19552 17952 19616
rect 18016 19552 18032 19616
rect 18096 19552 18112 19616
rect 18176 19552 18192 19616
rect 18256 19552 18262 19616
rect 17946 19551 18262 19552
rect 24761 19546 24827 19549
rect 26200 19546 27000 19576
rect 24761 19544 27000 19546
rect 24761 19488 24766 19544
rect 24822 19488 27000 19544
rect 24761 19486 27000 19488
rect 24761 19483 24827 19486
rect 26200 19456 27000 19486
rect 7005 19274 7071 19277
rect 13721 19276 13787 19277
rect 9622 19274 9628 19276
rect 7005 19272 9628 19274
rect 7005 19216 7010 19272
rect 7066 19216 9628 19272
rect 7005 19214 9628 19216
rect 7005 19211 7071 19214
rect 9622 19212 9628 19214
rect 9692 19212 9698 19276
rect 13670 19212 13676 19276
rect 13740 19274 13787 19276
rect 13740 19272 13832 19274
rect 13782 19216 13832 19272
rect 13740 19214 13832 19216
rect 13740 19212 13787 19214
rect 13721 19211 13787 19212
rect 2946 19072 3262 19073
rect 2946 19008 2952 19072
rect 3016 19008 3032 19072
rect 3096 19008 3112 19072
rect 3176 19008 3192 19072
rect 3256 19008 3262 19072
rect 2946 19007 3262 19008
rect 12946 19072 13262 19073
rect 12946 19008 12952 19072
rect 13016 19008 13032 19072
rect 13096 19008 13112 19072
rect 13176 19008 13192 19072
rect 13256 19008 13262 19072
rect 12946 19007 13262 19008
rect 22946 19072 23262 19073
rect 22946 19008 22952 19072
rect 23016 19008 23032 19072
rect 23096 19008 23112 19072
rect 23176 19008 23192 19072
rect 23256 19008 23262 19072
rect 22946 19007 23262 19008
rect 13537 18866 13603 18869
rect 15694 18866 15700 18868
rect 13537 18864 15700 18866
rect 13537 18808 13542 18864
rect 13598 18808 15700 18864
rect 13537 18806 15700 18808
rect 13537 18803 13603 18806
rect 15694 18804 15700 18806
rect 15764 18804 15770 18868
rect 0 18730 800 18760
rect 1301 18730 1367 18733
rect 17585 18732 17651 18733
rect 17534 18730 17540 18732
rect 0 18728 1367 18730
rect 0 18672 1306 18728
rect 1362 18672 1367 18728
rect 0 18670 1367 18672
rect 17494 18670 17540 18730
rect 17604 18728 17651 18732
rect 17646 18672 17651 18728
rect 0 18640 800 18670
rect 1301 18667 1367 18670
rect 17534 18668 17540 18670
rect 17604 18668 17651 18672
rect 17585 18667 17651 18668
rect 18321 18730 18387 18733
rect 18873 18730 18939 18733
rect 19926 18730 19932 18732
rect 18321 18728 19932 18730
rect 18321 18672 18326 18728
rect 18382 18672 18878 18728
rect 18934 18672 19932 18728
rect 18321 18670 19932 18672
rect 18321 18667 18387 18670
rect 18873 18667 18939 18670
rect 19926 18668 19932 18670
rect 19996 18668 20002 18732
rect 24669 18730 24735 18733
rect 26200 18730 27000 18760
rect 24669 18728 27000 18730
rect 24669 18672 24674 18728
rect 24730 18672 27000 18728
rect 24669 18670 27000 18672
rect 24669 18667 24735 18670
rect 26200 18640 27000 18670
rect 14733 18596 14799 18597
rect 14733 18594 14780 18596
rect 14688 18592 14780 18594
rect 14688 18536 14738 18592
rect 14688 18534 14780 18536
rect 14733 18532 14780 18534
rect 14844 18532 14850 18596
rect 14733 18531 14799 18532
rect 7946 18528 8262 18529
rect 7946 18464 7952 18528
rect 8016 18464 8032 18528
rect 8096 18464 8112 18528
rect 8176 18464 8192 18528
rect 8256 18464 8262 18528
rect 7946 18463 8262 18464
rect 17946 18528 18262 18529
rect 17946 18464 17952 18528
rect 18016 18464 18032 18528
rect 18096 18464 18112 18528
rect 18176 18464 18192 18528
rect 18256 18464 18262 18528
rect 17946 18463 18262 18464
rect 12014 18260 12020 18324
rect 12084 18322 12090 18324
rect 12341 18322 12407 18325
rect 12084 18320 12407 18322
rect 12084 18264 12346 18320
rect 12402 18264 12407 18320
rect 12084 18262 12407 18264
rect 12084 18260 12090 18262
rect 12341 18259 12407 18262
rect 2946 17984 3262 17985
rect 2946 17920 2952 17984
rect 3016 17920 3032 17984
rect 3096 17920 3112 17984
rect 3176 17920 3192 17984
rect 3256 17920 3262 17984
rect 2946 17919 3262 17920
rect 12946 17984 13262 17985
rect 12946 17920 12952 17984
rect 13016 17920 13032 17984
rect 13096 17920 13112 17984
rect 13176 17920 13192 17984
rect 13256 17920 13262 17984
rect 12946 17919 13262 17920
rect 22946 17984 23262 17985
rect 22946 17920 22952 17984
rect 23016 17920 23032 17984
rect 23096 17920 23112 17984
rect 23176 17920 23192 17984
rect 23256 17920 23262 17984
rect 22946 17919 23262 17920
rect 23381 17914 23447 17917
rect 26200 17914 27000 17944
rect 23381 17912 27000 17914
rect 23381 17856 23386 17912
rect 23442 17856 27000 17912
rect 23381 17854 27000 17856
rect 23381 17851 23447 17854
rect 26200 17824 27000 17854
rect 7946 17440 8262 17441
rect 7946 17376 7952 17440
rect 8016 17376 8032 17440
rect 8096 17376 8112 17440
rect 8176 17376 8192 17440
rect 8256 17376 8262 17440
rect 7946 17375 8262 17376
rect 17946 17440 18262 17441
rect 17946 17376 17952 17440
rect 18016 17376 18032 17440
rect 18096 17376 18112 17440
rect 18176 17376 18192 17440
rect 18256 17376 18262 17440
rect 17946 17375 18262 17376
rect 24761 17098 24827 17101
rect 26200 17098 27000 17128
rect 24761 17096 27000 17098
rect 24761 17040 24766 17096
rect 24822 17040 27000 17096
rect 24761 17038 27000 17040
rect 24761 17035 24827 17038
rect 26200 17008 27000 17038
rect 2946 16896 3262 16897
rect 2946 16832 2952 16896
rect 3016 16832 3032 16896
rect 3096 16832 3112 16896
rect 3176 16832 3192 16896
rect 3256 16832 3262 16896
rect 2946 16831 3262 16832
rect 12946 16896 13262 16897
rect 12946 16832 12952 16896
rect 13016 16832 13032 16896
rect 13096 16832 13112 16896
rect 13176 16832 13192 16896
rect 13256 16832 13262 16896
rect 12946 16831 13262 16832
rect 22946 16896 23262 16897
rect 22946 16832 22952 16896
rect 23016 16832 23032 16896
rect 23096 16832 23112 16896
rect 23176 16832 23192 16896
rect 23256 16832 23262 16896
rect 22946 16831 23262 16832
rect 12433 16826 12499 16829
rect 12566 16826 12572 16828
rect 12433 16824 12572 16826
rect 12433 16768 12438 16824
rect 12494 16768 12572 16824
rect 12433 16766 12572 16768
rect 12433 16763 12499 16766
rect 12566 16764 12572 16766
rect 12636 16826 12642 16828
rect 12801 16826 12867 16829
rect 12636 16824 12867 16826
rect 12636 16768 12806 16824
rect 12862 16768 12867 16824
rect 12636 16766 12867 16768
rect 12636 16764 12642 16766
rect 12801 16763 12867 16766
rect 20713 16556 20779 16557
rect 20662 16554 20668 16556
rect 20622 16494 20668 16554
rect 20732 16552 20779 16556
rect 20774 16496 20779 16552
rect 20662 16492 20668 16494
rect 20732 16492 20779 16496
rect 20713 16491 20779 16492
rect 21081 16554 21147 16557
rect 21214 16554 21220 16556
rect 21081 16552 21220 16554
rect 21081 16496 21086 16552
rect 21142 16496 21220 16552
rect 21081 16494 21220 16496
rect 21081 16491 21147 16494
rect 21214 16492 21220 16494
rect 21284 16492 21290 16556
rect 7946 16352 8262 16353
rect 0 16282 800 16312
rect 7946 16288 7952 16352
rect 8016 16288 8032 16352
rect 8096 16288 8112 16352
rect 8176 16288 8192 16352
rect 8256 16288 8262 16352
rect 7946 16287 8262 16288
rect 17946 16352 18262 16353
rect 17946 16288 17952 16352
rect 18016 16288 18032 16352
rect 18096 16288 18112 16352
rect 18176 16288 18192 16352
rect 18256 16288 18262 16352
rect 17946 16287 18262 16288
rect 1301 16282 1367 16285
rect 16205 16284 16271 16285
rect 16205 16282 16252 16284
rect 0 16280 1367 16282
rect 0 16224 1306 16280
rect 1362 16224 1367 16280
rect 0 16222 1367 16224
rect 16160 16280 16252 16282
rect 16160 16224 16210 16280
rect 16160 16222 16252 16224
rect 0 16192 800 16222
rect 1301 16219 1367 16222
rect 16205 16220 16252 16222
rect 16316 16220 16322 16284
rect 24669 16282 24735 16285
rect 26200 16282 27000 16312
rect 24669 16280 27000 16282
rect 24669 16224 24674 16280
rect 24730 16224 27000 16280
rect 24669 16222 27000 16224
rect 16205 16219 16271 16220
rect 24669 16219 24735 16222
rect 26200 16192 27000 16222
rect 2946 15808 3262 15809
rect 2946 15744 2952 15808
rect 3016 15744 3032 15808
rect 3096 15744 3112 15808
rect 3176 15744 3192 15808
rect 3256 15744 3262 15808
rect 2946 15743 3262 15744
rect 12946 15808 13262 15809
rect 12946 15744 12952 15808
rect 13016 15744 13032 15808
rect 13096 15744 13112 15808
rect 13176 15744 13192 15808
rect 13256 15744 13262 15808
rect 12946 15743 13262 15744
rect 22946 15808 23262 15809
rect 22946 15744 22952 15808
rect 23016 15744 23032 15808
rect 23096 15744 23112 15808
rect 23176 15744 23192 15808
rect 23256 15744 23262 15808
rect 22946 15743 23262 15744
rect 15009 15740 15075 15741
rect 14958 15676 14964 15740
rect 15028 15738 15075 15740
rect 15028 15736 15120 15738
rect 15070 15680 15120 15736
rect 15028 15678 15120 15680
rect 15028 15676 15075 15678
rect 15009 15675 15075 15676
rect 24945 15466 25011 15469
rect 26200 15466 27000 15496
rect 24945 15464 27000 15466
rect 24945 15408 24950 15464
rect 25006 15408 27000 15464
rect 24945 15406 27000 15408
rect 24945 15403 25011 15406
rect 26200 15376 27000 15406
rect 7946 15264 8262 15265
rect 7946 15200 7952 15264
rect 8016 15200 8032 15264
rect 8096 15200 8112 15264
rect 8176 15200 8192 15264
rect 8256 15200 8262 15264
rect 7946 15199 8262 15200
rect 17946 15264 18262 15265
rect 17946 15200 17952 15264
rect 18016 15200 18032 15264
rect 18096 15200 18112 15264
rect 18176 15200 18192 15264
rect 18256 15200 18262 15264
rect 17946 15199 18262 15200
rect 14273 15194 14339 15197
rect 15878 15194 15884 15196
rect 14273 15192 15884 15194
rect 14273 15136 14278 15192
rect 14334 15136 15884 15192
rect 14273 15134 15884 15136
rect 14273 15131 14339 15134
rect 15878 15132 15884 15134
rect 15948 15132 15954 15196
rect 2946 14720 3262 14721
rect 2946 14656 2952 14720
rect 3016 14656 3032 14720
rect 3096 14656 3112 14720
rect 3176 14656 3192 14720
rect 3256 14656 3262 14720
rect 2946 14655 3262 14656
rect 12946 14720 13262 14721
rect 12946 14656 12952 14720
rect 13016 14656 13032 14720
rect 13096 14656 13112 14720
rect 13176 14656 13192 14720
rect 13256 14656 13262 14720
rect 12946 14655 13262 14656
rect 22946 14720 23262 14721
rect 22946 14656 22952 14720
rect 23016 14656 23032 14720
rect 23096 14656 23112 14720
rect 23176 14656 23192 14720
rect 23256 14656 23262 14720
rect 22946 14655 23262 14656
rect 25129 14650 25195 14653
rect 26200 14650 27000 14680
rect 25129 14648 27000 14650
rect 25129 14592 25134 14648
rect 25190 14592 27000 14648
rect 25129 14590 27000 14592
rect 25129 14587 25195 14590
rect 26200 14560 27000 14590
rect 18413 14516 18479 14517
rect 18413 14514 18460 14516
rect 18368 14512 18460 14514
rect 18368 14456 18418 14512
rect 18368 14454 18460 14456
rect 18413 14452 18460 14454
rect 18524 14452 18530 14516
rect 18413 14451 18479 14452
rect 7946 14176 8262 14177
rect 7946 14112 7952 14176
rect 8016 14112 8032 14176
rect 8096 14112 8112 14176
rect 8176 14112 8192 14176
rect 8256 14112 8262 14176
rect 7946 14111 8262 14112
rect 17946 14176 18262 14177
rect 17946 14112 17952 14176
rect 18016 14112 18032 14176
rect 18096 14112 18112 14176
rect 18176 14112 18192 14176
rect 18256 14112 18262 14176
rect 17946 14111 18262 14112
rect 14917 14106 14983 14109
rect 17350 14106 17356 14108
rect 14917 14104 17356 14106
rect 14917 14048 14922 14104
rect 14978 14048 17356 14104
rect 14917 14046 17356 14048
rect 14917 14043 14983 14046
rect 17350 14044 17356 14046
rect 17420 14044 17426 14108
rect 0 13834 800 13864
rect 1301 13834 1367 13837
rect 0 13832 1367 13834
rect 0 13776 1306 13832
rect 1362 13776 1367 13832
rect 0 13774 1367 13776
rect 0 13744 800 13774
rect 1301 13771 1367 13774
rect 24761 13834 24827 13837
rect 26200 13834 27000 13864
rect 24761 13832 27000 13834
rect 24761 13776 24766 13832
rect 24822 13776 27000 13832
rect 24761 13774 27000 13776
rect 24761 13771 24827 13774
rect 26200 13744 27000 13774
rect 2946 13632 3262 13633
rect 2946 13568 2952 13632
rect 3016 13568 3032 13632
rect 3096 13568 3112 13632
rect 3176 13568 3192 13632
rect 3256 13568 3262 13632
rect 2946 13567 3262 13568
rect 12946 13632 13262 13633
rect 12946 13568 12952 13632
rect 13016 13568 13032 13632
rect 13096 13568 13112 13632
rect 13176 13568 13192 13632
rect 13256 13568 13262 13632
rect 12946 13567 13262 13568
rect 22946 13632 23262 13633
rect 22946 13568 22952 13632
rect 23016 13568 23032 13632
rect 23096 13568 23112 13632
rect 23176 13568 23192 13632
rect 23256 13568 23262 13632
rect 22946 13567 23262 13568
rect 13353 13154 13419 13157
rect 13670 13154 13676 13156
rect 13353 13152 13676 13154
rect 13353 13096 13358 13152
rect 13414 13096 13676 13152
rect 13353 13094 13676 13096
rect 13353 13091 13419 13094
rect 13670 13092 13676 13094
rect 13740 13092 13746 13156
rect 7946 13088 8262 13089
rect 7946 13024 7952 13088
rect 8016 13024 8032 13088
rect 8096 13024 8112 13088
rect 8176 13024 8192 13088
rect 8256 13024 8262 13088
rect 7946 13023 8262 13024
rect 17946 13088 18262 13089
rect 17946 13024 17952 13088
rect 18016 13024 18032 13088
rect 18096 13024 18112 13088
rect 18176 13024 18192 13088
rect 18256 13024 18262 13088
rect 17946 13023 18262 13024
rect 24945 13018 25011 13021
rect 26200 13018 27000 13048
rect 24945 13016 27000 13018
rect 24945 12960 24950 13016
rect 25006 12960 27000 13016
rect 24945 12958 27000 12960
rect 24945 12955 25011 12958
rect 26200 12928 27000 12958
rect 2946 12544 3262 12545
rect 2946 12480 2952 12544
rect 3016 12480 3032 12544
rect 3096 12480 3112 12544
rect 3176 12480 3192 12544
rect 3256 12480 3262 12544
rect 2946 12479 3262 12480
rect 12946 12544 13262 12545
rect 12946 12480 12952 12544
rect 13016 12480 13032 12544
rect 13096 12480 13112 12544
rect 13176 12480 13192 12544
rect 13256 12480 13262 12544
rect 12946 12479 13262 12480
rect 22946 12544 23262 12545
rect 22946 12480 22952 12544
rect 23016 12480 23032 12544
rect 23096 12480 23112 12544
rect 23176 12480 23192 12544
rect 23256 12480 23262 12544
rect 22946 12479 23262 12480
rect 25129 12202 25195 12205
rect 26200 12202 27000 12232
rect 25129 12200 27000 12202
rect 25129 12144 25134 12200
rect 25190 12144 27000 12200
rect 25129 12142 27000 12144
rect 25129 12139 25195 12142
rect 26200 12112 27000 12142
rect 7946 12000 8262 12001
rect 7946 11936 7952 12000
rect 8016 11936 8032 12000
rect 8096 11936 8112 12000
rect 8176 11936 8192 12000
rect 8256 11936 8262 12000
rect 7946 11935 8262 11936
rect 17946 12000 18262 12001
rect 17946 11936 17952 12000
rect 18016 11936 18032 12000
rect 18096 11936 18112 12000
rect 18176 11936 18192 12000
rect 18256 11936 18262 12000
rect 17946 11935 18262 11936
rect 2946 11456 3262 11457
rect 0 11386 800 11416
rect 2946 11392 2952 11456
rect 3016 11392 3032 11456
rect 3096 11392 3112 11456
rect 3176 11392 3192 11456
rect 3256 11392 3262 11456
rect 2946 11391 3262 11392
rect 12946 11456 13262 11457
rect 12946 11392 12952 11456
rect 13016 11392 13032 11456
rect 13096 11392 13112 11456
rect 13176 11392 13192 11456
rect 13256 11392 13262 11456
rect 12946 11391 13262 11392
rect 22946 11456 23262 11457
rect 22946 11392 22952 11456
rect 23016 11392 23032 11456
rect 23096 11392 23112 11456
rect 23176 11392 23192 11456
rect 23256 11392 23262 11456
rect 22946 11391 23262 11392
rect 2773 11386 2839 11389
rect 0 11384 2839 11386
rect 0 11328 2778 11384
rect 2834 11328 2839 11384
rect 0 11326 2839 11328
rect 0 11296 800 11326
rect 2773 11323 2839 11326
rect 24761 11386 24827 11389
rect 26200 11386 27000 11416
rect 24761 11384 27000 11386
rect 24761 11328 24766 11384
rect 24822 11328 27000 11384
rect 24761 11326 27000 11328
rect 24761 11323 24827 11326
rect 26200 11296 27000 11326
rect 15878 11188 15884 11252
rect 15948 11250 15954 11252
rect 16021 11250 16087 11253
rect 15948 11248 16087 11250
rect 15948 11192 16026 11248
rect 16082 11192 16087 11248
rect 15948 11190 16087 11192
rect 15948 11188 15954 11190
rect 16021 11187 16087 11190
rect 7946 10912 8262 10913
rect 7946 10848 7952 10912
rect 8016 10848 8032 10912
rect 8096 10848 8112 10912
rect 8176 10848 8192 10912
rect 8256 10848 8262 10912
rect 7946 10847 8262 10848
rect 17946 10912 18262 10913
rect 17946 10848 17952 10912
rect 18016 10848 18032 10912
rect 18096 10848 18112 10912
rect 18176 10848 18192 10912
rect 18256 10848 18262 10912
rect 17946 10847 18262 10848
rect 24669 10570 24735 10573
rect 26200 10570 27000 10600
rect 24669 10568 27000 10570
rect 24669 10512 24674 10568
rect 24730 10512 27000 10568
rect 24669 10510 27000 10512
rect 24669 10507 24735 10510
rect 26200 10480 27000 10510
rect 2946 10368 3262 10369
rect 2946 10304 2952 10368
rect 3016 10304 3032 10368
rect 3096 10304 3112 10368
rect 3176 10304 3192 10368
rect 3256 10304 3262 10368
rect 2946 10303 3262 10304
rect 12946 10368 13262 10369
rect 12946 10304 12952 10368
rect 13016 10304 13032 10368
rect 13096 10304 13112 10368
rect 13176 10304 13192 10368
rect 13256 10304 13262 10368
rect 12946 10303 13262 10304
rect 22946 10368 23262 10369
rect 22946 10304 22952 10368
rect 23016 10304 23032 10368
rect 23096 10304 23112 10368
rect 23176 10304 23192 10368
rect 23256 10304 23262 10368
rect 22946 10303 23262 10304
rect 7946 9824 8262 9825
rect 7946 9760 7952 9824
rect 8016 9760 8032 9824
rect 8096 9760 8112 9824
rect 8176 9760 8192 9824
rect 8256 9760 8262 9824
rect 7946 9759 8262 9760
rect 17946 9824 18262 9825
rect 17946 9760 17952 9824
rect 18016 9760 18032 9824
rect 18096 9760 18112 9824
rect 18176 9760 18192 9824
rect 18256 9760 18262 9824
rect 17946 9759 18262 9760
rect 24945 9754 25011 9757
rect 26200 9754 27000 9784
rect 24945 9752 27000 9754
rect 24945 9696 24950 9752
rect 25006 9696 27000 9752
rect 24945 9694 27000 9696
rect 24945 9691 25011 9694
rect 26200 9664 27000 9694
rect 2946 9280 3262 9281
rect 2946 9216 2952 9280
rect 3016 9216 3032 9280
rect 3096 9216 3112 9280
rect 3176 9216 3192 9280
rect 3256 9216 3262 9280
rect 2946 9215 3262 9216
rect 12946 9280 13262 9281
rect 12946 9216 12952 9280
rect 13016 9216 13032 9280
rect 13096 9216 13112 9280
rect 13176 9216 13192 9280
rect 13256 9216 13262 9280
rect 12946 9215 13262 9216
rect 22946 9280 23262 9281
rect 22946 9216 22952 9280
rect 23016 9216 23032 9280
rect 23096 9216 23112 9280
rect 23176 9216 23192 9280
rect 23256 9216 23262 9280
rect 22946 9215 23262 9216
rect 0 8938 800 8968
rect 2865 8938 2931 8941
rect 0 8936 2931 8938
rect 0 8880 2870 8936
rect 2926 8880 2931 8936
rect 0 8878 2931 8880
rect 0 8848 800 8878
rect 2865 8875 2931 8878
rect 25129 8938 25195 8941
rect 26200 8938 27000 8968
rect 25129 8936 27000 8938
rect 25129 8880 25134 8936
rect 25190 8880 27000 8936
rect 25129 8878 27000 8880
rect 25129 8875 25195 8878
rect 26200 8848 27000 8878
rect 7946 8736 8262 8737
rect 7946 8672 7952 8736
rect 8016 8672 8032 8736
rect 8096 8672 8112 8736
rect 8176 8672 8192 8736
rect 8256 8672 8262 8736
rect 7946 8671 8262 8672
rect 17946 8736 18262 8737
rect 17946 8672 17952 8736
rect 18016 8672 18032 8736
rect 18096 8672 18112 8736
rect 18176 8672 18192 8736
rect 18256 8672 18262 8736
rect 17946 8671 18262 8672
rect 2946 8192 3262 8193
rect 2946 8128 2952 8192
rect 3016 8128 3032 8192
rect 3096 8128 3112 8192
rect 3176 8128 3192 8192
rect 3256 8128 3262 8192
rect 2946 8127 3262 8128
rect 12946 8192 13262 8193
rect 12946 8128 12952 8192
rect 13016 8128 13032 8192
rect 13096 8128 13112 8192
rect 13176 8128 13192 8192
rect 13256 8128 13262 8192
rect 12946 8127 13262 8128
rect 22946 8192 23262 8193
rect 22946 8128 22952 8192
rect 23016 8128 23032 8192
rect 23096 8128 23112 8192
rect 23176 8128 23192 8192
rect 23256 8128 23262 8192
rect 22946 8127 23262 8128
rect 25129 8122 25195 8125
rect 26200 8122 27000 8152
rect 25129 8120 27000 8122
rect 25129 8064 25134 8120
rect 25190 8064 27000 8120
rect 25129 8062 27000 8064
rect 25129 8059 25195 8062
rect 26200 8032 27000 8062
rect 11053 7986 11119 7989
rect 14774 7986 14780 7988
rect 11053 7984 14780 7986
rect 11053 7928 11058 7984
rect 11114 7928 14780 7984
rect 11053 7926 14780 7928
rect 11053 7923 11119 7926
rect 14774 7924 14780 7926
rect 14844 7924 14850 7988
rect 7946 7648 8262 7649
rect 7946 7584 7952 7648
rect 8016 7584 8032 7648
rect 8096 7584 8112 7648
rect 8176 7584 8192 7648
rect 8256 7584 8262 7648
rect 7946 7583 8262 7584
rect 17946 7648 18262 7649
rect 17946 7584 17952 7648
rect 18016 7584 18032 7648
rect 18096 7584 18112 7648
rect 18176 7584 18192 7648
rect 18256 7584 18262 7648
rect 17946 7583 18262 7584
rect 24761 7306 24827 7309
rect 26200 7306 27000 7336
rect 24761 7304 27000 7306
rect 24761 7248 24766 7304
rect 24822 7248 27000 7304
rect 24761 7246 27000 7248
rect 24761 7243 24827 7246
rect 26200 7216 27000 7246
rect 2946 7104 3262 7105
rect 2946 7040 2952 7104
rect 3016 7040 3032 7104
rect 3096 7040 3112 7104
rect 3176 7040 3192 7104
rect 3256 7040 3262 7104
rect 2946 7039 3262 7040
rect 12946 7104 13262 7105
rect 12946 7040 12952 7104
rect 13016 7040 13032 7104
rect 13096 7040 13112 7104
rect 13176 7040 13192 7104
rect 13256 7040 13262 7104
rect 12946 7039 13262 7040
rect 22946 7104 23262 7105
rect 22946 7040 22952 7104
rect 23016 7040 23032 7104
rect 23096 7040 23112 7104
rect 23176 7040 23192 7104
rect 23256 7040 23262 7104
rect 22946 7039 23262 7040
rect 7946 6560 8262 6561
rect 0 6490 800 6520
rect 7946 6496 7952 6560
rect 8016 6496 8032 6560
rect 8096 6496 8112 6560
rect 8176 6496 8192 6560
rect 8256 6496 8262 6560
rect 7946 6495 8262 6496
rect 17946 6560 18262 6561
rect 17946 6496 17952 6560
rect 18016 6496 18032 6560
rect 18096 6496 18112 6560
rect 18176 6496 18192 6560
rect 18256 6496 18262 6560
rect 17946 6495 18262 6496
rect 3049 6490 3115 6493
rect 0 6488 3115 6490
rect 0 6432 3054 6488
rect 3110 6432 3115 6488
rect 0 6430 3115 6432
rect 0 6400 800 6430
rect 3049 6427 3115 6430
rect 25773 6490 25839 6493
rect 26200 6490 27000 6520
rect 25773 6488 27000 6490
rect 25773 6432 25778 6488
rect 25834 6432 27000 6488
rect 25773 6430 27000 6432
rect 25773 6427 25839 6430
rect 26200 6400 27000 6430
rect 2946 6016 3262 6017
rect 2946 5952 2952 6016
rect 3016 5952 3032 6016
rect 3096 5952 3112 6016
rect 3176 5952 3192 6016
rect 3256 5952 3262 6016
rect 2946 5951 3262 5952
rect 12946 6016 13262 6017
rect 12946 5952 12952 6016
rect 13016 5952 13032 6016
rect 13096 5952 13112 6016
rect 13176 5952 13192 6016
rect 13256 5952 13262 6016
rect 12946 5951 13262 5952
rect 22946 6016 23262 6017
rect 22946 5952 22952 6016
rect 23016 5952 23032 6016
rect 23096 5952 23112 6016
rect 23176 5952 23192 6016
rect 23256 5952 23262 6016
rect 22946 5951 23262 5952
rect 24761 5674 24827 5677
rect 26200 5674 27000 5704
rect 24761 5672 27000 5674
rect 24761 5616 24766 5672
rect 24822 5616 27000 5672
rect 24761 5614 27000 5616
rect 24761 5611 24827 5614
rect 26200 5584 27000 5614
rect 7946 5472 8262 5473
rect 7946 5408 7952 5472
rect 8016 5408 8032 5472
rect 8096 5408 8112 5472
rect 8176 5408 8192 5472
rect 8256 5408 8262 5472
rect 7946 5407 8262 5408
rect 17946 5472 18262 5473
rect 17946 5408 17952 5472
rect 18016 5408 18032 5472
rect 18096 5408 18112 5472
rect 18176 5408 18192 5472
rect 18256 5408 18262 5472
rect 17946 5407 18262 5408
rect 2946 4928 3262 4929
rect 2946 4864 2952 4928
rect 3016 4864 3032 4928
rect 3096 4864 3112 4928
rect 3176 4864 3192 4928
rect 3256 4864 3262 4928
rect 2946 4863 3262 4864
rect 12946 4928 13262 4929
rect 12946 4864 12952 4928
rect 13016 4864 13032 4928
rect 13096 4864 13112 4928
rect 13176 4864 13192 4928
rect 13256 4864 13262 4928
rect 12946 4863 13262 4864
rect 22946 4928 23262 4929
rect 22946 4864 22952 4928
rect 23016 4864 23032 4928
rect 23096 4864 23112 4928
rect 23176 4864 23192 4928
rect 23256 4864 23262 4928
rect 22946 4863 23262 4864
rect 23381 4858 23447 4861
rect 26200 4858 27000 4888
rect 23381 4856 27000 4858
rect 23381 4800 23386 4856
rect 23442 4800 27000 4856
rect 23381 4798 27000 4800
rect 23381 4795 23447 4798
rect 26200 4768 27000 4798
rect 7946 4384 8262 4385
rect 7946 4320 7952 4384
rect 8016 4320 8032 4384
rect 8096 4320 8112 4384
rect 8176 4320 8192 4384
rect 8256 4320 8262 4384
rect 7946 4319 8262 4320
rect 17946 4384 18262 4385
rect 17946 4320 17952 4384
rect 18016 4320 18032 4384
rect 18096 4320 18112 4384
rect 18176 4320 18192 4384
rect 18256 4320 18262 4384
rect 17946 4319 18262 4320
rect 8477 4178 8543 4181
rect 10174 4178 10180 4180
rect 8477 4176 10180 4178
rect 8477 4120 8482 4176
rect 8538 4120 10180 4176
rect 8477 4118 10180 4120
rect 8477 4115 8543 4118
rect 10174 4116 10180 4118
rect 10244 4116 10250 4180
rect 0 4042 800 4072
rect 2865 4042 2931 4045
rect 0 4040 2931 4042
rect 0 3984 2870 4040
rect 2926 3984 2931 4040
rect 0 3982 2931 3984
rect 0 3952 800 3982
rect 2865 3979 2931 3982
rect 22093 4042 22159 4045
rect 26200 4042 27000 4072
rect 22093 4040 27000 4042
rect 22093 3984 22098 4040
rect 22154 3984 27000 4040
rect 22093 3982 27000 3984
rect 22093 3979 22159 3982
rect 26200 3952 27000 3982
rect 2946 3840 3262 3841
rect 2946 3776 2952 3840
rect 3016 3776 3032 3840
rect 3096 3776 3112 3840
rect 3176 3776 3192 3840
rect 3256 3776 3262 3840
rect 2946 3775 3262 3776
rect 12946 3840 13262 3841
rect 12946 3776 12952 3840
rect 13016 3776 13032 3840
rect 13096 3776 13112 3840
rect 13176 3776 13192 3840
rect 13256 3776 13262 3840
rect 12946 3775 13262 3776
rect 22946 3840 23262 3841
rect 22946 3776 22952 3840
rect 23016 3776 23032 3840
rect 23096 3776 23112 3840
rect 23176 3776 23192 3840
rect 23256 3776 23262 3840
rect 22946 3775 23262 3776
rect 16798 3436 16804 3500
rect 16868 3498 16874 3500
rect 23749 3498 23815 3501
rect 16868 3496 23815 3498
rect 16868 3440 23754 3496
rect 23810 3440 23815 3496
rect 16868 3438 23815 3440
rect 16868 3436 16874 3438
rect 23749 3435 23815 3438
rect 7946 3296 8262 3297
rect 7946 3232 7952 3296
rect 8016 3232 8032 3296
rect 8096 3232 8112 3296
rect 8176 3232 8192 3296
rect 8256 3232 8262 3296
rect 7946 3231 8262 3232
rect 17946 3296 18262 3297
rect 17946 3232 17952 3296
rect 18016 3232 18032 3296
rect 18096 3232 18112 3296
rect 18176 3232 18192 3296
rect 18256 3232 18262 3296
rect 17946 3231 18262 3232
rect 11881 3226 11947 3229
rect 12014 3226 12020 3228
rect 11881 3224 12020 3226
rect 11881 3168 11886 3224
rect 11942 3168 12020 3224
rect 11881 3166 12020 3168
rect 11881 3163 11947 3166
rect 12014 3164 12020 3166
rect 12084 3164 12090 3228
rect 22737 3226 22803 3229
rect 26200 3226 27000 3256
rect 22737 3224 27000 3226
rect 22737 3168 22742 3224
rect 22798 3168 27000 3224
rect 22737 3166 27000 3168
rect 22737 3163 22803 3166
rect 26200 3136 27000 3166
rect 2946 2752 3262 2753
rect 2946 2688 2952 2752
rect 3016 2688 3032 2752
rect 3096 2688 3112 2752
rect 3176 2688 3192 2752
rect 3256 2688 3262 2752
rect 2946 2687 3262 2688
rect 12946 2752 13262 2753
rect 12946 2688 12952 2752
rect 13016 2688 13032 2752
rect 13096 2688 13112 2752
rect 13176 2688 13192 2752
rect 13256 2688 13262 2752
rect 12946 2687 13262 2688
rect 22946 2752 23262 2753
rect 22946 2688 22952 2752
rect 23016 2688 23032 2752
rect 23096 2688 23112 2752
rect 23176 2688 23192 2752
rect 23256 2688 23262 2752
rect 22946 2687 23262 2688
rect 21633 2410 21699 2413
rect 26200 2410 27000 2440
rect 21633 2408 27000 2410
rect 21633 2352 21638 2408
rect 21694 2352 27000 2408
rect 21633 2350 27000 2352
rect 21633 2347 21699 2350
rect 26200 2320 27000 2350
rect 7946 2208 8262 2209
rect 7946 2144 7952 2208
rect 8016 2144 8032 2208
rect 8096 2144 8112 2208
rect 8176 2144 8192 2208
rect 8256 2144 8262 2208
rect 7946 2143 8262 2144
rect 17946 2208 18262 2209
rect 17946 2144 17952 2208
rect 18016 2144 18032 2208
rect 18096 2144 18112 2208
rect 18176 2144 18192 2208
rect 18256 2144 18262 2208
rect 17946 2143 18262 2144
rect 0 1594 800 1624
rect 2865 1594 2931 1597
rect 0 1592 2931 1594
rect 0 1536 2870 1592
rect 2926 1536 2931 1592
rect 0 1534 2931 1536
rect 0 1504 800 1534
rect 2865 1531 2931 1534
rect 25313 1594 25379 1597
rect 26200 1594 27000 1624
rect 25313 1592 27000 1594
rect 25313 1536 25318 1592
rect 25374 1536 27000 1592
rect 25313 1534 27000 1536
rect 25313 1531 25379 1534
rect 26200 1504 27000 1534
rect 24945 778 25011 781
rect 26200 778 27000 808
rect 24945 776 27000 778
rect 24945 720 24950 776
rect 25006 720 27000 776
rect 24945 718 27000 720
rect 24945 715 25011 718
rect 26200 688 27000 718
<< via3 >>
rect 7952 54428 8016 54432
rect 7952 54372 7956 54428
rect 7956 54372 8012 54428
rect 8012 54372 8016 54428
rect 7952 54368 8016 54372
rect 8032 54428 8096 54432
rect 8032 54372 8036 54428
rect 8036 54372 8092 54428
rect 8092 54372 8096 54428
rect 8032 54368 8096 54372
rect 8112 54428 8176 54432
rect 8112 54372 8116 54428
rect 8116 54372 8172 54428
rect 8172 54372 8176 54428
rect 8112 54368 8176 54372
rect 8192 54428 8256 54432
rect 8192 54372 8196 54428
rect 8196 54372 8252 54428
rect 8252 54372 8256 54428
rect 8192 54368 8256 54372
rect 17952 54428 18016 54432
rect 17952 54372 17956 54428
rect 17956 54372 18012 54428
rect 18012 54372 18016 54428
rect 17952 54368 18016 54372
rect 18032 54428 18096 54432
rect 18032 54372 18036 54428
rect 18036 54372 18092 54428
rect 18092 54372 18096 54428
rect 18032 54368 18096 54372
rect 18112 54428 18176 54432
rect 18112 54372 18116 54428
rect 18116 54372 18172 54428
rect 18172 54372 18176 54428
rect 18112 54368 18176 54372
rect 18192 54428 18256 54432
rect 18192 54372 18196 54428
rect 18196 54372 18252 54428
rect 18252 54372 18256 54428
rect 18192 54368 18256 54372
rect 15884 53892 15948 53956
rect 22324 53952 22388 53956
rect 22324 53896 22374 53952
rect 22374 53896 22388 53952
rect 22324 53892 22388 53896
rect 2952 53884 3016 53888
rect 2952 53828 2956 53884
rect 2956 53828 3012 53884
rect 3012 53828 3016 53884
rect 2952 53824 3016 53828
rect 3032 53884 3096 53888
rect 3032 53828 3036 53884
rect 3036 53828 3092 53884
rect 3092 53828 3096 53884
rect 3032 53824 3096 53828
rect 3112 53884 3176 53888
rect 3112 53828 3116 53884
rect 3116 53828 3172 53884
rect 3172 53828 3176 53884
rect 3112 53824 3176 53828
rect 3192 53884 3256 53888
rect 3192 53828 3196 53884
rect 3196 53828 3252 53884
rect 3252 53828 3256 53884
rect 3192 53824 3256 53828
rect 12952 53884 13016 53888
rect 12952 53828 12956 53884
rect 12956 53828 13012 53884
rect 13012 53828 13016 53884
rect 12952 53824 13016 53828
rect 13032 53884 13096 53888
rect 13032 53828 13036 53884
rect 13036 53828 13092 53884
rect 13092 53828 13096 53884
rect 13032 53824 13096 53828
rect 13112 53884 13176 53888
rect 13112 53828 13116 53884
rect 13116 53828 13172 53884
rect 13172 53828 13176 53884
rect 13112 53824 13176 53828
rect 13192 53884 13256 53888
rect 13192 53828 13196 53884
rect 13196 53828 13252 53884
rect 13252 53828 13256 53884
rect 13192 53824 13256 53828
rect 22952 53884 23016 53888
rect 22952 53828 22956 53884
rect 22956 53828 23012 53884
rect 23012 53828 23016 53884
rect 22952 53824 23016 53828
rect 23032 53884 23096 53888
rect 23032 53828 23036 53884
rect 23036 53828 23092 53884
rect 23092 53828 23096 53884
rect 23032 53824 23096 53828
rect 23112 53884 23176 53888
rect 23112 53828 23116 53884
rect 23116 53828 23172 53884
rect 23172 53828 23176 53884
rect 23112 53824 23176 53828
rect 23192 53884 23256 53888
rect 23192 53828 23196 53884
rect 23196 53828 23252 53884
rect 23252 53828 23256 53884
rect 23192 53824 23256 53828
rect 7952 53340 8016 53344
rect 7952 53284 7956 53340
rect 7956 53284 8012 53340
rect 8012 53284 8016 53340
rect 7952 53280 8016 53284
rect 8032 53340 8096 53344
rect 8032 53284 8036 53340
rect 8036 53284 8092 53340
rect 8092 53284 8096 53340
rect 8032 53280 8096 53284
rect 8112 53340 8176 53344
rect 8112 53284 8116 53340
rect 8116 53284 8172 53340
rect 8172 53284 8176 53340
rect 8112 53280 8176 53284
rect 8192 53340 8256 53344
rect 8192 53284 8196 53340
rect 8196 53284 8252 53340
rect 8252 53284 8256 53340
rect 8192 53280 8256 53284
rect 17952 53340 18016 53344
rect 17952 53284 17956 53340
rect 17956 53284 18012 53340
rect 18012 53284 18016 53340
rect 17952 53280 18016 53284
rect 18032 53340 18096 53344
rect 18032 53284 18036 53340
rect 18036 53284 18092 53340
rect 18092 53284 18096 53340
rect 18032 53280 18096 53284
rect 18112 53340 18176 53344
rect 18112 53284 18116 53340
rect 18116 53284 18172 53340
rect 18172 53284 18176 53340
rect 18112 53280 18176 53284
rect 18192 53340 18256 53344
rect 18192 53284 18196 53340
rect 18196 53284 18252 53340
rect 18252 53284 18256 53340
rect 18192 53280 18256 53284
rect 22508 53212 22572 53276
rect 21036 52940 21100 53004
rect 2952 52796 3016 52800
rect 2952 52740 2956 52796
rect 2956 52740 3012 52796
rect 3012 52740 3016 52796
rect 2952 52736 3016 52740
rect 3032 52796 3096 52800
rect 3032 52740 3036 52796
rect 3036 52740 3092 52796
rect 3092 52740 3096 52796
rect 3032 52736 3096 52740
rect 3112 52796 3176 52800
rect 3112 52740 3116 52796
rect 3116 52740 3172 52796
rect 3172 52740 3176 52796
rect 3112 52736 3176 52740
rect 3192 52796 3256 52800
rect 3192 52740 3196 52796
rect 3196 52740 3252 52796
rect 3252 52740 3256 52796
rect 3192 52736 3256 52740
rect 12952 52796 13016 52800
rect 12952 52740 12956 52796
rect 12956 52740 13012 52796
rect 13012 52740 13016 52796
rect 12952 52736 13016 52740
rect 13032 52796 13096 52800
rect 13032 52740 13036 52796
rect 13036 52740 13092 52796
rect 13092 52740 13096 52796
rect 13032 52736 13096 52740
rect 13112 52796 13176 52800
rect 13112 52740 13116 52796
rect 13116 52740 13172 52796
rect 13172 52740 13176 52796
rect 13112 52736 13176 52740
rect 13192 52796 13256 52800
rect 13192 52740 13196 52796
rect 13196 52740 13252 52796
rect 13252 52740 13256 52796
rect 13192 52736 13256 52740
rect 22952 52796 23016 52800
rect 22952 52740 22956 52796
rect 22956 52740 23012 52796
rect 23012 52740 23016 52796
rect 22952 52736 23016 52740
rect 23032 52796 23096 52800
rect 23032 52740 23036 52796
rect 23036 52740 23092 52796
rect 23092 52740 23096 52796
rect 23032 52736 23096 52740
rect 23112 52796 23176 52800
rect 23112 52740 23116 52796
rect 23116 52740 23172 52796
rect 23172 52740 23176 52796
rect 23112 52736 23176 52740
rect 23192 52796 23256 52800
rect 23192 52740 23196 52796
rect 23196 52740 23252 52796
rect 23252 52740 23256 52796
rect 23192 52736 23256 52740
rect 13860 52532 13924 52596
rect 14044 52592 14108 52596
rect 14044 52536 14058 52592
rect 14058 52536 14108 52592
rect 14044 52532 14108 52536
rect 15332 52532 15396 52596
rect 17724 52532 17788 52596
rect 7952 52252 8016 52256
rect 7952 52196 7956 52252
rect 7956 52196 8012 52252
rect 8012 52196 8016 52252
rect 7952 52192 8016 52196
rect 8032 52252 8096 52256
rect 8032 52196 8036 52252
rect 8036 52196 8092 52252
rect 8092 52196 8096 52252
rect 8032 52192 8096 52196
rect 8112 52252 8176 52256
rect 8112 52196 8116 52252
rect 8116 52196 8172 52252
rect 8172 52196 8176 52252
rect 8112 52192 8176 52196
rect 8192 52252 8256 52256
rect 8192 52196 8196 52252
rect 8196 52196 8252 52252
rect 8252 52196 8256 52252
rect 8192 52192 8256 52196
rect 17952 52252 18016 52256
rect 17952 52196 17956 52252
rect 17956 52196 18012 52252
rect 18012 52196 18016 52252
rect 17952 52192 18016 52196
rect 18032 52252 18096 52256
rect 18032 52196 18036 52252
rect 18036 52196 18092 52252
rect 18092 52196 18096 52252
rect 18032 52192 18096 52196
rect 18112 52252 18176 52256
rect 18112 52196 18116 52252
rect 18116 52196 18172 52252
rect 18172 52196 18176 52252
rect 18112 52192 18176 52196
rect 18192 52252 18256 52256
rect 18192 52196 18196 52252
rect 18196 52196 18252 52252
rect 18252 52196 18256 52252
rect 18192 52192 18256 52196
rect 2952 51708 3016 51712
rect 2952 51652 2956 51708
rect 2956 51652 3012 51708
rect 3012 51652 3016 51708
rect 2952 51648 3016 51652
rect 3032 51708 3096 51712
rect 3032 51652 3036 51708
rect 3036 51652 3092 51708
rect 3092 51652 3096 51708
rect 3032 51648 3096 51652
rect 3112 51708 3176 51712
rect 3112 51652 3116 51708
rect 3116 51652 3172 51708
rect 3172 51652 3176 51708
rect 3112 51648 3176 51652
rect 3192 51708 3256 51712
rect 3192 51652 3196 51708
rect 3196 51652 3252 51708
rect 3252 51652 3256 51708
rect 3192 51648 3256 51652
rect 12952 51708 13016 51712
rect 12952 51652 12956 51708
rect 12956 51652 13012 51708
rect 13012 51652 13016 51708
rect 12952 51648 13016 51652
rect 13032 51708 13096 51712
rect 13032 51652 13036 51708
rect 13036 51652 13092 51708
rect 13092 51652 13096 51708
rect 13032 51648 13096 51652
rect 13112 51708 13176 51712
rect 13112 51652 13116 51708
rect 13116 51652 13172 51708
rect 13172 51652 13176 51708
rect 13112 51648 13176 51652
rect 13192 51708 13256 51712
rect 13192 51652 13196 51708
rect 13196 51652 13252 51708
rect 13252 51652 13256 51708
rect 13192 51648 13256 51652
rect 22952 51708 23016 51712
rect 22952 51652 22956 51708
rect 22956 51652 23012 51708
rect 23012 51652 23016 51708
rect 22952 51648 23016 51652
rect 23032 51708 23096 51712
rect 23032 51652 23036 51708
rect 23036 51652 23092 51708
rect 23092 51652 23096 51708
rect 23032 51648 23096 51652
rect 23112 51708 23176 51712
rect 23112 51652 23116 51708
rect 23116 51652 23172 51708
rect 23172 51652 23176 51708
rect 23112 51648 23176 51652
rect 23192 51708 23256 51712
rect 23192 51652 23196 51708
rect 23196 51652 23252 51708
rect 23252 51652 23256 51708
rect 23192 51648 23256 51652
rect 7952 51164 8016 51168
rect 7952 51108 7956 51164
rect 7956 51108 8012 51164
rect 8012 51108 8016 51164
rect 7952 51104 8016 51108
rect 8032 51164 8096 51168
rect 8032 51108 8036 51164
rect 8036 51108 8092 51164
rect 8092 51108 8096 51164
rect 8032 51104 8096 51108
rect 8112 51164 8176 51168
rect 8112 51108 8116 51164
rect 8116 51108 8172 51164
rect 8172 51108 8176 51164
rect 8112 51104 8176 51108
rect 8192 51164 8256 51168
rect 8192 51108 8196 51164
rect 8196 51108 8252 51164
rect 8252 51108 8256 51164
rect 8192 51104 8256 51108
rect 17952 51164 18016 51168
rect 17952 51108 17956 51164
rect 17956 51108 18012 51164
rect 18012 51108 18016 51164
rect 17952 51104 18016 51108
rect 18032 51164 18096 51168
rect 18032 51108 18036 51164
rect 18036 51108 18092 51164
rect 18092 51108 18096 51164
rect 18032 51104 18096 51108
rect 18112 51164 18176 51168
rect 18112 51108 18116 51164
rect 18116 51108 18172 51164
rect 18172 51108 18176 51164
rect 18112 51104 18176 51108
rect 18192 51164 18256 51168
rect 18192 51108 18196 51164
rect 18196 51108 18252 51164
rect 18252 51108 18256 51164
rect 18192 51104 18256 51108
rect 2952 50620 3016 50624
rect 2952 50564 2956 50620
rect 2956 50564 3012 50620
rect 3012 50564 3016 50620
rect 2952 50560 3016 50564
rect 3032 50620 3096 50624
rect 3032 50564 3036 50620
rect 3036 50564 3092 50620
rect 3092 50564 3096 50620
rect 3032 50560 3096 50564
rect 3112 50620 3176 50624
rect 3112 50564 3116 50620
rect 3116 50564 3172 50620
rect 3172 50564 3176 50620
rect 3112 50560 3176 50564
rect 3192 50620 3256 50624
rect 3192 50564 3196 50620
rect 3196 50564 3252 50620
rect 3252 50564 3256 50620
rect 3192 50560 3256 50564
rect 12952 50620 13016 50624
rect 12952 50564 12956 50620
rect 12956 50564 13012 50620
rect 13012 50564 13016 50620
rect 12952 50560 13016 50564
rect 13032 50620 13096 50624
rect 13032 50564 13036 50620
rect 13036 50564 13092 50620
rect 13092 50564 13096 50620
rect 13032 50560 13096 50564
rect 13112 50620 13176 50624
rect 13112 50564 13116 50620
rect 13116 50564 13172 50620
rect 13172 50564 13176 50620
rect 13112 50560 13176 50564
rect 13192 50620 13256 50624
rect 13192 50564 13196 50620
rect 13196 50564 13252 50620
rect 13252 50564 13256 50620
rect 13192 50560 13256 50564
rect 22952 50620 23016 50624
rect 22952 50564 22956 50620
rect 22956 50564 23012 50620
rect 23012 50564 23016 50620
rect 22952 50560 23016 50564
rect 23032 50620 23096 50624
rect 23032 50564 23036 50620
rect 23036 50564 23092 50620
rect 23092 50564 23096 50620
rect 23032 50560 23096 50564
rect 23112 50620 23176 50624
rect 23112 50564 23116 50620
rect 23116 50564 23172 50620
rect 23172 50564 23176 50620
rect 23112 50560 23176 50564
rect 23192 50620 23256 50624
rect 23192 50564 23196 50620
rect 23196 50564 23252 50620
rect 23252 50564 23256 50620
rect 23192 50560 23256 50564
rect 7952 50076 8016 50080
rect 7952 50020 7956 50076
rect 7956 50020 8012 50076
rect 8012 50020 8016 50076
rect 7952 50016 8016 50020
rect 8032 50076 8096 50080
rect 8032 50020 8036 50076
rect 8036 50020 8092 50076
rect 8092 50020 8096 50076
rect 8032 50016 8096 50020
rect 8112 50076 8176 50080
rect 8112 50020 8116 50076
rect 8116 50020 8172 50076
rect 8172 50020 8176 50076
rect 8112 50016 8176 50020
rect 8192 50076 8256 50080
rect 8192 50020 8196 50076
rect 8196 50020 8252 50076
rect 8252 50020 8256 50076
rect 8192 50016 8256 50020
rect 17952 50076 18016 50080
rect 17952 50020 17956 50076
rect 17956 50020 18012 50076
rect 18012 50020 18016 50076
rect 17952 50016 18016 50020
rect 18032 50076 18096 50080
rect 18032 50020 18036 50076
rect 18036 50020 18092 50076
rect 18092 50020 18096 50076
rect 18032 50016 18096 50020
rect 18112 50076 18176 50080
rect 18112 50020 18116 50076
rect 18116 50020 18172 50076
rect 18172 50020 18176 50076
rect 18112 50016 18176 50020
rect 18192 50076 18256 50080
rect 18192 50020 18196 50076
rect 18196 50020 18252 50076
rect 18252 50020 18256 50076
rect 18192 50016 18256 50020
rect 2952 49532 3016 49536
rect 2952 49476 2956 49532
rect 2956 49476 3012 49532
rect 3012 49476 3016 49532
rect 2952 49472 3016 49476
rect 3032 49532 3096 49536
rect 3032 49476 3036 49532
rect 3036 49476 3092 49532
rect 3092 49476 3096 49532
rect 3032 49472 3096 49476
rect 3112 49532 3176 49536
rect 3112 49476 3116 49532
rect 3116 49476 3172 49532
rect 3172 49476 3176 49532
rect 3112 49472 3176 49476
rect 3192 49532 3256 49536
rect 3192 49476 3196 49532
rect 3196 49476 3252 49532
rect 3252 49476 3256 49532
rect 3192 49472 3256 49476
rect 12952 49532 13016 49536
rect 12952 49476 12956 49532
rect 12956 49476 13012 49532
rect 13012 49476 13016 49532
rect 12952 49472 13016 49476
rect 13032 49532 13096 49536
rect 13032 49476 13036 49532
rect 13036 49476 13092 49532
rect 13092 49476 13096 49532
rect 13032 49472 13096 49476
rect 13112 49532 13176 49536
rect 13112 49476 13116 49532
rect 13116 49476 13172 49532
rect 13172 49476 13176 49532
rect 13112 49472 13176 49476
rect 13192 49532 13256 49536
rect 13192 49476 13196 49532
rect 13196 49476 13252 49532
rect 13252 49476 13256 49532
rect 13192 49472 13256 49476
rect 22952 49532 23016 49536
rect 22952 49476 22956 49532
rect 22956 49476 23012 49532
rect 23012 49476 23016 49532
rect 22952 49472 23016 49476
rect 23032 49532 23096 49536
rect 23032 49476 23036 49532
rect 23036 49476 23092 49532
rect 23092 49476 23096 49532
rect 23032 49472 23096 49476
rect 23112 49532 23176 49536
rect 23112 49476 23116 49532
rect 23116 49476 23172 49532
rect 23172 49476 23176 49532
rect 23112 49472 23176 49476
rect 23192 49532 23256 49536
rect 23192 49476 23196 49532
rect 23196 49476 23252 49532
rect 23252 49476 23256 49532
rect 23192 49472 23256 49476
rect 7952 48988 8016 48992
rect 7952 48932 7956 48988
rect 7956 48932 8012 48988
rect 8012 48932 8016 48988
rect 7952 48928 8016 48932
rect 8032 48988 8096 48992
rect 8032 48932 8036 48988
rect 8036 48932 8092 48988
rect 8092 48932 8096 48988
rect 8032 48928 8096 48932
rect 8112 48988 8176 48992
rect 8112 48932 8116 48988
rect 8116 48932 8172 48988
rect 8172 48932 8176 48988
rect 8112 48928 8176 48932
rect 8192 48988 8256 48992
rect 8192 48932 8196 48988
rect 8196 48932 8252 48988
rect 8252 48932 8256 48988
rect 8192 48928 8256 48932
rect 17952 48988 18016 48992
rect 17952 48932 17956 48988
rect 17956 48932 18012 48988
rect 18012 48932 18016 48988
rect 17952 48928 18016 48932
rect 18032 48988 18096 48992
rect 18032 48932 18036 48988
rect 18036 48932 18092 48988
rect 18092 48932 18096 48988
rect 18032 48928 18096 48932
rect 18112 48988 18176 48992
rect 18112 48932 18116 48988
rect 18116 48932 18172 48988
rect 18172 48932 18176 48988
rect 18112 48928 18176 48932
rect 18192 48988 18256 48992
rect 18192 48932 18196 48988
rect 18196 48932 18252 48988
rect 18252 48932 18256 48988
rect 18192 48928 18256 48932
rect 2952 48444 3016 48448
rect 2952 48388 2956 48444
rect 2956 48388 3012 48444
rect 3012 48388 3016 48444
rect 2952 48384 3016 48388
rect 3032 48444 3096 48448
rect 3032 48388 3036 48444
rect 3036 48388 3092 48444
rect 3092 48388 3096 48444
rect 3032 48384 3096 48388
rect 3112 48444 3176 48448
rect 3112 48388 3116 48444
rect 3116 48388 3172 48444
rect 3172 48388 3176 48444
rect 3112 48384 3176 48388
rect 3192 48444 3256 48448
rect 3192 48388 3196 48444
rect 3196 48388 3252 48444
rect 3252 48388 3256 48444
rect 3192 48384 3256 48388
rect 12952 48444 13016 48448
rect 12952 48388 12956 48444
rect 12956 48388 13012 48444
rect 13012 48388 13016 48444
rect 12952 48384 13016 48388
rect 13032 48444 13096 48448
rect 13032 48388 13036 48444
rect 13036 48388 13092 48444
rect 13092 48388 13096 48444
rect 13032 48384 13096 48388
rect 13112 48444 13176 48448
rect 13112 48388 13116 48444
rect 13116 48388 13172 48444
rect 13172 48388 13176 48444
rect 13112 48384 13176 48388
rect 13192 48444 13256 48448
rect 13192 48388 13196 48444
rect 13196 48388 13252 48444
rect 13252 48388 13256 48444
rect 13192 48384 13256 48388
rect 22952 48444 23016 48448
rect 22952 48388 22956 48444
rect 22956 48388 23012 48444
rect 23012 48388 23016 48444
rect 22952 48384 23016 48388
rect 23032 48444 23096 48448
rect 23032 48388 23036 48444
rect 23036 48388 23092 48444
rect 23092 48388 23096 48444
rect 23032 48384 23096 48388
rect 23112 48444 23176 48448
rect 23112 48388 23116 48444
rect 23116 48388 23172 48444
rect 23172 48388 23176 48444
rect 23112 48384 23176 48388
rect 23192 48444 23256 48448
rect 23192 48388 23196 48444
rect 23196 48388 23252 48444
rect 23252 48388 23256 48444
rect 23192 48384 23256 48388
rect 7952 47900 8016 47904
rect 7952 47844 7956 47900
rect 7956 47844 8012 47900
rect 8012 47844 8016 47900
rect 7952 47840 8016 47844
rect 8032 47900 8096 47904
rect 8032 47844 8036 47900
rect 8036 47844 8092 47900
rect 8092 47844 8096 47900
rect 8032 47840 8096 47844
rect 8112 47900 8176 47904
rect 8112 47844 8116 47900
rect 8116 47844 8172 47900
rect 8172 47844 8176 47900
rect 8112 47840 8176 47844
rect 8192 47900 8256 47904
rect 8192 47844 8196 47900
rect 8196 47844 8252 47900
rect 8252 47844 8256 47900
rect 8192 47840 8256 47844
rect 17952 47900 18016 47904
rect 17952 47844 17956 47900
rect 17956 47844 18012 47900
rect 18012 47844 18016 47900
rect 17952 47840 18016 47844
rect 18032 47900 18096 47904
rect 18032 47844 18036 47900
rect 18036 47844 18092 47900
rect 18092 47844 18096 47900
rect 18032 47840 18096 47844
rect 18112 47900 18176 47904
rect 18112 47844 18116 47900
rect 18116 47844 18172 47900
rect 18172 47844 18176 47900
rect 18112 47840 18176 47844
rect 18192 47900 18256 47904
rect 18192 47844 18196 47900
rect 18196 47844 18252 47900
rect 18252 47844 18256 47900
rect 18192 47840 18256 47844
rect 2952 47356 3016 47360
rect 2952 47300 2956 47356
rect 2956 47300 3012 47356
rect 3012 47300 3016 47356
rect 2952 47296 3016 47300
rect 3032 47356 3096 47360
rect 3032 47300 3036 47356
rect 3036 47300 3092 47356
rect 3092 47300 3096 47356
rect 3032 47296 3096 47300
rect 3112 47356 3176 47360
rect 3112 47300 3116 47356
rect 3116 47300 3172 47356
rect 3172 47300 3176 47356
rect 3112 47296 3176 47300
rect 3192 47356 3256 47360
rect 3192 47300 3196 47356
rect 3196 47300 3252 47356
rect 3252 47300 3256 47356
rect 3192 47296 3256 47300
rect 12952 47356 13016 47360
rect 12952 47300 12956 47356
rect 12956 47300 13012 47356
rect 13012 47300 13016 47356
rect 12952 47296 13016 47300
rect 13032 47356 13096 47360
rect 13032 47300 13036 47356
rect 13036 47300 13092 47356
rect 13092 47300 13096 47356
rect 13032 47296 13096 47300
rect 13112 47356 13176 47360
rect 13112 47300 13116 47356
rect 13116 47300 13172 47356
rect 13172 47300 13176 47356
rect 13112 47296 13176 47300
rect 13192 47356 13256 47360
rect 13192 47300 13196 47356
rect 13196 47300 13252 47356
rect 13252 47300 13256 47356
rect 13192 47296 13256 47300
rect 22952 47356 23016 47360
rect 22952 47300 22956 47356
rect 22956 47300 23012 47356
rect 23012 47300 23016 47356
rect 22952 47296 23016 47300
rect 23032 47356 23096 47360
rect 23032 47300 23036 47356
rect 23036 47300 23092 47356
rect 23092 47300 23096 47356
rect 23032 47296 23096 47300
rect 23112 47356 23176 47360
rect 23112 47300 23116 47356
rect 23116 47300 23172 47356
rect 23172 47300 23176 47356
rect 23112 47296 23176 47300
rect 23192 47356 23256 47360
rect 23192 47300 23196 47356
rect 23196 47300 23252 47356
rect 23252 47300 23256 47356
rect 23192 47296 23256 47300
rect 19196 46956 19260 47020
rect 7952 46812 8016 46816
rect 7952 46756 7956 46812
rect 7956 46756 8012 46812
rect 8012 46756 8016 46812
rect 7952 46752 8016 46756
rect 8032 46812 8096 46816
rect 8032 46756 8036 46812
rect 8036 46756 8092 46812
rect 8092 46756 8096 46812
rect 8032 46752 8096 46756
rect 8112 46812 8176 46816
rect 8112 46756 8116 46812
rect 8116 46756 8172 46812
rect 8172 46756 8176 46812
rect 8112 46752 8176 46756
rect 8192 46812 8256 46816
rect 8192 46756 8196 46812
rect 8196 46756 8252 46812
rect 8252 46756 8256 46812
rect 8192 46752 8256 46756
rect 17952 46812 18016 46816
rect 17952 46756 17956 46812
rect 17956 46756 18012 46812
rect 18012 46756 18016 46812
rect 17952 46752 18016 46756
rect 18032 46812 18096 46816
rect 18032 46756 18036 46812
rect 18036 46756 18092 46812
rect 18092 46756 18096 46812
rect 18032 46752 18096 46756
rect 18112 46812 18176 46816
rect 18112 46756 18116 46812
rect 18116 46756 18172 46812
rect 18172 46756 18176 46812
rect 18112 46752 18176 46756
rect 18192 46812 18256 46816
rect 18192 46756 18196 46812
rect 18196 46756 18252 46812
rect 18252 46756 18256 46812
rect 18192 46752 18256 46756
rect 20116 46684 20180 46748
rect 19932 46548 19996 46612
rect 2952 46268 3016 46272
rect 2952 46212 2956 46268
rect 2956 46212 3012 46268
rect 3012 46212 3016 46268
rect 2952 46208 3016 46212
rect 3032 46268 3096 46272
rect 3032 46212 3036 46268
rect 3036 46212 3092 46268
rect 3092 46212 3096 46268
rect 3032 46208 3096 46212
rect 3112 46268 3176 46272
rect 3112 46212 3116 46268
rect 3116 46212 3172 46268
rect 3172 46212 3176 46268
rect 3112 46208 3176 46212
rect 3192 46268 3256 46272
rect 3192 46212 3196 46268
rect 3196 46212 3252 46268
rect 3252 46212 3256 46268
rect 3192 46208 3256 46212
rect 12952 46268 13016 46272
rect 12952 46212 12956 46268
rect 12956 46212 13012 46268
rect 13012 46212 13016 46268
rect 12952 46208 13016 46212
rect 13032 46268 13096 46272
rect 13032 46212 13036 46268
rect 13036 46212 13092 46268
rect 13092 46212 13096 46268
rect 13032 46208 13096 46212
rect 13112 46268 13176 46272
rect 13112 46212 13116 46268
rect 13116 46212 13172 46268
rect 13172 46212 13176 46268
rect 13112 46208 13176 46212
rect 13192 46268 13256 46272
rect 13192 46212 13196 46268
rect 13196 46212 13252 46268
rect 13252 46212 13256 46268
rect 13192 46208 13256 46212
rect 22952 46268 23016 46272
rect 22952 46212 22956 46268
rect 22956 46212 23012 46268
rect 23012 46212 23016 46268
rect 22952 46208 23016 46212
rect 23032 46268 23096 46272
rect 23032 46212 23036 46268
rect 23036 46212 23092 46268
rect 23092 46212 23096 46268
rect 23032 46208 23096 46212
rect 23112 46268 23176 46272
rect 23112 46212 23116 46268
rect 23116 46212 23172 46268
rect 23172 46212 23176 46268
rect 23112 46208 23176 46212
rect 23192 46268 23256 46272
rect 23192 46212 23196 46268
rect 23196 46212 23252 46268
rect 23252 46212 23256 46268
rect 23192 46208 23256 46212
rect 21956 45928 22020 45932
rect 21956 45872 22006 45928
rect 22006 45872 22020 45928
rect 21956 45868 22020 45872
rect 7952 45724 8016 45728
rect 7952 45668 7956 45724
rect 7956 45668 8012 45724
rect 8012 45668 8016 45724
rect 7952 45664 8016 45668
rect 8032 45724 8096 45728
rect 8032 45668 8036 45724
rect 8036 45668 8092 45724
rect 8092 45668 8096 45724
rect 8032 45664 8096 45668
rect 8112 45724 8176 45728
rect 8112 45668 8116 45724
rect 8116 45668 8172 45724
rect 8172 45668 8176 45724
rect 8112 45664 8176 45668
rect 8192 45724 8256 45728
rect 8192 45668 8196 45724
rect 8196 45668 8252 45724
rect 8252 45668 8256 45724
rect 8192 45664 8256 45668
rect 17952 45724 18016 45728
rect 17952 45668 17956 45724
rect 17956 45668 18012 45724
rect 18012 45668 18016 45724
rect 17952 45664 18016 45668
rect 18032 45724 18096 45728
rect 18032 45668 18036 45724
rect 18036 45668 18092 45724
rect 18092 45668 18096 45724
rect 18032 45664 18096 45668
rect 18112 45724 18176 45728
rect 18112 45668 18116 45724
rect 18116 45668 18172 45724
rect 18172 45668 18176 45724
rect 18112 45664 18176 45668
rect 18192 45724 18256 45728
rect 18192 45668 18196 45724
rect 18196 45668 18252 45724
rect 18252 45668 18256 45724
rect 18192 45664 18256 45668
rect 24716 45656 24780 45660
rect 24716 45600 24766 45656
rect 24766 45600 24780 45656
rect 24716 45596 24780 45600
rect 11284 45324 11348 45388
rect 2952 45180 3016 45184
rect 2952 45124 2956 45180
rect 2956 45124 3012 45180
rect 3012 45124 3016 45180
rect 2952 45120 3016 45124
rect 3032 45180 3096 45184
rect 3032 45124 3036 45180
rect 3036 45124 3092 45180
rect 3092 45124 3096 45180
rect 3032 45120 3096 45124
rect 3112 45180 3176 45184
rect 3112 45124 3116 45180
rect 3116 45124 3172 45180
rect 3172 45124 3176 45180
rect 3112 45120 3176 45124
rect 3192 45180 3256 45184
rect 3192 45124 3196 45180
rect 3196 45124 3252 45180
rect 3252 45124 3256 45180
rect 3192 45120 3256 45124
rect 12952 45180 13016 45184
rect 12952 45124 12956 45180
rect 12956 45124 13012 45180
rect 13012 45124 13016 45180
rect 12952 45120 13016 45124
rect 13032 45180 13096 45184
rect 13032 45124 13036 45180
rect 13036 45124 13092 45180
rect 13092 45124 13096 45180
rect 13032 45120 13096 45124
rect 13112 45180 13176 45184
rect 13112 45124 13116 45180
rect 13116 45124 13172 45180
rect 13172 45124 13176 45180
rect 13112 45120 13176 45124
rect 13192 45180 13256 45184
rect 13192 45124 13196 45180
rect 13196 45124 13252 45180
rect 13252 45124 13256 45180
rect 13192 45120 13256 45124
rect 22952 45180 23016 45184
rect 22952 45124 22956 45180
rect 22956 45124 23012 45180
rect 23012 45124 23016 45180
rect 22952 45120 23016 45124
rect 23032 45180 23096 45184
rect 23032 45124 23036 45180
rect 23036 45124 23092 45180
rect 23092 45124 23096 45180
rect 23032 45120 23096 45124
rect 23112 45180 23176 45184
rect 23112 45124 23116 45180
rect 23116 45124 23172 45180
rect 23172 45124 23176 45180
rect 23112 45120 23176 45124
rect 23192 45180 23256 45184
rect 23192 45124 23196 45180
rect 23196 45124 23252 45180
rect 23252 45124 23256 45180
rect 23192 45120 23256 45124
rect 9812 44704 9876 44708
rect 9812 44648 9826 44704
rect 9826 44648 9876 44704
rect 9812 44644 9876 44648
rect 11468 44644 11532 44708
rect 18460 44644 18524 44708
rect 7952 44636 8016 44640
rect 7952 44580 7956 44636
rect 7956 44580 8012 44636
rect 8012 44580 8016 44636
rect 7952 44576 8016 44580
rect 8032 44636 8096 44640
rect 8032 44580 8036 44636
rect 8036 44580 8092 44636
rect 8092 44580 8096 44636
rect 8032 44576 8096 44580
rect 8112 44636 8176 44640
rect 8112 44580 8116 44636
rect 8116 44580 8172 44636
rect 8172 44580 8176 44636
rect 8112 44576 8176 44580
rect 8192 44636 8256 44640
rect 8192 44580 8196 44636
rect 8196 44580 8252 44636
rect 8252 44580 8256 44636
rect 8192 44576 8256 44580
rect 17952 44636 18016 44640
rect 17952 44580 17956 44636
rect 17956 44580 18012 44636
rect 18012 44580 18016 44636
rect 17952 44576 18016 44580
rect 18032 44636 18096 44640
rect 18032 44580 18036 44636
rect 18036 44580 18092 44636
rect 18092 44580 18096 44636
rect 18032 44576 18096 44580
rect 18112 44636 18176 44640
rect 18112 44580 18116 44636
rect 18116 44580 18172 44636
rect 18172 44580 18176 44636
rect 18112 44576 18176 44580
rect 18192 44636 18256 44640
rect 18192 44580 18196 44636
rect 18196 44580 18252 44636
rect 18252 44580 18256 44636
rect 18192 44576 18256 44580
rect 10364 44236 10428 44300
rect 11652 44296 11716 44300
rect 11652 44240 11666 44296
rect 11666 44240 11716 44296
rect 11652 44236 11716 44240
rect 24532 44236 24596 44300
rect 2952 44092 3016 44096
rect 2952 44036 2956 44092
rect 2956 44036 3012 44092
rect 3012 44036 3016 44092
rect 2952 44032 3016 44036
rect 3032 44092 3096 44096
rect 3032 44036 3036 44092
rect 3036 44036 3092 44092
rect 3092 44036 3096 44092
rect 3032 44032 3096 44036
rect 3112 44092 3176 44096
rect 3112 44036 3116 44092
rect 3116 44036 3172 44092
rect 3172 44036 3176 44092
rect 3112 44032 3176 44036
rect 3192 44092 3256 44096
rect 3192 44036 3196 44092
rect 3196 44036 3252 44092
rect 3252 44036 3256 44092
rect 3192 44032 3256 44036
rect 12952 44092 13016 44096
rect 12952 44036 12956 44092
rect 12956 44036 13012 44092
rect 13012 44036 13016 44092
rect 12952 44032 13016 44036
rect 13032 44092 13096 44096
rect 13032 44036 13036 44092
rect 13036 44036 13092 44092
rect 13092 44036 13096 44092
rect 13032 44032 13096 44036
rect 13112 44092 13176 44096
rect 13112 44036 13116 44092
rect 13116 44036 13172 44092
rect 13172 44036 13176 44092
rect 13112 44032 13176 44036
rect 13192 44092 13256 44096
rect 13192 44036 13196 44092
rect 13196 44036 13252 44092
rect 13252 44036 13256 44092
rect 13192 44032 13256 44036
rect 22952 44092 23016 44096
rect 22952 44036 22956 44092
rect 22956 44036 23012 44092
rect 23012 44036 23016 44092
rect 22952 44032 23016 44036
rect 23032 44092 23096 44096
rect 23032 44036 23036 44092
rect 23036 44036 23092 44092
rect 23092 44036 23096 44092
rect 23032 44032 23096 44036
rect 23112 44092 23176 44096
rect 23112 44036 23116 44092
rect 23116 44036 23172 44092
rect 23172 44036 23176 44092
rect 23112 44032 23176 44036
rect 23192 44092 23256 44096
rect 23192 44036 23196 44092
rect 23196 44036 23252 44092
rect 23252 44036 23256 44092
rect 23192 44032 23256 44036
rect 7952 43548 8016 43552
rect 7952 43492 7956 43548
rect 7956 43492 8012 43548
rect 8012 43492 8016 43548
rect 7952 43488 8016 43492
rect 8032 43548 8096 43552
rect 8032 43492 8036 43548
rect 8036 43492 8092 43548
rect 8092 43492 8096 43548
rect 8032 43488 8096 43492
rect 8112 43548 8176 43552
rect 8112 43492 8116 43548
rect 8116 43492 8172 43548
rect 8172 43492 8176 43548
rect 8112 43488 8176 43492
rect 8192 43548 8256 43552
rect 8192 43492 8196 43548
rect 8196 43492 8252 43548
rect 8252 43492 8256 43548
rect 8192 43488 8256 43492
rect 17952 43548 18016 43552
rect 17952 43492 17956 43548
rect 17956 43492 18012 43548
rect 18012 43492 18016 43548
rect 17952 43488 18016 43492
rect 18032 43548 18096 43552
rect 18032 43492 18036 43548
rect 18036 43492 18092 43548
rect 18092 43492 18096 43548
rect 18032 43488 18096 43492
rect 18112 43548 18176 43552
rect 18112 43492 18116 43548
rect 18116 43492 18172 43548
rect 18172 43492 18176 43548
rect 18112 43488 18176 43492
rect 18192 43548 18256 43552
rect 18192 43492 18196 43548
rect 18196 43492 18252 43548
rect 18252 43492 18256 43548
rect 18192 43488 18256 43492
rect 17356 43148 17420 43212
rect 2952 43004 3016 43008
rect 2952 42948 2956 43004
rect 2956 42948 3012 43004
rect 3012 42948 3016 43004
rect 2952 42944 3016 42948
rect 3032 43004 3096 43008
rect 3032 42948 3036 43004
rect 3036 42948 3092 43004
rect 3092 42948 3096 43004
rect 3032 42944 3096 42948
rect 3112 43004 3176 43008
rect 3112 42948 3116 43004
rect 3116 42948 3172 43004
rect 3172 42948 3176 43004
rect 3112 42944 3176 42948
rect 3192 43004 3256 43008
rect 3192 42948 3196 43004
rect 3196 42948 3252 43004
rect 3252 42948 3256 43004
rect 3192 42944 3256 42948
rect 12952 43004 13016 43008
rect 12952 42948 12956 43004
rect 12956 42948 13012 43004
rect 13012 42948 13016 43004
rect 12952 42944 13016 42948
rect 13032 43004 13096 43008
rect 13032 42948 13036 43004
rect 13036 42948 13092 43004
rect 13092 42948 13096 43004
rect 13032 42944 13096 42948
rect 13112 43004 13176 43008
rect 13112 42948 13116 43004
rect 13116 42948 13172 43004
rect 13172 42948 13176 43004
rect 13112 42944 13176 42948
rect 13192 43004 13256 43008
rect 13192 42948 13196 43004
rect 13196 42948 13252 43004
rect 13252 42948 13256 43004
rect 13192 42944 13256 42948
rect 22952 43004 23016 43008
rect 22952 42948 22956 43004
rect 22956 42948 23012 43004
rect 23012 42948 23016 43004
rect 22952 42944 23016 42948
rect 23032 43004 23096 43008
rect 23032 42948 23036 43004
rect 23036 42948 23092 43004
rect 23092 42948 23096 43004
rect 23032 42944 23096 42948
rect 23112 43004 23176 43008
rect 23112 42948 23116 43004
rect 23116 42948 23172 43004
rect 23172 42948 23176 43004
rect 23112 42944 23176 42948
rect 23192 43004 23256 43008
rect 23192 42948 23196 43004
rect 23196 42948 23252 43004
rect 23252 42948 23256 43004
rect 23192 42944 23256 42948
rect 7952 42460 8016 42464
rect 7952 42404 7956 42460
rect 7956 42404 8012 42460
rect 8012 42404 8016 42460
rect 7952 42400 8016 42404
rect 8032 42460 8096 42464
rect 8032 42404 8036 42460
rect 8036 42404 8092 42460
rect 8092 42404 8096 42460
rect 8032 42400 8096 42404
rect 8112 42460 8176 42464
rect 8112 42404 8116 42460
rect 8116 42404 8172 42460
rect 8172 42404 8176 42460
rect 8112 42400 8176 42404
rect 8192 42460 8256 42464
rect 8192 42404 8196 42460
rect 8196 42404 8252 42460
rect 8252 42404 8256 42460
rect 8192 42400 8256 42404
rect 17952 42460 18016 42464
rect 17952 42404 17956 42460
rect 17956 42404 18012 42460
rect 18012 42404 18016 42460
rect 17952 42400 18016 42404
rect 18032 42460 18096 42464
rect 18032 42404 18036 42460
rect 18036 42404 18092 42460
rect 18092 42404 18096 42460
rect 18032 42400 18096 42404
rect 18112 42460 18176 42464
rect 18112 42404 18116 42460
rect 18116 42404 18172 42460
rect 18172 42404 18176 42460
rect 18112 42400 18176 42404
rect 18192 42460 18256 42464
rect 18192 42404 18196 42460
rect 18196 42404 18252 42460
rect 18252 42404 18256 42460
rect 18192 42400 18256 42404
rect 2952 41916 3016 41920
rect 2952 41860 2956 41916
rect 2956 41860 3012 41916
rect 3012 41860 3016 41916
rect 2952 41856 3016 41860
rect 3032 41916 3096 41920
rect 3032 41860 3036 41916
rect 3036 41860 3092 41916
rect 3092 41860 3096 41916
rect 3032 41856 3096 41860
rect 3112 41916 3176 41920
rect 3112 41860 3116 41916
rect 3116 41860 3172 41916
rect 3172 41860 3176 41916
rect 3112 41856 3176 41860
rect 3192 41916 3256 41920
rect 3192 41860 3196 41916
rect 3196 41860 3252 41916
rect 3252 41860 3256 41916
rect 3192 41856 3256 41860
rect 12952 41916 13016 41920
rect 12952 41860 12956 41916
rect 12956 41860 13012 41916
rect 13012 41860 13016 41916
rect 12952 41856 13016 41860
rect 13032 41916 13096 41920
rect 13032 41860 13036 41916
rect 13036 41860 13092 41916
rect 13092 41860 13096 41916
rect 13032 41856 13096 41860
rect 13112 41916 13176 41920
rect 13112 41860 13116 41916
rect 13116 41860 13172 41916
rect 13172 41860 13176 41916
rect 13112 41856 13176 41860
rect 13192 41916 13256 41920
rect 13192 41860 13196 41916
rect 13196 41860 13252 41916
rect 13252 41860 13256 41916
rect 13192 41856 13256 41860
rect 22952 41916 23016 41920
rect 22952 41860 22956 41916
rect 22956 41860 23012 41916
rect 23012 41860 23016 41916
rect 22952 41856 23016 41860
rect 23032 41916 23096 41920
rect 23032 41860 23036 41916
rect 23036 41860 23092 41916
rect 23092 41860 23096 41916
rect 23032 41856 23096 41860
rect 23112 41916 23176 41920
rect 23112 41860 23116 41916
rect 23116 41860 23172 41916
rect 23172 41860 23176 41916
rect 23112 41856 23176 41860
rect 23192 41916 23256 41920
rect 23192 41860 23196 41916
rect 23196 41860 23252 41916
rect 23252 41860 23256 41916
rect 23192 41856 23256 41860
rect 7952 41372 8016 41376
rect 7952 41316 7956 41372
rect 7956 41316 8012 41372
rect 8012 41316 8016 41372
rect 7952 41312 8016 41316
rect 8032 41372 8096 41376
rect 8032 41316 8036 41372
rect 8036 41316 8092 41372
rect 8092 41316 8096 41372
rect 8032 41312 8096 41316
rect 8112 41372 8176 41376
rect 8112 41316 8116 41372
rect 8116 41316 8172 41372
rect 8172 41316 8176 41372
rect 8112 41312 8176 41316
rect 8192 41372 8256 41376
rect 8192 41316 8196 41372
rect 8196 41316 8252 41372
rect 8252 41316 8256 41372
rect 8192 41312 8256 41316
rect 17952 41372 18016 41376
rect 17952 41316 17956 41372
rect 17956 41316 18012 41372
rect 18012 41316 18016 41372
rect 17952 41312 18016 41316
rect 18032 41372 18096 41376
rect 18032 41316 18036 41372
rect 18036 41316 18092 41372
rect 18092 41316 18096 41372
rect 18032 41312 18096 41316
rect 18112 41372 18176 41376
rect 18112 41316 18116 41372
rect 18116 41316 18172 41372
rect 18172 41316 18176 41372
rect 18112 41312 18176 41316
rect 18192 41372 18256 41376
rect 18192 41316 18196 41372
rect 18196 41316 18252 41372
rect 18252 41316 18256 41372
rect 18192 41312 18256 41316
rect 22692 41380 22756 41444
rect 2952 40828 3016 40832
rect 2952 40772 2956 40828
rect 2956 40772 3012 40828
rect 3012 40772 3016 40828
rect 2952 40768 3016 40772
rect 3032 40828 3096 40832
rect 3032 40772 3036 40828
rect 3036 40772 3092 40828
rect 3092 40772 3096 40828
rect 3032 40768 3096 40772
rect 3112 40828 3176 40832
rect 3112 40772 3116 40828
rect 3116 40772 3172 40828
rect 3172 40772 3176 40828
rect 3112 40768 3176 40772
rect 3192 40828 3256 40832
rect 3192 40772 3196 40828
rect 3196 40772 3252 40828
rect 3252 40772 3256 40828
rect 3192 40768 3256 40772
rect 12952 40828 13016 40832
rect 12952 40772 12956 40828
rect 12956 40772 13012 40828
rect 13012 40772 13016 40828
rect 12952 40768 13016 40772
rect 13032 40828 13096 40832
rect 13032 40772 13036 40828
rect 13036 40772 13092 40828
rect 13092 40772 13096 40828
rect 13032 40768 13096 40772
rect 13112 40828 13176 40832
rect 13112 40772 13116 40828
rect 13116 40772 13172 40828
rect 13172 40772 13176 40828
rect 13112 40768 13176 40772
rect 13192 40828 13256 40832
rect 13192 40772 13196 40828
rect 13196 40772 13252 40828
rect 13252 40772 13256 40828
rect 13192 40768 13256 40772
rect 22952 40828 23016 40832
rect 22952 40772 22956 40828
rect 22956 40772 23012 40828
rect 23012 40772 23016 40828
rect 22952 40768 23016 40772
rect 23032 40828 23096 40832
rect 23032 40772 23036 40828
rect 23036 40772 23092 40828
rect 23092 40772 23096 40828
rect 23032 40768 23096 40772
rect 23112 40828 23176 40832
rect 23112 40772 23116 40828
rect 23116 40772 23172 40828
rect 23172 40772 23176 40828
rect 23112 40768 23176 40772
rect 23192 40828 23256 40832
rect 23192 40772 23196 40828
rect 23196 40772 23252 40828
rect 23252 40772 23256 40828
rect 23192 40768 23256 40772
rect 17724 40564 17788 40628
rect 7952 40284 8016 40288
rect 7952 40228 7956 40284
rect 7956 40228 8012 40284
rect 8012 40228 8016 40284
rect 7952 40224 8016 40228
rect 8032 40284 8096 40288
rect 8032 40228 8036 40284
rect 8036 40228 8092 40284
rect 8092 40228 8096 40284
rect 8032 40224 8096 40228
rect 8112 40284 8176 40288
rect 8112 40228 8116 40284
rect 8116 40228 8172 40284
rect 8172 40228 8176 40284
rect 8112 40224 8176 40228
rect 8192 40284 8256 40288
rect 8192 40228 8196 40284
rect 8196 40228 8252 40284
rect 8252 40228 8256 40284
rect 8192 40224 8256 40228
rect 17952 40284 18016 40288
rect 17952 40228 17956 40284
rect 17956 40228 18012 40284
rect 18012 40228 18016 40284
rect 17952 40224 18016 40228
rect 18032 40284 18096 40288
rect 18032 40228 18036 40284
rect 18036 40228 18092 40284
rect 18092 40228 18096 40284
rect 18032 40224 18096 40228
rect 18112 40284 18176 40288
rect 18112 40228 18116 40284
rect 18116 40228 18172 40284
rect 18172 40228 18176 40284
rect 18112 40224 18176 40228
rect 18192 40284 18256 40288
rect 18192 40228 18196 40284
rect 18196 40228 18252 40284
rect 18252 40228 18256 40284
rect 18192 40224 18256 40228
rect 22508 40156 22572 40220
rect 22140 40020 22204 40084
rect 22324 40020 22388 40084
rect 23428 40020 23492 40084
rect 2952 39740 3016 39744
rect 2952 39684 2956 39740
rect 2956 39684 3012 39740
rect 3012 39684 3016 39740
rect 2952 39680 3016 39684
rect 3032 39740 3096 39744
rect 3032 39684 3036 39740
rect 3036 39684 3092 39740
rect 3092 39684 3096 39740
rect 3032 39680 3096 39684
rect 3112 39740 3176 39744
rect 3112 39684 3116 39740
rect 3116 39684 3172 39740
rect 3172 39684 3176 39740
rect 3112 39680 3176 39684
rect 3192 39740 3256 39744
rect 3192 39684 3196 39740
rect 3196 39684 3252 39740
rect 3252 39684 3256 39740
rect 3192 39680 3256 39684
rect 12952 39740 13016 39744
rect 12952 39684 12956 39740
rect 12956 39684 13012 39740
rect 13012 39684 13016 39740
rect 12952 39680 13016 39684
rect 13032 39740 13096 39744
rect 13032 39684 13036 39740
rect 13036 39684 13092 39740
rect 13092 39684 13096 39740
rect 13032 39680 13096 39684
rect 13112 39740 13176 39744
rect 13112 39684 13116 39740
rect 13116 39684 13172 39740
rect 13172 39684 13176 39740
rect 13112 39680 13176 39684
rect 13192 39740 13256 39744
rect 13192 39684 13196 39740
rect 13196 39684 13252 39740
rect 13252 39684 13256 39740
rect 13192 39680 13256 39684
rect 22952 39740 23016 39744
rect 22952 39684 22956 39740
rect 22956 39684 23012 39740
rect 23012 39684 23016 39740
rect 22952 39680 23016 39684
rect 23032 39740 23096 39744
rect 23032 39684 23036 39740
rect 23036 39684 23092 39740
rect 23092 39684 23096 39740
rect 23032 39680 23096 39684
rect 23112 39740 23176 39744
rect 23112 39684 23116 39740
rect 23116 39684 23172 39740
rect 23172 39684 23176 39740
rect 23112 39680 23176 39684
rect 23192 39740 23256 39744
rect 23192 39684 23196 39740
rect 23196 39684 23252 39740
rect 23252 39684 23256 39740
rect 23192 39680 23256 39684
rect 7952 39196 8016 39200
rect 7952 39140 7956 39196
rect 7956 39140 8012 39196
rect 8012 39140 8016 39196
rect 7952 39136 8016 39140
rect 8032 39196 8096 39200
rect 8032 39140 8036 39196
rect 8036 39140 8092 39196
rect 8092 39140 8096 39196
rect 8032 39136 8096 39140
rect 8112 39196 8176 39200
rect 8112 39140 8116 39196
rect 8116 39140 8172 39196
rect 8172 39140 8176 39196
rect 8112 39136 8176 39140
rect 8192 39196 8256 39200
rect 8192 39140 8196 39196
rect 8196 39140 8252 39196
rect 8252 39140 8256 39196
rect 8192 39136 8256 39140
rect 17952 39196 18016 39200
rect 17952 39140 17956 39196
rect 17956 39140 18012 39196
rect 18012 39140 18016 39196
rect 17952 39136 18016 39140
rect 18032 39196 18096 39200
rect 18032 39140 18036 39196
rect 18036 39140 18092 39196
rect 18092 39140 18096 39196
rect 18032 39136 18096 39140
rect 18112 39196 18176 39200
rect 18112 39140 18116 39196
rect 18116 39140 18172 39196
rect 18172 39140 18176 39196
rect 18112 39136 18176 39140
rect 18192 39196 18256 39200
rect 18192 39140 18196 39196
rect 18196 39140 18252 39196
rect 18252 39140 18256 39196
rect 18192 39136 18256 39140
rect 16068 38660 16132 38724
rect 2952 38652 3016 38656
rect 2952 38596 2956 38652
rect 2956 38596 3012 38652
rect 3012 38596 3016 38652
rect 2952 38592 3016 38596
rect 3032 38652 3096 38656
rect 3032 38596 3036 38652
rect 3036 38596 3092 38652
rect 3092 38596 3096 38652
rect 3032 38592 3096 38596
rect 3112 38652 3176 38656
rect 3112 38596 3116 38652
rect 3116 38596 3172 38652
rect 3172 38596 3176 38652
rect 3112 38592 3176 38596
rect 3192 38652 3256 38656
rect 3192 38596 3196 38652
rect 3196 38596 3252 38652
rect 3252 38596 3256 38652
rect 3192 38592 3256 38596
rect 12952 38652 13016 38656
rect 12952 38596 12956 38652
rect 12956 38596 13012 38652
rect 13012 38596 13016 38652
rect 12952 38592 13016 38596
rect 13032 38652 13096 38656
rect 13032 38596 13036 38652
rect 13036 38596 13092 38652
rect 13092 38596 13096 38652
rect 13032 38592 13096 38596
rect 13112 38652 13176 38656
rect 13112 38596 13116 38652
rect 13116 38596 13172 38652
rect 13172 38596 13176 38652
rect 13112 38592 13176 38596
rect 13192 38652 13256 38656
rect 13192 38596 13196 38652
rect 13196 38596 13252 38652
rect 13252 38596 13256 38652
rect 13192 38592 13256 38596
rect 22952 38652 23016 38656
rect 22952 38596 22956 38652
rect 22956 38596 23012 38652
rect 23012 38596 23016 38652
rect 22952 38592 23016 38596
rect 23032 38652 23096 38656
rect 23032 38596 23036 38652
rect 23036 38596 23092 38652
rect 23092 38596 23096 38652
rect 23032 38592 23096 38596
rect 23112 38652 23176 38656
rect 23112 38596 23116 38652
rect 23116 38596 23172 38652
rect 23172 38596 23176 38652
rect 23112 38592 23176 38596
rect 23192 38652 23256 38656
rect 23192 38596 23196 38652
rect 23196 38596 23252 38652
rect 23252 38596 23256 38652
rect 23192 38592 23256 38596
rect 21588 38388 21652 38452
rect 12572 38312 12636 38316
rect 12572 38256 12622 38312
rect 12622 38256 12636 38312
rect 12572 38252 12636 38256
rect 7952 38108 8016 38112
rect 7952 38052 7956 38108
rect 7956 38052 8012 38108
rect 8012 38052 8016 38108
rect 7952 38048 8016 38052
rect 8032 38108 8096 38112
rect 8032 38052 8036 38108
rect 8036 38052 8092 38108
rect 8092 38052 8096 38108
rect 8032 38048 8096 38052
rect 8112 38108 8176 38112
rect 8112 38052 8116 38108
rect 8116 38052 8172 38108
rect 8172 38052 8176 38108
rect 8112 38048 8176 38052
rect 8192 38108 8256 38112
rect 8192 38052 8196 38108
rect 8196 38052 8252 38108
rect 8252 38052 8256 38108
rect 8192 38048 8256 38052
rect 17952 38108 18016 38112
rect 17952 38052 17956 38108
rect 17956 38052 18012 38108
rect 18012 38052 18016 38108
rect 17952 38048 18016 38052
rect 18032 38108 18096 38112
rect 18032 38052 18036 38108
rect 18036 38052 18092 38108
rect 18092 38052 18096 38108
rect 18032 38048 18096 38052
rect 18112 38108 18176 38112
rect 18112 38052 18116 38108
rect 18116 38052 18172 38108
rect 18172 38052 18176 38108
rect 18112 38048 18176 38052
rect 18192 38108 18256 38112
rect 18192 38052 18196 38108
rect 18196 38052 18252 38108
rect 18252 38052 18256 38108
rect 18192 38048 18256 38052
rect 22692 38040 22756 38044
rect 22692 37984 22706 38040
rect 22706 37984 22756 38040
rect 22692 37980 22756 37984
rect 2952 37564 3016 37568
rect 2952 37508 2956 37564
rect 2956 37508 3012 37564
rect 3012 37508 3016 37564
rect 2952 37504 3016 37508
rect 3032 37564 3096 37568
rect 3032 37508 3036 37564
rect 3036 37508 3092 37564
rect 3092 37508 3096 37564
rect 3032 37504 3096 37508
rect 3112 37564 3176 37568
rect 3112 37508 3116 37564
rect 3116 37508 3172 37564
rect 3172 37508 3176 37564
rect 3112 37504 3176 37508
rect 3192 37564 3256 37568
rect 3192 37508 3196 37564
rect 3196 37508 3252 37564
rect 3252 37508 3256 37564
rect 3192 37504 3256 37508
rect 12952 37564 13016 37568
rect 12952 37508 12956 37564
rect 12956 37508 13012 37564
rect 13012 37508 13016 37564
rect 12952 37504 13016 37508
rect 13032 37564 13096 37568
rect 13032 37508 13036 37564
rect 13036 37508 13092 37564
rect 13092 37508 13096 37564
rect 13032 37504 13096 37508
rect 13112 37564 13176 37568
rect 13112 37508 13116 37564
rect 13116 37508 13172 37564
rect 13172 37508 13176 37564
rect 13112 37504 13176 37508
rect 13192 37564 13256 37568
rect 13192 37508 13196 37564
rect 13196 37508 13252 37564
rect 13252 37508 13256 37564
rect 13192 37504 13256 37508
rect 22952 37564 23016 37568
rect 22952 37508 22956 37564
rect 22956 37508 23012 37564
rect 23012 37508 23016 37564
rect 22952 37504 23016 37508
rect 23032 37564 23096 37568
rect 23032 37508 23036 37564
rect 23036 37508 23092 37564
rect 23092 37508 23096 37564
rect 23032 37504 23096 37508
rect 23112 37564 23176 37568
rect 23112 37508 23116 37564
rect 23116 37508 23172 37564
rect 23172 37508 23176 37564
rect 23112 37504 23176 37508
rect 23192 37564 23256 37568
rect 23192 37508 23196 37564
rect 23196 37508 23252 37564
rect 23252 37508 23256 37564
rect 23192 37504 23256 37508
rect 19380 37360 19444 37364
rect 19380 37304 19394 37360
rect 19394 37304 19444 37360
rect 19380 37300 19444 37304
rect 7952 37020 8016 37024
rect 7952 36964 7956 37020
rect 7956 36964 8012 37020
rect 8012 36964 8016 37020
rect 7952 36960 8016 36964
rect 8032 37020 8096 37024
rect 8032 36964 8036 37020
rect 8036 36964 8092 37020
rect 8092 36964 8096 37020
rect 8032 36960 8096 36964
rect 8112 37020 8176 37024
rect 8112 36964 8116 37020
rect 8116 36964 8172 37020
rect 8172 36964 8176 37020
rect 8112 36960 8176 36964
rect 8192 37020 8256 37024
rect 8192 36964 8196 37020
rect 8196 36964 8252 37020
rect 8252 36964 8256 37020
rect 8192 36960 8256 36964
rect 17952 37020 18016 37024
rect 17952 36964 17956 37020
rect 17956 36964 18012 37020
rect 18012 36964 18016 37020
rect 17952 36960 18016 36964
rect 18032 37020 18096 37024
rect 18032 36964 18036 37020
rect 18036 36964 18092 37020
rect 18092 36964 18096 37020
rect 18032 36960 18096 36964
rect 18112 37020 18176 37024
rect 18112 36964 18116 37020
rect 18116 36964 18172 37020
rect 18172 36964 18176 37020
rect 18112 36960 18176 36964
rect 18192 37020 18256 37024
rect 18192 36964 18196 37020
rect 18196 36964 18252 37020
rect 18252 36964 18256 37020
rect 18192 36960 18256 36964
rect 9812 36756 9876 36820
rect 21036 36544 21100 36548
rect 21036 36488 21086 36544
rect 21086 36488 21100 36544
rect 21036 36484 21100 36488
rect 2952 36476 3016 36480
rect 2952 36420 2956 36476
rect 2956 36420 3012 36476
rect 3012 36420 3016 36476
rect 2952 36416 3016 36420
rect 3032 36476 3096 36480
rect 3032 36420 3036 36476
rect 3036 36420 3092 36476
rect 3092 36420 3096 36476
rect 3032 36416 3096 36420
rect 3112 36476 3176 36480
rect 3112 36420 3116 36476
rect 3116 36420 3172 36476
rect 3172 36420 3176 36476
rect 3112 36416 3176 36420
rect 3192 36476 3256 36480
rect 3192 36420 3196 36476
rect 3196 36420 3252 36476
rect 3252 36420 3256 36476
rect 3192 36416 3256 36420
rect 12952 36476 13016 36480
rect 12952 36420 12956 36476
rect 12956 36420 13012 36476
rect 13012 36420 13016 36476
rect 12952 36416 13016 36420
rect 13032 36476 13096 36480
rect 13032 36420 13036 36476
rect 13036 36420 13092 36476
rect 13092 36420 13096 36476
rect 13032 36416 13096 36420
rect 13112 36476 13176 36480
rect 13112 36420 13116 36476
rect 13116 36420 13172 36476
rect 13172 36420 13176 36476
rect 13112 36416 13176 36420
rect 13192 36476 13256 36480
rect 13192 36420 13196 36476
rect 13196 36420 13252 36476
rect 13252 36420 13256 36476
rect 13192 36416 13256 36420
rect 22952 36476 23016 36480
rect 22952 36420 22956 36476
rect 22956 36420 23012 36476
rect 23012 36420 23016 36476
rect 22952 36416 23016 36420
rect 23032 36476 23096 36480
rect 23032 36420 23036 36476
rect 23036 36420 23092 36476
rect 23092 36420 23096 36476
rect 23032 36416 23096 36420
rect 23112 36476 23176 36480
rect 23112 36420 23116 36476
rect 23116 36420 23172 36476
rect 23172 36420 23176 36476
rect 23112 36416 23176 36420
rect 23192 36476 23256 36480
rect 23192 36420 23196 36476
rect 23196 36420 23252 36476
rect 23252 36420 23256 36476
rect 23192 36416 23256 36420
rect 11284 36408 11348 36412
rect 11284 36352 11298 36408
rect 11298 36352 11348 36408
rect 11284 36348 11348 36352
rect 14780 35940 14844 36004
rect 7952 35932 8016 35936
rect 7952 35876 7956 35932
rect 7956 35876 8012 35932
rect 8012 35876 8016 35932
rect 7952 35872 8016 35876
rect 8032 35932 8096 35936
rect 8032 35876 8036 35932
rect 8036 35876 8092 35932
rect 8092 35876 8096 35932
rect 8032 35872 8096 35876
rect 8112 35932 8176 35936
rect 8112 35876 8116 35932
rect 8116 35876 8172 35932
rect 8172 35876 8176 35932
rect 8112 35872 8176 35876
rect 8192 35932 8256 35936
rect 8192 35876 8196 35932
rect 8196 35876 8252 35932
rect 8252 35876 8256 35932
rect 8192 35872 8256 35876
rect 17952 35932 18016 35936
rect 17952 35876 17956 35932
rect 17956 35876 18012 35932
rect 18012 35876 18016 35932
rect 17952 35872 18016 35876
rect 18032 35932 18096 35936
rect 18032 35876 18036 35932
rect 18036 35876 18092 35932
rect 18092 35876 18096 35932
rect 18032 35872 18096 35876
rect 18112 35932 18176 35936
rect 18112 35876 18116 35932
rect 18116 35876 18172 35932
rect 18172 35876 18176 35932
rect 18112 35872 18176 35876
rect 18192 35932 18256 35936
rect 18192 35876 18196 35932
rect 18196 35876 18252 35932
rect 18252 35876 18256 35932
rect 18192 35872 18256 35876
rect 2952 35388 3016 35392
rect 2952 35332 2956 35388
rect 2956 35332 3012 35388
rect 3012 35332 3016 35388
rect 2952 35328 3016 35332
rect 3032 35388 3096 35392
rect 3032 35332 3036 35388
rect 3036 35332 3092 35388
rect 3092 35332 3096 35388
rect 3032 35328 3096 35332
rect 3112 35388 3176 35392
rect 3112 35332 3116 35388
rect 3116 35332 3172 35388
rect 3172 35332 3176 35388
rect 3112 35328 3176 35332
rect 3192 35388 3256 35392
rect 3192 35332 3196 35388
rect 3196 35332 3252 35388
rect 3252 35332 3256 35388
rect 3192 35328 3256 35332
rect 12952 35388 13016 35392
rect 12952 35332 12956 35388
rect 12956 35332 13012 35388
rect 13012 35332 13016 35388
rect 12952 35328 13016 35332
rect 13032 35388 13096 35392
rect 13032 35332 13036 35388
rect 13036 35332 13092 35388
rect 13092 35332 13096 35388
rect 13032 35328 13096 35332
rect 13112 35388 13176 35392
rect 13112 35332 13116 35388
rect 13116 35332 13172 35388
rect 13172 35332 13176 35388
rect 13112 35328 13176 35332
rect 13192 35388 13256 35392
rect 13192 35332 13196 35388
rect 13196 35332 13252 35388
rect 13252 35332 13256 35388
rect 13192 35328 13256 35332
rect 22952 35388 23016 35392
rect 22952 35332 22956 35388
rect 22956 35332 23012 35388
rect 23012 35332 23016 35388
rect 22952 35328 23016 35332
rect 23032 35388 23096 35392
rect 23032 35332 23036 35388
rect 23036 35332 23092 35388
rect 23092 35332 23096 35388
rect 23032 35328 23096 35332
rect 23112 35388 23176 35392
rect 23112 35332 23116 35388
rect 23116 35332 23172 35388
rect 23172 35332 23176 35388
rect 23112 35328 23176 35332
rect 23192 35388 23256 35392
rect 23192 35332 23196 35388
rect 23196 35332 23252 35388
rect 23252 35332 23256 35388
rect 23192 35328 23256 35332
rect 24532 35124 24596 35188
rect 7952 34844 8016 34848
rect 7952 34788 7956 34844
rect 7956 34788 8012 34844
rect 8012 34788 8016 34844
rect 7952 34784 8016 34788
rect 8032 34844 8096 34848
rect 8032 34788 8036 34844
rect 8036 34788 8092 34844
rect 8092 34788 8096 34844
rect 8032 34784 8096 34788
rect 8112 34844 8176 34848
rect 8112 34788 8116 34844
rect 8116 34788 8172 34844
rect 8172 34788 8176 34844
rect 8112 34784 8176 34788
rect 8192 34844 8256 34848
rect 8192 34788 8196 34844
rect 8196 34788 8252 34844
rect 8252 34788 8256 34844
rect 8192 34784 8256 34788
rect 17952 34844 18016 34848
rect 17952 34788 17956 34844
rect 17956 34788 18012 34844
rect 18012 34788 18016 34844
rect 17952 34784 18016 34788
rect 18032 34844 18096 34848
rect 18032 34788 18036 34844
rect 18036 34788 18092 34844
rect 18092 34788 18096 34844
rect 18032 34784 18096 34788
rect 18112 34844 18176 34848
rect 18112 34788 18116 34844
rect 18116 34788 18172 34844
rect 18172 34788 18176 34844
rect 18112 34784 18176 34788
rect 18192 34844 18256 34848
rect 18192 34788 18196 34844
rect 18196 34788 18252 34844
rect 18252 34788 18256 34844
rect 18192 34784 18256 34788
rect 2952 34300 3016 34304
rect 2952 34244 2956 34300
rect 2956 34244 3012 34300
rect 3012 34244 3016 34300
rect 2952 34240 3016 34244
rect 3032 34300 3096 34304
rect 3032 34244 3036 34300
rect 3036 34244 3092 34300
rect 3092 34244 3096 34300
rect 3032 34240 3096 34244
rect 3112 34300 3176 34304
rect 3112 34244 3116 34300
rect 3116 34244 3172 34300
rect 3172 34244 3176 34300
rect 3112 34240 3176 34244
rect 3192 34300 3256 34304
rect 3192 34244 3196 34300
rect 3196 34244 3252 34300
rect 3252 34244 3256 34300
rect 3192 34240 3256 34244
rect 12952 34300 13016 34304
rect 12952 34244 12956 34300
rect 12956 34244 13012 34300
rect 13012 34244 13016 34300
rect 12952 34240 13016 34244
rect 13032 34300 13096 34304
rect 13032 34244 13036 34300
rect 13036 34244 13092 34300
rect 13092 34244 13096 34300
rect 13032 34240 13096 34244
rect 13112 34300 13176 34304
rect 13112 34244 13116 34300
rect 13116 34244 13172 34300
rect 13172 34244 13176 34300
rect 13112 34240 13176 34244
rect 13192 34300 13256 34304
rect 13192 34244 13196 34300
rect 13196 34244 13252 34300
rect 13252 34244 13256 34300
rect 13192 34240 13256 34244
rect 22952 34300 23016 34304
rect 22952 34244 22956 34300
rect 22956 34244 23012 34300
rect 23012 34244 23016 34300
rect 22952 34240 23016 34244
rect 23032 34300 23096 34304
rect 23032 34244 23036 34300
rect 23036 34244 23092 34300
rect 23092 34244 23096 34300
rect 23032 34240 23096 34244
rect 23112 34300 23176 34304
rect 23112 34244 23116 34300
rect 23116 34244 23172 34300
rect 23172 34244 23176 34300
rect 23112 34240 23176 34244
rect 23192 34300 23256 34304
rect 23192 34244 23196 34300
rect 23196 34244 23252 34300
rect 23252 34244 23256 34300
rect 23192 34240 23256 34244
rect 7952 33756 8016 33760
rect 7952 33700 7956 33756
rect 7956 33700 8012 33756
rect 8012 33700 8016 33756
rect 7952 33696 8016 33700
rect 8032 33756 8096 33760
rect 8032 33700 8036 33756
rect 8036 33700 8092 33756
rect 8092 33700 8096 33756
rect 8032 33696 8096 33700
rect 8112 33756 8176 33760
rect 8112 33700 8116 33756
rect 8116 33700 8172 33756
rect 8172 33700 8176 33756
rect 8112 33696 8176 33700
rect 8192 33756 8256 33760
rect 8192 33700 8196 33756
rect 8196 33700 8252 33756
rect 8252 33700 8256 33756
rect 8192 33696 8256 33700
rect 17952 33756 18016 33760
rect 17952 33700 17956 33756
rect 17956 33700 18012 33756
rect 18012 33700 18016 33756
rect 17952 33696 18016 33700
rect 18032 33756 18096 33760
rect 18032 33700 18036 33756
rect 18036 33700 18092 33756
rect 18092 33700 18096 33756
rect 18032 33696 18096 33700
rect 18112 33756 18176 33760
rect 18112 33700 18116 33756
rect 18116 33700 18172 33756
rect 18172 33700 18176 33756
rect 18112 33696 18176 33700
rect 18192 33756 18256 33760
rect 18192 33700 18196 33756
rect 18196 33700 18252 33756
rect 18252 33700 18256 33756
rect 18192 33696 18256 33700
rect 24716 33356 24780 33420
rect 12572 33280 12636 33284
rect 12572 33224 12586 33280
rect 12586 33224 12636 33280
rect 12572 33220 12636 33224
rect 2952 33212 3016 33216
rect 2952 33156 2956 33212
rect 2956 33156 3012 33212
rect 3012 33156 3016 33212
rect 2952 33152 3016 33156
rect 3032 33212 3096 33216
rect 3032 33156 3036 33212
rect 3036 33156 3092 33212
rect 3092 33156 3096 33212
rect 3032 33152 3096 33156
rect 3112 33212 3176 33216
rect 3112 33156 3116 33212
rect 3116 33156 3172 33212
rect 3172 33156 3176 33212
rect 3112 33152 3176 33156
rect 3192 33212 3256 33216
rect 3192 33156 3196 33212
rect 3196 33156 3252 33212
rect 3252 33156 3256 33212
rect 3192 33152 3256 33156
rect 12952 33212 13016 33216
rect 12952 33156 12956 33212
rect 12956 33156 13012 33212
rect 13012 33156 13016 33212
rect 12952 33152 13016 33156
rect 13032 33212 13096 33216
rect 13032 33156 13036 33212
rect 13036 33156 13092 33212
rect 13092 33156 13096 33212
rect 13032 33152 13096 33156
rect 13112 33212 13176 33216
rect 13112 33156 13116 33212
rect 13116 33156 13172 33212
rect 13172 33156 13176 33212
rect 13112 33152 13176 33156
rect 13192 33212 13256 33216
rect 13192 33156 13196 33212
rect 13196 33156 13252 33212
rect 13252 33156 13256 33212
rect 13192 33152 13256 33156
rect 22952 33212 23016 33216
rect 22952 33156 22956 33212
rect 22956 33156 23012 33212
rect 23012 33156 23016 33212
rect 22952 33152 23016 33156
rect 23032 33212 23096 33216
rect 23032 33156 23036 33212
rect 23036 33156 23092 33212
rect 23092 33156 23096 33212
rect 23032 33152 23096 33156
rect 23112 33212 23176 33216
rect 23112 33156 23116 33212
rect 23116 33156 23172 33212
rect 23172 33156 23176 33212
rect 23112 33152 23176 33156
rect 23192 33212 23256 33216
rect 23192 33156 23196 33212
rect 23196 33156 23252 33212
rect 23252 33156 23256 33212
rect 23192 33152 23256 33156
rect 19196 33084 19260 33148
rect 22140 33144 22204 33148
rect 22140 33088 22190 33144
rect 22190 33088 22204 33144
rect 22140 33084 22204 33088
rect 11468 32948 11532 33012
rect 23428 32948 23492 33012
rect 13860 32812 13924 32876
rect 7952 32668 8016 32672
rect 7952 32612 7956 32668
rect 7956 32612 8012 32668
rect 8012 32612 8016 32668
rect 7952 32608 8016 32612
rect 8032 32668 8096 32672
rect 8032 32612 8036 32668
rect 8036 32612 8092 32668
rect 8092 32612 8096 32668
rect 8032 32608 8096 32612
rect 8112 32668 8176 32672
rect 8112 32612 8116 32668
rect 8116 32612 8172 32668
rect 8172 32612 8176 32668
rect 8112 32608 8176 32612
rect 8192 32668 8256 32672
rect 8192 32612 8196 32668
rect 8196 32612 8252 32668
rect 8252 32612 8256 32668
rect 8192 32608 8256 32612
rect 17952 32668 18016 32672
rect 17952 32612 17956 32668
rect 17956 32612 18012 32668
rect 18012 32612 18016 32668
rect 17952 32608 18016 32612
rect 18032 32668 18096 32672
rect 18032 32612 18036 32668
rect 18036 32612 18092 32668
rect 18092 32612 18096 32668
rect 18032 32608 18096 32612
rect 18112 32668 18176 32672
rect 18112 32612 18116 32668
rect 18116 32612 18172 32668
rect 18172 32612 18176 32668
rect 18112 32608 18176 32612
rect 18192 32668 18256 32672
rect 18192 32612 18196 32668
rect 18196 32612 18252 32668
rect 18252 32612 18256 32668
rect 18192 32608 18256 32612
rect 11652 32540 11716 32604
rect 2952 32124 3016 32128
rect 2952 32068 2956 32124
rect 2956 32068 3012 32124
rect 3012 32068 3016 32124
rect 2952 32064 3016 32068
rect 3032 32124 3096 32128
rect 3032 32068 3036 32124
rect 3036 32068 3092 32124
rect 3092 32068 3096 32124
rect 3032 32064 3096 32068
rect 3112 32124 3176 32128
rect 3112 32068 3116 32124
rect 3116 32068 3172 32124
rect 3172 32068 3176 32124
rect 3112 32064 3176 32068
rect 3192 32124 3256 32128
rect 3192 32068 3196 32124
rect 3196 32068 3252 32124
rect 3252 32068 3256 32124
rect 3192 32064 3256 32068
rect 12952 32124 13016 32128
rect 12952 32068 12956 32124
rect 12956 32068 13012 32124
rect 13012 32068 13016 32124
rect 12952 32064 13016 32068
rect 13032 32124 13096 32128
rect 13032 32068 13036 32124
rect 13036 32068 13092 32124
rect 13092 32068 13096 32124
rect 13032 32064 13096 32068
rect 13112 32124 13176 32128
rect 13112 32068 13116 32124
rect 13116 32068 13172 32124
rect 13172 32068 13176 32124
rect 13112 32064 13176 32068
rect 13192 32124 13256 32128
rect 13192 32068 13196 32124
rect 13196 32068 13252 32124
rect 13252 32068 13256 32124
rect 13192 32064 13256 32068
rect 22952 32124 23016 32128
rect 22952 32068 22956 32124
rect 22956 32068 23012 32124
rect 23012 32068 23016 32124
rect 22952 32064 23016 32068
rect 23032 32124 23096 32128
rect 23032 32068 23036 32124
rect 23036 32068 23092 32124
rect 23092 32068 23096 32124
rect 23032 32064 23096 32068
rect 23112 32124 23176 32128
rect 23112 32068 23116 32124
rect 23116 32068 23172 32124
rect 23172 32068 23176 32124
rect 23112 32064 23176 32068
rect 23192 32124 23256 32128
rect 23192 32068 23196 32124
rect 23196 32068 23252 32124
rect 23252 32068 23256 32124
rect 23192 32064 23256 32068
rect 21588 32056 21652 32060
rect 21588 32000 21602 32056
rect 21602 32000 21652 32056
rect 21588 31996 21652 32000
rect 20116 31860 20180 31924
rect 21036 31724 21100 31788
rect 7952 31580 8016 31584
rect 7952 31524 7956 31580
rect 7956 31524 8012 31580
rect 8012 31524 8016 31580
rect 7952 31520 8016 31524
rect 8032 31580 8096 31584
rect 8032 31524 8036 31580
rect 8036 31524 8092 31580
rect 8092 31524 8096 31580
rect 8032 31520 8096 31524
rect 8112 31580 8176 31584
rect 8112 31524 8116 31580
rect 8116 31524 8172 31580
rect 8172 31524 8176 31580
rect 8112 31520 8176 31524
rect 8192 31580 8256 31584
rect 8192 31524 8196 31580
rect 8196 31524 8252 31580
rect 8252 31524 8256 31580
rect 8192 31520 8256 31524
rect 17952 31580 18016 31584
rect 17952 31524 17956 31580
rect 17956 31524 18012 31580
rect 18012 31524 18016 31580
rect 17952 31520 18016 31524
rect 18032 31580 18096 31584
rect 18032 31524 18036 31580
rect 18036 31524 18092 31580
rect 18092 31524 18096 31580
rect 18032 31520 18096 31524
rect 18112 31580 18176 31584
rect 18112 31524 18116 31580
rect 18116 31524 18172 31580
rect 18172 31524 18176 31580
rect 18112 31520 18176 31524
rect 18192 31580 18256 31584
rect 18192 31524 18196 31580
rect 18196 31524 18252 31580
rect 18252 31524 18256 31580
rect 18192 31520 18256 31524
rect 2952 31036 3016 31040
rect 2952 30980 2956 31036
rect 2956 30980 3012 31036
rect 3012 30980 3016 31036
rect 2952 30976 3016 30980
rect 3032 31036 3096 31040
rect 3032 30980 3036 31036
rect 3036 30980 3092 31036
rect 3092 30980 3096 31036
rect 3032 30976 3096 30980
rect 3112 31036 3176 31040
rect 3112 30980 3116 31036
rect 3116 30980 3172 31036
rect 3172 30980 3176 31036
rect 3112 30976 3176 30980
rect 3192 31036 3256 31040
rect 3192 30980 3196 31036
rect 3196 30980 3252 31036
rect 3252 30980 3256 31036
rect 3192 30976 3256 30980
rect 12952 31036 13016 31040
rect 12952 30980 12956 31036
rect 12956 30980 13012 31036
rect 13012 30980 13016 31036
rect 12952 30976 13016 30980
rect 13032 31036 13096 31040
rect 13032 30980 13036 31036
rect 13036 30980 13092 31036
rect 13092 30980 13096 31036
rect 13032 30976 13096 30980
rect 13112 31036 13176 31040
rect 13112 30980 13116 31036
rect 13116 30980 13172 31036
rect 13172 30980 13176 31036
rect 13112 30976 13176 30980
rect 13192 31036 13256 31040
rect 13192 30980 13196 31036
rect 13196 30980 13252 31036
rect 13252 30980 13256 31036
rect 13192 30976 13256 30980
rect 22952 31036 23016 31040
rect 22952 30980 22956 31036
rect 22956 30980 23012 31036
rect 23012 30980 23016 31036
rect 22952 30976 23016 30980
rect 23032 31036 23096 31040
rect 23032 30980 23036 31036
rect 23036 30980 23092 31036
rect 23092 30980 23096 31036
rect 23032 30976 23096 30980
rect 23112 31036 23176 31040
rect 23112 30980 23116 31036
rect 23116 30980 23172 31036
rect 23172 30980 23176 31036
rect 23112 30976 23176 30980
rect 23192 31036 23256 31040
rect 23192 30980 23196 31036
rect 23196 30980 23252 31036
rect 23252 30980 23256 31036
rect 23192 30976 23256 30980
rect 10364 30772 10428 30836
rect 19380 30772 19444 30836
rect 15332 30560 15396 30564
rect 15332 30504 15382 30560
rect 15382 30504 15396 30560
rect 15332 30500 15396 30504
rect 19932 30560 19996 30564
rect 19932 30504 19946 30560
rect 19946 30504 19996 30560
rect 19932 30500 19996 30504
rect 7952 30492 8016 30496
rect 7952 30436 7956 30492
rect 7956 30436 8012 30492
rect 8012 30436 8016 30492
rect 7952 30432 8016 30436
rect 8032 30492 8096 30496
rect 8032 30436 8036 30492
rect 8036 30436 8092 30492
rect 8092 30436 8096 30492
rect 8032 30432 8096 30436
rect 8112 30492 8176 30496
rect 8112 30436 8116 30492
rect 8116 30436 8172 30492
rect 8172 30436 8176 30492
rect 8112 30432 8176 30436
rect 8192 30492 8256 30496
rect 8192 30436 8196 30492
rect 8196 30436 8252 30492
rect 8252 30436 8256 30492
rect 8192 30432 8256 30436
rect 17952 30492 18016 30496
rect 17952 30436 17956 30492
rect 17956 30436 18012 30492
rect 18012 30436 18016 30492
rect 17952 30432 18016 30436
rect 18032 30492 18096 30496
rect 18032 30436 18036 30492
rect 18036 30436 18092 30492
rect 18092 30436 18096 30492
rect 18032 30432 18096 30436
rect 18112 30492 18176 30496
rect 18112 30436 18116 30492
rect 18116 30436 18172 30492
rect 18172 30436 18176 30492
rect 18112 30432 18176 30436
rect 18192 30492 18256 30496
rect 18192 30436 18196 30492
rect 18196 30436 18252 30492
rect 18252 30436 18256 30492
rect 18192 30432 18256 30436
rect 18460 29956 18524 30020
rect 19748 30016 19812 30020
rect 19748 29960 19798 30016
rect 19798 29960 19812 30016
rect 19748 29956 19812 29960
rect 2952 29948 3016 29952
rect 2952 29892 2956 29948
rect 2956 29892 3012 29948
rect 3012 29892 3016 29948
rect 2952 29888 3016 29892
rect 3032 29948 3096 29952
rect 3032 29892 3036 29948
rect 3036 29892 3092 29948
rect 3092 29892 3096 29948
rect 3032 29888 3096 29892
rect 3112 29948 3176 29952
rect 3112 29892 3116 29948
rect 3116 29892 3172 29948
rect 3172 29892 3176 29948
rect 3112 29888 3176 29892
rect 3192 29948 3256 29952
rect 3192 29892 3196 29948
rect 3196 29892 3252 29948
rect 3252 29892 3256 29948
rect 3192 29888 3256 29892
rect 12952 29948 13016 29952
rect 12952 29892 12956 29948
rect 12956 29892 13012 29948
rect 13012 29892 13016 29948
rect 12952 29888 13016 29892
rect 13032 29948 13096 29952
rect 13032 29892 13036 29948
rect 13036 29892 13092 29948
rect 13092 29892 13096 29948
rect 13032 29888 13096 29892
rect 13112 29948 13176 29952
rect 13112 29892 13116 29948
rect 13116 29892 13172 29948
rect 13172 29892 13176 29948
rect 13112 29888 13176 29892
rect 13192 29948 13256 29952
rect 13192 29892 13196 29948
rect 13196 29892 13252 29948
rect 13252 29892 13256 29948
rect 13192 29888 13256 29892
rect 22952 29948 23016 29952
rect 22952 29892 22956 29948
rect 22956 29892 23012 29948
rect 23012 29892 23016 29948
rect 22952 29888 23016 29892
rect 23032 29948 23096 29952
rect 23032 29892 23036 29948
rect 23036 29892 23092 29948
rect 23092 29892 23096 29948
rect 23032 29888 23096 29892
rect 23112 29948 23176 29952
rect 23112 29892 23116 29948
rect 23116 29892 23172 29948
rect 23172 29892 23176 29948
rect 23112 29888 23176 29892
rect 23192 29948 23256 29952
rect 23192 29892 23196 29948
rect 23196 29892 23252 29948
rect 23252 29892 23256 29948
rect 23192 29888 23256 29892
rect 16804 29472 16868 29476
rect 16804 29416 16818 29472
rect 16818 29416 16868 29472
rect 16804 29412 16868 29416
rect 7952 29404 8016 29408
rect 7952 29348 7956 29404
rect 7956 29348 8012 29404
rect 8012 29348 8016 29404
rect 7952 29344 8016 29348
rect 8032 29404 8096 29408
rect 8032 29348 8036 29404
rect 8036 29348 8092 29404
rect 8092 29348 8096 29404
rect 8032 29344 8096 29348
rect 8112 29404 8176 29408
rect 8112 29348 8116 29404
rect 8116 29348 8172 29404
rect 8172 29348 8176 29404
rect 8112 29344 8176 29348
rect 8192 29404 8256 29408
rect 8192 29348 8196 29404
rect 8196 29348 8252 29404
rect 8252 29348 8256 29404
rect 8192 29344 8256 29348
rect 17952 29404 18016 29408
rect 17952 29348 17956 29404
rect 17956 29348 18012 29404
rect 18012 29348 18016 29404
rect 17952 29344 18016 29348
rect 18032 29404 18096 29408
rect 18032 29348 18036 29404
rect 18036 29348 18092 29404
rect 18092 29348 18096 29404
rect 18032 29344 18096 29348
rect 18112 29404 18176 29408
rect 18112 29348 18116 29404
rect 18116 29348 18172 29404
rect 18172 29348 18176 29404
rect 18112 29344 18176 29348
rect 18192 29404 18256 29408
rect 18192 29348 18196 29404
rect 18196 29348 18252 29404
rect 18252 29348 18256 29404
rect 18192 29344 18256 29348
rect 15884 29276 15948 29340
rect 15332 29004 15396 29068
rect 16252 29004 16316 29068
rect 2952 28860 3016 28864
rect 2952 28804 2956 28860
rect 2956 28804 3012 28860
rect 3012 28804 3016 28860
rect 2952 28800 3016 28804
rect 3032 28860 3096 28864
rect 3032 28804 3036 28860
rect 3036 28804 3092 28860
rect 3092 28804 3096 28860
rect 3032 28800 3096 28804
rect 3112 28860 3176 28864
rect 3112 28804 3116 28860
rect 3116 28804 3172 28860
rect 3172 28804 3176 28860
rect 3112 28800 3176 28804
rect 3192 28860 3256 28864
rect 3192 28804 3196 28860
rect 3196 28804 3252 28860
rect 3252 28804 3256 28860
rect 3192 28800 3256 28804
rect 12952 28860 13016 28864
rect 12952 28804 12956 28860
rect 12956 28804 13012 28860
rect 13012 28804 13016 28860
rect 12952 28800 13016 28804
rect 13032 28860 13096 28864
rect 13032 28804 13036 28860
rect 13036 28804 13092 28860
rect 13092 28804 13096 28860
rect 13032 28800 13096 28804
rect 13112 28860 13176 28864
rect 13112 28804 13116 28860
rect 13116 28804 13172 28860
rect 13172 28804 13176 28860
rect 13112 28800 13176 28804
rect 13192 28860 13256 28864
rect 13192 28804 13196 28860
rect 13196 28804 13252 28860
rect 13252 28804 13256 28860
rect 13192 28800 13256 28804
rect 22952 28860 23016 28864
rect 22952 28804 22956 28860
rect 22956 28804 23012 28860
rect 23012 28804 23016 28860
rect 22952 28800 23016 28804
rect 23032 28860 23096 28864
rect 23032 28804 23036 28860
rect 23036 28804 23092 28860
rect 23092 28804 23096 28860
rect 23032 28800 23096 28804
rect 23112 28860 23176 28864
rect 23112 28804 23116 28860
rect 23116 28804 23172 28860
rect 23172 28804 23176 28860
rect 23112 28800 23176 28804
rect 23192 28860 23256 28864
rect 23192 28804 23196 28860
rect 23196 28804 23252 28860
rect 23252 28804 23256 28860
rect 23192 28800 23256 28804
rect 17356 28384 17420 28388
rect 17356 28328 17370 28384
rect 17370 28328 17420 28384
rect 17356 28324 17420 28328
rect 17540 28324 17604 28388
rect 7952 28316 8016 28320
rect 7952 28260 7956 28316
rect 7956 28260 8012 28316
rect 8012 28260 8016 28316
rect 7952 28256 8016 28260
rect 8032 28316 8096 28320
rect 8032 28260 8036 28316
rect 8036 28260 8092 28316
rect 8092 28260 8096 28316
rect 8032 28256 8096 28260
rect 8112 28316 8176 28320
rect 8112 28260 8116 28316
rect 8116 28260 8172 28316
rect 8172 28260 8176 28316
rect 8112 28256 8176 28260
rect 8192 28316 8256 28320
rect 8192 28260 8196 28316
rect 8196 28260 8252 28316
rect 8252 28260 8256 28316
rect 8192 28256 8256 28260
rect 17952 28316 18016 28320
rect 17952 28260 17956 28316
rect 17956 28260 18012 28316
rect 18012 28260 18016 28316
rect 17952 28256 18016 28260
rect 18032 28316 18096 28320
rect 18032 28260 18036 28316
rect 18036 28260 18092 28316
rect 18092 28260 18096 28316
rect 18032 28256 18096 28260
rect 18112 28316 18176 28320
rect 18112 28260 18116 28316
rect 18116 28260 18172 28316
rect 18172 28260 18176 28316
rect 18112 28256 18176 28260
rect 18192 28316 18256 28320
rect 18192 28260 18196 28316
rect 18196 28260 18252 28316
rect 18252 28260 18256 28316
rect 18192 28256 18256 28260
rect 15700 28188 15764 28252
rect 17724 28248 17788 28252
rect 17724 28192 17738 28248
rect 17738 28192 17788 28248
rect 17724 28188 17788 28192
rect 2952 27772 3016 27776
rect 2952 27716 2956 27772
rect 2956 27716 3012 27772
rect 3012 27716 3016 27772
rect 2952 27712 3016 27716
rect 3032 27772 3096 27776
rect 3032 27716 3036 27772
rect 3036 27716 3092 27772
rect 3092 27716 3096 27772
rect 3032 27712 3096 27716
rect 3112 27772 3176 27776
rect 3112 27716 3116 27772
rect 3116 27716 3172 27772
rect 3172 27716 3176 27772
rect 3112 27712 3176 27716
rect 3192 27772 3256 27776
rect 3192 27716 3196 27772
rect 3196 27716 3252 27772
rect 3252 27716 3256 27772
rect 3192 27712 3256 27716
rect 12952 27772 13016 27776
rect 12952 27716 12956 27772
rect 12956 27716 13012 27772
rect 13012 27716 13016 27772
rect 12952 27712 13016 27716
rect 13032 27772 13096 27776
rect 13032 27716 13036 27772
rect 13036 27716 13092 27772
rect 13092 27716 13096 27772
rect 13032 27712 13096 27716
rect 13112 27772 13176 27776
rect 13112 27716 13116 27772
rect 13116 27716 13172 27772
rect 13172 27716 13176 27772
rect 13112 27712 13176 27716
rect 13192 27772 13256 27776
rect 13192 27716 13196 27772
rect 13196 27716 13252 27772
rect 13252 27716 13256 27772
rect 13192 27712 13256 27716
rect 22952 27772 23016 27776
rect 22952 27716 22956 27772
rect 22956 27716 23012 27772
rect 23012 27716 23016 27772
rect 22952 27712 23016 27716
rect 23032 27772 23096 27776
rect 23032 27716 23036 27772
rect 23036 27716 23092 27772
rect 23092 27716 23096 27772
rect 23032 27712 23096 27716
rect 23112 27772 23176 27776
rect 23112 27716 23116 27772
rect 23116 27716 23172 27772
rect 23172 27716 23176 27772
rect 23112 27712 23176 27716
rect 23192 27772 23256 27776
rect 23192 27716 23196 27772
rect 23196 27716 23252 27772
rect 23252 27716 23256 27772
rect 23192 27712 23256 27716
rect 7952 27228 8016 27232
rect 7952 27172 7956 27228
rect 7956 27172 8012 27228
rect 8012 27172 8016 27228
rect 7952 27168 8016 27172
rect 8032 27228 8096 27232
rect 8032 27172 8036 27228
rect 8036 27172 8092 27228
rect 8092 27172 8096 27228
rect 8032 27168 8096 27172
rect 8112 27228 8176 27232
rect 8112 27172 8116 27228
rect 8116 27172 8172 27228
rect 8172 27172 8176 27228
rect 8112 27168 8176 27172
rect 8192 27228 8256 27232
rect 8192 27172 8196 27228
rect 8196 27172 8252 27228
rect 8252 27172 8256 27228
rect 8192 27168 8256 27172
rect 17952 27228 18016 27232
rect 17952 27172 17956 27228
rect 17956 27172 18012 27228
rect 18012 27172 18016 27228
rect 17952 27168 18016 27172
rect 18032 27228 18096 27232
rect 18032 27172 18036 27228
rect 18036 27172 18092 27228
rect 18092 27172 18096 27228
rect 18032 27168 18096 27172
rect 18112 27228 18176 27232
rect 18112 27172 18116 27228
rect 18116 27172 18172 27228
rect 18172 27172 18176 27228
rect 18112 27168 18176 27172
rect 18192 27228 18256 27232
rect 18192 27172 18196 27228
rect 18196 27172 18252 27228
rect 18252 27172 18256 27228
rect 18192 27168 18256 27172
rect 21956 27100 22020 27164
rect 19748 26828 19812 26892
rect 14044 26692 14108 26756
rect 14964 26692 15028 26756
rect 2952 26684 3016 26688
rect 2952 26628 2956 26684
rect 2956 26628 3012 26684
rect 3012 26628 3016 26684
rect 2952 26624 3016 26628
rect 3032 26684 3096 26688
rect 3032 26628 3036 26684
rect 3036 26628 3092 26684
rect 3092 26628 3096 26684
rect 3032 26624 3096 26628
rect 3112 26684 3176 26688
rect 3112 26628 3116 26684
rect 3116 26628 3172 26684
rect 3172 26628 3176 26684
rect 3112 26624 3176 26628
rect 3192 26684 3256 26688
rect 3192 26628 3196 26684
rect 3196 26628 3252 26684
rect 3252 26628 3256 26684
rect 3192 26624 3256 26628
rect 12952 26684 13016 26688
rect 12952 26628 12956 26684
rect 12956 26628 13012 26684
rect 13012 26628 13016 26684
rect 12952 26624 13016 26628
rect 13032 26684 13096 26688
rect 13032 26628 13036 26684
rect 13036 26628 13092 26684
rect 13092 26628 13096 26684
rect 13032 26624 13096 26628
rect 13112 26684 13176 26688
rect 13112 26628 13116 26684
rect 13116 26628 13172 26684
rect 13172 26628 13176 26684
rect 13112 26624 13176 26628
rect 13192 26684 13256 26688
rect 13192 26628 13196 26684
rect 13196 26628 13252 26684
rect 13252 26628 13256 26684
rect 13192 26624 13256 26628
rect 22952 26684 23016 26688
rect 22952 26628 22956 26684
rect 22956 26628 23012 26684
rect 23012 26628 23016 26684
rect 22952 26624 23016 26628
rect 23032 26684 23096 26688
rect 23032 26628 23036 26684
rect 23036 26628 23092 26684
rect 23092 26628 23096 26684
rect 23032 26624 23096 26628
rect 23112 26684 23176 26688
rect 23112 26628 23116 26684
rect 23116 26628 23172 26684
rect 23172 26628 23176 26684
rect 23112 26624 23176 26628
rect 23192 26684 23256 26688
rect 23192 26628 23196 26684
rect 23196 26628 23252 26684
rect 23252 26628 23256 26684
rect 23192 26624 23256 26628
rect 21036 26556 21100 26620
rect 7952 26140 8016 26144
rect 7952 26084 7956 26140
rect 7956 26084 8012 26140
rect 8012 26084 8016 26140
rect 7952 26080 8016 26084
rect 8032 26140 8096 26144
rect 8032 26084 8036 26140
rect 8036 26084 8092 26140
rect 8092 26084 8096 26140
rect 8032 26080 8096 26084
rect 8112 26140 8176 26144
rect 8112 26084 8116 26140
rect 8116 26084 8172 26140
rect 8172 26084 8176 26140
rect 8112 26080 8176 26084
rect 8192 26140 8256 26144
rect 8192 26084 8196 26140
rect 8196 26084 8252 26140
rect 8252 26084 8256 26140
rect 8192 26080 8256 26084
rect 17952 26140 18016 26144
rect 17952 26084 17956 26140
rect 17956 26084 18012 26140
rect 18012 26084 18016 26140
rect 17952 26080 18016 26084
rect 18032 26140 18096 26144
rect 18032 26084 18036 26140
rect 18036 26084 18092 26140
rect 18092 26084 18096 26140
rect 18032 26080 18096 26084
rect 18112 26140 18176 26144
rect 18112 26084 18116 26140
rect 18116 26084 18172 26140
rect 18172 26084 18176 26140
rect 18112 26080 18176 26084
rect 18192 26140 18256 26144
rect 18192 26084 18196 26140
rect 18196 26084 18252 26140
rect 18252 26084 18256 26140
rect 18192 26080 18256 26084
rect 2952 25596 3016 25600
rect 2952 25540 2956 25596
rect 2956 25540 3012 25596
rect 3012 25540 3016 25596
rect 2952 25536 3016 25540
rect 3032 25596 3096 25600
rect 3032 25540 3036 25596
rect 3036 25540 3092 25596
rect 3092 25540 3096 25596
rect 3032 25536 3096 25540
rect 3112 25596 3176 25600
rect 3112 25540 3116 25596
rect 3116 25540 3172 25596
rect 3172 25540 3176 25596
rect 3112 25536 3176 25540
rect 3192 25596 3256 25600
rect 3192 25540 3196 25596
rect 3196 25540 3252 25596
rect 3252 25540 3256 25596
rect 3192 25536 3256 25540
rect 12952 25596 13016 25600
rect 12952 25540 12956 25596
rect 12956 25540 13012 25596
rect 13012 25540 13016 25596
rect 12952 25536 13016 25540
rect 13032 25596 13096 25600
rect 13032 25540 13036 25596
rect 13036 25540 13092 25596
rect 13092 25540 13096 25596
rect 13032 25536 13096 25540
rect 13112 25596 13176 25600
rect 13112 25540 13116 25596
rect 13116 25540 13172 25596
rect 13172 25540 13176 25596
rect 13112 25536 13176 25540
rect 13192 25596 13256 25600
rect 13192 25540 13196 25596
rect 13196 25540 13252 25596
rect 13252 25540 13256 25596
rect 13192 25536 13256 25540
rect 22952 25596 23016 25600
rect 22952 25540 22956 25596
rect 22956 25540 23012 25596
rect 23012 25540 23016 25596
rect 22952 25536 23016 25540
rect 23032 25596 23096 25600
rect 23032 25540 23036 25596
rect 23036 25540 23092 25596
rect 23092 25540 23096 25596
rect 23032 25536 23096 25540
rect 23112 25596 23176 25600
rect 23112 25540 23116 25596
rect 23116 25540 23172 25596
rect 23172 25540 23176 25596
rect 23112 25536 23176 25540
rect 23192 25596 23256 25600
rect 23192 25540 23196 25596
rect 23196 25540 23252 25596
rect 23252 25540 23256 25596
rect 23192 25536 23256 25540
rect 7952 25052 8016 25056
rect 7952 24996 7956 25052
rect 7956 24996 8012 25052
rect 8012 24996 8016 25052
rect 7952 24992 8016 24996
rect 8032 25052 8096 25056
rect 8032 24996 8036 25052
rect 8036 24996 8092 25052
rect 8092 24996 8096 25052
rect 8032 24992 8096 24996
rect 8112 25052 8176 25056
rect 8112 24996 8116 25052
rect 8116 24996 8172 25052
rect 8172 24996 8176 25052
rect 8112 24992 8176 24996
rect 8192 25052 8256 25056
rect 8192 24996 8196 25052
rect 8196 24996 8252 25052
rect 8252 24996 8256 25052
rect 8192 24992 8256 24996
rect 17952 25052 18016 25056
rect 17952 24996 17956 25052
rect 17956 24996 18012 25052
rect 18012 24996 18016 25052
rect 17952 24992 18016 24996
rect 18032 25052 18096 25056
rect 18032 24996 18036 25052
rect 18036 24996 18092 25052
rect 18092 24996 18096 25052
rect 18032 24992 18096 24996
rect 18112 25052 18176 25056
rect 18112 24996 18116 25052
rect 18116 24996 18172 25052
rect 18172 24996 18176 25052
rect 18112 24992 18176 24996
rect 18192 25052 18256 25056
rect 18192 24996 18196 25052
rect 18196 24996 18252 25052
rect 18252 24996 18256 25052
rect 18192 24992 18256 24996
rect 9628 24788 9692 24852
rect 2952 24508 3016 24512
rect 2952 24452 2956 24508
rect 2956 24452 3012 24508
rect 3012 24452 3016 24508
rect 2952 24448 3016 24452
rect 3032 24508 3096 24512
rect 3032 24452 3036 24508
rect 3036 24452 3092 24508
rect 3092 24452 3096 24508
rect 3032 24448 3096 24452
rect 3112 24508 3176 24512
rect 3112 24452 3116 24508
rect 3116 24452 3172 24508
rect 3172 24452 3176 24508
rect 3112 24448 3176 24452
rect 3192 24508 3256 24512
rect 3192 24452 3196 24508
rect 3196 24452 3252 24508
rect 3252 24452 3256 24508
rect 3192 24448 3256 24452
rect 12952 24508 13016 24512
rect 12952 24452 12956 24508
rect 12956 24452 13012 24508
rect 13012 24452 13016 24508
rect 12952 24448 13016 24452
rect 13032 24508 13096 24512
rect 13032 24452 13036 24508
rect 13036 24452 13092 24508
rect 13092 24452 13096 24508
rect 13032 24448 13096 24452
rect 13112 24508 13176 24512
rect 13112 24452 13116 24508
rect 13116 24452 13172 24508
rect 13172 24452 13176 24508
rect 13112 24448 13176 24452
rect 13192 24508 13256 24512
rect 13192 24452 13196 24508
rect 13196 24452 13252 24508
rect 13252 24452 13256 24508
rect 13192 24448 13256 24452
rect 22952 24508 23016 24512
rect 22952 24452 22956 24508
rect 22956 24452 23012 24508
rect 23012 24452 23016 24508
rect 22952 24448 23016 24452
rect 23032 24508 23096 24512
rect 23032 24452 23036 24508
rect 23036 24452 23092 24508
rect 23092 24452 23096 24508
rect 23032 24448 23096 24452
rect 23112 24508 23176 24512
rect 23112 24452 23116 24508
rect 23116 24452 23172 24508
rect 23172 24452 23176 24508
rect 23112 24448 23176 24452
rect 23192 24508 23256 24512
rect 23192 24452 23196 24508
rect 23196 24452 23252 24508
rect 23252 24452 23256 24508
rect 23192 24448 23256 24452
rect 7952 23964 8016 23968
rect 7952 23908 7956 23964
rect 7956 23908 8012 23964
rect 8012 23908 8016 23964
rect 7952 23904 8016 23908
rect 8032 23964 8096 23968
rect 8032 23908 8036 23964
rect 8036 23908 8092 23964
rect 8092 23908 8096 23964
rect 8032 23904 8096 23908
rect 8112 23964 8176 23968
rect 8112 23908 8116 23964
rect 8116 23908 8172 23964
rect 8172 23908 8176 23964
rect 8112 23904 8176 23908
rect 8192 23964 8256 23968
rect 8192 23908 8196 23964
rect 8196 23908 8252 23964
rect 8252 23908 8256 23964
rect 8192 23904 8256 23908
rect 17952 23964 18016 23968
rect 17952 23908 17956 23964
rect 17956 23908 18012 23964
rect 18012 23908 18016 23964
rect 17952 23904 18016 23908
rect 18032 23964 18096 23968
rect 18032 23908 18036 23964
rect 18036 23908 18092 23964
rect 18092 23908 18096 23964
rect 18032 23904 18096 23908
rect 18112 23964 18176 23968
rect 18112 23908 18116 23964
rect 18116 23908 18172 23964
rect 18172 23908 18176 23964
rect 18112 23904 18176 23908
rect 18192 23964 18256 23968
rect 18192 23908 18196 23964
rect 18196 23908 18252 23964
rect 18252 23908 18256 23964
rect 18192 23904 18256 23908
rect 18460 23700 18524 23764
rect 2952 23420 3016 23424
rect 2952 23364 2956 23420
rect 2956 23364 3012 23420
rect 3012 23364 3016 23420
rect 2952 23360 3016 23364
rect 3032 23420 3096 23424
rect 3032 23364 3036 23420
rect 3036 23364 3092 23420
rect 3092 23364 3096 23420
rect 3032 23360 3096 23364
rect 3112 23420 3176 23424
rect 3112 23364 3116 23420
rect 3116 23364 3172 23420
rect 3172 23364 3176 23420
rect 3112 23360 3176 23364
rect 3192 23420 3256 23424
rect 3192 23364 3196 23420
rect 3196 23364 3252 23420
rect 3252 23364 3256 23420
rect 3192 23360 3256 23364
rect 12952 23420 13016 23424
rect 12952 23364 12956 23420
rect 12956 23364 13012 23420
rect 13012 23364 13016 23420
rect 12952 23360 13016 23364
rect 13032 23420 13096 23424
rect 13032 23364 13036 23420
rect 13036 23364 13092 23420
rect 13092 23364 13096 23420
rect 13032 23360 13096 23364
rect 13112 23420 13176 23424
rect 13112 23364 13116 23420
rect 13116 23364 13172 23420
rect 13172 23364 13176 23420
rect 13112 23360 13176 23364
rect 13192 23420 13256 23424
rect 13192 23364 13196 23420
rect 13196 23364 13252 23420
rect 13252 23364 13256 23420
rect 13192 23360 13256 23364
rect 22952 23420 23016 23424
rect 22952 23364 22956 23420
rect 22956 23364 23012 23420
rect 23012 23364 23016 23420
rect 22952 23360 23016 23364
rect 23032 23420 23096 23424
rect 23032 23364 23036 23420
rect 23036 23364 23092 23420
rect 23092 23364 23096 23420
rect 23032 23360 23096 23364
rect 23112 23420 23176 23424
rect 23112 23364 23116 23420
rect 23116 23364 23172 23420
rect 23172 23364 23176 23420
rect 23112 23360 23176 23364
rect 23192 23420 23256 23424
rect 23192 23364 23196 23420
rect 23196 23364 23252 23420
rect 23252 23364 23256 23420
rect 23192 23360 23256 23364
rect 7952 22876 8016 22880
rect 7952 22820 7956 22876
rect 7956 22820 8012 22876
rect 8012 22820 8016 22876
rect 7952 22816 8016 22820
rect 8032 22876 8096 22880
rect 8032 22820 8036 22876
rect 8036 22820 8092 22876
rect 8092 22820 8096 22876
rect 8032 22816 8096 22820
rect 8112 22876 8176 22880
rect 8112 22820 8116 22876
rect 8116 22820 8172 22876
rect 8172 22820 8176 22876
rect 8112 22816 8176 22820
rect 8192 22876 8256 22880
rect 8192 22820 8196 22876
rect 8196 22820 8252 22876
rect 8252 22820 8256 22876
rect 8192 22816 8256 22820
rect 17952 22876 18016 22880
rect 17952 22820 17956 22876
rect 17956 22820 18012 22876
rect 18012 22820 18016 22876
rect 17952 22816 18016 22820
rect 18032 22876 18096 22880
rect 18032 22820 18036 22876
rect 18036 22820 18092 22876
rect 18092 22820 18096 22876
rect 18032 22816 18096 22820
rect 18112 22876 18176 22880
rect 18112 22820 18116 22876
rect 18116 22820 18172 22876
rect 18172 22820 18176 22876
rect 18112 22816 18176 22820
rect 18192 22876 18256 22880
rect 18192 22820 18196 22876
rect 18196 22820 18252 22876
rect 18252 22820 18256 22876
rect 18192 22816 18256 22820
rect 2952 22332 3016 22336
rect 2952 22276 2956 22332
rect 2956 22276 3012 22332
rect 3012 22276 3016 22332
rect 2952 22272 3016 22276
rect 3032 22332 3096 22336
rect 3032 22276 3036 22332
rect 3036 22276 3092 22332
rect 3092 22276 3096 22332
rect 3032 22272 3096 22276
rect 3112 22332 3176 22336
rect 3112 22276 3116 22332
rect 3116 22276 3172 22332
rect 3172 22276 3176 22332
rect 3112 22272 3176 22276
rect 3192 22332 3256 22336
rect 3192 22276 3196 22332
rect 3196 22276 3252 22332
rect 3252 22276 3256 22332
rect 3192 22272 3256 22276
rect 12952 22332 13016 22336
rect 12952 22276 12956 22332
rect 12956 22276 13012 22332
rect 13012 22276 13016 22332
rect 12952 22272 13016 22276
rect 13032 22332 13096 22336
rect 13032 22276 13036 22332
rect 13036 22276 13092 22332
rect 13092 22276 13096 22332
rect 13032 22272 13096 22276
rect 13112 22332 13176 22336
rect 13112 22276 13116 22332
rect 13116 22276 13172 22332
rect 13172 22276 13176 22332
rect 13112 22272 13176 22276
rect 13192 22332 13256 22336
rect 13192 22276 13196 22332
rect 13196 22276 13252 22332
rect 13252 22276 13256 22332
rect 13192 22272 13256 22276
rect 22952 22332 23016 22336
rect 22952 22276 22956 22332
rect 22956 22276 23012 22332
rect 23012 22276 23016 22332
rect 22952 22272 23016 22276
rect 23032 22332 23096 22336
rect 23032 22276 23036 22332
rect 23036 22276 23092 22332
rect 23092 22276 23096 22332
rect 23032 22272 23096 22276
rect 23112 22332 23176 22336
rect 23112 22276 23116 22332
rect 23116 22276 23172 22332
rect 23172 22276 23176 22332
rect 23112 22272 23176 22276
rect 23192 22332 23256 22336
rect 23192 22276 23196 22332
rect 23196 22276 23252 22332
rect 23252 22276 23256 22332
rect 23192 22272 23256 22276
rect 21220 22204 21284 22268
rect 7952 21788 8016 21792
rect 7952 21732 7956 21788
rect 7956 21732 8012 21788
rect 8012 21732 8016 21788
rect 7952 21728 8016 21732
rect 8032 21788 8096 21792
rect 8032 21732 8036 21788
rect 8036 21732 8092 21788
rect 8092 21732 8096 21788
rect 8032 21728 8096 21732
rect 8112 21788 8176 21792
rect 8112 21732 8116 21788
rect 8116 21732 8172 21788
rect 8172 21732 8176 21788
rect 8112 21728 8176 21732
rect 8192 21788 8256 21792
rect 8192 21732 8196 21788
rect 8196 21732 8252 21788
rect 8252 21732 8256 21788
rect 8192 21728 8256 21732
rect 17952 21788 18016 21792
rect 17952 21732 17956 21788
rect 17956 21732 18012 21788
rect 18012 21732 18016 21788
rect 17952 21728 18016 21732
rect 18032 21788 18096 21792
rect 18032 21732 18036 21788
rect 18036 21732 18092 21788
rect 18092 21732 18096 21788
rect 18032 21728 18096 21732
rect 18112 21788 18176 21792
rect 18112 21732 18116 21788
rect 18116 21732 18172 21788
rect 18172 21732 18176 21788
rect 18112 21728 18176 21732
rect 18192 21788 18256 21792
rect 18192 21732 18196 21788
rect 18196 21732 18252 21788
rect 18252 21732 18256 21788
rect 18192 21728 18256 21732
rect 2952 21244 3016 21248
rect 2952 21188 2956 21244
rect 2956 21188 3012 21244
rect 3012 21188 3016 21244
rect 2952 21184 3016 21188
rect 3032 21244 3096 21248
rect 3032 21188 3036 21244
rect 3036 21188 3092 21244
rect 3092 21188 3096 21244
rect 3032 21184 3096 21188
rect 3112 21244 3176 21248
rect 3112 21188 3116 21244
rect 3116 21188 3172 21244
rect 3172 21188 3176 21244
rect 3112 21184 3176 21188
rect 3192 21244 3256 21248
rect 3192 21188 3196 21244
rect 3196 21188 3252 21244
rect 3252 21188 3256 21244
rect 3192 21184 3256 21188
rect 12952 21244 13016 21248
rect 12952 21188 12956 21244
rect 12956 21188 13012 21244
rect 13012 21188 13016 21244
rect 12952 21184 13016 21188
rect 13032 21244 13096 21248
rect 13032 21188 13036 21244
rect 13036 21188 13092 21244
rect 13092 21188 13096 21244
rect 13032 21184 13096 21188
rect 13112 21244 13176 21248
rect 13112 21188 13116 21244
rect 13116 21188 13172 21244
rect 13172 21188 13176 21244
rect 13112 21184 13176 21188
rect 13192 21244 13256 21248
rect 13192 21188 13196 21244
rect 13196 21188 13252 21244
rect 13252 21188 13256 21244
rect 13192 21184 13256 21188
rect 22952 21244 23016 21248
rect 22952 21188 22956 21244
rect 22956 21188 23012 21244
rect 23012 21188 23016 21244
rect 22952 21184 23016 21188
rect 23032 21244 23096 21248
rect 23032 21188 23036 21244
rect 23036 21188 23092 21244
rect 23092 21188 23096 21244
rect 23032 21184 23096 21188
rect 23112 21244 23176 21248
rect 23112 21188 23116 21244
rect 23116 21188 23172 21244
rect 23172 21188 23176 21244
rect 23112 21184 23176 21188
rect 23192 21244 23256 21248
rect 23192 21188 23196 21244
rect 23196 21188 23252 21244
rect 23252 21188 23256 21244
rect 23192 21184 23256 21188
rect 16068 21116 16132 21180
rect 7952 20700 8016 20704
rect 7952 20644 7956 20700
rect 7956 20644 8012 20700
rect 8012 20644 8016 20700
rect 7952 20640 8016 20644
rect 8032 20700 8096 20704
rect 8032 20644 8036 20700
rect 8036 20644 8092 20700
rect 8092 20644 8096 20700
rect 8032 20640 8096 20644
rect 8112 20700 8176 20704
rect 8112 20644 8116 20700
rect 8116 20644 8172 20700
rect 8172 20644 8176 20700
rect 8112 20640 8176 20644
rect 8192 20700 8256 20704
rect 8192 20644 8196 20700
rect 8196 20644 8252 20700
rect 8252 20644 8256 20700
rect 8192 20640 8256 20644
rect 17952 20700 18016 20704
rect 17952 20644 17956 20700
rect 17956 20644 18012 20700
rect 18012 20644 18016 20700
rect 17952 20640 18016 20644
rect 18032 20700 18096 20704
rect 18032 20644 18036 20700
rect 18036 20644 18092 20700
rect 18092 20644 18096 20700
rect 18032 20640 18096 20644
rect 18112 20700 18176 20704
rect 18112 20644 18116 20700
rect 18116 20644 18172 20700
rect 18172 20644 18176 20700
rect 18112 20640 18176 20644
rect 18192 20700 18256 20704
rect 18192 20644 18196 20700
rect 18196 20644 18252 20700
rect 18252 20644 18256 20700
rect 18192 20640 18256 20644
rect 20668 20436 20732 20500
rect 2952 20156 3016 20160
rect 2952 20100 2956 20156
rect 2956 20100 3012 20156
rect 3012 20100 3016 20156
rect 2952 20096 3016 20100
rect 3032 20156 3096 20160
rect 3032 20100 3036 20156
rect 3036 20100 3092 20156
rect 3092 20100 3096 20156
rect 3032 20096 3096 20100
rect 3112 20156 3176 20160
rect 3112 20100 3116 20156
rect 3116 20100 3172 20156
rect 3172 20100 3176 20156
rect 3112 20096 3176 20100
rect 3192 20156 3256 20160
rect 3192 20100 3196 20156
rect 3196 20100 3252 20156
rect 3252 20100 3256 20156
rect 3192 20096 3256 20100
rect 12952 20156 13016 20160
rect 12952 20100 12956 20156
rect 12956 20100 13012 20156
rect 13012 20100 13016 20156
rect 12952 20096 13016 20100
rect 13032 20156 13096 20160
rect 13032 20100 13036 20156
rect 13036 20100 13092 20156
rect 13092 20100 13096 20156
rect 13032 20096 13096 20100
rect 13112 20156 13176 20160
rect 13112 20100 13116 20156
rect 13116 20100 13172 20156
rect 13172 20100 13176 20156
rect 13112 20096 13176 20100
rect 13192 20156 13256 20160
rect 13192 20100 13196 20156
rect 13196 20100 13252 20156
rect 13252 20100 13256 20156
rect 13192 20096 13256 20100
rect 22952 20156 23016 20160
rect 22952 20100 22956 20156
rect 22956 20100 23012 20156
rect 23012 20100 23016 20156
rect 22952 20096 23016 20100
rect 23032 20156 23096 20160
rect 23032 20100 23036 20156
rect 23036 20100 23092 20156
rect 23092 20100 23096 20156
rect 23032 20096 23096 20100
rect 23112 20156 23176 20160
rect 23112 20100 23116 20156
rect 23116 20100 23172 20156
rect 23172 20100 23176 20156
rect 23112 20096 23176 20100
rect 23192 20156 23256 20160
rect 23192 20100 23196 20156
rect 23196 20100 23252 20156
rect 23252 20100 23256 20156
rect 23192 20096 23256 20100
rect 7952 19612 8016 19616
rect 7952 19556 7956 19612
rect 7956 19556 8012 19612
rect 8012 19556 8016 19612
rect 7952 19552 8016 19556
rect 8032 19612 8096 19616
rect 8032 19556 8036 19612
rect 8036 19556 8092 19612
rect 8092 19556 8096 19612
rect 8032 19552 8096 19556
rect 8112 19612 8176 19616
rect 8112 19556 8116 19612
rect 8116 19556 8172 19612
rect 8172 19556 8176 19612
rect 8112 19552 8176 19556
rect 8192 19612 8256 19616
rect 8192 19556 8196 19612
rect 8196 19556 8252 19612
rect 8252 19556 8256 19612
rect 8192 19552 8256 19556
rect 17952 19612 18016 19616
rect 17952 19556 17956 19612
rect 17956 19556 18012 19612
rect 18012 19556 18016 19612
rect 17952 19552 18016 19556
rect 18032 19612 18096 19616
rect 18032 19556 18036 19612
rect 18036 19556 18092 19612
rect 18092 19556 18096 19612
rect 18032 19552 18096 19556
rect 18112 19612 18176 19616
rect 18112 19556 18116 19612
rect 18116 19556 18172 19612
rect 18172 19556 18176 19612
rect 18112 19552 18176 19556
rect 18192 19612 18256 19616
rect 18192 19556 18196 19612
rect 18196 19556 18252 19612
rect 18252 19556 18256 19612
rect 18192 19552 18256 19556
rect 9628 19212 9692 19276
rect 13676 19272 13740 19276
rect 13676 19216 13726 19272
rect 13726 19216 13740 19272
rect 13676 19212 13740 19216
rect 2952 19068 3016 19072
rect 2952 19012 2956 19068
rect 2956 19012 3012 19068
rect 3012 19012 3016 19068
rect 2952 19008 3016 19012
rect 3032 19068 3096 19072
rect 3032 19012 3036 19068
rect 3036 19012 3092 19068
rect 3092 19012 3096 19068
rect 3032 19008 3096 19012
rect 3112 19068 3176 19072
rect 3112 19012 3116 19068
rect 3116 19012 3172 19068
rect 3172 19012 3176 19068
rect 3112 19008 3176 19012
rect 3192 19068 3256 19072
rect 3192 19012 3196 19068
rect 3196 19012 3252 19068
rect 3252 19012 3256 19068
rect 3192 19008 3256 19012
rect 12952 19068 13016 19072
rect 12952 19012 12956 19068
rect 12956 19012 13012 19068
rect 13012 19012 13016 19068
rect 12952 19008 13016 19012
rect 13032 19068 13096 19072
rect 13032 19012 13036 19068
rect 13036 19012 13092 19068
rect 13092 19012 13096 19068
rect 13032 19008 13096 19012
rect 13112 19068 13176 19072
rect 13112 19012 13116 19068
rect 13116 19012 13172 19068
rect 13172 19012 13176 19068
rect 13112 19008 13176 19012
rect 13192 19068 13256 19072
rect 13192 19012 13196 19068
rect 13196 19012 13252 19068
rect 13252 19012 13256 19068
rect 13192 19008 13256 19012
rect 22952 19068 23016 19072
rect 22952 19012 22956 19068
rect 22956 19012 23012 19068
rect 23012 19012 23016 19068
rect 22952 19008 23016 19012
rect 23032 19068 23096 19072
rect 23032 19012 23036 19068
rect 23036 19012 23092 19068
rect 23092 19012 23096 19068
rect 23032 19008 23096 19012
rect 23112 19068 23176 19072
rect 23112 19012 23116 19068
rect 23116 19012 23172 19068
rect 23172 19012 23176 19068
rect 23112 19008 23176 19012
rect 23192 19068 23256 19072
rect 23192 19012 23196 19068
rect 23196 19012 23252 19068
rect 23252 19012 23256 19068
rect 23192 19008 23256 19012
rect 15700 18804 15764 18868
rect 17540 18728 17604 18732
rect 17540 18672 17590 18728
rect 17590 18672 17604 18728
rect 17540 18668 17604 18672
rect 19932 18668 19996 18732
rect 14780 18592 14844 18596
rect 14780 18536 14794 18592
rect 14794 18536 14844 18592
rect 14780 18532 14844 18536
rect 7952 18524 8016 18528
rect 7952 18468 7956 18524
rect 7956 18468 8012 18524
rect 8012 18468 8016 18524
rect 7952 18464 8016 18468
rect 8032 18524 8096 18528
rect 8032 18468 8036 18524
rect 8036 18468 8092 18524
rect 8092 18468 8096 18524
rect 8032 18464 8096 18468
rect 8112 18524 8176 18528
rect 8112 18468 8116 18524
rect 8116 18468 8172 18524
rect 8172 18468 8176 18524
rect 8112 18464 8176 18468
rect 8192 18524 8256 18528
rect 8192 18468 8196 18524
rect 8196 18468 8252 18524
rect 8252 18468 8256 18524
rect 8192 18464 8256 18468
rect 17952 18524 18016 18528
rect 17952 18468 17956 18524
rect 17956 18468 18012 18524
rect 18012 18468 18016 18524
rect 17952 18464 18016 18468
rect 18032 18524 18096 18528
rect 18032 18468 18036 18524
rect 18036 18468 18092 18524
rect 18092 18468 18096 18524
rect 18032 18464 18096 18468
rect 18112 18524 18176 18528
rect 18112 18468 18116 18524
rect 18116 18468 18172 18524
rect 18172 18468 18176 18524
rect 18112 18464 18176 18468
rect 18192 18524 18256 18528
rect 18192 18468 18196 18524
rect 18196 18468 18252 18524
rect 18252 18468 18256 18524
rect 18192 18464 18256 18468
rect 12020 18260 12084 18324
rect 2952 17980 3016 17984
rect 2952 17924 2956 17980
rect 2956 17924 3012 17980
rect 3012 17924 3016 17980
rect 2952 17920 3016 17924
rect 3032 17980 3096 17984
rect 3032 17924 3036 17980
rect 3036 17924 3092 17980
rect 3092 17924 3096 17980
rect 3032 17920 3096 17924
rect 3112 17980 3176 17984
rect 3112 17924 3116 17980
rect 3116 17924 3172 17980
rect 3172 17924 3176 17980
rect 3112 17920 3176 17924
rect 3192 17980 3256 17984
rect 3192 17924 3196 17980
rect 3196 17924 3252 17980
rect 3252 17924 3256 17980
rect 3192 17920 3256 17924
rect 12952 17980 13016 17984
rect 12952 17924 12956 17980
rect 12956 17924 13012 17980
rect 13012 17924 13016 17980
rect 12952 17920 13016 17924
rect 13032 17980 13096 17984
rect 13032 17924 13036 17980
rect 13036 17924 13092 17980
rect 13092 17924 13096 17980
rect 13032 17920 13096 17924
rect 13112 17980 13176 17984
rect 13112 17924 13116 17980
rect 13116 17924 13172 17980
rect 13172 17924 13176 17980
rect 13112 17920 13176 17924
rect 13192 17980 13256 17984
rect 13192 17924 13196 17980
rect 13196 17924 13252 17980
rect 13252 17924 13256 17980
rect 13192 17920 13256 17924
rect 22952 17980 23016 17984
rect 22952 17924 22956 17980
rect 22956 17924 23012 17980
rect 23012 17924 23016 17980
rect 22952 17920 23016 17924
rect 23032 17980 23096 17984
rect 23032 17924 23036 17980
rect 23036 17924 23092 17980
rect 23092 17924 23096 17980
rect 23032 17920 23096 17924
rect 23112 17980 23176 17984
rect 23112 17924 23116 17980
rect 23116 17924 23172 17980
rect 23172 17924 23176 17980
rect 23112 17920 23176 17924
rect 23192 17980 23256 17984
rect 23192 17924 23196 17980
rect 23196 17924 23252 17980
rect 23252 17924 23256 17980
rect 23192 17920 23256 17924
rect 7952 17436 8016 17440
rect 7952 17380 7956 17436
rect 7956 17380 8012 17436
rect 8012 17380 8016 17436
rect 7952 17376 8016 17380
rect 8032 17436 8096 17440
rect 8032 17380 8036 17436
rect 8036 17380 8092 17436
rect 8092 17380 8096 17436
rect 8032 17376 8096 17380
rect 8112 17436 8176 17440
rect 8112 17380 8116 17436
rect 8116 17380 8172 17436
rect 8172 17380 8176 17436
rect 8112 17376 8176 17380
rect 8192 17436 8256 17440
rect 8192 17380 8196 17436
rect 8196 17380 8252 17436
rect 8252 17380 8256 17436
rect 8192 17376 8256 17380
rect 17952 17436 18016 17440
rect 17952 17380 17956 17436
rect 17956 17380 18012 17436
rect 18012 17380 18016 17436
rect 17952 17376 18016 17380
rect 18032 17436 18096 17440
rect 18032 17380 18036 17436
rect 18036 17380 18092 17436
rect 18092 17380 18096 17436
rect 18032 17376 18096 17380
rect 18112 17436 18176 17440
rect 18112 17380 18116 17436
rect 18116 17380 18172 17436
rect 18172 17380 18176 17436
rect 18112 17376 18176 17380
rect 18192 17436 18256 17440
rect 18192 17380 18196 17436
rect 18196 17380 18252 17436
rect 18252 17380 18256 17436
rect 18192 17376 18256 17380
rect 2952 16892 3016 16896
rect 2952 16836 2956 16892
rect 2956 16836 3012 16892
rect 3012 16836 3016 16892
rect 2952 16832 3016 16836
rect 3032 16892 3096 16896
rect 3032 16836 3036 16892
rect 3036 16836 3092 16892
rect 3092 16836 3096 16892
rect 3032 16832 3096 16836
rect 3112 16892 3176 16896
rect 3112 16836 3116 16892
rect 3116 16836 3172 16892
rect 3172 16836 3176 16892
rect 3112 16832 3176 16836
rect 3192 16892 3256 16896
rect 3192 16836 3196 16892
rect 3196 16836 3252 16892
rect 3252 16836 3256 16892
rect 3192 16832 3256 16836
rect 12952 16892 13016 16896
rect 12952 16836 12956 16892
rect 12956 16836 13012 16892
rect 13012 16836 13016 16892
rect 12952 16832 13016 16836
rect 13032 16892 13096 16896
rect 13032 16836 13036 16892
rect 13036 16836 13092 16892
rect 13092 16836 13096 16892
rect 13032 16832 13096 16836
rect 13112 16892 13176 16896
rect 13112 16836 13116 16892
rect 13116 16836 13172 16892
rect 13172 16836 13176 16892
rect 13112 16832 13176 16836
rect 13192 16892 13256 16896
rect 13192 16836 13196 16892
rect 13196 16836 13252 16892
rect 13252 16836 13256 16892
rect 13192 16832 13256 16836
rect 22952 16892 23016 16896
rect 22952 16836 22956 16892
rect 22956 16836 23012 16892
rect 23012 16836 23016 16892
rect 22952 16832 23016 16836
rect 23032 16892 23096 16896
rect 23032 16836 23036 16892
rect 23036 16836 23092 16892
rect 23092 16836 23096 16892
rect 23032 16832 23096 16836
rect 23112 16892 23176 16896
rect 23112 16836 23116 16892
rect 23116 16836 23172 16892
rect 23172 16836 23176 16892
rect 23112 16832 23176 16836
rect 23192 16892 23256 16896
rect 23192 16836 23196 16892
rect 23196 16836 23252 16892
rect 23252 16836 23256 16892
rect 23192 16832 23256 16836
rect 12572 16764 12636 16828
rect 20668 16552 20732 16556
rect 20668 16496 20718 16552
rect 20718 16496 20732 16552
rect 20668 16492 20732 16496
rect 21220 16492 21284 16556
rect 7952 16348 8016 16352
rect 7952 16292 7956 16348
rect 7956 16292 8012 16348
rect 8012 16292 8016 16348
rect 7952 16288 8016 16292
rect 8032 16348 8096 16352
rect 8032 16292 8036 16348
rect 8036 16292 8092 16348
rect 8092 16292 8096 16348
rect 8032 16288 8096 16292
rect 8112 16348 8176 16352
rect 8112 16292 8116 16348
rect 8116 16292 8172 16348
rect 8172 16292 8176 16348
rect 8112 16288 8176 16292
rect 8192 16348 8256 16352
rect 8192 16292 8196 16348
rect 8196 16292 8252 16348
rect 8252 16292 8256 16348
rect 8192 16288 8256 16292
rect 17952 16348 18016 16352
rect 17952 16292 17956 16348
rect 17956 16292 18012 16348
rect 18012 16292 18016 16348
rect 17952 16288 18016 16292
rect 18032 16348 18096 16352
rect 18032 16292 18036 16348
rect 18036 16292 18092 16348
rect 18092 16292 18096 16348
rect 18032 16288 18096 16292
rect 18112 16348 18176 16352
rect 18112 16292 18116 16348
rect 18116 16292 18172 16348
rect 18172 16292 18176 16348
rect 18112 16288 18176 16292
rect 18192 16348 18256 16352
rect 18192 16292 18196 16348
rect 18196 16292 18252 16348
rect 18252 16292 18256 16348
rect 18192 16288 18256 16292
rect 16252 16280 16316 16284
rect 16252 16224 16266 16280
rect 16266 16224 16316 16280
rect 16252 16220 16316 16224
rect 2952 15804 3016 15808
rect 2952 15748 2956 15804
rect 2956 15748 3012 15804
rect 3012 15748 3016 15804
rect 2952 15744 3016 15748
rect 3032 15804 3096 15808
rect 3032 15748 3036 15804
rect 3036 15748 3092 15804
rect 3092 15748 3096 15804
rect 3032 15744 3096 15748
rect 3112 15804 3176 15808
rect 3112 15748 3116 15804
rect 3116 15748 3172 15804
rect 3172 15748 3176 15804
rect 3112 15744 3176 15748
rect 3192 15804 3256 15808
rect 3192 15748 3196 15804
rect 3196 15748 3252 15804
rect 3252 15748 3256 15804
rect 3192 15744 3256 15748
rect 12952 15804 13016 15808
rect 12952 15748 12956 15804
rect 12956 15748 13012 15804
rect 13012 15748 13016 15804
rect 12952 15744 13016 15748
rect 13032 15804 13096 15808
rect 13032 15748 13036 15804
rect 13036 15748 13092 15804
rect 13092 15748 13096 15804
rect 13032 15744 13096 15748
rect 13112 15804 13176 15808
rect 13112 15748 13116 15804
rect 13116 15748 13172 15804
rect 13172 15748 13176 15804
rect 13112 15744 13176 15748
rect 13192 15804 13256 15808
rect 13192 15748 13196 15804
rect 13196 15748 13252 15804
rect 13252 15748 13256 15804
rect 13192 15744 13256 15748
rect 22952 15804 23016 15808
rect 22952 15748 22956 15804
rect 22956 15748 23012 15804
rect 23012 15748 23016 15804
rect 22952 15744 23016 15748
rect 23032 15804 23096 15808
rect 23032 15748 23036 15804
rect 23036 15748 23092 15804
rect 23092 15748 23096 15804
rect 23032 15744 23096 15748
rect 23112 15804 23176 15808
rect 23112 15748 23116 15804
rect 23116 15748 23172 15804
rect 23172 15748 23176 15804
rect 23112 15744 23176 15748
rect 23192 15804 23256 15808
rect 23192 15748 23196 15804
rect 23196 15748 23252 15804
rect 23252 15748 23256 15804
rect 23192 15744 23256 15748
rect 14964 15736 15028 15740
rect 14964 15680 15014 15736
rect 15014 15680 15028 15736
rect 14964 15676 15028 15680
rect 7952 15260 8016 15264
rect 7952 15204 7956 15260
rect 7956 15204 8012 15260
rect 8012 15204 8016 15260
rect 7952 15200 8016 15204
rect 8032 15260 8096 15264
rect 8032 15204 8036 15260
rect 8036 15204 8092 15260
rect 8092 15204 8096 15260
rect 8032 15200 8096 15204
rect 8112 15260 8176 15264
rect 8112 15204 8116 15260
rect 8116 15204 8172 15260
rect 8172 15204 8176 15260
rect 8112 15200 8176 15204
rect 8192 15260 8256 15264
rect 8192 15204 8196 15260
rect 8196 15204 8252 15260
rect 8252 15204 8256 15260
rect 8192 15200 8256 15204
rect 17952 15260 18016 15264
rect 17952 15204 17956 15260
rect 17956 15204 18012 15260
rect 18012 15204 18016 15260
rect 17952 15200 18016 15204
rect 18032 15260 18096 15264
rect 18032 15204 18036 15260
rect 18036 15204 18092 15260
rect 18092 15204 18096 15260
rect 18032 15200 18096 15204
rect 18112 15260 18176 15264
rect 18112 15204 18116 15260
rect 18116 15204 18172 15260
rect 18172 15204 18176 15260
rect 18112 15200 18176 15204
rect 18192 15260 18256 15264
rect 18192 15204 18196 15260
rect 18196 15204 18252 15260
rect 18252 15204 18256 15260
rect 18192 15200 18256 15204
rect 15884 15132 15948 15196
rect 2952 14716 3016 14720
rect 2952 14660 2956 14716
rect 2956 14660 3012 14716
rect 3012 14660 3016 14716
rect 2952 14656 3016 14660
rect 3032 14716 3096 14720
rect 3032 14660 3036 14716
rect 3036 14660 3092 14716
rect 3092 14660 3096 14716
rect 3032 14656 3096 14660
rect 3112 14716 3176 14720
rect 3112 14660 3116 14716
rect 3116 14660 3172 14716
rect 3172 14660 3176 14716
rect 3112 14656 3176 14660
rect 3192 14716 3256 14720
rect 3192 14660 3196 14716
rect 3196 14660 3252 14716
rect 3252 14660 3256 14716
rect 3192 14656 3256 14660
rect 12952 14716 13016 14720
rect 12952 14660 12956 14716
rect 12956 14660 13012 14716
rect 13012 14660 13016 14716
rect 12952 14656 13016 14660
rect 13032 14716 13096 14720
rect 13032 14660 13036 14716
rect 13036 14660 13092 14716
rect 13092 14660 13096 14716
rect 13032 14656 13096 14660
rect 13112 14716 13176 14720
rect 13112 14660 13116 14716
rect 13116 14660 13172 14716
rect 13172 14660 13176 14716
rect 13112 14656 13176 14660
rect 13192 14716 13256 14720
rect 13192 14660 13196 14716
rect 13196 14660 13252 14716
rect 13252 14660 13256 14716
rect 13192 14656 13256 14660
rect 22952 14716 23016 14720
rect 22952 14660 22956 14716
rect 22956 14660 23012 14716
rect 23012 14660 23016 14716
rect 22952 14656 23016 14660
rect 23032 14716 23096 14720
rect 23032 14660 23036 14716
rect 23036 14660 23092 14716
rect 23092 14660 23096 14716
rect 23032 14656 23096 14660
rect 23112 14716 23176 14720
rect 23112 14660 23116 14716
rect 23116 14660 23172 14716
rect 23172 14660 23176 14716
rect 23112 14656 23176 14660
rect 23192 14716 23256 14720
rect 23192 14660 23196 14716
rect 23196 14660 23252 14716
rect 23252 14660 23256 14716
rect 23192 14656 23256 14660
rect 18460 14512 18524 14516
rect 18460 14456 18474 14512
rect 18474 14456 18524 14512
rect 18460 14452 18524 14456
rect 7952 14172 8016 14176
rect 7952 14116 7956 14172
rect 7956 14116 8012 14172
rect 8012 14116 8016 14172
rect 7952 14112 8016 14116
rect 8032 14172 8096 14176
rect 8032 14116 8036 14172
rect 8036 14116 8092 14172
rect 8092 14116 8096 14172
rect 8032 14112 8096 14116
rect 8112 14172 8176 14176
rect 8112 14116 8116 14172
rect 8116 14116 8172 14172
rect 8172 14116 8176 14172
rect 8112 14112 8176 14116
rect 8192 14172 8256 14176
rect 8192 14116 8196 14172
rect 8196 14116 8252 14172
rect 8252 14116 8256 14172
rect 8192 14112 8256 14116
rect 17952 14172 18016 14176
rect 17952 14116 17956 14172
rect 17956 14116 18012 14172
rect 18012 14116 18016 14172
rect 17952 14112 18016 14116
rect 18032 14172 18096 14176
rect 18032 14116 18036 14172
rect 18036 14116 18092 14172
rect 18092 14116 18096 14172
rect 18032 14112 18096 14116
rect 18112 14172 18176 14176
rect 18112 14116 18116 14172
rect 18116 14116 18172 14172
rect 18172 14116 18176 14172
rect 18112 14112 18176 14116
rect 18192 14172 18256 14176
rect 18192 14116 18196 14172
rect 18196 14116 18252 14172
rect 18252 14116 18256 14172
rect 18192 14112 18256 14116
rect 17356 14044 17420 14108
rect 2952 13628 3016 13632
rect 2952 13572 2956 13628
rect 2956 13572 3012 13628
rect 3012 13572 3016 13628
rect 2952 13568 3016 13572
rect 3032 13628 3096 13632
rect 3032 13572 3036 13628
rect 3036 13572 3092 13628
rect 3092 13572 3096 13628
rect 3032 13568 3096 13572
rect 3112 13628 3176 13632
rect 3112 13572 3116 13628
rect 3116 13572 3172 13628
rect 3172 13572 3176 13628
rect 3112 13568 3176 13572
rect 3192 13628 3256 13632
rect 3192 13572 3196 13628
rect 3196 13572 3252 13628
rect 3252 13572 3256 13628
rect 3192 13568 3256 13572
rect 12952 13628 13016 13632
rect 12952 13572 12956 13628
rect 12956 13572 13012 13628
rect 13012 13572 13016 13628
rect 12952 13568 13016 13572
rect 13032 13628 13096 13632
rect 13032 13572 13036 13628
rect 13036 13572 13092 13628
rect 13092 13572 13096 13628
rect 13032 13568 13096 13572
rect 13112 13628 13176 13632
rect 13112 13572 13116 13628
rect 13116 13572 13172 13628
rect 13172 13572 13176 13628
rect 13112 13568 13176 13572
rect 13192 13628 13256 13632
rect 13192 13572 13196 13628
rect 13196 13572 13252 13628
rect 13252 13572 13256 13628
rect 13192 13568 13256 13572
rect 22952 13628 23016 13632
rect 22952 13572 22956 13628
rect 22956 13572 23012 13628
rect 23012 13572 23016 13628
rect 22952 13568 23016 13572
rect 23032 13628 23096 13632
rect 23032 13572 23036 13628
rect 23036 13572 23092 13628
rect 23092 13572 23096 13628
rect 23032 13568 23096 13572
rect 23112 13628 23176 13632
rect 23112 13572 23116 13628
rect 23116 13572 23172 13628
rect 23172 13572 23176 13628
rect 23112 13568 23176 13572
rect 23192 13628 23256 13632
rect 23192 13572 23196 13628
rect 23196 13572 23252 13628
rect 23252 13572 23256 13628
rect 23192 13568 23256 13572
rect 13676 13092 13740 13156
rect 7952 13084 8016 13088
rect 7952 13028 7956 13084
rect 7956 13028 8012 13084
rect 8012 13028 8016 13084
rect 7952 13024 8016 13028
rect 8032 13084 8096 13088
rect 8032 13028 8036 13084
rect 8036 13028 8092 13084
rect 8092 13028 8096 13084
rect 8032 13024 8096 13028
rect 8112 13084 8176 13088
rect 8112 13028 8116 13084
rect 8116 13028 8172 13084
rect 8172 13028 8176 13084
rect 8112 13024 8176 13028
rect 8192 13084 8256 13088
rect 8192 13028 8196 13084
rect 8196 13028 8252 13084
rect 8252 13028 8256 13084
rect 8192 13024 8256 13028
rect 17952 13084 18016 13088
rect 17952 13028 17956 13084
rect 17956 13028 18012 13084
rect 18012 13028 18016 13084
rect 17952 13024 18016 13028
rect 18032 13084 18096 13088
rect 18032 13028 18036 13084
rect 18036 13028 18092 13084
rect 18092 13028 18096 13084
rect 18032 13024 18096 13028
rect 18112 13084 18176 13088
rect 18112 13028 18116 13084
rect 18116 13028 18172 13084
rect 18172 13028 18176 13084
rect 18112 13024 18176 13028
rect 18192 13084 18256 13088
rect 18192 13028 18196 13084
rect 18196 13028 18252 13084
rect 18252 13028 18256 13084
rect 18192 13024 18256 13028
rect 2952 12540 3016 12544
rect 2952 12484 2956 12540
rect 2956 12484 3012 12540
rect 3012 12484 3016 12540
rect 2952 12480 3016 12484
rect 3032 12540 3096 12544
rect 3032 12484 3036 12540
rect 3036 12484 3092 12540
rect 3092 12484 3096 12540
rect 3032 12480 3096 12484
rect 3112 12540 3176 12544
rect 3112 12484 3116 12540
rect 3116 12484 3172 12540
rect 3172 12484 3176 12540
rect 3112 12480 3176 12484
rect 3192 12540 3256 12544
rect 3192 12484 3196 12540
rect 3196 12484 3252 12540
rect 3252 12484 3256 12540
rect 3192 12480 3256 12484
rect 12952 12540 13016 12544
rect 12952 12484 12956 12540
rect 12956 12484 13012 12540
rect 13012 12484 13016 12540
rect 12952 12480 13016 12484
rect 13032 12540 13096 12544
rect 13032 12484 13036 12540
rect 13036 12484 13092 12540
rect 13092 12484 13096 12540
rect 13032 12480 13096 12484
rect 13112 12540 13176 12544
rect 13112 12484 13116 12540
rect 13116 12484 13172 12540
rect 13172 12484 13176 12540
rect 13112 12480 13176 12484
rect 13192 12540 13256 12544
rect 13192 12484 13196 12540
rect 13196 12484 13252 12540
rect 13252 12484 13256 12540
rect 13192 12480 13256 12484
rect 22952 12540 23016 12544
rect 22952 12484 22956 12540
rect 22956 12484 23012 12540
rect 23012 12484 23016 12540
rect 22952 12480 23016 12484
rect 23032 12540 23096 12544
rect 23032 12484 23036 12540
rect 23036 12484 23092 12540
rect 23092 12484 23096 12540
rect 23032 12480 23096 12484
rect 23112 12540 23176 12544
rect 23112 12484 23116 12540
rect 23116 12484 23172 12540
rect 23172 12484 23176 12540
rect 23112 12480 23176 12484
rect 23192 12540 23256 12544
rect 23192 12484 23196 12540
rect 23196 12484 23252 12540
rect 23252 12484 23256 12540
rect 23192 12480 23256 12484
rect 7952 11996 8016 12000
rect 7952 11940 7956 11996
rect 7956 11940 8012 11996
rect 8012 11940 8016 11996
rect 7952 11936 8016 11940
rect 8032 11996 8096 12000
rect 8032 11940 8036 11996
rect 8036 11940 8092 11996
rect 8092 11940 8096 11996
rect 8032 11936 8096 11940
rect 8112 11996 8176 12000
rect 8112 11940 8116 11996
rect 8116 11940 8172 11996
rect 8172 11940 8176 11996
rect 8112 11936 8176 11940
rect 8192 11996 8256 12000
rect 8192 11940 8196 11996
rect 8196 11940 8252 11996
rect 8252 11940 8256 11996
rect 8192 11936 8256 11940
rect 17952 11996 18016 12000
rect 17952 11940 17956 11996
rect 17956 11940 18012 11996
rect 18012 11940 18016 11996
rect 17952 11936 18016 11940
rect 18032 11996 18096 12000
rect 18032 11940 18036 11996
rect 18036 11940 18092 11996
rect 18092 11940 18096 11996
rect 18032 11936 18096 11940
rect 18112 11996 18176 12000
rect 18112 11940 18116 11996
rect 18116 11940 18172 11996
rect 18172 11940 18176 11996
rect 18112 11936 18176 11940
rect 18192 11996 18256 12000
rect 18192 11940 18196 11996
rect 18196 11940 18252 11996
rect 18252 11940 18256 11996
rect 18192 11936 18256 11940
rect 2952 11452 3016 11456
rect 2952 11396 2956 11452
rect 2956 11396 3012 11452
rect 3012 11396 3016 11452
rect 2952 11392 3016 11396
rect 3032 11452 3096 11456
rect 3032 11396 3036 11452
rect 3036 11396 3092 11452
rect 3092 11396 3096 11452
rect 3032 11392 3096 11396
rect 3112 11452 3176 11456
rect 3112 11396 3116 11452
rect 3116 11396 3172 11452
rect 3172 11396 3176 11452
rect 3112 11392 3176 11396
rect 3192 11452 3256 11456
rect 3192 11396 3196 11452
rect 3196 11396 3252 11452
rect 3252 11396 3256 11452
rect 3192 11392 3256 11396
rect 12952 11452 13016 11456
rect 12952 11396 12956 11452
rect 12956 11396 13012 11452
rect 13012 11396 13016 11452
rect 12952 11392 13016 11396
rect 13032 11452 13096 11456
rect 13032 11396 13036 11452
rect 13036 11396 13092 11452
rect 13092 11396 13096 11452
rect 13032 11392 13096 11396
rect 13112 11452 13176 11456
rect 13112 11396 13116 11452
rect 13116 11396 13172 11452
rect 13172 11396 13176 11452
rect 13112 11392 13176 11396
rect 13192 11452 13256 11456
rect 13192 11396 13196 11452
rect 13196 11396 13252 11452
rect 13252 11396 13256 11452
rect 13192 11392 13256 11396
rect 22952 11452 23016 11456
rect 22952 11396 22956 11452
rect 22956 11396 23012 11452
rect 23012 11396 23016 11452
rect 22952 11392 23016 11396
rect 23032 11452 23096 11456
rect 23032 11396 23036 11452
rect 23036 11396 23092 11452
rect 23092 11396 23096 11452
rect 23032 11392 23096 11396
rect 23112 11452 23176 11456
rect 23112 11396 23116 11452
rect 23116 11396 23172 11452
rect 23172 11396 23176 11452
rect 23112 11392 23176 11396
rect 23192 11452 23256 11456
rect 23192 11396 23196 11452
rect 23196 11396 23252 11452
rect 23252 11396 23256 11452
rect 23192 11392 23256 11396
rect 15884 11188 15948 11252
rect 7952 10908 8016 10912
rect 7952 10852 7956 10908
rect 7956 10852 8012 10908
rect 8012 10852 8016 10908
rect 7952 10848 8016 10852
rect 8032 10908 8096 10912
rect 8032 10852 8036 10908
rect 8036 10852 8092 10908
rect 8092 10852 8096 10908
rect 8032 10848 8096 10852
rect 8112 10908 8176 10912
rect 8112 10852 8116 10908
rect 8116 10852 8172 10908
rect 8172 10852 8176 10908
rect 8112 10848 8176 10852
rect 8192 10908 8256 10912
rect 8192 10852 8196 10908
rect 8196 10852 8252 10908
rect 8252 10852 8256 10908
rect 8192 10848 8256 10852
rect 17952 10908 18016 10912
rect 17952 10852 17956 10908
rect 17956 10852 18012 10908
rect 18012 10852 18016 10908
rect 17952 10848 18016 10852
rect 18032 10908 18096 10912
rect 18032 10852 18036 10908
rect 18036 10852 18092 10908
rect 18092 10852 18096 10908
rect 18032 10848 18096 10852
rect 18112 10908 18176 10912
rect 18112 10852 18116 10908
rect 18116 10852 18172 10908
rect 18172 10852 18176 10908
rect 18112 10848 18176 10852
rect 18192 10908 18256 10912
rect 18192 10852 18196 10908
rect 18196 10852 18252 10908
rect 18252 10852 18256 10908
rect 18192 10848 18256 10852
rect 2952 10364 3016 10368
rect 2952 10308 2956 10364
rect 2956 10308 3012 10364
rect 3012 10308 3016 10364
rect 2952 10304 3016 10308
rect 3032 10364 3096 10368
rect 3032 10308 3036 10364
rect 3036 10308 3092 10364
rect 3092 10308 3096 10364
rect 3032 10304 3096 10308
rect 3112 10364 3176 10368
rect 3112 10308 3116 10364
rect 3116 10308 3172 10364
rect 3172 10308 3176 10364
rect 3112 10304 3176 10308
rect 3192 10364 3256 10368
rect 3192 10308 3196 10364
rect 3196 10308 3252 10364
rect 3252 10308 3256 10364
rect 3192 10304 3256 10308
rect 12952 10364 13016 10368
rect 12952 10308 12956 10364
rect 12956 10308 13012 10364
rect 13012 10308 13016 10364
rect 12952 10304 13016 10308
rect 13032 10364 13096 10368
rect 13032 10308 13036 10364
rect 13036 10308 13092 10364
rect 13092 10308 13096 10364
rect 13032 10304 13096 10308
rect 13112 10364 13176 10368
rect 13112 10308 13116 10364
rect 13116 10308 13172 10364
rect 13172 10308 13176 10364
rect 13112 10304 13176 10308
rect 13192 10364 13256 10368
rect 13192 10308 13196 10364
rect 13196 10308 13252 10364
rect 13252 10308 13256 10364
rect 13192 10304 13256 10308
rect 22952 10364 23016 10368
rect 22952 10308 22956 10364
rect 22956 10308 23012 10364
rect 23012 10308 23016 10364
rect 22952 10304 23016 10308
rect 23032 10364 23096 10368
rect 23032 10308 23036 10364
rect 23036 10308 23092 10364
rect 23092 10308 23096 10364
rect 23032 10304 23096 10308
rect 23112 10364 23176 10368
rect 23112 10308 23116 10364
rect 23116 10308 23172 10364
rect 23172 10308 23176 10364
rect 23112 10304 23176 10308
rect 23192 10364 23256 10368
rect 23192 10308 23196 10364
rect 23196 10308 23252 10364
rect 23252 10308 23256 10364
rect 23192 10304 23256 10308
rect 7952 9820 8016 9824
rect 7952 9764 7956 9820
rect 7956 9764 8012 9820
rect 8012 9764 8016 9820
rect 7952 9760 8016 9764
rect 8032 9820 8096 9824
rect 8032 9764 8036 9820
rect 8036 9764 8092 9820
rect 8092 9764 8096 9820
rect 8032 9760 8096 9764
rect 8112 9820 8176 9824
rect 8112 9764 8116 9820
rect 8116 9764 8172 9820
rect 8172 9764 8176 9820
rect 8112 9760 8176 9764
rect 8192 9820 8256 9824
rect 8192 9764 8196 9820
rect 8196 9764 8252 9820
rect 8252 9764 8256 9820
rect 8192 9760 8256 9764
rect 17952 9820 18016 9824
rect 17952 9764 17956 9820
rect 17956 9764 18012 9820
rect 18012 9764 18016 9820
rect 17952 9760 18016 9764
rect 18032 9820 18096 9824
rect 18032 9764 18036 9820
rect 18036 9764 18092 9820
rect 18092 9764 18096 9820
rect 18032 9760 18096 9764
rect 18112 9820 18176 9824
rect 18112 9764 18116 9820
rect 18116 9764 18172 9820
rect 18172 9764 18176 9820
rect 18112 9760 18176 9764
rect 18192 9820 18256 9824
rect 18192 9764 18196 9820
rect 18196 9764 18252 9820
rect 18252 9764 18256 9820
rect 18192 9760 18256 9764
rect 2952 9276 3016 9280
rect 2952 9220 2956 9276
rect 2956 9220 3012 9276
rect 3012 9220 3016 9276
rect 2952 9216 3016 9220
rect 3032 9276 3096 9280
rect 3032 9220 3036 9276
rect 3036 9220 3092 9276
rect 3092 9220 3096 9276
rect 3032 9216 3096 9220
rect 3112 9276 3176 9280
rect 3112 9220 3116 9276
rect 3116 9220 3172 9276
rect 3172 9220 3176 9276
rect 3112 9216 3176 9220
rect 3192 9276 3256 9280
rect 3192 9220 3196 9276
rect 3196 9220 3252 9276
rect 3252 9220 3256 9276
rect 3192 9216 3256 9220
rect 12952 9276 13016 9280
rect 12952 9220 12956 9276
rect 12956 9220 13012 9276
rect 13012 9220 13016 9276
rect 12952 9216 13016 9220
rect 13032 9276 13096 9280
rect 13032 9220 13036 9276
rect 13036 9220 13092 9276
rect 13092 9220 13096 9276
rect 13032 9216 13096 9220
rect 13112 9276 13176 9280
rect 13112 9220 13116 9276
rect 13116 9220 13172 9276
rect 13172 9220 13176 9276
rect 13112 9216 13176 9220
rect 13192 9276 13256 9280
rect 13192 9220 13196 9276
rect 13196 9220 13252 9276
rect 13252 9220 13256 9276
rect 13192 9216 13256 9220
rect 22952 9276 23016 9280
rect 22952 9220 22956 9276
rect 22956 9220 23012 9276
rect 23012 9220 23016 9276
rect 22952 9216 23016 9220
rect 23032 9276 23096 9280
rect 23032 9220 23036 9276
rect 23036 9220 23092 9276
rect 23092 9220 23096 9276
rect 23032 9216 23096 9220
rect 23112 9276 23176 9280
rect 23112 9220 23116 9276
rect 23116 9220 23172 9276
rect 23172 9220 23176 9276
rect 23112 9216 23176 9220
rect 23192 9276 23256 9280
rect 23192 9220 23196 9276
rect 23196 9220 23252 9276
rect 23252 9220 23256 9276
rect 23192 9216 23256 9220
rect 7952 8732 8016 8736
rect 7952 8676 7956 8732
rect 7956 8676 8012 8732
rect 8012 8676 8016 8732
rect 7952 8672 8016 8676
rect 8032 8732 8096 8736
rect 8032 8676 8036 8732
rect 8036 8676 8092 8732
rect 8092 8676 8096 8732
rect 8032 8672 8096 8676
rect 8112 8732 8176 8736
rect 8112 8676 8116 8732
rect 8116 8676 8172 8732
rect 8172 8676 8176 8732
rect 8112 8672 8176 8676
rect 8192 8732 8256 8736
rect 8192 8676 8196 8732
rect 8196 8676 8252 8732
rect 8252 8676 8256 8732
rect 8192 8672 8256 8676
rect 17952 8732 18016 8736
rect 17952 8676 17956 8732
rect 17956 8676 18012 8732
rect 18012 8676 18016 8732
rect 17952 8672 18016 8676
rect 18032 8732 18096 8736
rect 18032 8676 18036 8732
rect 18036 8676 18092 8732
rect 18092 8676 18096 8732
rect 18032 8672 18096 8676
rect 18112 8732 18176 8736
rect 18112 8676 18116 8732
rect 18116 8676 18172 8732
rect 18172 8676 18176 8732
rect 18112 8672 18176 8676
rect 18192 8732 18256 8736
rect 18192 8676 18196 8732
rect 18196 8676 18252 8732
rect 18252 8676 18256 8732
rect 18192 8672 18256 8676
rect 2952 8188 3016 8192
rect 2952 8132 2956 8188
rect 2956 8132 3012 8188
rect 3012 8132 3016 8188
rect 2952 8128 3016 8132
rect 3032 8188 3096 8192
rect 3032 8132 3036 8188
rect 3036 8132 3092 8188
rect 3092 8132 3096 8188
rect 3032 8128 3096 8132
rect 3112 8188 3176 8192
rect 3112 8132 3116 8188
rect 3116 8132 3172 8188
rect 3172 8132 3176 8188
rect 3112 8128 3176 8132
rect 3192 8188 3256 8192
rect 3192 8132 3196 8188
rect 3196 8132 3252 8188
rect 3252 8132 3256 8188
rect 3192 8128 3256 8132
rect 12952 8188 13016 8192
rect 12952 8132 12956 8188
rect 12956 8132 13012 8188
rect 13012 8132 13016 8188
rect 12952 8128 13016 8132
rect 13032 8188 13096 8192
rect 13032 8132 13036 8188
rect 13036 8132 13092 8188
rect 13092 8132 13096 8188
rect 13032 8128 13096 8132
rect 13112 8188 13176 8192
rect 13112 8132 13116 8188
rect 13116 8132 13172 8188
rect 13172 8132 13176 8188
rect 13112 8128 13176 8132
rect 13192 8188 13256 8192
rect 13192 8132 13196 8188
rect 13196 8132 13252 8188
rect 13252 8132 13256 8188
rect 13192 8128 13256 8132
rect 22952 8188 23016 8192
rect 22952 8132 22956 8188
rect 22956 8132 23012 8188
rect 23012 8132 23016 8188
rect 22952 8128 23016 8132
rect 23032 8188 23096 8192
rect 23032 8132 23036 8188
rect 23036 8132 23092 8188
rect 23092 8132 23096 8188
rect 23032 8128 23096 8132
rect 23112 8188 23176 8192
rect 23112 8132 23116 8188
rect 23116 8132 23172 8188
rect 23172 8132 23176 8188
rect 23112 8128 23176 8132
rect 23192 8188 23256 8192
rect 23192 8132 23196 8188
rect 23196 8132 23252 8188
rect 23252 8132 23256 8188
rect 23192 8128 23256 8132
rect 14780 7924 14844 7988
rect 7952 7644 8016 7648
rect 7952 7588 7956 7644
rect 7956 7588 8012 7644
rect 8012 7588 8016 7644
rect 7952 7584 8016 7588
rect 8032 7644 8096 7648
rect 8032 7588 8036 7644
rect 8036 7588 8092 7644
rect 8092 7588 8096 7644
rect 8032 7584 8096 7588
rect 8112 7644 8176 7648
rect 8112 7588 8116 7644
rect 8116 7588 8172 7644
rect 8172 7588 8176 7644
rect 8112 7584 8176 7588
rect 8192 7644 8256 7648
rect 8192 7588 8196 7644
rect 8196 7588 8252 7644
rect 8252 7588 8256 7644
rect 8192 7584 8256 7588
rect 17952 7644 18016 7648
rect 17952 7588 17956 7644
rect 17956 7588 18012 7644
rect 18012 7588 18016 7644
rect 17952 7584 18016 7588
rect 18032 7644 18096 7648
rect 18032 7588 18036 7644
rect 18036 7588 18092 7644
rect 18092 7588 18096 7644
rect 18032 7584 18096 7588
rect 18112 7644 18176 7648
rect 18112 7588 18116 7644
rect 18116 7588 18172 7644
rect 18172 7588 18176 7644
rect 18112 7584 18176 7588
rect 18192 7644 18256 7648
rect 18192 7588 18196 7644
rect 18196 7588 18252 7644
rect 18252 7588 18256 7644
rect 18192 7584 18256 7588
rect 2952 7100 3016 7104
rect 2952 7044 2956 7100
rect 2956 7044 3012 7100
rect 3012 7044 3016 7100
rect 2952 7040 3016 7044
rect 3032 7100 3096 7104
rect 3032 7044 3036 7100
rect 3036 7044 3092 7100
rect 3092 7044 3096 7100
rect 3032 7040 3096 7044
rect 3112 7100 3176 7104
rect 3112 7044 3116 7100
rect 3116 7044 3172 7100
rect 3172 7044 3176 7100
rect 3112 7040 3176 7044
rect 3192 7100 3256 7104
rect 3192 7044 3196 7100
rect 3196 7044 3252 7100
rect 3252 7044 3256 7100
rect 3192 7040 3256 7044
rect 12952 7100 13016 7104
rect 12952 7044 12956 7100
rect 12956 7044 13012 7100
rect 13012 7044 13016 7100
rect 12952 7040 13016 7044
rect 13032 7100 13096 7104
rect 13032 7044 13036 7100
rect 13036 7044 13092 7100
rect 13092 7044 13096 7100
rect 13032 7040 13096 7044
rect 13112 7100 13176 7104
rect 13112 7044 13116 7100
rect 13116 7044 13172 7100
rect 13172 7044 13176 7100
rect 13112 7040 13176 7044
rect 13192 7100 13256 7104
rect 13192 7044 13196 7100
rect 13196 7044 13252 7100
rect 13252 7044 13256 7100
rect 13192 7040 13256 7044
rect 22952 7100 23016 7104
rect 22952 7044 22956 7100
rect 22956 7044 23012 7100
rect 23012 7044 23016 7100
rect 22952 7040 23016 7044
rect 23032 7100 23096 7104
rect 23032 7044 23036 7100
rect 23036 7044 23092 7100
rect 23092 7044 23096 7100
rect 23032 7040 23096 7044
rect 23112 7100 23176 7104
rect 23112 7044 23116 7100
rect 23116 7044 23172 7100
rect 23172 7044 23176 7100
rect 23112 7040 23176 7044
rect 23192 7100 23256 7104
rect 23192 7044 23196 7100
rect 23196 7044 23252 7100
rect 23252 7044 23256 7100
rect 23192 7040 23256 7044
rect 7952 6556 8016 6560
rect 7952 6500 7956 6556
rect 7956 6500 8012 6556
rect 8012 6500 8016 6556
rect 7952 6496 8016 6500
rect 8032 6556 8096 6560
rect 8032 6500 8036 6556
rect 8036 6500 8092 6556
rect 8092 6500 8096 6556
rect 8032 6496 8096 6500
rect 8112 6556 8176 6560
rect 8112 6500 8116 6556
rect 8116 6500 8172 6556
rect 8172 6500 8176 6556
rect 8112 6496 8176 6500
rect 8192 6556 8256 6560
rect 8192 6500 8196 6556
rect 8196 6500 8252 6556
rect 8252 6500 8256 6556
rect 8192 6496 8256 6500
rect 17952 6556 18016 6560
rect 17952 6500 17956 6556
rect 17956 6500 18012 6556
rect 18012 6500 18016 6556
rect 17952 6496 18016 6500
rect 18032 6556 18096 6560
rect 18032 6500 18036 6556
rect 18036 6500 18092 6556
rect 18092 6500 18096 6556
rect 18032 6496 18096 6500
rect 18112 6556 18176 6560
rect 18112 6500 18116 6556
rect 18116 6500 18172 6556
rect 18172 6500 18176 6556
rect 18112 6496 18176 6500
rect 18192 6556 18256 6560
rect 18192 6500 18196 6556
rect 18196 6500 18252 6556
rect 18252 6500 18256 6556
rect 18192 6496 18256 6500
rect 2952 6012 3016 6016
rect 2952 5956 2956 6012
rect 2956 5956 3012 6012
rect 3012 5956 3016 6012
rect 2952 5952 3016 5956
rect 3032 6012 3096 6016
rect 3032 5956 3036 6012
rect 3036 5956 3092 6012
rect 3092 5956 3096 6012
rect 3032 5952 3096 5956
rect 3112 6012 3176 6016
rect 3112 5956 3116 6012
rect 3116 5956 3172 6012
rect 3172 5956 3176 6012
rect 3112 5952 3176 5956
rect 3192 6012 3256 6016
rect 3192 5956 3196 6012
rect 3196 5956 3252 6012
rect 3252 5956 3256 6012
rect 3192 5952 3256 5956
rect 12952 6012 13016 6016
rect 12952 5956 12956 6012
rect 12956 5956 13012 6012
rect 13012 5956 13016 6012
rect 12952 5952 13016 5956
rect 13032 6012 13096 6016
rect 13032 5956 13036 6012
rect 13036 5956 13092 6012
rect 13092 5956 13096 6012
rect 13032 5952 13096 5956
rect 13112 6012 13176 6016
rect 13112 5956 13116 6012
rect 13116 5956 13172 6012
rect 13172 5956 13176 6012
rect 13112 5952 13176 5956
rect 13192 6012 13256 6016
rect 13192 5956 13196 6012
rect 13196 5956 13252 6012
rect 13252 5956 13256 6012
rect 13192 5952 13256 5956
rect 22952 6012 23016 6016
rect 22952 5956 22956 6012
rect 22956 5956 23012 6012
rect 23012 5956 23016 6012
rect 22952 5952 23016 5956
rect 23032 6012 23096 6016
rect 23032 5956 23036 6012
rect 23036 5956 23092 6012
rect 23092 5956 23096 6012
rect 23032 5952 23096 5956
rect 23112 6012 23176 6016
rect 23112 5956 23116 6012
rect 23116 5956 23172 6012
rect 23172 5956 23176 6012
rect 23112 5952 23176 5956
rect 23192 6012 23256 6016
rect 23192 5956 23196 6012
rect 23196 5956 23252 6012
rect 23252 5956 23256 6012
rect 23192 5952 23256 5956
rect 7952 5468 8016 5472
rect 7952 5412 7956 5468
rect 7956 5412 8012 5468
rect 8012 5412 8016 5468
rect 7952 5408 8016 5412
rect 8032 5468 8096 5472
rect 8032 5412 8036 5468
rect 8036 5412 8092 5468
rect 8092 5412 8096 5468
rect 8032 5408 8096 5412
rect 8112 5468 8176 5472
rect 8112 5412 8116 5468
rect 8116 5412 8172 5468
rect 8172 5412 8176 5468
rect 8112 5408 8176 5412
rect 8192 5468 8256 5472
rect 8192 5412 8196 5468
rect 8196 5412 8252 5468
rect 8252 5412 8256 5468
rect 8192 5408 8256 5412
rect 17952 5468 18016 5472
rect 17952 5412 17956 5468
rect 17956 5412 18012 5468
rect 18012 5412 18016 5468
rect 17952 5408 18016 5412
rect 18032 5468 18096 5472
rect 18032 5412 18036 5468
rect 18036 5412 18092 5468
rect 18092 5412 18096 5468
rect 18032 5408 18096 5412
rect 18112 5468 18176 5472
rect 18112 5412 18116 5468
rect 18116 5412 18172 5468
rect 18172 5412 18176 5468
rect 18112 5408 18176 5412
rect 18192 5468 18256 5472
rect 18192 5412 18196 5468
rect 18196 5412 18252 5468
rect 18252 5412 18256 5468
rect 18192 5408 18256 5412
rect 2952 4924 3016 4928
rect 2952 4868 2956 4924
rect 2956 4868 3012 4924
rect 3012 4868 3016 4924
rect 2952 4864 3016 4868
rect 3032 4924 3096 4928
rect 3032 4868 3036 4924
rect 3036 4868 3092 4924
rect 3092 4868 3096 4924
rect 3032 4864 3096 4868
rect 3112 4924 3176 4928
rect 3112 4868 3116 4924
rect 3116 4868 3172 4924
rect 3172 4868 3176 4924
rect 3112 4864 3176 4868
rect 3192 4924 3256 4928
rect 3192 4868 3196 4924
rect 3196 4868 3252 4924
rect 3252 4868 3256 4924
rect 3192 4864 3256 4868
rect 12952 4924 13016 4928
rect 12952 4868 12956 4924
rect 12956 4868 13012 4924
rect 13012 4868 13016 4924
rect 12952 4864 13016 4868
rect 13032 4924 13096 4928
rect 13032 4868 13036 4924
rect 13036 4868 13092 4924
rect 13092 4868 13096 4924
rect 13032 4864 13096 4868
rect 13112 4924 13176 4928
rect 13112 4868 13116 4924
rect 13116 4868 13172 4924
rect 13172 4868 13176 4924
rect 13112 4864 13176 4868
rect 13192 4924 13256 4928
rect 13192 4868 13196 4924
rect 13196 4868 13252 4924
rect 13252 4868 13256 4924
rect 13192 4864 13256 4868
rect 22952 4924 23016 4928
rect 22952 4868 22956 4924
rect 22956 4868 23012 4924
rect 23012 4868 23016 4924
rect 22952 4864 23016 4868
rect 23032 4924 23096 4928
rect 23032 4868 23036 4924
rect 23036 4868 23092 4924
rect 23092 4868 23096 4924
rect 23032 4864 23096 4868
rect 23112 4924 23176 4928
rect 23112 4868 23116 4924
rect 23116 4868 23172 4924
rect 23172 4868 23176 4924
rect 23112 4864 23176 4868
rect 23192 4924 23256 4928
rect 23192 4868 23196 4924
rect 23196 4868 23252 4924
rect 23252 4868 23256 4924
rect 23192 4864 23256 4868
rect 7952 4380 8016 4384
rect 7952 4324 7956 4380
rect 7956 4324 8012 4380
rect 8012 4324 8016 4380
rect 7952 4320 8016 4324
rect 8032 4380 8096 4384
rect 8032 4324 8036 4380
rect 8036 4324 8092 4380
rect 8092 4324 8096 4380
rect 8032 4320 8096 4324
rect 8112 4380 8176 4384
rect 8112 4324 8116 4380
rect 8116 4324 8172 4380
rect 8172 4324 8176 4380
rect 8112 4320 8176 4324
rect 8192 4380 8256 4384
rect 8192 4324 8196 4380
rect 8196 4324 8252 4380
rect 8252 4324 8256 4380
rect 8192 4320 8256 4324
rect 17952 4380 18016 4384
rect 17952 4324 17956 4380
rect 17956 4324 18012 4380
rect 18012 4324 18016 4380
rect 17952 4320 18016 4324
rect 18032 4380 18096 4384
rect 18032 4324 18036 4380
rect 18036 4324 18092 4380
rect 18092 4324 18096 4380
rect 18032 4320 18096 4324
rect 18112 4380 18176 4384
rect 18112 4324 18116 4380
rect 18116 4324 18172 4380
rect 18172 4324 18176 4380
rect 18112 4320 18176 4324
rect 18192 4380 18256 4384
rect 18192 4324 18196 4380
rect 18196 4324 18252 4380
rect 18252 4324 18256 4380
rect 18192 4320 18256 4324
rect 10180 4116 10244 4180
rect 2952 3836 3016 3840
rect 2952 3780 2956 3836
rect 2956 3780 3012 3836
rect 3012 3780 3016 3836
rect 2952 3776 3016 3780
rect 3032 3836 3096 3840
rect 3032 3780 3036 3836
rect 3036 3780 3092 3836
rect 3092 3780 3096 3836
rect 3032 3776 3096 3780
rect 3112 3836 3176 3840
rect 3112 3780 3116 3836
rect 3116 3780 3172 3836
rect 3172 3780 3176 3836
rect 3112 3776 3176 3780
rect 3192 3836 3256 3840
rect 3192 3780 3196 3836
rect 3196 3780 3252 3836
rect 3252 3780 3256 3836
rect 3192 3776 3256 3780
rect 12952 3836 13016 3840
rect 12952 3780 12956 3836
rect 12956 3780 13012 3836
rect 13012 3780 13016 3836
rect 12952 3776 13016 3780
rect 13032 3836 13096 3840
rect 13032 3780 13036 3836
rect 13036 3780 13092 3836
rect 13092 3780 13096 3836
rect 13032 3776 13096 3780
rect 13112 3836 13176 3840
rect 13112 3780 13116 3836
rect 13116 3780 13172 3836
rect 13172 3780 13176 3836
rect 13112 3776 13176 3780
rect 13192 3836 13256 3840
rect 13192 3780 13196 3836
rect 13196 3780 13252 3836
rect 13252 3780 13256 3836
rect 13192 3776 13256 3780
rect 22952 3836 23016 3840
rect 22952 3780 22956 3836
rect 22956 3780 23012 3836
rect 23012 3780 23016 3836
rect 22952 3776 23016 3780
rect 23032 3836 23096 3840
rect 23032 3780 23036 3836
rect 23036 3780 23092 3836
rect 23092 3780 23096 3836
rect 23032 3776 23096 3780
rect 23112 3836 23176 3840
rect 23112 3780 23116 3836
rect 23116 3780 23172 3836
rect 23172 3780 23176 3836
rect 23112 3776 23176 3780
rect 23192 3836 23256 3840
rect 23192 3780 23196 3836
rect 23196 3780 23252 3836
rect 23252 3780 23256 3836
rect 23192 3776 23256 3780
rect 16804 3436 16868 3500
rect 7952 3292 8016 3296
rect 7952 3236 7956 3292
rect 7956 3236 8012 3292
rect 8012 3236 8016 3292
rect 7952 3232 8016 3236
rect 8032 3292 8096 3296
rect 8032 3236 8036 3292
rect 8036 3236 8092 3292
rect 8092 3236 8096 3292
rect 8032 3232 8096 3236
rect 8112 3292 8176 3296
rect 8112 3236 8116 3292
rect 8116 3236 8172 3292
rect 8172 3236 8176 3292
rect 8112 3232 8176 3236
rect 8192 3292 8256 3296
rect 8192 3236 8196 3292
rect 8196 3236 8252 3292
rect 8252 3236 8256 3292
rect 8192 3232 8256 3236
rect 17952 3292 18016 3296
rect 17952 3236 17956 3292
rect 17956 3236 18012 3292
rect 18012 3236 18016 3292
rect 17952 3232 18016 3236
rect 18032 3292 18096 3296
rect 18032 3236 18036 3292
rect 18036 3236 18092 3292
rect 18092 3236 18096 3292
rect 18032 3232 18096 3236
rect 18112 3292 18176 3296
rect 18112 3236 18116 3292
rect 18116 3236 18172 3292
rect 18172 3236 18176 3292
rect 18112 3232 18176 3236
rect 18192 3292 18256 3296
rect 18192 3236 18196 3292
rect 18196 3236 18252 3292
rect 18252 3236 18256 3292
rect 18192 3232 18256 3236
rect 12020 3164 12084 3228
rect 2952 2748 3016 2752
rect 2952 2692 2956 2748
rect 2956 2692 3012 2748
rect 3012 2692 3016 2748
rect 2952 2688 3016 2692
rect 3032 2748 3096 2752
rect 3032 2692 3036 2748
rect 3036 2692 3092 2748
rect 3092 2692 3096 2748
rect 3032 2688 3096 2692
rect 3112 2748 3176 2752
rect 3112 2692 3116 2748
rect 3116 2692 3172 2748
rect 3172 2692 3176 2748
rect 3112 2688 3176 2692
rect 3192 2748 3256 2752
rect 3192 2692 3196 2748
rect 3196 2692 3252 2748
rect 3252 2692 3256 2748
rect 3192 2688 3256 2692
rect 12952 2748 13016 2752
rect 12952 2692 12956 2748
rect 12956 2692 13012 2748
rect 13012 2692 13016 2748
rect 12952 2688 13016 2692
rect 13032 2748 13096 2752
rect 13032 2692 13036 2748
rect 13036 2692 13092 2748
rect 13092 2692 13096 2748
rect 13032 2688 13096 2692
rect 13112 2748 13176 2752
rect 13112 2692 13116 2748
rect 13116 2692 13172 2748
rect 13172 2692 13176 2748
rect 13112 2688 13176 2692
rect 13192 2748 13256 2752
rect 13192 2692 13196 2748
rect 13196 2692 13252 2748
rect 13252 2692 13256 2748
rect 13192 2688 13256 2692
rect 22952 2748 23016 2752
rect 22952 2692 22956 2748
rect 22956 2692 23012 2748
rect 23012 2692 23016 2748
rect 22952 2688 23016 2692
rect 23032 2748 23096 2752
rect 23032 2692 23036 2748
rect 23036 2692 23092 2748
rect 23092 2692 23096 2748
rect 23032 2688 23096 2692
rect 23112 2748 23176 2752
rect 23112 2692 23116 2748
rect 23116 2692 23172 2748
rect 23172 2692 23176 2748
rect 23112 2688 23176 2692
rect 23192 2748 23256 2752
rect 23192 2692 23196 2748
rect 23196 2692 23252 2748
rect 23252 2692 23256 2748
rect 23192 2688 23256 2692
rect 7952 2204 8016 2208
rect 7952 2148 7956 2204
rect 7956 2148 8012 2204
rect 8012 2148 8016 2204
rect 7952 2144 8016 2148
rect 8032 2204 8096 2208
rect 8032 2148 8036 2204
rect 8036 2148 8092 2204
rect 8092 2148 8096 2204
rect 8032 2144 8096 2148
rect 8112 2204 8176 2208
rect 8112 2148 8116 2204
rect 8116 2148 8172 2204
rect 8172 2148 8176 2204
rect 8112 2144 8176 2148
rect 8192 2204 8256 2208
rect 8192 2148 8196 2204
rect 8196 2148 8252 2204
rect 8252 2148 8256 2204
rect 8192 2144 8256 2148
rect 17952 2204 18016 2208
rect 17952 2148 17956 2204
rect 17956 2148 18012 2204
rect 18012 2148 18016 2204
rect 17952 2144 18016 2148
rect 18032 2204 18096 2208
rect 18032 2148 18036 2204
rect 18036 2148 18092 2204
rect 18092 2148 18096 2204
rect 18032 2144 18096 2148
rect 18112 2204 18176 2208
rect 18112 2148 18116 2204
rect 18116 2148 18172 2204
rect 18172 2148 18176 2204
rect 18112 2144 18176 2148
rect 18192 2204 18256 2208
rect 18192 2148 18196 2204
rect 18196 2148 18252 2204
rect 18252 2148 18256 2204
rect 18192 2144 18256 2148
<< metal4 >>
rect 2944 53888 3264 54448
rect 2944 53824 2952 53888
rect 3016 53824 3032 53888
rect 3096 53824 3112 53888
rect 3176 53824 3192 53888
rect 3256 53824 3264 53888
rect 2944 52800 3264 53824
rect 2944 52736 2952 52800
rect 3016 52736 3032 52800
rect 3096 52736 3112 52800
rect 3176 52736 3192 52800
rect 3256 52736 3264 52800
rect 2944 51712 3264 52736
rect 2944 51648 2952 51712
rect 3016 51648 3032 51712
rect 3096 51648 3112 51712
rect 3176 51648 3192 51712
rect 3256 51648 3264 51712
rect 2944 50624 3264 51648
rect 2944 50560 2952 50624
rect 3016 50560 3032 50624
rect 3096 50560 3112 50624
rect 3176 50560 3192 50624
rect 3256 50560 3264 50624
rect 2944 49536 3264 50560
rect 2944 49472 2952 49536
rect 3016 49472 3032 49536
rect 3096 49472 3112 49536
rect 3176 49472 3192 49536
rect 3256 49472 3264 49536
rect 2944 48448 3264 49472
rect 2944 48384 2952 48448
rect 3016 48384 3032 48448
rect 3096 48384 3112 48448
rect 3176 48384 3192 48448
rect 3256 48384 3264 48448
rect 2944 47360 3264 48384
rect 2944 47296 2952 47360
rect 3016 47296 3032 47360
rect 3096 47296 3112 47360
rect 3176 47296 3192 47360
rect 3256 47296 3264 47360
rect 2944 46272 3264 47296
rect 2944 46208 2952 46272
rect 3016 46208 3032 46272
rect 3096 46208 3112 46272
rect 3176 46208 3192 46272
rect 3256 46208 3264 46272
rect 2944 45184 3264 46208
rect 2944 45120 2952 45184
rect 3016 45120 3032 45184
rect 3096 45120 3112 45184
rect 3176 45120 3192 45184
rect 3256 45120 3264 45184
rect 2944 44096 3264 45120
rect 2944 44032 2952 44096
rect 3016 44032 3032 44096
rect 3096 44032 3112 44096
rect 3176 44032 3192 44096
rect 3256 44032 3264 44096
rect 2944 43008 3264 44032
rect 2944 42944 2952 43008
rect 3016 42944 3032 43008
rect 3096 42944 3112 43008
rect 3176 42944 3192 43008
rect 3256 42944 3264 43008
rect 2944 41920 3264 42944
rect 2944 41856 2952 41920
rect 3016 41856 3032 41920
rect 3096 41856 3112 41920
rect 3176 41856 3192 41920
rect 3256 41856 3264 41920
rect 2944 40832 3264 41856
rect 2944 40768 2952 40832
rect 3016 40768 3032 40832
rect 3096 40768 3112 40832
rect 3176 40768 3192 40832
rect 3256 40768 3264 40832
rect 2944 39744 3264 40768
rect 2944 39680 2952 39744
rect 3016 39680 3032 39744
rect 3096 39680 3112 39744
rect 3176 39680 3192 39744
rect 3256 39680 3264 39744
rect 2944 38656 3264 39680
rect 2944 38592 2952 38656
rect 3016 38592 3032 38656
rect 3096 38592 3112 38656
rect 3176 38592 3192 38656
rect 3256 38592 3264 38656
rect 2944 37568 3264 38592
rect 2944 37504 2952 37568
rect 3016 37504 3032 37568
rect 3096 37504 3112 37568
rect 3176 37504 3192 37568
rect 3256 37504 3264 37568
rect 2944 36480 3264 37504
rect 2944 36416 2952 36480
rect 3016 36416 3032 36480
rect 3096 36416 3112 36480
rect 3176 36416 3192 36480
rect 3256 36416 3264 36480
rect 2944 35392 3264 36416
rect 2944 35328 2952 35392
rect 3016 35328 3032 35392
rect 3096 35328 3112 35392
rect 3176 35328 3192 35392
rect 3256 35328 3264 35392
rect 2944 34304 3264 35328
rect 2944 34240 2952 34304
rect 3016 34240 3032 34304
rect 3096 34240 3112 34304
rect 3176 34240 3192 34304
rect 3256 34240 3264 34304
rect 2944 33216 3264 34240
rect 2944 33152 2952 33216
rect 3016 33152 3032 33216
rect 3096 33152 3112 33216
rect 3176 33152 3192 33216
rect 3256 33152 3264 33216
rect 2944 32128 3264 33152
rect 2944 32064 2952 32128
rect 3016 32064 3032 32128
rect 3096 32064 3112 32128
rect 3176 32064 3192 32128
rect 3256 32064 3264 32128
rect 2944 31040 3264 32064
rect 2944 30976 2952 31040
rect 3016 30976 3032 31040
rect 3096 30976 3112 31040
rect 3176 30976 3192 31040
rect 3256 30976 3264 31040
rect 2944 29952 3264 30976
rect 2944 29888 2952 29952
rect 3016 29888 3032 29952
rect 3096 29888 3112 29952
rect 3176 29888 3192 29952
rect 3256 29888 3264 29952
rect 2944 28864 3264 29888
rect 2944 28800 2952 28864
rect 3016 28800 3032 28864
rect 3096 28800 3112 28864
rect 3176 28800 3192 28864
rect 3256 28800 3264 28864
rect 2944 27776 3264 28800
rect 2944 27712 2952 27776
rect 3016 27712 3032 27776
rect 3096 27712 3112 27776
rect 3176 27712 3192 27776
rect 3256 27712 3264 27776
rect 2944 26688 3264 27712
rect 2944 26624 2952 26688
rect 3016 26624 3032 26688
rect 3096 26624 3112 26688
rect 3176 26624 3192 26688
rect 3256 26624 3264 26688
rect 2944 25600 3264 26624
rect 2944 25536 2952 25600
rect 3016 25536 3032 25600
rect 3096 25536 3112 25600
rect 3176 25536 3192 25600
rect 3256 25536 3264 25600
rect 2944 24512 3264 25536
rect 2944 24448 2952 24512
rect 3016 24448 3032 24512
rect 3096 24448 3112 24512
rect 3176 24448 3192 24512
rect 3256 24448 3264 24512
rect 2944 23424 3264 24448
rect 2944 23360 2952 23424
rect 3016 23360 3032 23424
rect 3096 23360 3112 23424
rect 3176 23360 3192 23424
rect 3256 23360 3264 23424
rect 2944 22336 3264 23360
rect 2944 22272 2952 22336
rect 3016 22272 3032 22336
rect 3096 22272 3112 22336
rect 3176 22272 3192 22336
rect 3256 22272 3264 22336
rect 2944 21248 3264 22272
rect 2944 21184 2952 21248
rect 3016 21184 3032 21248
rect 3096 21184 3112 21248
rect 3176 21184 3192 21248
rect 3256 21184 3264 21248
rect 2944 20160 3264 21184
rect 2944 20096 2952 20160
rect 3016 20096 3032 20160
rect 3096 20096 3112 20160
rect 3176 20096 3192 20160
rect 3256 20096 3264 20160
rect 2944 19072 3264 20096
rect 2944 19008 2952 19072
rect 3016 19008 3032 19072
rect 3096 19008 3112 19072
rect 3176 19008 3192 19072
rect 3256 19008 3264 19072
rect 2944 17984 3264 19008
rect 2944 17920 2952 17984
rect 3016 17920 3032 17984
rect 3096 17920 3112 17984
rect 3176 17920 3192 17984
rect 3256 17920 3264 17984
rect 2944 16896 3264 17920
rect 2944 16832 2952 16896
rect 3016 16832 3032 16896
rect 3096 16832 3112 16896
rect 3176 16832 3192 16896
rect 3256 16832 3264 16896
rect 2944 15808 3264 16832
rect 2944 15744 2952 15808
rect 3016 15744 3032 15808
rect 3096 15744 3112 15808
rect 3176 15744 3192 15808
rect 3256 15744 3264 15808
rect 2944 14720 3264 15744
rect 2944 14656 2952 14720
rect 3016 14656 3032 14720
rect 3096 14656 3112 14720
rect 3176 14656 3192 14720
rect 3256 14656 3264 14720
rect 2944 13632 3264 14656
rect 2944 13568 2952 13632
rect 3016 13568 3032 13632
rect 3096 13568 3112 13632
rect 3176 13568 3192 13632
rect 3256 13568 3264 13632
rect 2944 12544 3264 13568
rect 2944 12480 2952 12544
rect 3016 12480 3032 12544
rect 3096 12480 3112 12544
rect 3176 12480 3192 12544
rect 3256 12480 3264 12544
rect 2944 11456 3264 12480
rect 2944 11392 2952 11456
rect 3016 11392 3032 11456
rect 3096 11392 3112 11456
rect 3176 11392 3192 11456
rect 3256 11392 3264 11456
rect 2944 10368 3264 11392
rect 2944 10304 2952 10368
rect 3016 10304 3032 10368
rect 3096 10304 3112 10368
rect 3176 10304 3192 10368
rect 3256 10304 3264 10368
rect 2944 9280 3264 10304
rect 2944 9216 2952 9280
rect 3016 9216 3032 9280
rect 3096 9216 3112 9280
rect 3176 9216 3192 9280
rect 3256 9216 3264 9280
rect 2944 8192 3264 9216
rect 2944 8128 2952 8192
rect 3016 8128 3032 8192
rect 3096 8128 3112 8192
rect 3176 8128 3192 8192
rect 3256 8128 3264 8192
rect 2944 7104 3264 8128
rect 2944 7040 2952 7104
rect 3016 7040 3032 7104
rect 3096 7040 3112 7104
rect 3176 7040 3192 7104
rect 3256 7040 3264 7104
rect 2944 6016 3264 7040
rect 2944 5952 2952 6016
rect 3016 5952 3032 6016
rect 3096 5952 3112 6016
rect 3176 5952 3192 6016
rect 3256 5952 3264 6016
rect 2944 4928 3264 5952
rect 2944 4864 2952 4928
rect 3016 4864 3032 4928
rect 3096 4864 3112 4928
rect 3176 4864 3192 4928
rect 3256 4864 3264 4928
rect 2944 3840 3264 4864
rect 2944 3776 2952 3840
rect 3016 3776 3032 3840
rect 3096 3776 3112 3840
rect 3176 3776 3192 3840
rect 3256 3776 3264 3840
rect 2944 2752 3264 3776
rect 2944 2688 2952 2752
rect 3016 2688 3032 2752
rect 3096 2688 3112 2752
rect 3176 2688 3192 2752
rect 3256 2688 3264 2752
rect 2944 2128 3264 2688
rect 7944 54432 8264 54448
rect 7944 54368 7952 54432
rect 8016 54368 8032 54432
rect 8096 54368 8112 54432
rect 8176 54368 8192 54432
rect 8256 54368 8264 54432
rect 7944 53344 8264 54368
rect 7944 53280 7952 53344
rect 8016 53280 8032 53344
rect 8096 53280 8112 53344
rect 8176 53280 8192 53344
rect 8256 53280 8264 53344
rect 7944 52256 8264 53280
rect 7944 52192 7952 52256
rect 8016 52192 8032 52256
rect 8096 52192 8112 52256
rect 8176 52192 8192 52256
rect 8256 52192 8264 52256
rect 7944 51168 8264 52192
rect 7944 51104 7952 51168
rect 8016 51104 8032 51168
rect 8096 51104 8112 51168
rect 8176 51104 8192 51168
rect 8256 51104 8264 51168
rect 7944 50080 8264 51104
rect 7944 50016 7952 50080
rect 8016 50016 8032 50080
rect 8096 50016 8112 50080
rect 8176 50016 8192 50080
rect 8256 50016 8264 50080
rect 7944 48992 8264 50016
rect 7944 48928 7952 48992
rect 8016 48928 8032 48992
rect 8096 48928 8112 48992
rect 8176 48928 8192 48992
rect 8256 48928 8264 48992
rect 7944 47904 8264 48928
rect 7944 47840 7952 47904
rect 8016 47840 8032 47904
rect 8096 47840 8112 47904
rect 8176 47840 8192 47904
rect 8256 47840 8264 47904
rect 7944 46816 8264 47840
rect 7944 46752 7952 46816
rect 8016 46752 8032 46816
rect 8096 46752 8112 46816
rect 8176 46752 8192 46816
rect 8256 46752 8264 46816
rect 7944 45728 8264 46752
rect 7944 45664 7952 45728
rect 8016 45664 8032 45728
rect 8096 45664 8112 45728
rect 8176 45664 8192 45728
rect 8256 45664 8264 45728
rect 7944 44640 8264 45664
rect 12944 53888 13264 54448
rect 17944 54432 18264 54448
rect 17944 54368 17952 54432
rect 18016 54368 18032 54432
rect 18096 54368 18112 54432
rect 18176 54368 18192 54432
rect 18256 54368 18264 54432
rect 15883 53956 15949 53957
rect 15883 53892 15884 53956
rect 15948 53892 15949 53956
rect 15883 53891 15949 53892
rect 12944 53824 12952 53888
rect 13016 53824 13032 53888
rect 13096 53824 13112 53888
rect 13176 53824 13192 53888
rect 13256 53824 13264 53888
rect 12944 52800 13264 53824
rect 12944 52736 12952 52800
rect 13016 52736 13032 52800
rect 13096 52736 13112 52800
rect 13176 52736 13192 52800
rect 13256 52736 13264 52800
rect 12944 51712 13264 52736
rect 13859 52596 13925 52597
rect 13859 52532 13860 52596
rect 13924 52532 13925 52596
rect 13859 52531 13925 52532
rect 14043 52596 14109 52597
rect 14043 52532 14044 52596
rect 14108 52532 14109 52596
rect 14043 52531 14109 52532
rect 15331 52596 15397 52597
rect 15331 52532 15332 52596
rect 15396 52532 15397 52596
rect 15331 52531 15397 52532
rect 12944 51648 12952 51712
rect 13016 51648 13032 51712
rect 13096 51648 13112 51712
rect 13176 51648 13192 51712
rect 13256 51648 13264 51712
rect 12944 50624 13264 51648
rect 12944 50560 12952 50624
rect 13016 50560 13032 50624
rect 13096 50560 13112 50624
rect 13176 50560 13192 50624
rect 13256 50560 13264 50624
rect 12944 49536 13264 50560
rect 12944 49472 12952 49536
rect 13016 49472 13032 49536
rect 13096 49472 13112 49536
rect 13176 49472 13192 49536
rect 13256 49472 13264 49536
rect 12944 48448 13264 49472
rect 12944 48384 12952 48448
rect 13016 48384 13032 48448
rect 13096 48384 13112 48448
rect 13176 48384 13192 48448
rect 13256 48384 13264 48448
rect 12944 47360 13264 48384
rect 12944 47296 12952 47360
rect 13016 47296 13032 47360
rect 13096 47296 13112 47360
rect 13176 47296 13192 47360
rect 13256 47296 13264 47360
rect 12944 46272 13264 47296
rect 12944 46208 12952 46272
rect 13016 46208 13032 46272
rect 13096 46208 13112 46272
rect 13176 46208 13192 46272
rect 13256 46208 13264 46272
rect 11283 45388 11349 45389
rect 11283 45324 11284 45388
rect 11348 45324 11349 45388
rect 11283 45323 11349 45324
rect 9811 44708 9877 44709
rect 9811 44644 9812 44708
rect 9876 44644 9877 44708
rect 9811 44643 9877 44644
rect 7944 44576 7952 44640
rect 8016 44576 8032 44640
rect 8096 44576 8112 44640
rect 8176 44576 8192 44640
rect 8256 44576 8264 44640
rect 7944 43552 8264 44576
rect 7944 43488 7952 43552
rect 8016 43488 8032 43552
rect 8096 43488 8112 43552
rect 8176 43488 8192 43552
rect 8256 43488 8264 43552
rect 7944 42464 8264 43488
rect 7944 42400 7952 42464
rect 8016 42400 8032 42464
rect 8096 42400 8112 42464
rect 8176 42400 8192 42464
rect 8256 42400 8264 42464
rect 7944 41376 8264 42400
rect 7944 41312 7952 41376
rect 8016 41312 8032 41376
rect 8096 41312 8112 41376
rect 8176 41312 8192 41376
rect 8256 41312 8264 41376
rect 7944 40288 8264 41312
rect 7944 40224 7952 40288
rect 8016 40224 8032 40288
rect 8096 40224 8112 40288
rect 8176 40224 8192 40288
rect 8256 40224 8264 40288
rect 7944 39200 8264 40224
rect 7944 39136 7952 39200
rect 8016 39136 8032 39200
rect 8096 39136 8112 39200
rect 8176 39136 8192 39200
rect 8256 39136 8264 39200
rect 7944 38112 8264 39136
rect 7944 38048 7952 38112
rect 8016 38048 8032 38112
rect 8096 38048 8112 38112
rect 8176 38048 8192 38112
rect 8256 38048 8264 38112
rect 7944 37024 8264 38048
rect 7944 36960 7952 37024
rect 8016 36960 8032 37024
rect 8096 36960 8112 37024
rect 8176 36960 8192 37024
rect 8256 36960 8264 37024
rect 7944 35936 8264 36960
rect 9814 36821 9874 44643
rect 10363 44300 10429 44301
rect 10363 44236 10364 44300
rect 10428 44236 10429 44300
rect 10363 44235 10429 44236
rect 9811 36820 9877 36821
rect 9811 36756 9812 36820
rect 9876 36756 9877 36820
rect 9811 36755 9877 36756
rect 7944 35872 7952 35936
rect 8016 35872 8032 35936
rect 8096 35872 8112 35936
rect 8176 35872 8192 35936
rect 8256 35872 8264 35936
rect 7944 34848 8264 35872
rect 7944 34784 7952 34848
rect 8016 34784 8032 34848
rect 8096 34784 8112 34848
rect 8176 34784 8192 34848
rect 8256 34784 8264 34848
rect 7944 33760 8264 34784
rect 7944 33696 7952 33760
rect 8016 33696 8032 33760
rect 8096 33696 8112 33760
rect 8176 33696 8192 33760
rect 8256 33696 8264 33760
rect 7944 32672 8264 33696
rect 7944 32608 7952 32672
rect 8016 32608 8032 32672
rect 8096 32608 8112 32672
rect 8176 32608 8192 32672
rect 8256 32608 8264 32672
rect 7944 31584 8264 32608
rect 7944 31520 7952 31584
rect 8016 31520 8032 31584
rect 8096 31520 8112 31584
rect 8176 31520 8192 31584
rect 8256 31520 8264 31584
rect 7944 30496 8264 31520
rect 10366 30837 10426 44235
rect 11286 36413 11346 45323
rect 12944 45184 13264 46208
rect 12944 45120 12952 45184
rect 13016 45120 13032 45184
rect 13096 45120 13112 45184
rect 13176 45120 13192 45184
rect 13256 45120 13264 45184
rect 11467 44708 11533 44709
rect 11467 44644 11468 44708
rect 11532 44644 11533 44708
rect 11467 44643 11533 44644
rect 11283 36412 11349 36413
rect 11283 36348 11284 36412
rect 11348 36348 11349 36412
rect 11283 36347 11349 36348
rect 11470 33013 11530 44643
rect 11651 44300 11717 44301
rect 11651 44236 11652 44300
rect 11716 44236 11717 44300
rect 11651 44235 11717 44236
rect 11467 33012 11533 33013
rect 11467 32948 11468 33012
rect 11532 32948 11533 33012
rect 11467 32947 11533 32948
rect 11654 32605 11714 44235
rect 12944 44096 13264 45120
rect 12944 44032 12952 44096
rect 13016 44032 13032 44096
rect 13096 44032 13112 44096
rect 13176 44032 13192 44096
rect 13256 44032 13264 44096
rect 12944 43008 13264 44032
rect 12944 42944 12952 43008
rect 13016 42944 13032 43008
rect 13096 42944 13112 43008
rect 13176 42944 13192 43008
rect 13256 42944 13264 43008
rect 12944 41920 13264 42944
rect 12944 41856 12952 41920
rect 13016 41856 13032 41920
rect 13096 41856 13112 41920
rect 13176 41856 13192 41920
rect 13256 41856 13264 41920
rect 12944 40832 13264 41856
rect 12944 40768 12952 40832
rect 13016 40768 13032 40832
rect 13096 40768 13112 40832
rect 13176 40768 13192 40832
rect 13256 40768 13264 40832
rect 12944 39744 13264 40768
rect 12944 39680 12952 39744
rect 13016 39680 13032 39744
rect 13096 39680 13112 39744
rect 13176 39680 13192 39744
rect 13256 39680 13264 39744
rect 12944 38656 13264 39680
rect 12944 38592 12952 38656
rect 13016 38592 13032 38656
rect 13096 38592 13112 38656
rect 13176 38592 13192 38656
rect 13256 38592 13264 38656
rect 12571 38316 12637 38317
rect 12571 38252 12572 38316
rect 12636 38252 12637 38316
rect 12571 38251 12637 38252
rect 12574 33285 12634 38251
rect 12944 37568 13264 38592
rect 12944 37504 12952 37568
rect 13016 37504 13032 37568
rect 13096 37504 13112 37568
rect 13176 37504 13192 37568
rect 13256 37504 13264 37568
rect 12944 36480 13264 37504
rect 12944 36416 12952 36480
rect 13016 36416 13032 36480
rect 13096 36416 13112 36480
rect 13176 36416 13192 36480
rect 13256 36416 13264 36480
rect 12944 35392 13264 36416
rect 12944 35328 12952 35392
rect 13016 35328 13032 35392
rect 13096 35328 13112 35392
rect 13176 35328 13192 35392
rect 13256 35328 13264 35392
rect 12944 34304 13264 35328
rect 12944 34240 12952 34304
rect 13016 34240 13032 34304
rect 13096 34240 13112 34304
rect 13176 34240 13192 34304
rect 13256 34240 13264 34304
rect 12571 33284 12637 33285
rect 12571 33220 12572 33284
rect 12636 33220 12637 33284
rect 12571 33219 12637 33220
rect 11651 32604 11717 32605
rect 11651 32540 11652 32604
rect 11716 32540 11717 32604
rect 11651 32539 11717 32540
rect 10363 30836 10429 30837
rect 10363 30772 10364 30836
rect 10428 30772 10429 30836
rect 10363 30771 10429 30772
rect 7944 30432 7952 30496
rect 8016 30432 8032 30496
rect 8096 30432 8112 30496
rect 8176 30432 8192 30496
rect 8256 30432 8264 30496
rect 7944 29408 8264 30432
rect 7944 29344 7952 29408
rect 8016 29344 8032 29408
rect 8096 29344 8112 29408
rect 8176 29344 8192 29408
rect 8256 29344 8264 29408
rect 7944 28320 8264 29344
rect 10366 29010 10426 30771
rect 7944 28256 7952 28320
rect 8016 28256 8032 28320
rect 8096 28256 8112 28320
rect 8176 28256 8192 28320
rect 8256 28256 8264 28320
rect 7944 27232 8264 28256
rect 7944 27168 7952 27232
rect 8016 27168 8032 27232
rect 8096 27168 8112 27232
rect 8176 27168 8192 27232
rect 8256 27168 8264 27232
rect 7944 26144 8264 27168
rect 7944 26080 7952 26144
rect 8016 26080 8032 26144
rect 8096 26080 8112 26144
rect 8176 26080 8192 26144
rect 8256 26080 8264 26144
rect 7944 25056 8264 26080
rect 7944 24992 7952 25056
rect 8016 24992 8032 25056
rect 8096 24992 8112 25056
rect 8176 24992 8192 25056
rect 8256 24992 8264 25056
rect 7944 23968 8264 24992
rect 10182 28950 10426 29010
rect 9627 24852 9693 24853
rect 9627 24788 9628 24852
rect 9692 24788 9693 24852
rect 9627 24787 9693 24788
rect 7944 23904 7952 23968
rect 8016 23904 8032 23968
rect 8096 23904 8112 23968
rect 8176 23904 8192 23968
rect 8256 23904 8264 23968
rect 7944 22880 8264 23904
rect 7944 22816 7952 22880
rect 8016 22816 8032 22880
rect 8096 22816 8112 22880
rect 8176 22816 8192 22880
rect 8256 22816 8264 22880
rect 7944 21792 8264 22816
rect 7944 21728 7952 21792
rect 8016 21728 8032 21792
rect 8096 21728 8112 21792
rect 8176 21728 8192 21792
rect 8256 21728 8264 21792
rect 7944 20704 8264 21728
rect 7944 20640 7952 20704
rect 8016 20640 8032 20704
rect 8096 20640 8112 20704
rect 8176 20640 8192 20704
rect 8256 20640 8264 20704
rect 7944 19616 8264 20640
rect 7944 19552 7952 19616
rect 8016 19552 8032 19616
rect 8096 19552 8112 19616
rect 8176 19552 8192 19616
rect 8256 19552 8264 19616
rect 7944 18528 8264 19552
rect 9630 19277 9690 24787
rect 9627 19276 9693 19277
rect 9627 19212 9628 19276
rect 9692 19212 9693 19276
rect 9627 19211 9693 19212
rect 7944 18464 7952 18528
rect 8016 18464 8032 18528
rect 8096 18464 8112 18528
rect 8176 18464 8192 18528
rect 8256 18464 8264 18528
rect 7944 17440 8264 18464
rect 7944 17376 7952 17440
rect 8016 17376 8032 17440
rect 8096 17376 8112 17440
rect 8176 17376 8192 17440
rect 8256 17376 8264 17440
rect 7944 16352 8264 17376
rect 7944 16288 7952 16352
rect 8016 16288 8032 16352
rect 8096 16288 8112 16352
rect 8176 16288 8192 16352
rect 8256 16288 8264 16352
rect 7944 15264 8264 16288
rect 7944 15200 7952 15264
rect 8016 15200 8032 15264
rect 8096 15200 8112 15264
rect 8176 15200 8192 15264
rect 8256 15200 8264 15264
rect 7944 14176 8264 15200
rect 7944 14112 7952 14176
rect 8016 14112 8032 14176
rect 8096 14112 8112 14176
rect 8176 14112 8192 14176
rect 8256 14112 8264 14176
rect 7944 13088 8264 14112
rect 7944 13024 7952 13088
rect 8016 13024 8032 13088
rect 8096 13024 8112 13088
rect 8176 13024 8192 13088
rect 8256 13024 8264 13088
rect 7944 12000 8264 13024
rect 7944 11936 7952 12000
rect 8016 11936 8032 12000
rect 8096 11936 8112 12000
rect 8176 11936 8192 12000
rect 8256 11936 8264 12000
rect 7944 10912 8264 11936
rect 7944 10848 7952 10912
rect 8016 10848 8032 10912
rect 8096 10848 8112 10912
rect 8176 10848 8192 10912
rect 8256 10848 8264 10912
rect 7944 9824 8264 10848
rect 7944 9760 7952 9824
rect 8016 9760 8032 9824
rect 8096 9760 8112 9824
rect 8176 9760 8192 9824
rect 8256 9760 8264 9824
rect 7944 8736 8264 9760
rect 7944 8672 7952 8736
rect 8016 8672 8032 8736
rect 8096 8672 8112 8736
rect 8176 8672 8192 8736
rect 8256 8672 8264 8736
rect 7944 7648 8264 8672
rect 7944 7584 7952 7648
rect 8016 7584 8032 7648
rect 8096 7584 8112 7648
rect 8176 7584 8192 7648
rect 8256 7584 8264 7648
rect 7944 6560 8264 7584
rect 7944 6496 7952 6560
rect 8016 6496 8032 6560
rect 8096 6496 8112 6560
rect 8176 6496 8192 6560
rect 8256 6496 8264 6560
rect 7944 5472 8264 6496
rect 7944 5408 7952 5472
rect 8016 5408 8032 5472
rect 8096 5408 8112 5472
rect 8176 5408 8192 5472
rect 8256 5408 8264 5472
rect 7944 4384 8264 5408
rect 7944 4320 7952 4384
rect 8016 4320 8032 4384
rect 8096 4320 8112 4384
rect 8176 4320 8192 4384
rect 8256 4320 8264 4384
rect 7944 3296 8264 4320
rect 10182 4181 10242 28950
rect 12019 18324 12085 18325
rect 12019 18260 12020 18324
rect 12084 18260 12085 18324
rect 12019 18259 12085 18260
rect 10179 4180 10245 4181
rect 10179 4116 10180 4180
rect 10244 4116 10245 4180
rect 10179 4115 10245 4116
rect 7944 3232 7952 3296
rect 8016 3232 8032 3296
rect 8096 3232 8112 3296
rect 8176 3232 8192 3296
rect 8256 3232 8264 3296
rect 7944 2208 8264 3232
rect 12022 3229 12082 18259
rect 12574 16829 12634 33219
rect 12944 33216 13264 34240
rect 12944 33152 12952 33216
rect 13016 33152 13032 33216
rect 13096 33152 13112 33216
rect 13176 33152 13192 33216
rect 13256 33152 13264 33216
rect 12944 32128 13264 33152
rect 13862 32877 13922 52531
rect 13859 32876 13925 32877
rect 13859 32812 13860 32876
rect 13924 32812 13925 32876
rect 13859 32811 13925 32812
rect 12944 32064 12952 32128
rect 13016 32064 13032 32128
rect 13096 32064 13112 32128
rect 13176 32064 13192 32128
rect 13256 32064 13264 32128
rect 12944 31040 13264 32064
rect 12944 30976 12952 31040
rect 13016 30976 13032 31040
rect 13096 30976 13112 31040
rect 13176 30976 13192 31040
rect 13256 30976 13264 31040
rect 12944 29952 13264 30976
rect 12944 29888 12952 29952
rect 13016 29888 13032 29952
rect 13096 29888 13112 29952
rect 13176 29888 13192 29952
rect 13256 29888 13264 29952
rect 12944 28864 13264 29888
rect 12944 28800 12952 28864
rect 13016 28800 13032 28864
rect 13096 28800 13112 28864
rect 13176 28800 13192 28864
rect 13256 28800 13264 28864
rect 12944 27776 13264 28800
rect 12944 27712 12952 27776
rect 13016 27712 13032 27776
rect 13096 27712 13112 27776
rect 13176 27712 13192 27776
rect 13256 27712 13264 27776
rect 12944 26688 13264 27712
rect 14046 26757 14106 52531
rect 14779 36004 14845 36005
rect 14779 35940 14780 36004
rect 14844 35940 14845 36004
rect 14779 35939 14845 35940
rect 14043 26756 14109 26757
rect 14043 26692 14044 26756
rect 14108 26692 14109 26756
rect 14043 26691 14109 26692
rect 12944 26624 12952 26688
rect 13016 26624 13032 26688
rect 13096 26624 13112 26688
rect 13176 26624 13192 26688
rect 13256 26624 13264 26688
rect 12944 25600 13264 26624
rect 12944 25536 12952 25600
rect 13016 25536 13032 25600
rect 13096 25536 13112 25600
rect 13176 25536 13192 25600
rect 13256 25536 13264 25600
rect 12944 24512 13264 25536
rect 12944 24448 12952 24512
rect 13016 24448 13032 24512
rect 13096 24448 13112 24512
rect 13176 24448 13192 24512
rect 13256 24448 13264 24512
rect 12944 23424 13264 24448
rect 12944 23360 12952 23424
rect 13016 23360 13032 23424
rect 13096 23360 13112 23424
rect 13176 23360 13192 23424
rect 13256 23360 13264 23424
rect 12944 22336 13264 23360
rect 12944 22272 12952 22336
rect 13016 22272 13032 22336
rect 13096 22272 13112 22336
rect 13176 22272 13192 22336
rect 13256 22272 13264 22336
rect 12944 21248 13264 22272
rect 12944 21184 12952 21248
rect 13016 21184 13032 21248
rect 13096 21184 13112 21248
rect 13176 21184 13192 21248
rect 13256 21184 13264 21248
rect 12944 20160 13264 21184
rect 12944 20096 12952 20160
rect 13016 20096 13032 20160
rect 13096 20096 13112 20160
rect 13176 20096 13192 20160
rect 13256 20096 13264 20160
rect 12944 19072 13264 20096
rect 13675 19276 13741 19277
rect 13675 19212 13676 19276
rect 13740 19212 13741 19276
rect 13675 19211 13741 19212
rect 12944 19008 12952 19072
rect 13016 19008 13032 19072
rect 13096 19008 13112 19072
rect 13176 19008 13192 19072
rect 13256 19008 13264 19072
rect 12944 17984 13264 19008
rect 12944 17920 12952 17984
rect 13016 17920 13032 17984
rect 13096 17920 13112 17984
rect 13176 17920 13192 17984
rect 13256 17920 13264 17984
rect 12944 16896 13264 17920
rect 12944 16832 12952 16896
rect 13016 16832 13032 16896
rect 13096 16832 13112 16896
rect 13176 16832 13192 16896
rect 13256 16832 13264 16896
rect 12571 16828 12637 16829
rect 12571 16764 12572 16828
rect 12636 16764 12637 16828
rect 12571 16763 12637 16764
rect 12944 15808 13264 16832
rect 12944 15744 12952 15808
rect 13016 15744 13032 15808
rect 13096 15744 13112 15808
rect 13176 15744 13192 15808
rect 13256 15744 13264 15808
rect 12944 14720 13264 15744
rect 12944 14656 12952 14720
rect 13016 14656 13032 14720
rect 13096 14656 13112 14720
rect 13176 14656 13192 14720
rect 13256 14656 13264 14720
rect 12944 13632 13264 14656
rect 12944 13568 12952 13632
rect 13016 13568 13032 13632
rect 13096 13568 13112 13632
rect 13176 13568 13192 13632
rect 13256 13568 13264 13632
rect 12944 12544 13264 13568
rect 13678 13157 13738 19211
rect 14782 18597 14842 35939
rect 15334 30565 15394 52531
rect 15331 30564 15397 30565
rect 15331 30500 15332 30564
rect 15396 30500 15397 30564
rect 15331 30499 15397 30500
rect 15334 29069 15394 30499
rect 15886 29341 15946 53891
rect 17944 53344 18264 54368
rect 22323 53956 22389 53957
rect 22323 53892 22324 53956
rect 22388 53892 22389 53956
rect 22323 53891 22389 53892
rect 17944 53280 17952 53344
rect 18016 53280 18032 53344
rect 18096 53280 18112 53344
rect 18176 53280 18192 53344
rect 18256 53280 18264 53344
rect 17723 52596 17789 52597
rect 17723 52532 17724 52596
rect 17788 52532 17789 52596
rect 17723 52531 17789 52532
rect 17355 43212 17421 43213
rect 17355 43148 17356 43212
rect 17420 43148 17421 43212
rect 17355 43147 17421 43148
rect 16067 38724 16133 38725
rect 16067 38660 16068 38724
rect 16132 38660 16133 38724
rect 16067 38659 16133 38660
rect 15883 29340 15949 29341
rect 15883 29276 15884 29340
rect 15948 29276 15949 29340
rect 15883 29275 15949 29276
rect 15331 29068 15397 29069
rect 15331 29004 15332 29068
rect 15396 29004 15397 29068
rect 15331 29003 15397 29004
rect 15699 28252 15765 28253
rect 15699 28188 15700 28252
rect 15764 28188 15765 28252
rect 15699 28187 15765 28188
rect 14963 26756 15029 26757
rect 14963 26692 14964 26756
rect 15028 26692 15029 26756
rect 14963 26691 15029 26692
rect 14779 18596 14845 18597
rect 14779 18532 14780 18596
rect 14844 18532 14845 18596
rect 14779 18531 14845 18532
rect 13675 13156 13741 13157
rect 13675 13092 13676 13156
rect 13740 13092 13741 13156
rect 13675 13091 13741 13092
rect 12944 12480 12952 12544
rect 13016 12480 13032 12544
rect 13096 12480 13112 12544
rect 13176 12480 13192 12544
rect 13256 12480 13264 12544
rect 12944 11456 13264 12480
rect 12944 11392 12952 11456
rect 13016 11392 13032 11456
rect 13096 11392 13112 11456
rect 13176 11392 13192 11456
rect 13256 11392 13264 11456
rect 12944 10368 13264 11392
rect 12944 10304 12952 10368
rect 13016 10304 13032 10368
rect 13096 10304 13112 10368
rect 13176 10304 13192 10368
rect 13256 10304 13264 10368
rect 12944 9280 13264 10304
rect 12944 9216 12952 9280
rect 13016 9216 13032 9280
rect 13096 9216 13112 9280
rect 13176 9216 13192 9280
rect 13256 9216 13264 9280
rect 12944 8192 13264 9216
rect 12944 8128 12952 8192
rect 13016 8128 13032 8192
rect 13096 8128 13112 8192
rect 13176 8128 13192 8192
rect 13256 8128 13264 8192
rect 12944 7104 13264 8128
rect 14782 7989 14842 18531
rect 14966 15741 15026 26691
rect 15702 18869 15762 28187
rect 16070 21181 16130 38659
rect 17358 31770 17418 43147
rect 17726 40629 17786 52531
rect 17944 52256 18264 53280
rect 21035 53004 21101 53005
rect 21035 52940 21036 53004
rect 21100 52940 21101 53004
rect 21035 52939 21101 52940
rect 17944 52192 17952 52256
rect 18016 52192 18032 52256
rect 18096 52192 18112 52256
rect 18176 52192 18192 52256
rect 18256 52192 18264 52256
rect 17944 51168 18264 52192
rect 17944 51104 17952 51168
rect 18016 51104 18032 51168
rect 18096 51104 18112 51168
rect 18176 51104 18192 51168
rect 18256 51104 18264 51168
rect 17944 50080 18264 51104
rect 17944 50016 17952 50080
rect 18016 50016 18032 50080
rect 18096 50016 18112 50080
rect 18176 50016 18192 50080
rect 18256 50016 18264 50080
rect 17944 48992 18264 50016
rect 17944 48928 17952 48992
rect 18016 48928 18032 48992
rect 18096 48928 18112 48992
rect 18176 48928 18192 48992
rect 18256 48928 18264 48992
rect 17944 47904 18264 48928
rect 17944 47840 17952 47904
rect 18016 47840 18032 47904
rect 18096 47840 18112 47904
rect 18176 47840 18192 47904
rect 18256 47840 18264 47904
rect 17944 46816 18264 47840
rect 19195 47020 19261 47021
rect 19195 46956 19196 47020
rect 19260 46956 19261 47020
rect 19195 46955 19261 46956
rect 17944 46752 17952 46816
rect 18016 46752 18032 46816
rect 18096 46752 18112 46816
rect 18176 46752 18192 46816
rect 18256 46752 18264 46816
rect 17944 45728 18264 46752
rect 17944 45664 17952 45728
rect 18016 45664 18032 45728
rect 18096 45664 18112 45728
rect 18176 45664 18192 45728
rect 18256 45664 18264 45728
rect 17944 44640 18264 45664
rect 18459 44708 18525 44709
rect 18459 44644 18460 44708
rect 18524 44644 18525 44708
rect 18459 44643 18525 44644
rect 17944 44576 17952 44640
rect 18016 44576 18032 44640
rect 18096 44576 18112 44640
rect 18176 44576 18192 44640
rect 18256 44576 18264 44640
rect 17944 43552 18264 44576
rect 17944 43488 17952 43552
rect 18016 43488 18032 43552
rect 18096 43488 18112 43552
rect 18176 43488 18192 43552
rect 18256 43488 18264 43552
rect 17944 42464 18264 43488
rect 17944 42400 17952 42464
rect 18016 42400 18032 42464
rect 18096 42400 18112 42464
rect 18176 42400 18192 42464
rect 18256 42400 18264 42464
rect 17944 41376 18264 42400
rect 17944 41312 17952 41376
rect 18016 41312 18032 41376
rect 18096 41312 18112 41376
rect 18176 41312 18192 41376
rect 18256 41312 18264 41376
rect 17723 40628 17789 40629
rect 17723 40564 17724 40628
rect 17788 40564 17789 40628
rect 17723 40563 17789 40564
rect 17358 31710 17602 31770
rect 16803 29476 16869 29477
rect 16803 29412 16804 29476
rect 16868 29412 16869 29476
rect 16803 29411 16869 29412
rect 16251 29068 16317 29069
rect 16251 29004 16252 29068
rect 16316 29004 16317 29068
rect 16251 29003 16317 29004
rect 16067 21180 16133 21181
rect 16067 21116 16068 21180
rect 16132 21116 16133 21180
rect 16067 21115 16133 21116
rect 15699 18868 15765 18869
rect 15699 18804 15700 18868
rect 15764 18804 15765 18868
rect 15699 18803 15765 18804
rect 16254 16285 16314 29003
rect 16251 16284 16317 16285
rect 16251 16220 16252 16284
rect 16316 16220 16317 16284
rect 16251 16219 16317 16220
rect 14963 15740 15029 15741
rect 14963 15676 14964 15740
rect 15028 15676 15029 15740
rect 14963 15675 15029 15676
rect 15883 15196 15949 15197
rect 15883 15132 15884 15196
rect 15948 15132 15949 15196
rect 15883 15131 15949 15132
rect 15886 11253 15946 15131
rect 15883 11252 15949 11253
rect 15883 11188 15884 11252
rect 15948 11188 15949 11252
rect 15883 11187 15949 11188
rect 14779 7988 14845 7989
rect 14779 7924 14780 7988
rect 14844 7924 14845 7988
rect 14779 7923 14845 7924
rect 12944 7040 12952 7104
rect 13016 7040 13032 7104
rect 13096 7040 13112 7104
rect 13176 7040 13192 7104
rect 13256 7040 13264 7104
rect 12944 6016 13264 7040
rect 12944 5952 12952 6016
rect 13016 5952 13032 6016
rect 13096 5952 13112 6016
rect 13176 5952 13192 6016
rect 13256 5952 13264 6016
rect 12944 4928 13264 5952
rect 12944 4864 12952 4928
rect 13016 4864 13032 4928
rect 13096 4864 13112 4928
rect 13176 4864 13192 4928
rect 13256 4864 13264 4928
rect 12944 3840 13264 4864
rect 12944 3776 12952 3840
rect 13016 3776 13032 3840
rect 13096 3776 13112 3840
rect 13176 3776 13192 3840
rect 13256 3776 13264 3840
rect 12019 3228 12085 3229
rect 12019 3164 12020 3228
rect 12084 3164 12085 3228
rect 12019 3163 12085 3164
rect 7944 2144 7952 2208
rect 8016 2144 8032 2208
rect 8096 2144 8112 2208
rect 8176 2144 8192 2208
rect 8256 2144 8264 2208
rect 7944 2128 8264 2144
rect 12944 2752 13264 3776
rect 16806 3501 16866 29411
rect 17542 28389 17602 31710
rect 17355 28388 17421 28389
rect 17355 28324 17356 28388
rect 17420 28324 17421 28388
rect 17355 28323 17421 28324
rect 17539 28388 17605 28389
rect 17539 28324 17540 28388
rect 17604 28324 17605 28388
rect 17539 28323 17605 28324
rect 17358 14109 17418 28323
rect 17542 18733 17602 28323
rect 17726 28253 17786 40563
rect 17944 40288 18264 41312
rect 17944 40224 17952 40288
rect 18016 40224 18032 40288
rect 18096 40224 18112 40288
rect 18176 40224 18192 40288
rect 18256 40224 18264 40288
rect 17944 39200 18264 40224
rect 17944 39136 17952 39200
rect 18016 39136 18032 39200
rect 18096 39136 18112 39200
rect 18176 39136 18192 39200
rect 18256 39136 18264 39200
rect 17944 38112 18264 39136
rect 17944 38048 17952 38112
rect 18016 38048 18032 38112
rect 18096 38048 18112 38112
rect 18176 38048 18192 38112
rect 18256 38048 18264 38112
rect 17944 37024 18264 38048
rect 17944 36960 17952 37024
rect 18016 36960 18032 37024
rect 18096 36960 18112 37024
rect 18176 36960 18192 37024
rect 18256 36960 18264 37024
rect 17944 35936 18264 36960
rect 17944 35872 17952 35936
rect 18016 35872 18032 35936
rect 18096 35872 18112 35936
rect 18176 35872 18192 35936
rect 18256 35872 18264 35936
rect 17944 34848 18264 35872
rect 17944 34784 17952 34848
rect 18016 34784 18032 34848
rect 18096 34784 18112 34848
rect 18176 34784 18192 34848
rect 18256 34784 18264 34848
rect 17944 33760 18264 34784
rect 17944 33696 17952 33760
rect 18016 33696 18032 33760
rect 18096 33696 18112 33760
rect 18176 33696 18192 33760
rect 18256 33696 18264 33760
rect 17944 32672 18264 33696
rect 17944 32608 17952 32672
rect 18016 32608 18032 32672
rect 18096 32608 18112 32672
rect 18176 32608 18192 32672
rect 18256 32608 18264 32672
rect 17944 31584 18264 32608
rect 17944 31520 17952 31584
rect 18016 31520 18032 31584
rect 18096 31520 18112 31584
rect 18176 31520 18192 31584
rect 18256 31520 18264 31584
rect 17944 30496 18264 31520
rect 17944 30432 17952 30496
rect 18016 30432 18032 30496
rect 18096 30432 18112 30496
rect 18176 30432 18192 30496
rect 18256 30432 18264 30496
rect 17944 29408 18264 30432
rect 18462 30021 18522 44643
rect 19198 33149 19258 46955
rect 20115 46748 20181 46749
rect 20115 46684 20116 46748
rect 20180 46684 20181 46748
rect 20115 46683 20181 46684
rect 19931 46612 19997 46613
rect 19931 46548 19932 46612
rect 19996 46548 19997 46612
rect 19931 46547 19997 46548
rect 19379 37364 19445 37365
rect 19379 37300 19380 37364
rect 19444 37300 19445 37364
rect 19379 37299 19445 37300
rect 19195 33148 19261 33149
rect 19195 33084 19196 33148
rect 19260 33084 19261 33148
rect 19195 33083 19261 33084
rect 19382 30837 19442 37299
rect 19379 30836 19445 30837
rect 19379 30772 19380 30836
rect 19444 30772 19445 30836
rect 19379 30771 19445 30772
rect 19934 30565 19994 46547
rect 20118 31925 20178 46683
rect 21038 36549 21098 52939
rect 21955 45932 22021 45933
rect 21955 45868 21956 45932
rect 22020 45868 22021 45932
rect 21955 45867 22021 45868
rect 21587 38452 21653 38453
rect 21587 38388 21588 38452
rect 21652 38388 21653 38452
rect 21587 38387 21653 38388
rect 21035 36548 21101 36549
rect 21035 36484 21036 36548
rect 21100 36484 21101 36548
rect 21035 36483 21101 36484
rect 20115 31924 20181 31925
rect 20115 31860 20116 31924
rect 20180 31860 20181 31924
rect 20115 31859 20181 31860
rect 21038 31789 21098 36483
rect 21590 32061 21650 38387
rect 21587 32060 21653 32061
rect 21587 31996 21588 32060
rect 21652 31996 21653 32060
rect 21587 31995 21653 31996
rect 21035 31788 21101 31789
rect 21035 31724 21036 31788
rect 21100 31724 21101 31788
rect 21035 31723 21101 31724
rect 19931 30564 19997 30565
rect 19931 30500 19932 30564
rect 19996 30500 19997 30564
rect 19931 30499 19997 30500
rect 18459 30020 18525 30021
rect 18459 29956 18460 30020
rect 18524 29956 18525 30020
rect 18459 29955 18525 29956
rect 19747 30020 19813 30021
rect 19747 29956 19748 30020
rect 19812 29956 19813 30020
rect 19747 29955 19813 29956
rect 17944 29344 17952 29408
rect 18016 29344 18032 29408
rect 18096 29344 18112 29408
rect 18176 29344 18192 29408
rect 18256 29344 18264 29408
rect 17944 28320 18264 29344
rect 17944 28256 17952 28320
rect 18016 28256 18032 28320
rect 18096 28256 18112 28320
rect 18176 28256 18192 28320
rect 18256 28256 18264 28320
rect 17723 28252 17789 28253
rect 17723 28188 17724 28252
rect 17788 28188 17789 28252
rect 17723 28187 17789 28188
rect 17944 27232 18264 28256
rect 17944 27168 17952 27232
rect 18016 27168 18032 27232
rect 18096 27168 18112 27232
rect 18176 27168 18192 27232
rect 18256 27168 18264 27232
rect 17944 26144 18264 27168
rect 17944 26080 17952 26144
rect 18016 26080 18032 26144
rect 18096 26080 18112 26144
rect 18176 26080 18192 26144
rect 18256 26080 18264 26144
rect 17944 25056 18264 26080
rect 17944 24992 17952 25056
rect 18016 24992 18032 25056
rect 18096 24992 18112 25056
rect 18176 24992 18192 25056
rect 18256 24992 18264 25056
rect 17944 23968 18264 24992
rect 17944 23904 17952 23968
rect 18016 23904 18032 23968
rect 18096 23904 18112 23968
rect 18176 23904 18192 23968
rect 18256 23904 18264 23968
rect 17944 22880 18264 23904
rect 18462 23765 18522 29955
rect 19750 26893 19810 29955
rect 19747 26892 19813 26893
rect 19747 26828 19748 26892
rect 19812 26828 19813 26892
rect 19747 26827 19813 26828
rect 18459 23764 18525 23765
rect 18459 23700 18460 23764
rect 18524 23700 18525 23764
rect 18459 23699 18525 23700
rect 17944 22816 17952 22880
rect 18016 22816 18032 22880
rect 18096 22816 18112 22880
rect 18176 22816 18192 22880
rect 18256 22816 18264 22880
rect 17944 21792 18264 22816
rect 17944 21728 17952 21792
rect 18016 21728 18032 21792
rect 18096 21728 18112 21792
rect 18176 21728 18192 21792
rect 18256 21728 18264 21792
rect 17944 20704 18264 21728
rect 17944 20640 17952 20704
rect 18016 20640 18032 20704
rect 18096 20640 18112 20704
rect 18176 20640 18192 20704
rect 18256 20640 18264 20704
rect 17944 19616 18264 20640
rect 17944 19552 17952 19616
rect 18016 19552 18032 19616
rect 18096 19552 18112 19616
rect 18176 19552 18192 19616
rect 18256 19552 18264 19616
rect 17539 18732 17605 18733
rect 17539 18668 17540 18732
rect 17604 18668 17605 18732
rect 17539 18667 17605 18668
rect 17944 18528 18264 19552
rect 17944 18464 17952 18528
rect 18016 18464 18032 18528
rect 18096 18464 18112 18528
rect 18176 18464 18192 18528
rect 18256 18464 18264 18528
rect 17944 17440 18264 18464
rect 17944 17376 17952 17440
rect 18016 17376 18032 17440
rect 18096 17376 18112 17440
rect 18176 17376 18192 17440
rect 18256 17376 18264 17440
rect 17944 16352 18264 17376
rect 17944 16288 17952 16352
rect 18016 16288 18032 16352
rect 18096 16288 18112 16352
rect 18176 16288 18192 16352
rect 18256 16288 18264 16352
rect 17944 15264 18264 16288
rect 17944 15200 17952 15264
rect 18016 15200 18032 15264
rect 18096 15200 18112 15264
rect 18176 15200 18192 15264
rect 18256 15200 18264 15264
rect 17944 14176 18264 15200
rect 18462 14517 18522 23699
rect 19934 18733 19994 30499
rect 21038 26621 21098 31723
rect 21958 27165 22018 45867
rect 22326 40085 22386 53891
rect 22944 53888 23264 54448
rect 22944 53824 22952 53888
rect 23016 53824 23032 53888
rect 23096 53824 23112 53888
rect 23176 53824 23192 53888
rect 23256 53824 23264 53888
rect 22507 53276 22573 53277
rect 22507 53212 22508 53276
rect 22572 53212 22573 53276
rect 22507 53211 22573 53212
rect 22510 40221 22570 53211
rect 22944 52800 23264 53824
rect 22944 52736 22952 52800
rect 23016 52736 23032 52800
rect 23096 52736 23112 52800
rect 23176 52736 23192 52800
rect 23256 52736 23264 52800
rect 22944 51712 23264 52736
rect 22944 51648 22952 51712
rect 23016 51648 23032 51712
rect 23096 51648 23112 51712
rect 23176 51648 23192 51712
rect 23256 51648 23264 51712
rect 22944 50624 23264 51648
rect 22944 50560 22952 50624
rect 23016 50560 23032 50624
rect 23096 50560 23112 50624
rect 23176 50560 23192 50624
rect 23256 50560 23264 50624
rect 22944 49536 23264 50560
rect 22944 49472 22952 49536
rect 23016 49472 23032 49536
rect 23096 49472 23112 49536
rect 23176 49472 23192 49536
rect 23256 49472 23264 49536
rect 22944 48448 23264 49472
rect 22944 48384 22952 48448
rect 23016 48384 23032 48448
rect 23096 48384 23112 48448
rect 23176 48384 23192 48448
rect 23256 48384 23264 48448
rect 22944 47360 23264 48384
rect 22944 47296 22952 47360
rect 23016 47296 23032 47360
rect 23096 47296 23112 47360
rect 23176 47296 23192 47360
rect 23256 47296 23264 47360
rect 22944 46272 23264 47296
rect 22944 46208 22952 46272
rect 23016 46208 23032 46272
rect 23096 46208 23112 46272
rect 23176 46208 23192 46272
rect 23256 46208 23264 46272
rect 22944 45184 23264 46208
rect 24715 45660 24781 45661
rect 24715 45596 24716 45660
rect 24780 45596 24781 45660
rect 24715 45595 24781 45596
rect 22944 45120 22952 45184
rect 23016 45120 23032 45184
rect 23096 45120 23112 45184
rect 23176 45120 23192 45184
rect 23256 45120 23264 45184
rect 22944 44096 23264 45120
rect 24531 44300 24597 44301
rect 24531 44236 24532 44300
rect 24596 44236 24597 44300
rect 24531 44235 24597 44236
rect 22944 44032 22952 44096
rect 23016 44032 23032 44096
rect 23096 44032 23112 44096
rect 23176 44032 23192 44096
rect 23256 44032 23264 44096
rect 22944 43008 23264 44032
rect 22944 42944 22952 43008
rect 23016 42944 23032 43008
rect 23096 42944 23112 43008
rect 23176 42944 23192 43008
rect 23256 42944 23264 43008
rect 22944 41920 23264 42944
rect 22944 41856 22952 41920
rect 23016 41856 23032 41920
rect 23096 41856 23112 41920
rect 23176 41856 23192 41920
rect 23256 41856 23264 41920
rect 22691 41444 22757 41445
rect 22691 41380 22692 41444
rect 22756 41380 22757 41444
rect 22691 41379 22757 41380
rect 22507 40220 22573 40221
rect 22507 40156 22508 40220
rect 22572 40156 22573 40220
rect 22507 40155 22573 40156
rect 22139 40084 22205 40085
rect 22139 40020 22140 40084
rect 22204 40020 22205 40084
rect 22139 40019 22205 40020
rect 22323 40084 22389 40085
rect 22323 40020 22324 40084
rect 22388 40020 22389 40084
rect 22323 40019 22389 40020
rect 22142 33149 22202 40019
rect 22694 38045 22754 41379
rect 22944 40832 23264 41856
rect 22944 40768 22952 40832
rect 23016 40768 23032 40832
rect 23096 40768 23112 40832
rect 23176 40768 23192 40832
rect 23256 40768 23264 40832
rect 22944 39744 23264 40768
rect 23427 40084 23493 40085
rect 23427 40020 23428 40084
rect 23492 40020 23493 40084
rect 23427 40019 23493 40020
rect 22944 39680 22952 39744
rect 23016 39680 23032 39744
rect 23096 39680 23112 39744
rect 23176 39680 23192 39744
rect 23256 39680 23264 39744
rect 22944 38656 23264 39680
rect 22944 38592 22952 38656
rect 23016 38592 23032 38656
rect 23096 38592 23112 38656
rect 23176 38592 23192 38656
rect 23256 38592 23264 38656
rect 22691 38044 22757 38045
rect 22691 37980 22692 38044
rect 22756 37980 22757 38044
rect 22691 37979 22757 37980
rect 22944 37568 23264 38592
rect 22944 37504 22952 37568
rect 23016 37504 23032 37568
rect 23096 37504 23112 37568
rect 23176 37504 23192 37568
rect 23256 37504 23264 37568
rect 22944 36480 23264 37504
rect 22944 36416 22952 36480
rect 23016 36416 23032 36480
rect 23096 36416 23112 36480
rect 23176 36416 23192 36480
rect 23256 36416 23264 36480
rect 22944 35392 23264 36416
rect 22944 35328 22952 35392
rect 23016 35328 23032 35392
rect 23096 35328 23112 35392
rect 23176 35328 23192 35392
rect 23256 35328 23264 35392
rect 22944 34304 23264 35328
rect 22944 34240 22952 34304
rect 23016 34240 23032 34304
rect 23096 34240 23112 34304
rect 23176 34240 23192 34304
rect 23256 34240 23264 34304
rect 22944 33216 23264 34240
rect 22944 33152 22952 33216
rect 23016 33152 23032 33216
rect 23096 33152 23112 33216
rect 23176 33152 23192 33216
rect 23256 33152 23264 33216
rect 22139 33148 22205 33149
rect 22139 33084 22140 33148
rect 22204 33084 22205 33148
rect 22139 33083 22205 33084
rect 22944 32128 23264 33152
rect 23430 33013 23490 40019
rect 24534 35189 24594 44235
rect 24531 35188 24597 35189
rect 24531 35124 24532 35188
rect 24596 35124 24597 35188
rect 24531 35123 24597 35124
rect 24718 33421 24778 45595
rect 24715 33420 24781 33421
rect 24715 33356 24716 33420
rect 24780 33356 24781 33420
rect 24715 33355 24781 33356
rect 23427 33012 23493 33013
rect 23427 32948 23428 33012
rect 23492 32948 23493 33012
rect 23427 32947 23493 32948
rect 22944 32064 22952 32128
rect 23016 32064 23032 32128
rect 23096 32064 23112 32128
rect 23176 32064 23192 32128
rect 23256 32064 23264 32128
rect 22944 31040 23264 32064
rect 22944 30976 22952 31040
rect 23016 30976 23032 31040
rect 23096 30976 23112 31040
rect 23176 30976 23192 31040
rect 23256 30976 23264 31040
rect 22944 29952 23264 30976
rect 22944 29888 22952 29952
rect 23016 29888 23032 29952
rect 23096 29888 23112 29952
rect 23176 29888 23192 29952
rect 23256 29888 23264 29952
rect 22944 28864 23264 29888
rect 22944 28800 22952 28864
rect 23016 28800 23032 28864
rect 23096 28800 23112 28864
rect 23176 28800 23192 28864
rect 23256 28800 23264 28864
rect 22944 27776 23264 28800
rect 22944 27712 22952 27776
rect 23016 27712 23032 27776
rect 23096 27712 23112 27776
rect 23176 27712 23192 27776
rect 23256 27712 23264 27776
rect 21955 27164 22021 27165
rect 21955 27100 21956 27164
rect 22020 27100 22021 27164
rect 21955 27099 22021 27100
rect 22944 26688 23264 27712
rect 22944 26624 22952 26688
rect 23016 26624 23032 26688
rect 23096 26624 23112 26688
rect 23176 26624 23192 26688
rect 23256 26624 23264 26688
rect 21035 26620 21101 26621
rect 21035 26556 21036 26620
rect 21100 26556 21101 26620
rect 21035 26555 21101 26556
rect 22944 25600 23264 26624
rect 22944 25536 22952 25600
rect 23016 25536 23032 25600
rect 23096 25536 23112 25600
rect 23176 25536 23192 25600
rect 23256 25536 23264 25600
rect 22944 24512 23264 25536
rect 22944 24448 22952 24512
rect 23016 24448 23032 24512
rect 23096 24448 23112 24512
rect 23176 24448 23192 24512
rect 23256 24448 23264 24512
rect 22944 23424 23264 24448
rect 22944 23360 22952 23424
rect 23016 23360 23032 23424
rect 23096 23360 23112 23424
rect 23176 23360 23192 23424
rect 23256 23360 23264 23424
rect 22944 22336 23264 23360
rect 22944 22272 22952 22336
rect 23016 22272 23032 22336
rect 23096 22272 23112 22336
rect 23176 22272 23192 22336
rect 23256 22272 23264 22336
rect 21219 22268 21285 22269
rect 21219 22204 21220 22268
rect 21284 22204 21285 22268
rect 21219 22203 21285 22204
rect 20667 20500 20733 20501
rect 20667 20436 20668 20500
rect 20732 20436 20733 20500
rect 20667 20435 20733 20436
rect 19931 18732 19997 18733
rect 19931 18668 19932 18732
rect 19996 18668 19997 18732
rect 19931 18667 19997 18668
rect 20670 16557 20730 20435
rect 21222 16557 21282 22203
rect 22944 21248 23264 22272
rect 22944 21184 22952 21248
rect 23016 21184 23032 21248
rect 23096 21184 23112 21248
rect 23176 21184 23192 21248
rect 23256 21184 23264 21248
rect 22944 20160 23264 21184
rect 22944 20096 22952 20160
rect 23016 20096 23032 20160
rect 23096 20096 23112 20160
rect 23176 20096 23192 20160
rect 23256 20096 23264 20160
rect 22944 19072 23264 20096
rect 22944 19008 22952 19072
rect 23016 19008 23032 19072
rect 23096 19008 23112 19072
rect 23176 19008 23192 19072
rect 23256 19008 23264 19072
rect 22944 17984 23264 19008
rect 22944 17920 22952 17984
rect 23016 17920 23032 17984
rect 23096 17920 23112 17984
rect 23176 17920 23192 17984
rect 23256 17920 23264 17984
rect 22944 16896 23264 17920
rect 22944 16832 22952 16896
rect 23016 16832 23032 16896
rect 23096 16832 23112 16896
rect 23176 16832 23192 16896
rect 23256 16832 23264 16896
rect 20667 16556 20733 16557
rect 20667 16492 20668 16556
rect 20732 16492 20733 16556
rect 20667 16491 20733 16492
rect 21219 16556 21285 16557
rect 21219 16492 21220 16556
rect 21284 16492 21285 16556
rect 21219 16491 21285 16492
rect 22944 15808 23264 16832
rect 22944 15744 22952 15808
rect 23016 15744 23032 15808
rect 23096 15744 23112 15808
rect 23176 15744 23192 15808
rect 23256 15744 23264 15808
rect 22944 14720 23264 15744
rect 22944 14656 22952 14720
rect 23016 14656 23032 14720
rect 23096 14656 23112 14720
rect 23176 14656 23192 14720
rect 23256 14656 23264 14720
rect 18459 14516 18525 14517
rect 18459 14452 18460 14516
rect 18524 14452 18525 14516
rect 18459 14451 18525 14452
rect 17944 14112 17952 14176
rect 18016 14112 18032 14176
rect 18096 14112 18112 14176
rect 18176 14112 18192 14176
rect 18256 14112 18264 14176
rect 17355 14108 17421 14109
rect 17355 14044 17356 14108
rect 17420 14044 17421 14108
rect 17355 14043 17421 14044
rect 17944 13088 18264 14112
rect 17944 13024 17952 13088
rect 18016 13024 18032 13088
rect 18096 13024 18112 13088
rect 18176 13024 18192 13088
rect 18256 13024 18264 13088
rect 17944 12000 18264 13024
rect 17944 11936 17952 12000
rect 18016 11936 18032 12000
rect 18096 11936 18112 12000
rect 18176 11936 18192 12000
rect 18256 11936 18264 12000
rect 17944 10912 18264 11936
rect 17944 10848 17952 10912
rect 18016 10848 18032 10912
rect 18096 10848 18112 10912
rect 18176 10848 18192 10912
rect 18256 10848 18264 10912
rect 17944 9824 18264 10848
rect 17944 9760 17952 9824
rect 18016 9760 18032 9824
rect 18096 9760 18112 9824
rect 18176 9760 18192 9824
rect 18256 9760 18264 9824
rect 17944 8736 18264 9760
rect 17944 8672 17952 8736
rect 18016 8672 18032 8736
rect 18096 8672 18112 8736
rect 18176 8672 18192 8736
rect 18256 8672 18264 8736
rect 17944 7648 18264 8672
rect 17944 7584 17952 7648
rect 18016 7584 18032 7648
rect 18096 7584 18112 7648
rect 18176 7584 18192 7648
rect 18256 7584 18264 7648
rect 17944 6560 18264 7584
rect 17944 6496 17952 6560
rect 18016 6496 18032 6560
rect 18096 6496 18112 6560
rect 18176 6496 18192 6560
rect 18256 6496 18264 6560
rect 17944 5472 18264 6496
rect 17944 5408 17952 5472
rect 18016 5408 18032 5472
rect 18096 5408 18112 5472
rect 18176 5408 18192 5472
rect 18256 5408 18264 5472
rect 17944 4384 18264 5408
rect 17944 4320 17952 4384
rect 18016 4320 18032 4384
rect 18096 4320 18112 4384
rect 18176 4320 18192 4384
rect 18256 4320 18264 4384
rect 16803 3500 16869 3501
rect 16803 3436 16804 3500
rect 16868 3436 16869 3500
rect 16803 3435 16869 3436
rect 12944 2688 12952 2752
rect 13016 2688 13032 2752
rect 13096 2688 13112 2752
rect 13176 2688 13192 2752
rect 13256 2688 13264 2752
rect 12944 2128 13264 2688
rect 17944 3296 18264 4320
rect 17944 3232 17952 3296
rect 18016 3232 18032 3296
rect 18096 3232 18112 3296
rect 18176 3232 18192 3296
rect 18256 3232 18264 3296
rect 17944 2208 18264 3232
rect 17944 2144 17952 2208
rect 18016 2144 18032 2208
rect 18096 2144 18112 2208
rect 18176 2144 18192 2208
rect 18256 2144 18264 2208
rect 17944 2128 18264 2144
rect 22944 13632 23264 14656
rect 22944 13568 22952 13632
rect 23016 13568 23032 13632
rect 23096 13568 23112 13632
rect 23176 13568 23192 13632
rect 23256 13568 23264 13632
rect 22944 12544 23264 13568
rect 22944 12480 22952 12544
rect 23016 12480 23032 12544
rect 23096 12480 23112 12544
rect 23176 12480 23192 12544
rect 23256 12480 23264 12544
rect 22944 11456 23264 12480
rect 22944 11392 22952 11456
rect 23016 11392 23032 11456
rect 23096 11392 23112 11456
rect 23176 11392 23192 11456
rect 23256 11392 23264 11456
rect 22944 10368 23264 11392
rect 22944 10304 22952 10368
rect 23016 10304 23032 10368
rect 23096 10304 23112 10368
rect 23176 10304 23192 10368
rect 23256 10304 23264 10368
rect 22944 9280 23264 10304
rect 22944 9216 22952 9280
rect 23016 9216 23032 9280
rect 23096 9216 23112 9280
rect 23176 9216 23192 9280
rect 23256 9216 23264 9280
rect 22944 8192 23264 9216
rect 22944 8128 22952 8192
rect 23016 8128 23032 8192
rect 23096 8128 23112 8192
rect 23176 8128 23192 8192
rect 23256 8128 23264 8192
rect 22944 7104 23264 8128
rect 22944 7040 22952 7104
rect 23016 7040 23032 7104
rect 23096 7040 23112 7104
rect 23176 7040 23192 7104
rect 23256 7040 23264 7104
rect 22944 6016 23264 7040
rect 22944 5952 22952 6016
rect 23016 5952 23032 6016
rect 23096 5952 23112 6016
rect 23176 5952 23192 6016
rect 23256 5952 23264 6016
rect 22944 4928 23264 5952
rect 22944 4864 22952 4928
rect 23016 4864 23032 4928
rect 23096 4864 23112 4928
rect 23176 4864 23192 4928
rect 23256 4864 23264 4928
rect 22944 3840 23264 4864
rect 22944 3776 22952 3840
rect 23016 3776 23032 3840
rect 23096 3776 23112 3840
rect 23176 3776 23192 3840
rect 23256 3776 23264 3840
rect 22944 2752 23264 3776
rect 22944 2688 22952 2752
rect 23016 2688 23032 2752
rect 23096 2688 23112 2752
rect 23176 2688 23192 2752
rect 23256 2688 23264 2752
rect 22944 2128 23264 2688
use sky130_fd_sc_hd__clkbuf_2  _109_ pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1679235063
transform 1 0 24564 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _110_
timestamp 1679235063
transform 1 0 24564 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _111_ pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1679235063
transform 1 0 23184 0 1 4352
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_1  _112_ pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1679235063
transform 1 0 24656 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  _113_
timestamp 1679235063
transform 1 0 23736 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  _114_
timestamp 1679235063
transform 1 0 24656 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _115_
timestamp 1679235063
transform 1 0 23184 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  _116_
timestamp 1679235063
transform 1 0 16008 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  _117_
timestamp 1679235063
transform 1 0 23184 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _118_
timestamp 1679235063
transform 1 0 22448 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  _119_
timestamp 1679235063
transform 1 0 21620 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _120_
timestamp 1679235063
transform 1 0 23184 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _121_
timestamp 1679235063
transform 1 0 22448 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _122_
timestamp 1679235063
transform 1 0 20240 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _123_
timestamp 1679235063
transform 1 0 23092 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _124_
timestamp 1679235063
transform 1 0 20976 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _125_
timestamp 1679235063
transform 1 0 20332 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _126_
timestamp 1679235063
transform 1 0 24564 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _127_
timestamp 1679235063
transform 1 0 24564 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _128_
timestamp 1679235063
transform 1 0 25024 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _129_
timestamp 1679235063
transform 1 0 23736 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _130_
timestamp 1679235063
transform 1 0 24564 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _131_
timestamp 1679235063
transform 1 0 24564 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _132_
timestamp 1679235063
transform 1 0 23736 0 1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _133_
timestamp 1679235063
transform 1 0 24564 0 -1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _134_
timestamp 1679235063
transform 1 0 24564 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  _135_
timestamp 1679235063
transform 1 0 24656 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  _136_
timestamp 1679235063
transform 1 0 24564 0 -1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  _137_
timestamp 1679235063
transform 1 0 24564 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  _138_
timestamp 1679235063
transform 1 0 14260 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _139_
timestamp 1679235063
transform 1 0 14444 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _140_
timestamp 1679235063
transform 1 0 13432 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _141_
timestamp 1679235063
transform 1 0 11868 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _142_
timestamp 1679235063
transform 1 0 14260 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _143_
timestamp 1679235063
transform 1 0 14260 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _144_
timestamp 1679235063
transform 1 0 15548 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _145_
timestamp 1679235063
transform 1 0 16744 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _146_
timestamp 1679235063
transform 1 0 15916 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _147_
timestamp 1679235063
transform 1 0 15364 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _148_
timestamp 1679235063
transform 1 0 16836 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _149_
timestamp 1679235063
transform 1 0 14444 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _150_
timestamp 1679235063
transform 1 0 17572 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _151_
timestamp 1679235063
transform 1 0 17664 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _152_
timestamp 1679235063
transform 1 0 17480 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _153_
timestamp 1679235063
transform 1 0 16836 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _154_
timestamp 1679235063
transform 1 0 18308 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _155_
timestamp 1679235063
transform 1 0 18308 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _156_
timestamp 1679235063
transform 1 0 18584 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _157_
timestamp 1679235063
transform 1 0 20700 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _158_
timestamp 1679235063
transform 1 0 19412 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _159_
timestamp 1679235063
transform 1 0 20148 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _160_
timestamp 1679235063
transform 1 0 21988 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _161_
timestamp 1679235063
transform 1 0 18768 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _162_
timestamp 1679235063
transform 1 0 18400 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _163_
timestamp 1679235063
transform 1 0 20884 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _164_
timestamp 1679235063
transform 1 0 18768 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  _165_
timestamp 1679235063
transform 1 0 20424 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _166_
timestamp 1679235063
transform 1 0 20056 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  _167_
timestamp 1679235063
transform 1 0 19320 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _168_
timestamp 1679235063
transform 1 0 3404 0 -1 41344
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _169_
timestamp 1679235063
transform 1 0 4508 0 -1 41344
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _170_
timestamp 1679235063
transform 1 0 3956 0 1 41344
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _171_
timestamp 1679235063
transform 1 0 6716 0 -1 51136
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _172_
timestamp 1679235063
transform 1 0 4692 0 1 42432
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _173_
timestamp 1679235063
transform 1 0 4692 0 1 41344
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _174_
timestamp 1679235063
transform 1 0 5612 0 -1 42432
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _175_
timestamp 1679235063
transform 1 0 6808 0 -1 52224
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _176_
timestamp 1679235063
transform 1 0 6532 0 1 43520
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _177_
timestamp 1679235063
transform 1 0 6532 0 -1 44608
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _178_
timestamp 1679235063
transform 1 0 7268 0 -1 44608
box -38 -48 406 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _179_
timestamp 1679235063
transform 1 0 7452 0 -1 51136
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_2  _180_
timestamp 1679235063
transform 1 0 7636 0 1 44608
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _181_
timestamp 1679235063
transform 1 0 7912 0 1 45696
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _182_
timestamp 1679235063
transform 1 0 8832 0 -1 44608
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  _183_
timestamp 1679235063
transform 1 0 6808 0 1 50048
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  _184_
timestamp 1679235063
transform 1 0 9108 0 1 44608
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _185_
timestamp 1679235063
transform 1 0 8372 0 -1 43520
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _186_
timestamp 1679235063
transform 1 0 10120 0 -1 44608
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  _187_
timestamp 1679235063
transform 1 0 9200 0 1 50048
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  _188_
timestamp 1679235063
transform 1 0 10856 0 -1 44608
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _189_
timestamp 1679235063
transform 1 0 11040 0 1 44608
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _190_
timestamp 1679235063
transform 1 0 11684 0 -1 45696
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _191_
timestamp 1679235063
transform 1 0 9108 0 -1 50048
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _192_
timestamp 1679235063
transform 1 0 9292 0 -1 51136
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _193_
timestamp 1679235063
transform 1 0 12144 0 1 44608
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  _194_
timestamp 1679235063
transform 1 0 10212 0 1 51136
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _195_
timestamp 1679235063
transform 1 0 11684 0 -1 52224
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _196_
timestamp 1679235063
transform 1 0 12604 0 1 52224
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _197_
timestamp 1679235063
transform 1 0 12328 0 -1 52224
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  _198_
timestamp 1679235063
transform 1 0 2116 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _199_
timestamp 1679235063
transform 1 0 2024 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  _200_
timestamp 1679235063
transform 1 0 2024 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _201_
timestamp 1679235063
transform 1 0 2024 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_1 pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1679235063
transform 1 0 12604 0 -1 33728
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__138__A
timestamp 1679235063
transform 1 0 14812 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__139__A
timestamp 1679235063
transform 1 0 14996 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__140__A
timestamp 1679235063
transform 1 0 13800 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__141__A
timestamp 1679235063
transform 1 0 12420 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__142__A
timestamp 1679235063
transform 1 0 14812 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__143__A
timestamp 1679235063
transform 1 0 14812 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__144__A
timestamp 1679235063
transform 1 0 16100 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__146__A
timestamp 1679235063
transform 1 0 17112 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__147__A
timestamp 1679235063
transform 1 0 15916 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__148__A
timestamp 1679235063
transform 1 0 17204 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__150__A
timestamp 1679235063
transform 1 0 18124 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__151__A
timestamp 1679235063
transform 1 0 18860 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__152__A
timestamp 1679235063
transform 1 0 17940 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__154__A
timestamp 1679235063
transform 1 0 18860 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__155__A
timestamp 1679235063
transform 1 0 18860 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__156__A
timestamp 1679235063
transform 1 0 19228 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__158__A
timestamp 1679235063
transform 1 0 19872 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__159__A
timestamp 1679235063
transform 1 0 20700 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__160__A
timestamp 1679235063
transform 1 0 23184 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__163__A
timestamp 1679235063
transform 1 0 21252 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__168__A
timestamp 1679235063
transform 1 0 3956 0 -1 41344
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__169__A
timestamp 1679235063
transform 1 0 5060 0 -1 41344
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__170__A
timestamp 1679235063
transform 1 0 3496 0 1 41344
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__172__A
timestamp 1679235063
transform 1 0 5244 0 1 42432
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__173__A
timestamp 1679235063
transform 1 0 5244 0 1 41344
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__174__A
timestamp 1679235063
transform 1 0 5244 0 -1 42432
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__176__A
timestamp 1679235063
transform 1 0 7084 0 1 43520
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__177__A
timestamp 1679235063
transform 1 0 6348 0 1 44608
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__178__A
timestamp 1679235063
transform 1 0 7820 0 -1 44608
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__180__A
timestamp 1679235063
transform 1 0 7268 0 1 44608
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__181__A
timestamp 1679235063
transform 1 0 8464 0 1 45696
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__182__A
timestamp 1679235063
transform 1 0 9384 0 -1 44608
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__184__A
timestamp 1679235063
transform 1 0 9660 0 1 44608
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__185__A
timestamp 1679235063
transform 1 0 7360 0 -1 43520
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__186__A
timestamp 1679235063
transform 1 0 9752 0 -1 44608
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__188__A
timestamp 1679235063
transform 1 0 11500 0 -1 44608
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__189__A
timestamp 1679235063
transform 1 0 11592 0 1 44608
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__190__A
timestamp 1679235063
transform 1 0 12236 0 -1 45696
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__193__A
timestamp 1679235063
transform 1 0 12696 0 1 44608
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_cby_0__1_.cby_0__1_.mem_right_ipin_0.sky130_fd_sc_hd__dfrtp_1_0__RESET_B
timestamp 1679235063
transform 1 0 6348 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_cby_0__1_.cby_0__1_.mem_right_ipin_0.sky130_fd_sc_hd__dfrtp_1_1__D
timestamp 1679235063
transform 1 0 11408 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_cby_0__1_.cby_0__1_.mem_right_ipin_0.sky130_fd_sc_hd__dfrtp_1_1__RESET_B
timestamp 1679235063
transform 1 0 11224 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_cby_0__1_.cby_0__1_.mem_right_ipin_0.sky130_fd_sc_hd__dfrtp_1_2__RESET_B
timestamp 1679235063
transform 1 0 8280 0 1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_cby_0__1_.cby_0__1_.mem_right_ipin_0.sky130_fd_sc_hd__dfrtp_1_3__RESET_B
timestamp 1679235063
transform 1 0 8556 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_cby_0__1_.cby_0__1_.mem_right_ipin_1.sky130_fd_sc_hd__dfrtp_1_0__RESET_B
timestamp 1679235063
transform 1 0 10120 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_cby_0__1_.cby_0__1_.mem_right_ipin_1.sky130_fd_sc_hd__dfrtp_1_1__RESET_B
timestamp 1679235063
transform 1 0 13892 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_cby_0__1_.cby_0__1_.mem_right_ipin_1.sky130_fd_sc_hd__dfrtp_1_2__RESET_B
timestamp 1679235063
transform 1 0 10120 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_cby_0__1_.cby_0__1_.mem_right_ipin_1.sky130_fd_sc_hd__dfrtp_1_3__RESET_B
timestamp 1679235063
transform 1 0 7728 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_cby_0__1_.cby_0__1_.mem_right_ipin_2.sky130_fd_sc_hd__dfrtp_1_0__RESET_B
timestamp 1679235063
transform 1 0 10396 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_cby_0__1_.cby_0__1_.mem_right_ipin_2.sky130_fd_sc_hd__dfrtp_1_1__RESET_B
timestamp 1679235063
transform 1 0 12144 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_cby_0__1_.cby_0__1_.mem_right_ipin_2.sky130_fd_sc_hd__dfrtp_1_2__RESET_B
timestamp 1679235063
transform 1 0 8004 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_cby_0__1_.cby_0__1_.mem_right_ipin_2.sky130_fd_sc_hd__dfrtp_1_3__RESET_B
timestamp 1679235063
transform 1 0 6624 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_cby_0__1_.cby_0__1_.mem_right_ipin_3.sky130_fd_sc_hd__dfrtp_1_0__RESET_B
timestamp 1679235063
transform 1 0 8648 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_cby_0__1_.cby_0__1_.mem_right_ipin_3.sky130_fd_sc_hd__dfrtp_1_1__RESET_B
timestamp 1679235063
transform 1 0 10396 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_cby_0__1_.cby_0__1_.mem_right_ipin_3.sky130_fd_sc_hd__dfrtp_1_2__RESET_B
timestamp 1679235063
transform 1 0 7360 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_cby_0__1_.cby_0__1_.mem_right_ipin_3.sky130_fd_sc_hd__dfrtp_1_3__RESET_B
timestamp 1679235063
transform 1 0 6164 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_cby_0__1_.cby_0__1_.mux_right_ipin_0.mux_l1_in_0__A1
timestamp 1679235063
transform 1 0 12420 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_cby_0__1_.cby_0__1_.mux_right_ipin_0.mux_l1_in_0__S
timestamp 1679235063
transform 1 0 12604 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_cby_0__1_.cby_0__1_.mux_right_ipin_0.mux_l1_in_1__A1
timestamp 1679235063
transform 1 0 12420 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_cby_0__1_.cby_0__1_.mux_right_ipin_0.mux_l1_in_1__S
timestamp 1679235063
transform 1 0 12696 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_cby_0__1_.cby_0__1_.mux_right_ipin_0.mux_l1_in_2__A1
timestamp 1679235063
transform 1 0 14628 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_cby_0__1_.cby_0__1_.mux_right_ipin_0.mux_l1_in_2__S
timestamp 1679235063
transform 1 0 14444 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_cby_0__1_.cby_0__1_.mux_right_ipin_0.mux_l1_in_3__A0
timestamp 1679235063
transform 1 0 13340 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_cby_0__1_.cby_0__1_.mux_right_ipin_0.mux_l1_in_3__A1
timestamp 1679235063
transform 1 0 11592 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_cby_0__1_.cby_0__1_.mux_right_ipin_0.mux_l1_in_3__S
timestamp 1679235063
transform 1 0 11776 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_cby_0__1_.cby_0__1_.mux_right_ipin_0.mux_l1_in_4__A1
timestamp 1679235063
transform 1 0 10580 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_cby_0__1_.cby_0__1_.mux_right_ipin_0.mux_l1_in_4__S
timestamp 1679235063
transform 1 0 10212 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_cby_0__1_.cby_0__1_.mux_right_ipin_0.mux_l2_in_2__A0
timestamp 1679235063
transform 1 0 8648 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_cby_0__1_.cby_0__1_.mux_right_ipin_0.mux_l2_in_3__A1
timestamp 1679235063
transform 1 0 10304 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_cby_0__1_.cby_0__1_.mux_right_ipin_1.mux_l1_in_1__A0
timestamp 1679235063
transform 1 0 16100 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_cby_0__1_.cby_0__1_.mux_right_ipin_1.mux_l1_in_1__A1
timestamp 1679235063
transform 1 0 14720 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_cby_0__1_.cby_0__1_.mux_right_ipin_1.mux_l1_in_2__A0
timestamp 1679235063
transform 1 0 15548 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_cby_0__1_.cby_0__1_.mux_right_ipin_1.mux_l1_in_2__A1
timestamp 1679235063
transform 1 0 14076 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_cby_0__1_.cby_0__1_.mux_right_ipin_1.mux_l1_in_3__A0
timestamp 1679235063
transform 1 0 14996 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_cby_0__1_.cby_0__1_.mux_right_ipin_1.mux_l1_in_3__A1
timestamp 1679235063
transform 1 0 13800 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_cby_0__1_.cby_0__1_.mux_right_ipin_1.mux_l1_in_4__A0
timestamp 1679235063
transform 1 0 11960 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_cby_0__1_.cby_0__1_.mux_right_ipin_1.mux_l1_in_4__A1
timestamp 1679235063
transform 1 0 10764 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_cby_0__1_.cby_0__1_.mux_right_ipin_1.mux_l2_in_2__A0
timestamp 1679235063
transform 1 0 9200 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_cby_0__1_.cby_0__1_.mux_right_ipin_1.mux_l2_in_3__A1
timestamp 1679235063
transform 1 0 12696 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_cby_0__1_.cby_0__1_.mux_right_ipin_2.mux_l1_in_0__A1
timestamp 1679235063
transform 1 0 16376 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_cby_0__1_.cby_0__1_.mux_right_ipin_2.mux_l1_in_1__A1
timestamp 1679235063
transform 1 0 12972 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_cby_0__1_.cby_0__1_.mux_right_ipin_2.mux_l1_in_2__A0
timestamp 1679235063
transform 1 0 15272 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_cby_0__1_.cby_0__1_.mux_right_ipin_2.mux_l1_in_2__A1
timestamp 1679235063
transform 1 0 13892 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_cby_0__1_.cby_0__1_.mux_right_ipin_2.mux_l1_in_3__A1
timestamp 1679235063
transform 1 0 12880 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_cby_0__1_.cby_0__1_.mux_right_ipin_2.mux_l1_in_4__A0
timestamp 1679235063
transform 1 0 11592 0 1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_cby_0__1_.cby_0__1_.mux_right_ipin_2.mux_l1_in_4__A1
timestamp 1679235063
transform 1 0 10028 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_cby_0__1_.cby_0__1_.mux_right_ipin_2.mux_l2_in_2__A0
timestamp 1679235063
transform 1 0 9200 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_cby_0__1_.cby_0__1_.mux_right_ipin_2.mux_l2_in_3__A1
timestamp 1679235063
transform 1 0 10028 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_cby_0__1_.cby_0__1_.mux_right_ipin_3.mux_l1_in_0__A1
timestamp 1679235063
transform 1 0 12604 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_cby_0__1_.cby_0__1_.mux_right_ipin_3.mux_l1_in_1__A1
timestamp 1679235063
transform 1 0 12236 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_cby_0__1_.cby_0__1_.mux_right_ipin_3.mux_l1_in_2__A0
timestamp 1679235063
transform 1 0 14260 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_cby_0__1_.cby_0__1_.mux_right_ipin_3.mux_l1_in_2__A1
timestamp 1679235063
transform 1 0 12880 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_cby_0__1_.cby_0__1_.mux_right_ipin_3.mux_l1_in_3__A0
timestamp 1679235063
transform 1 0 12972 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_cby_0__1_.cby_0__1_.mux_right_ipin_3.mux_l1_in_3__A1
timestamp 1679235063
transform 1 0 11224 0 -1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_cby_0__1_.cby_0__1_.mux_right_ipin_3.mux_l1_in_4__A0
timestamp 1679235063
transform 1 0 10856 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_cby_0__1_.cby_0__1_.mux_right_ipin_3.mux_l1_in_4__A1
timestamp 1679235063
transform 1 0 10488 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_cby_0__1_.cby_0__1_.mux_right_ipin_3.mux_l2_in_2__A0
timestamp 1679235063
transform 1 0 9384 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_cby_0__1_.cby_0__1_.mux_right_ipin_3.mux_l2_in_3__A1
timestamp 1679235063
transform 1 0 10028 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_cby_0__1_.grid_io_left_left_0__1_.logical_tile_io_mode_io__0.logical_tile_io_mode_physical__iopad_0.io_0_.ISOL_EN_GATE_B_N
timestamp 1679235063
transform 1 0 3496 0 1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_cby_0__1_.grid_io_left_left_0__1_.logical_tile_io_mode_io__0.logical_tile_io_mode_physical__iopad_0.io_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_0__RESET_B
timestamp 1679235063
transform 1 0 5980 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_cby_0__1_.grid_io_left_left_0__1_.logical_tile_io_mode_io__1.logical_tile_io_mode_physical__iopad_0.io_0_.ISOL_EN_GATE_B_N
timestamp 1679235063
transform 1 0 2944 0 -1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_cby_0__1_.grid_io_left_left_0__1_.logical_tile_io_mode_io__1.logical_tile_io_mode_physical__iopad_0.io_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_0__RESET_B
timestamp 1679235063
transform 1 0 5980 0 -1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_cby_0__1_.grid_io_left_left_0__1_.logical_tile_io_mode_io__2.logical_tile_io_mode_physical__iopad_0.io_0_.ISOL_EN_GATE_B_N
timestamp 1679235063
transform 1 0 3956 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_cby_0__1_.grid_io_left_left_0__1_.logical_tile_io_mode_io__2.logical_tile_io_mode_physical__iopad_0.io_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_0__RESET_B
timestamp 1679235063
transform 1 0 5980 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_cby_0__1_.grid_io_left_left_0__1_.logical_tile_io_mode_io__3.logical_tile_io_mode_physical__iopad_0.io_0_.ISOL_EN_GATE_A
timestamp 1679235063
transform 1 0 7544 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_cby_0__1_.grid_io_left_left_0__1_.logical_tile_io_mode_io__3.logical_tile_io_mode_physical__iopad_0.io_0_.ISOL_EN_GATE_B_N
timestamp 1679235063
transform 1 0 6716 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_cby_0__1_.grid_io_left_left_0__1_.logical_tile_io_mode_io__3.logical_tile_io_mode_physical__iopad_0.io_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_0__RESET_B
timestamp 1679235063
transform 1 0 12328 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_0_prog_clk_A
timestamp 1679235063
transform 1 0 16652 0 1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_4_0_0_prog_clk_A
timestamp 1679235063
transform 1 0 10304 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_4_1_0_prog_clk_A
timestamp 1679235063
transform 1 0 12696 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_4_2_0_prog_clk_A
timestamp 1679235063
transform 1 0 9384 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_4_3_0_prog_clk_A
timestamp 1679235063
transform 1 0 11408 0 1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_4_4_0_prog_clk_A
timestamp 1679235063
transform 1 0 19228 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_4_5_0_prog_clk_A
timestamp 1679235063
transform 1 0 20056 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_4_6_0_prog_clk_A
timestamp 1679235063
transform 1 0 17664 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_4_7_0_prog_clk_A
timestamp 1679235063
transform 1 0 20516 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_4_8_0_prog_clk_A
timestamp 1679235063
transform 1 0 10304 0 -1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_4_9_0_prog_clk_A
timestamp 1679235063
transform 1 0 10948 0 1 35904
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_4_10_0_prog_clk_A
timestamp 1679235063
transform 1 0 10304 0 1 40256
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_4_11_0_prog_clk_A
timestamp 1679235063
transform 1 0 13064 0 -1 41344
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_4_12_0_prog_clk_A
timestamp 1679235063
transform 1 0 18584 0 1 38080
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_4_13_0_prog_clk_A
timestamp 1679235063
transform 1 0 20976 0 1 38080
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_4_14_0_prog_clk_A
timestamp 1679235063
transform 1 0 17572 0 1 42432
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_4_15_0_prog_clk_A
timestamp 1679235063
transform 1 0 20516 0 1 43520
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_hold107_A
timestamp 1679235063
transform 1 0 20332 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input1_A
timestamp 1679235063
transform 1 0 2024 0 -1 53312
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input2_A
timestamp 1679235063
transform 1 0 2024 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input3_A
timestamp 1679235063
transform 1 0 21804 0 -1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input4_A
timestamp 1679235063
transform 1 0 25208 0 1 33728
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input5_A
timestamp 1679235063
transform 1 0 24564 0 1 35904
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input6_A
timestamp 1679235063
transform 1 0 24748 0 1 35904
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input7_A
timestamp 1679235063
transform 1 0 23920 0 1 38080
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input8_A
timestamp 1679235063
transform 1 0 21804 0 -1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input9_A
timestamp 1679235063
transform 1 0 23000 0 -1 40256
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input10_A
timestamp 1679235063
transform 1 0 23460 0 1 40256
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input11_A
timestamp 1679235063
transform 1 0 22448 0 -1 41344
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input12_A
timestamp 1679235063
transform 1 0 24104 0 1 45696
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input13_A
timestamp 1679235063
transform 1 0 21804 0 -1 42432
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input14_A
timestamp 1679235063
transform 1 0 20884 0 -1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input15_A
timestamp 1679235063
transform 1 0 22816 0 1 42432
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input16_A
timestamp 1679235063
transform 1 0 23184 0 -1 43520
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input17_A
timestamp 1679235063
transform 1 0 24104 0 -1 46784
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input18_A
timestamp 1679235063
transform 1 0 25208 0 1 46784
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input19_A
timestamp 1679235063
transform 1 0 24380 0 1 46784
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input20_A
timestamp 1679235063
transform 1 0 25208 0 1 47872
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input21_A
timestamp 1679235063
transform 1 0 25392 0 1 47872
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input22_A
timestamp 1679235063
transform 1 0 24748 0 1 50048
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input23_A
timestamp 1679235063
transform 1 0 24748 0 1 48960
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input24_A
timestamp 1679235063
transform 1 0 24564 0 1 50048
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input25_A
timestamp 1679235063
transform 1 0 23552 0 -1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input26_A
timestamp 1679235063
transform 1 0 25116 0 -1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input27_A
timestamp 1679235063
transform 1 0 25392 0 -1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input28_A
timestamp 1679235063
transform 1 0 25208 0 -1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input29_A
timestamp 1679235063
transform 1 0 24748 0 1 30464
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input30_A
timestamp 1679235063
transform 1 0 24748 0 1 31552
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input31_A
timestamp 1679235063
transform 1 0 24748 0 1 32640
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input32_A
timestamp 1679235063
transform 1 0 24748 0 -1 32640
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input33_A
timestamp 1679235063
transform 1 0 2392 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input34_A
timestamp 1679235063
transform 1 0 4600 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input35_A
timestamp 1679235063
transform 1 0 6072 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input36_A
timestamp 1679235063
transform 1 0 6348 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input37_A
timestamp 1679235063
transform 1 0 6348 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input38_A
timestamp 1679235063
transform 1 0 7176 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input39_A
timestamp 1679235063
transform 1 0 6348 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input40_A
timestamp 1679235063
transform 1 0 6532 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input41_A
timestamp 1679235063
transform 1 0 7636 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input42_A
timestamp 1679235063
transform 1 0 7452 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input43_A
timestamp 1679235063
transform 1 0 8648 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input44_A
timestamp 1679235063
transform 1 0 2208 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input45_A
timestamp 1679235063
transform 1 0 9936 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input46_A
timestamp 1679235063
transform 1 0 9476 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input47_A
timestamp 1679235063
transform 1 0 9660 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input48_A
timestamp 1679235063
transform 1 0 9016 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input49_A
timestamp 1679235063
transform 1 0 11040 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input50_A
timestamp 1679235063
transform 1 0 10396 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input51_A
timestamp 1679235063
transform 1 0 10580 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input52_A
timestamp 1679235063
transform 1 0 11224 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input53_A
timestamp 1679235063
transform 1 0 14076 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input54_A
timestamp 1679235063
transform 1 0 9200 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input55_A
timestamp 1679235063
transform 1 0 1380 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input56_A
timestamp 1679235063
transform 1 0 2852 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input57_A
timestamp 1679235063
transform 1 0 3036 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input58_A
timestamp 1679235063
transform 1 0 3220 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input59_A
timestamp 1679235063
transform 1 0 3496 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input60_A
timestamp 1679235063
transform 1 0 4324 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input61_A
timestamp 1679235063
transform 1 0 5796 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input62_A
timestamp 1679235063
transform 1 0 4692 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input63_A
timestamp 1679235063
transform 1 0 14076 0 -1 54400
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input64_A
timestamp 1679235063
transform 1 0 16284 0 1 53312
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input65_A
timestamp 1679235063
transform 1 0 18860 0 -1 54400
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input66_A
timestamp 1679235063
transform 1 0 17204 0 -1 53312
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input67_A
timestamp 1679235063
transform 1 0 18860 0 1 53312
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input68_A
timestamp 1679235063
transform 1 0 18676 0 1 53312
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input69_A
timestamp 1679235063
transform 1 0 19688 0 -1 53312
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input70_A
timestamp 1679235063
transform 1 0 19320 0 -1 53312
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input71_A
timestamp 1679235063
transform 1 0 19504 0 -1 53312
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input72_A
timestamp 1679235063
transform 1 0 21436 0 -1 54400
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input73_A
timestamp 1679235063
transform 1 0 20700 0 1 53312
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input74_A
timestamp 1679235063
transform 1 0 13156 0 -1 52224
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input75_A
timestamp 1679235063
transform 1 0 20792 0 -1 53312
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input76_A
timestamp 1679235063
transform 1 0 21160 0 -1 53312
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input77_A
timestamp 1679235063
transform 1 0 20976 0 -1 53312
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input78_A
timestamp 1679235063
transform 1 0 23276 0 -1 54400
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input79_A
timestamp 1679235063
transform 1 0 21804 0 -1 53312
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input80_A
timestamp 1679235063
transform 1 0 22264 0 -1 53312
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input81_A
timestamp 1679235063
transform 1 0 22540 0 -1 53312
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input82_A
timestamp 1679235063
transform 1 0 24380 0 1 53312
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input83_A
timestamp 1679235063
transform 1 0 22908 0 -1 53312
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input84_A
timestamp 1679235063
transform 1 0 24380 0 -1 53312
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input85_A
timestamp 1679235063
transform 1 0 14076 0 1 52224
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input86_A
timestamp 1679235063
transform 1 0 14812 0 1 53312
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input87_A
timestamp 1679235063
transform 1 0 14904 0 -1 53312
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input88_A
timestamp 1679235063
transform 1 0 14444 0 -1 54400
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input89_A
timestamp 1679235063
transform 1 0 16100 0 -1 54400
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input90_A
timestamp 1679235063
transform 1 0 16100 0 1 53312
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input91_A
timestamp 1679235063
transform 1 0 16376 0 -1 53312
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input92_A
timestamp 1679235063
transform 1 0 16376 0 -1 54400
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input93_A
timestamp 1679235063
transform 1 0 2024 0 -1 33728
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input94_A
timestamp 1679235063
transform 1 0 2024 0 1 35904
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input95_A
timestamp 1679235063
transform 1 0 2024 0 1 38080
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input96_A
timestamp 1679235063
transform 1 0 2024 0 -1 41344
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input97_A
timestamp 1679235063
transform 1 0 2116 0 -1 43520
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input98_A
timestamp 1679235063
transform 1 0 25392 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input99_A
timestamp 1679235063
transform 1 0 24656 0 -1 51136
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input100_A
timestamp 1679235063
transform 1 0 25392 0 -1 52224
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input101_A
timestamp 1679235063
transform 1 0 24656 0 1 52224
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input102_A
timestamp 1679235063
transform 1 0 24656 0 -1 53312
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input103_A
timestamp 1679235063
transform 1 0 25208 0 -1 52224
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input104_A
timestamp 1679235063
transform 1 0 24472 0 1 52224
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input105_A
timestamp 1679235063
transform 1 0 24564 0 -1 54400
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input106_A
timestamp 1679235063
transform 1 0 24380 0 -1 54400
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output107_A
timestamp 1679235063
transform 1 0 17848 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output108_A
timestamp 1679235063
transform 1 0 3220 0 1 48960
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output141_A
timestamp 1679235063
transform 1 0 18492 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__1_.mem_bottom_track_1.sky130_fd_sc_hd__dfrtp_1_0__RESET_B
timestamp 1679235063
transform 1 0 21068 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__1_.mem_bottom_track_1.sky130_fd_sc_hd__dfrtp_1_1__RESET_B
timestamp 1679235063
transform 1 0 18952 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__1_.mem_bottom_track_1.sky130_fd_sc_hd__dfrtp_1_2__RESET_B
timestamp 1679235063
transform 1 0 20700 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__1_.mem_bottom_track_3.sky130_fd_sc_hd__dfrtp_1_0__RESET_B
timestamp 1679235063
transform 1 0 21436 0 1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__1_.mem_bottom_track_3.sky130_fd_sc_hd__dfrtp_1_1__RESET_B
timestamp 1679235063
transform 1 0 21804 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__1_.mem_bottom_track_3.sky130_fd_sc_hd__dfrtp_1_2__RESET_B
timestamp 1679235063
transform 1 0 21896 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__1_.mem_bottom_track_5.sky130_fd_sc_hd__dfrtp_1_0__RESET_B
timestamp 1679235063
transform 1 0 25116 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__1_.mem_bottom_track_5.sky130_fd_sc_hd__dfrtp_1_1__RESET_B
timestamp 1679235063
transform 1 0 25116 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__1_.mem_bottom_track_5.sky130_fd_sc_hd__dfrtp_1_2__RESET_B
timestamp 1679235063
transform 1 0 25208 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__1_.mem_bottom_track_7.sky130_fd_sc_hd__dfrtp_1_0__RESET_B
timestamp 1679235063
transform 1 0 25024 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__1_.mem_bottom_track_7.sky130_fd_sc_hd__dfrtp_1_1__RESET_B
timestamp 1679235063
transform 1 0 19228 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__1_.mem_bottom_track_7.sky130_fd_sc_hd__dfrtp_1_2__RESET_B
timestamp 1679235063
transform 1 0 18768 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__1_.mem_bottom_track_11.sky130_fd_sc_hd__dfrtp_1_0__RESET_B
timestamp 1679235063
transform 1 0 16652 0 -1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__1_.mem_bottom_track_11.sky130_fd_sc_hd__dfrtp_1_1__RESET_B
timestamp 1679235063
transform 1 0 14996 0 -1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__1_.mem_bottom_track_11.sky130_fd_sc_hd__dfrtp_1_2__RESET_B
timestamp 1679235063
transform 1 0 15272 0 -1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__1_.mem_bottom_track_13.sky130_fd_sc_hd__dfrtp_1_0__RESET_B
timestamp 1679235063
transform 1 0 18676 0 1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__1_.mem_bottom_track_13.sky130_fd_sc_hd__dfrtp_1_1__RESET_B
timestamp 1679235063
transform 1 0 21160 0 -1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__1_.mem_bottom_track_13.sky130_fd_sc_hd__dfrtp_1_2__RESET_B
timestamp 1679235063
transform 1 0 21988 0 -1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__1_.mem_bottom_track_21.sky130_fd_sc_hd__dfrtp_1_0__RESET_B
timestamp 1679235063
transform 1 0 25116 0 -1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__1_.mem_bottom_track_21.sky130_fd_sc_hd__dfrtp_1_1__RESET_B
timestamp 1679235063
transform 1 0 24104 0 -1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__1_.mem_bottom_track_21.sky130_fd_sc_hd__dfrtp_1_2__RESET_B
timestamp 1679235063
transform 1 0 25024 0 -1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__1_.mem_bottom_track_29.sky130_fd_sc_hd__dfrtp_1_0__RESET_B
timestamp 1679235063
transform 1 0 24104 0 -1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__1_.mem_bottom_track_29.sky130_fd_sc_hd__dfrtp_1_1__RESET_B
timestamp 1679235063
transform 1 0 18952 0 -1 30464
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__1_.mem_bottom_track_29.sky130_fd_sc_hd__dfrtp_1_2__RESET_B
timestamp 1679235063
transform 1 0 16652 0 -1 30464
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__1_.mem_bottom_track_37.sky130_fd_sc_hd__dfrtp_1_0__RESET_B
timestamp 1679235063
transform 1 0 18492 0 1 31552
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__1_.mem_bottom_track_37.sky130_fd_sc_hd__dfrtp_1_1__RESET_B
timestamp 1679235063
transform 1 0 16008 0 -1 33728
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__1_.mem_bottom_track_37.sky130_fd_sc_hd__dfrtp_1_2__RESET_B
timestamp 1679235063
transform 1 0 14628 0 -1 31552
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__1_.mem_bottom_track_45.sky130_fd_sc_hd__dfrtp_1_0__RESET_B
timestamp 1679235063
transform 1 0 17664 0 1 33728
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__1_.mem_bottom_track_45.sky130_fd_sc_hd__dfrtp_1_1__RESET_B
timestamp 1679235063
transform 1 0 21252 0 -1 35904
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__1_.mem_bottom_track_45.sky130_fd_sc_hd__dfrtp_1_2__RESET_B
timestamp 1679235063
transform 1 0 21528 0 -1 33728
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__1_.mem_bottom_track_53.sky130_fd_sc_hd__dfrtp_1_0__RESET_B
timestamp 1679235063
transform 1 0 17480 0 1 34816
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__1_.mem_bottom_track_53.sky130_fd_sc_hd__dfrtp_1_1__RESET_B
timestamp 1679235063
transform 1 0 11224 0 1 43520
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__1_.mem_right_track_0.sky130_fd_sc_hd__dfrtp_1_0__RESET_B
timestamp 1679235063
transform 1 0 20884 0 -1 35904
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__1_.mem_right_track_0.sky130_fd_sc_hd__dfrtp_1_1__RESET_B
timestamp 1679235063
transform 1 0 24748 0 -1 31552
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__1_.mem_right_track_0.sky130_fd_sc_hd__dfrtp_1_2__RESET_B
timestamp 1679235063
transform 1 0 25392 0 -1 30464
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__1_.mem_right_track_2.sky130_fd_sc_hd__dfrtp_1_0__RESET_B
timestamp 1679235063
transform 1 0 25392 0 1 33728
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__1_.mem_right_track_2.sky130_fd_sc_hd__dfrtp_1_1__RESET_B
timestamp 1679235063
transform 1 0 24656 0 1 43520
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__1_.mem_right_track_2.sky130_fd_sc_hd__dfrtp_1_2__RESET_B
timestamp 1679235063
transform 1 0 25392 0 1 46784
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__1_.mem_right_track_4.sky130_fd_sc_hd__dfrtp_1_0__RESET_B
timestamp 1679235063
transform 1 0 24472 0 1 43520
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__1_.mem_right_track_4.sky130_fd_sc_hd__dfrtp_1_1__RESET_B
timestamp 1679235063
transform 1 0 21988 0 -1 39168
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__1_.mem_right_track_4.sky130_fd_sc_hd__dfrtp_1_2__RESET_B
timestamp 1679235063
transform 1 0 24196 0 -1 34816
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__1_.mem_right_track_6.sky130_fd_sc_hd__dfrtp_1_0__RESET_B
timestamp 1679235063
transform 1 0 25300 0 -1 35904
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__1_.mem_right_track_6.sky130_fd_sc_hd__dfrtp_1_1__RESET_B
timestamp 1679235063
transform 1 0 24380 0 1 35904
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__1_.mem_right_track_6.sky130_fd_sc_hd__dfrtp_1_2__RESET_B
timestamp 1679235063
transform 1 0 21804 0 -1 39168
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__1_.mem_right_track_8.sky130_fd_sc_hd__dfrtp_1_0__RESET_B
timestamp 1679235063
transform 1 0 22816 0 -1 40256
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__1_.mem_right_track_8.sky130_fd_sc_hd__dfrtp_1_1__RESET_B
timestamp 1679235063
transform 1 0 24104 0 -1 45696
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__1_.mem_right_track_8.sky130_fd_sc_hd__dfrtp_1_2__RESET_B
timestamp 1679235063
transform 1 0 23920 0 1 45696
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__1_.mem_right_track_10.sky130_fd_sc_hd__dfrtp_1_0__RESET_B
timestamp 1679235063
transform 1 0 23736 0 1 45696
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__1_.mem_right_track_10.sky130_fd_sc_hd__dfrtp_1_1__RESET_B
timestamp 1679235063
transform 1 0 21988 0 -1 42432
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__1_.mem_right_track_10.sky130_fd_sc_hd__dfrtp_1_2__RESET_B
timestamp 1679235063
transform 1 0 20792 0 -1 42432
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__1_.mem_right_track_12.sky130_fd_sc_hd__dfrtp_1_0__RESET_B
timestamp 1679235063
transform 1 0 21712 0 1 44608
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__1_.mem_right_track_12.sky130_fd_sc_hd__dfrtp_1_1__RESET_B
timestamp 1679235063
transform 1 0 21528 0 1 45696
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__1_.mem_right_track_12.sky130_fd_sc_hd__dfrtp_1_2__RESET_B
timestamp 1679235063
transform 1 0 20332 0 1 43520
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__1_.mem_right_track_14.sky130_fd_sc_hd__dfrtp_1_0__RESET_B
timestamp 1679235063
transform 1 0 21436 0 -1 45696
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__1_.mem_right_track_14.sky130_fd_sc_hd__dfrtp_1_1__RESET_B
timestamp 1679235063
transform 1 0 18952 0 -1 46784
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__1_.mem_right_track_14.sky130_fd_sc_hd__dfrtp_1_2__RESET_B
timestamp 1679235063
transform 1 0 18676 0 1 43520
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__1_.mem_right_track_16.sky130_fd_sc_hd__dfrtp_1_0__RESET_B
timestamp 1679235063
transform 1 0 19136 0 -1 46784
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__1_.mem_right_track_16.sky130_fd_sc_hd__dfrtp_1_1__RESET_B
timestamp 1679235063
transform 1 0 17756 0 1 46784
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__1_.mem_right_track_16.sky130_fd_sc_hd__dfrtp_1_2__RESET_B
timestamp 1679235063
transform 1 0 17112 0 1 44608
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__1_.mem_right_track_18.sky130_fd_sc_hd__dfrtp_1_0__RESET_B
timestamp 1679235063
transform 1 0 16744 0 1 45696
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__1_.mem_right_track_18.sky130_fd_sc_hd__dfrtp_1_1__RESET_B
timestamp 1679235063
transform 1 0 16376 0 -1 45696
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__1_.mem_right_track_18.sky130_fd_sc_hd__dfrtp_1_2__RESET_B
timestamp 1679235063
transform 1 0 15824 0 -1 41344
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__1_.mem_right_track_20.sky130_fd_sc_hd__dfrtp_1_0__RESET_B
timestamp 1679235063
transform 1 0 14996 0 -1 40256
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__1_.mem_right_track_20.sky130_fd_sc_hd__dfrtp_1_1__RESET_B
timestamp 1679235063
transform 1 0 13892 0 -1 38080
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__1_.mem_right_track_20.sky130_fd_sc_hd__dfrtp_1_2__RESET_B
timestamp 1679235063
transform 1 0 13432 0 1 33728
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__1_.mem_right_track_22.sky130_fd_sc_hd__dfrtp_1_0__RESET_B
timestamp 1679235063
transform 1 0 13708 0 -1 35904
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__1_.mem_right_track_22.sky130_fd_sc_hd__dfrtp_1_1__RESET_B
timestamp 1679235063
transform 1 0 12328 0 1 34816
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__1_.mem_right_track_22.sky130_fd_sc_hd__dfrtp_1_2__RESET_B
timestamp 1679235063
transform 1 0 11500 0 -1 31552
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__1_.mem_right_track_24.sky130_fd_sc_hd__dfrtp_1_0__RESET_B
timestamp 1679235063
transform 1 0 11500 0 -1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__1_.mem_right_track_24.sky130_fd_sc_hd__dfrtp_1_1__RESET_B
timestamp 1679235063
transform 1 0 11040 0 1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__1_.mem_right_track_26.sky130_fd_sc_hd__dfrtp_1_0__RESET_B
timestamp 1679235063
transform 1 0 10948 0 -1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__1_.mem_right_track_26.sky130_fd_sc_hd__dfrtp_1_1__RESET_B
timestamp 1679235063
transform 1 0 9016 0 -1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__1_.mem_right_track_28.sky130_fd_sc_hd__dfrtp_1_0__RESET_B
timestamp 1679235063
transform 1 0 8556 0 -1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__1_.mem_right_track_28.sky130_fd_sc_hd__dfrtp_1_1__RESET_B
timestamp 1679235063
transform 1 0 8556 0 -1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__1_.mem_right_track_30.sky130_fd_sc_hd__dfrtp_1_0__RESET_B
timestamp 1679235063
transform 1 0 8464 0 1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__1_.mem_right_track_30.sky130_fd_sc_hd__dfrtp_1_1__RESET_B
timestamp 1679235063
transform 1 0 9476 0 -1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__1_.mem_right_track_32.sky130_fd_sc_hd__dfrtp_1_0__RESET_B
timestamp 1679235063
transform 1 0 11132 0 -1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__1_.mem_right_track_32.sky130_fd_sc_hd__dfrtp_1_1__RESET_B
timestamp 1679235063
transform 1 0 13156 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__1_.mem_right_track_34.sky130_fd_sc_hd__dfrtp_1_0__RESET_B
timestamp 1679235063
transform 1 0 15272 0 1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__1_.mem_right_track_34.sky130_fd_sc_hd__dfrtp_1_1__RESET_B
timestamp 1679235063
transform 1 0 16928 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__1_.mem_right_track_36.sky130_fd_sc_hd__dfrtp_1_0__RESET_B
timestamp 1679235063
transform 1 0 15088 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__1_.mem_right_track_36.sky130_fd_sc_hd__dfrtp_1_1__RESET_B
timestamp 1679235063
transform 1 0 13064 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__1_.mem_right_track_36.sky130_fd_sc_hd__dfrtp_1_2__RESET_B
timestamp 1679235063
transform 1 0 10856 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__1_.mem_right_track_38.sky130_fd_sc_hd__dfrtp_1_0__RESET_B
timestamp 1679235063
transform 1 0 11500 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__1_.mem_right_track_38.sky130_fd_sc_hd__dfrtp_1_1__RESET_B
timestamp 1679235063
transform 1 0 13800 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__1_.mem_right_track_40.sky130_fd_sc_hd__dfrtp_1_0__RESET_B
timestamp 1679235063
transform 1 0 16192 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__1_.mem_right_track_40.sky130_fd_sc_hd__dfrtp_1_1__RESET_B
timestamp 1679235063
transform 1 0 17388 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__1_.mem_right_track_44.sky130_fd_sc_hd__dfrtp_1_0__RESET_B
timestamp 1679235063
transform 1 0 17756 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__1_.mem_right_track_44.sky130_fd_sc_hd__dfrtp_1_1__RESET_B
timestamp 1679235063
transform 1 0 17480 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__1_.mem_right_track_46.sky130_fd_sc_hd__dfrtp_1_0__RESET_B
timestamp 1679235063
transform 1 0 18860 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__1_.mem_right_track_46.sky130_fd_sc_hd__dfrtp_1_1__RESET_B
timestamp 1679235063
transform 1 0 19872 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__1_.mem_right_track_48.sky130_fd_sc_hd__dfrtp_1_0__RESET_B
timestamp 1679235063
transform 1 0 21528 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__1_.mem_right_track_48.sky130_fd_sc_hd__dfrtp_1_1__RESET_B
timestamp 1679235063
transform 1 0 23920 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__1_.mem_right_track_50.sky130_fd_sc_hd__dfrtp_1_0__RESET_B
timestamp 1679235063
transform 1 0 24196 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__1_.mem_right_track_50.sky130_fd_sc_hd__dfrtp_1_1__RESET_B
timestamp 1679235063
transform 1 0 24012 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__1_.mem_right_track_52.sky130_fd_sc_hd__dfrtp_1_0__RESET_B
timestamp 1679235063
transform 1 0 23736 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__1_.mem_right_track_52.sky130_fd_sc_hd__dfrtp_1_1__RESET_B
timestamp 1679235063
transform 1 0 23000 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__1_.mem_right_track_54.sky130_fd_sc_hd__dfrtp_1_0__RESET_B
timestamp 1679235063
transform 1 0 22264 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__1_.mem_right_track_54.sky130_fd_sc_hd__dfrtp_1_1__RESET_B
timestamp 1679235063
transform 1 0 21068 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__1_.mem_right_track_56.sky130_fd_sc_hd__dfrtp_1_0__RESET_B
timestamp 1679235063
transform 1 0 20056 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__1_.mem_right_track_56.sky130_fd_sc_hd__dfrtp_1_1__RESET_B
timestamp 1679235063
transform 1 0 21436 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__1_.mem_top_track_0.sky130_fd_sc_hd__dfrtp_1_0__CLK
timestamp 1679235063
transform 1 0 6348 0 -1 50048
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__1_.mem_top_track_0.sky130_fd_sc_hd__dfrtp_1_0__RESET_B
timestamp 1679235063
transform 1 0 6532 0 -1 50048
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__1_.mem_top_track_0.sky130_fd_sc_hd__dfrtp_1_1__CLK
timestamp 1679235063
transform 1 0 11132 0 -1 45696
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__1_.mem_top_track_0.sky130_fd_sc_hd__dfrtp_1_1__D
timestamp 1679235063
transform 1 0 8740 0 -1 45696
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__1_.mem_top_track_0.sky130_fd_sc_hd__dfrtp_1_1__RESET_B
timestamp 1679235063
transform 1 0 11776 0 1 44608
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__1_.mem_top_track_0.sky130_fd_sc_hd__dfrtp_1_2__RESET_B
timestamp 1679235063
transform 1 0 11960 0 -1 47872
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__1_.mem_top_track_2.sky130_fd_sc_hd__dfrtp_1_0__RESET_B
timestamp 1679235063
transform 1 0 14076 0 1 45696
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__1_.mem_top_track_2.sky130_fd_sc_hd__dfrtp_1_1__RESET_B
timestamp 1679235063
transform 1 0 15088 0 -1 44608
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__1_.mem_top_track_2.sky130_fd_sc_hd__dfrtp_1_2__RESET_B
timestamp 1679235063
transform 1 0 14168 0 1 46784
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__1_.mem_top_track_4.sky130_fd_sc_hd__dfrtp_1_0__RESET_B
timestamp 1679235063
transform 1 0 15824 0 -1 43520
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__1_.mem_top_track_4.sky130_fd_sc_hd__dfrtp_1_1__D
timestamp 1679235063
transform 1 0 13432 0 1 39168
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__1_.mem_top_track_4.sky130_fd_sc_hd__dfrtp_1_1__RESET_B
timestamp 1679235063
transform 1 0 13248 0 1 39168
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__1_.mem_top_track_4.sky130_fd_sc_hd__dfrtp_1_2__CLK
timestamp 1679235063
transform 1 0 11040 0 -1 41344
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__1_.mem_top_track_4.sky130_fd_sc_hd__dfrtp_1_2__RESET_B
timestamp 1679235063
transform 1 0 11224 0 -1 41344
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__1_.mem_top_track_6.sky130_fd_sc_hd__dfrtp_1_0__RESET_B
timestamp 1679235063
transform 1 0 10764 0 1 40256
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__1_.mem_top_track_6.sky130_fd_sc_hd__dfrtp_1_1__D
timestamp 1679235063
transform 1 0 8648 0 -1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__1_.mem_top_track_6.sky130_fd_sc_hd__dfrtp_1_1__RESET_B
timestamp 1679235063
transform 1 0 8832 0 -1 38080
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__1_.mem_top_track_6.sky130_fd_sc_hd__dfrtp_1_2__CLK
timestamp 1679235063
transform 1 0 8648 0 1 38080
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__1_.mem_top_track_6.sky130_fd_sc_hd__dfrtp_1_2__RESET_B
timestamp 1679235063
transform 1 0 7268 0 -1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__1_.mem_top_track_10.sky130_fd_sc_hd__dfrtp_1_0__RESET_B
timestamp 1679235063
transform 1 0 9016 0 -1 38080
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__1_.mem_top_track_10.sky130_fd_sc_hd__dfrtp_1_1__D
timestamp 1679235063
transform 1 0 7084 0 -1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__1_.mem_top_track_10.sky130_fd_sc_hd__dfrtp_1_1__RESET_B
timestamp 1679235063
transform 1 0 7268 0 1 35904
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__1_.mem_top_track_10.sky130_fd_sc_hd__dfrtp_1_2__RESET_B
timestamp 1679235063
transform 1 0 6348 0 -1 35904
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__1_.mem_top_track_12.sky130_fd_sc_hd__dfrtp_1_0__RESET_B
timestamp 1679235063
transform 1 0 7360 0 -1 34816
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__1_.mem_top_track_12.sky130_fd_sc_hd__dfrtp_1_1__D
timestamp 1679235063
transform 1 0 8464 0 1 31552
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__1_.mem_top_track_12.sky130_fd_sc_hd__dfrtp_1_1__RESET_B
timestamp 1679235063
transform 1 0 8280 0 1 31552
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__1_.mem_top_track_12.sky130_fd_sc_hd__dfrtp_1_2__RESET_B
timestamp 1679235063
transform 1 0 7176 0 -1 33728
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__1_.mem_top_track_20.sky130_fd_sc_hd__dfrtp_1_0__RESET_B
timestamp 1679235063
transform 1 0 9752 0 -1 32640
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__1_.mem_top_track_20.sky130_fd_sc_hd__dfrtp_1_1__RESET_B
timestamp 1679235063
transform 1 0 11500 0 1 31552
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__1_.mem_top_track_20.sky130_fd_sc_hd__dfrtp_1_2__RESET_B
timestamp 1679235063
transform 1 0 9752 0 -1 34816
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__1_.mem_top_track_28.sky130_fd_sc_hd__dfrtp_1_0__RESET_B
timestamp 1679235063
transform 1 0 10120 0 -1 35904
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__1_.mem_top_track_28.sky130_fd_sc_hd__dfrtp_1_1__RESET_B
timestamp 1679235063
transform 1 0 8280 0 1 34816
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__1_.mem_top_track_28.sky130_fd_sc_hd__dfrtp_1_2__RESET_B
timestamp 1679235063
transform 1 0 6072 0 1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__1_.mem_top_track_36.sky130_fd_sc_hd__dfrtp_1_0__CLK
timestamp 1679235063
transform 1 0 8372 0 1 39168
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__1_.mem_top_track_36.sky130_fd_sc_hd__dfrtp_1_0__RESET_B
timestamp 1679235063
transform 1 0 8556 0 1 39168
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__1_.mem_top_track_36.sky130_fd_sc_hd__dfrtp_1_1__CLK
timestamp 1679235063
transform 1 0 8464 0 1 40256
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__1_.mem_top_track_36.sky130_fd_sc_hd__dfrtp_1_1__RESET_B
timestamp 1679235063
transform 1 0 8648 0 1 40256
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__1_.mem_top_track_36.sky130_fd_sc_hd__dfrtp_1_2__CLK
timestamp 1679235063
transform 1 0 8004 0 1 41344
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__1_.mem_top_track_36.sky130_fd_sc_hd__dfrtp_1_2__RESET_B
timestamp 1679235063
transform 1 0 8188 0 1 41344
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__1_.mem_top_track_44.sky130_fd_sc_hd__dfrtp_1_0__CLK
timestamp 1679235063
transform 1 0 10948 0 -1 42432
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__1_.mem_top_track_44.sky130_fd_sc_hd__dfrtp_1_0__RESET_B
timestamp 1679235063
transform 1 0 9384 0 1 42432
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__1_.mem_top_track_44.sky130_fd_sc_hd__dfrtp_1_1__RESET_B
timestamp 1679235063
transform 1 0 12880 0 1 42432
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__1_.mem_top_track_52.sky130_fd_sc_hd__dfrtp_1_0__RESET_B
timestamp 1679235063
transform 1 0 16744 0 1 42432
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__1_.mem_top_track_52.sky130_fd_sc_hd__dfrtp_1_1__RESET_B
timestamp 1679235063
transform 1 0 18952 0 -1 41344
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__1_.mem_top_track_52.sky130_fd_sc_hd__dfrtp_1_2__RESET_B
timestamp 1679235063
transform 1 0 18860 0 -1 39168
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__1_.mux_bottom_track_1.mux_l1_in_0__A0
timestamp 1679235063
transform 1 0 17020 0 -1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__1_.mux_bottom_track_1.mux_l1_in_0__A1
timestamp 1679235063
transform 1 0 18584 0 -1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__1_.mux_bottom_track_1.mux_l1_in_0__S
timestamp 1679235063
transform 1 0 18400 0 -1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__1_.mux_bottom_track_1.mux_l1_in_1__A0
timestamp 1679235063
transform 1 0 21436 0 -1 32640
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__1_.mux_bottom_track_1.mux_l1_in_1__A1
timestamp 1679235063
transform 1 0 19228 0 1 31552
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__1_.mux_bottom_track_1.mux_l1_in_1__S
timestamp 1679235063
transform 1 0 19412 0 1 31552
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__1_.mux_bottom_track_1.mux_l1_in_2__A0
timestamp 1679235063
transform 1 0 12420 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__1_.mux_bottom_track_1.mux_l1_in_2__A1
timestamp 1679235063
transform 1 0 13432 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__1_.mux_bottom_track_1.mux_l1_in_2__S
timestamp 1679235063
transform 1 0 14260 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__1_.mux_bottom_track_3.mux_l1_in_0__A0
timestamp 1679235063
transform 1 0 18952 0 1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__1_.mux_bottom_track_3.mux_l1_in_0__A1
timestamp 1679235063
transform 1 0 20332 0 -1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__1_.mux_bottom_track_3.mux_l1_in_1__A1
timestamp 1679235063
transform 1 0 20792 0 1 31552
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__1_.mux_bottom_track_3.mux_l2_in_1__A1
timestamp 1679235063
transform 1 0 16744 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__1_.mux_bottom_track_5.mux_l1_in_0__A0
timestamp 1679235063
transform 1 0 19412 0 -1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__1_.mux_bottom_track_5.mux_l1_in_0__A1
timestamp 1679235063
transform 1 0 20792 0 -1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__1_.mux_bottom_track_5.mux_l1_in_1__A1
timestamp 1679235063
transform 1 0 22816 0 1 30464
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__1_.mux_bottom_track_5.mux_l1_in_2__A0
timestamp 1679235063
transform 1 0 19596 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__1_.mux_bottom_track_7.mux_l1_in_0__A0
timestamp 1679235063
transform 1 0 17204 0 1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__1_.mux_bottom_track_7.mux_l1_in_0__A1
timestamp 1679235063
transform 1 0 17664 0 1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__1_.mux_bottom_track_7.mux_l1_in_1__A1
timestamp 1679235063
transform 1 0 20976 0 1 31552
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__1_.mux_bottom_track_7.mux_l1_in_2__A0
timestamp 1679235063
transform 1 0 16376 0 1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__1_.mux_bottom_track_7.mux_l1_in_3__A1
timestamp 1679235063
transform 1 0 14996 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__1_.mux_bottom_track_11.mux_l1_in_0__A0
timestamp 1679235063
transform 1 0 18676 0 1 31552
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__1_.mux_bottom_track_11.mux_l1_in_0__A1
timestamp 1679235063
transform 1 0 18860 0 1 31552
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__1_.mux_bottom_track_11.mux_l1_in_1__A1
timestamp 1679235063
transform 1 0 19412 0 -1 34816
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__1_.mux_bottom_track_11.mux_l1_in_2__A0
timestamp 1679235063
transform 1 0 14536 0 1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__1_.mux_bottom_track_11.mux_l1_in_3__A1
timestamp 1679235063
transform 1 0 12144 0 -1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__1_.mux_bottom_track_13.mux_l1_in_0__A0
timestamp 1679235063
transform 1 0 17020 0 -1 30464
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__1_.mux_bottom_track_13.mux_l1_in_0__A1
timestamp 1679235063
transform 1 0 18400 0 -1 30464
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__1_.mux_bottom_track_13.mux_l1_in_1__A1
timestamp 1679235063
transform 1 0 21804 0 1 33728
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__1_.mux_bottom_track_13.mux_l1_in_2__A0
timestamp 1679235063
transform 1 0 17848 0 1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__1_.mux_bottom_track_21.mux_l1_in_0__A0
timestamp 1679235063
transform 1 0 19228 0 -1 30464
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__1_.mux_bottom_track_21.mux_l1_in_0__A1
timestamp 1679235063
transform 1 0 20424 0 1 30464
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__1_.mux_bottom_track_21.mux_l1_in_1__A1
timestamp 1679235063
transform 1 0 23000 0 -1 34816
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__1_.mux_bottom_track_21.mux_l1_in_2__A0
timestamp 1679235063
transform 1 0 20424 0 1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__1_.mux_bottom_track_29.mux_l1_in_0__A0
timestamp 1679235063
transform 1 0 16376 0 -1 32640
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__1_.mux_bottom_track_29.mux_l1_in_0__A1
timestamp 1679235063
transform 1 0 17572 0 1 32640
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__1_.mux_bottom_track_29.mux_l1_in_1__A1
timestamp 1679235063
transform 1 0 21160 0 1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__1_.mux_bottom_track_29.mux_l1_in_2__A0
timestamp 1679235063
transform 1 0 17848 0 1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__1_.mux_bottom_track_37.mux_l1_in_0__A0
timestamp 1679235063
transform 1 0 18768 0 1 38080
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__1_.mux_bottom_track_37.mux_l1_in_0__A1
timestamp 1679235063
transform 1 0 18952 0 1 38080
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__1_.mux_bottom_track_37.mux_l2_in_1__A1
timestamp 1679235063
transform 1 0 11224 0 -1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__1_.mux_bottom_track_45.mux_l1_in_0__A1
timestamp 1679235063
transform 1 0 20424 0 1 39168
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__1_.mux_bottom_track_53.mux_l1_in_0__A1
timestamp 1679235063
transform 1 0 15916 0 -1 39168
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__1_.mux_bottom_track_53.mux_l2_in_0__S
timestamp 1679235063
transform 1 0 10948 0 1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__1_.mux_right_track_0.mux_l1_in_0__A0
timestamp 1679235063
transform 1 0 23184 0 1 32640
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__1_.mux_right_track_0.mux_l1_in_0__A1
timestamp 1679235063
transform 1 0 23000 0 1 32640
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__1_.mux_right_track_0.mux_l1_in_1__A0
timestamp 1679235063
transform 1 0 23552 0 1 32640
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__1_.mux_right_track_0.mux_l1_in_1__A1
timestamp 1679235063
transform 1 0 23368 0 1 32640
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__1_.mux_right_track_0.mux_l2_in_1__A1
timestamp 1679235063
transform 1 0 20700 0 1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__1_.mux_right_track_2.mux_l1_in_0__A0
timestamp 1679235063
transform 1 0 21896 0 1 45696
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__1_.mux_right_track_2.mux_l1_in_1__A0
timestamp 1679235063
transform 1 0 22356 0 -1 40256
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__1_.mux_right_track_2.mux_l1_in_1__A1
timestamp 1679235063
transform 1 0 22172 0 -1 40256
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__1_.mux_right_track_2.mux_l1_in_2__A0
timestamp 1679235063
transform 1 0 19596 0 -1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__1_.mux_right_track_2.mux_l1_in_2__A1
timestamp 1679235063
transform 1 0 20976 0 -1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__1_.mux_right_track_4.mux_l1_in_0__A0
timestamp 1679235063
transform 1 0 21896 0 -1 44608
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__1_.mux_right_track_4.mux_l1_in_1__A0
timestamp 1679235063
transform 1 0 24104 0 1 38080
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__1_.mux_right_track_4.mux_l1_in_1__A1
timestamp 1679235063
transform 1 0 23736 0 1 38080
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__1_.mux_right_track_4.mux_l2_in_1__A1
timestamp 1679235063
transform 1 0 19412 0 1 33728
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__1_.mux_right_track_6.mux_l1_in_0__A0
timestamp 1679235063
transform 1 0 23000 0 -1 43520
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__1_.mux_right_track_6.mux_l1_in_1__A0
timestamp 1679235063
transform 1 0 23184 0 -1 38080
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__1_.mux_right_track_6.mux_l1_in_1__A1
timestamp 1679235063
transform 1 0 23000 0 -1 38080
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__1_.mux_right_track_6.mux_l1_in_2__A0
timestamp 1679235063
transform 1 0 18952 0 1 32640
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__1_.mux_right_track_6.mux_l1_in_2__A1
timestamp 1679235063
transform 1 0 18768 0 1 32640
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__1_.mux_right_track_8.mux_l1_in_0__A0
timestamp 1679235063
transform 1 0 21528 0 -1 46784
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__1_.mux_right_track_8.mux_l1_in_1__A0
timestamp 1679235063
transform 1 0 22080 0 1 40256
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__1_.mux_right_track_8.mux_l1_in_1__A1
timestamp 1679235063
transform 1 0 21896 0 1 40256
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__1_.mux_right_track_8.mux_l1_in_2__A0
timestamp 1679235063
transform 1 0 19228 0 1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__1_.mux_right_track_8.mux_l1_in_2__A1
timestamp 1679235063
transform 1 0 20148 0 -1 38080
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__1_.mux_right_track_10.mux_l1_in_0__A0
timestamp 1679235063
transform 1 0 19320 0 1 44608
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__1_.mux_right_track_10.mux_l1_in_1__A0
timestamp 1679235063
transform 1 0 21988 0 -1 40256
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__1_.mux_right_track_10.mux_l1_in_1__A1
timestamp 1679235063
transform 1 0 21804 0 -1 40256
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__1_.mux_right_track_10.mux_l2_in_1__A1
timestamp 1679235063
transform 1 0 16008 0 -1 35904
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__1_.mux_right_track_12.mux_l1_in_0__A0
timestamp 1679235063
transform 1 0 19320 0 -1 46784
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__1_.mux_right_track_12.mux_l2_in_0__A0
timestamp 1679235063
transform 1 0 20332 0 -1 41344
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__1_.mux_right_track_12.mux_l2_in_1__A1
timestamp 1679235063
transform 1 0 16652 0 -1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__1_.mux_right_track_14.mux_l1_in_0__A0
timestamp 1679235063
transform 1 0 19044 0 -1 47872
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__1_.mux_right_track_14.mux_l2_in_0__A0
timestamp 1679235063
transform 1 0 19228 0 1 41344
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__1_.mux_right_track_14.mux_l2_in_1__A1
timestamp 1679235063
transform 1 0 15824 0 1 38080
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__1_.mux_right_track_16.mux_l1_in_0__A1
timestamp 1679235063
transform 1 0 19228 0 -1 47872
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__1_.mux_right_track_16.mux_l2_in_0__A0
timestamp 1679235063
transform 1 0 18216 0 1 43520
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__1_.mux_right_track_16.mux_l2_in_1__A1
timestamp 1679235063
transform 1 0 14076 0 1 39168
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__1_.mux_right_track_18.mux_l1_in_0__A1
timestamp 1679235063
transform 1 0 18032 0 1 47872
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__1_.mux_right_track_18.mux_l2_in_0__A0
timestamp 1679235063
transform 1 0 17388 0 1 41344
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__1_.mux_right_track_18.mux_l2_in_1__A1
timestamp 1679235063
transform 1 0 11500 0 -1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__1_.mux_right_track_20.mux_l1_in_0__A1
timestamp 1679235063
transform 1 0 16008 0 -1 43520
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__1_.mux_right_track_20.mux_l2_in_0__A0
timestamp 1679235063
transform 1 0 15456 0 -1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__1_.mux_right_track_20.mux_l2_in_1__A1
timestamp 1679235063
transform 1 0 11684 0 1 31552
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__1_.mux_right_track_22.mux_l1_in_0__A1
timestamp 1679235063
transform 1 0 13616 0 1 40256
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__1_.mux_right_track_22.mux_l2_in_0__A0
timestamp 1679235063
transform 1 0 14076 0 -1 34816
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__1_.mux_right_track_22.mux_l2_in_1__A1
timestamp 1679235063
transform 1 0 10028 0 -1 30464
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__1_.mux_right_track_24.mux_l1_in_0__A0
timestamp 1679235063
transform 1 0 15456 0 1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__1_.mux_right_track_24.mux_l1_in_0__A1
timestamp 1679235063
transform 1 0 15272 0 1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__1_.mux_right_track_24.mux_l1_in_1__A1
timestamp 1679235063
transform 1 0 10396 0 1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__1_.mux_right_track_26.mux_l1_in_0__A0
timestamp 1679235063
transform 1 0 15456 0 1 30464
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__1_.mux_right_track_26.mux_l1_in_0__A1
timestamp 1679235063
transform 1 0 15272 0 1 30464
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__1_.mux_right_track_26.mux_l1_in_1__A1
timestamp 1679235063
transform 1 0 8740 0 -1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__1_.mux_right_track_28.mux_l1_in_0__A0
timestamp 1679235063
transform 1 0 12972 0 -1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__1_.mux_right_track_28.mux_l1_in_0__A1
timestamp 1679235063
transform 1 0 12788 0 1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__1_.mux_right_track_28.mux_l1_in_1__A1
timestamp 1679235063
transform 1 0 7084 0 1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__1_.mux_right_track_30.mux_l1_in_0__A0
timestamp 1679235063
transform 1 0 13616 0 1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__1_.mux_right_track_30.mux_l1_in_0__A1
timestamp 1679235063
transform 1 0 13800 0 1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__1_.mux_right_track_30.mux_l1_in_1__A1
timestamp 1679235063
transform 1 0 7912 0 -1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__1_.mux_right_track_32.mux_l1_in_0__A0
timestamp 1679235063
transform 1 0 14076 0 1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__1_.mux_right_track_32.mux_l1_in_0__A1
timestamp 1679235063
transform 1 0 12604 0 1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__1_.mux_right_track_32.mux_l1_in_1__A1
timestamp 1679235063
transform 1 0 10488 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__1_.mux_right_track_34.mux_l1_in_0__A0
timestamp 1679235063
transform 1 0 17664 0 1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__1_.mux_right_track_34.mux_l1_in_0__A1
timestamp 1679235063
transform 1 0 16376 0 -1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__1_.mux_right_track_34.mux_l1_in_1__A1
timestamp 1679235063
transform 1 0 12236 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__1_.mux_right_track_36.mux_l1_in_0__A0
timestamp 1679235063
transform 1 0 14352 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__1_.mux_right_track_36.mux_l1_in_0__A1
timestamp 1679235063
transform 1 0 14536 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__1_.mux_right_track_36.mux_l2_in_0__A0
timestamp 1679235063
transform 1 0 8464 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__1_.mux_right_track_38.mux_l1_in_0__A0
timestamp 1679235063
transform 1 0 12052 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__1_.mux_right_track_38.mux_l1_in_0__A1
timestamp 1679235063
transform 1 0 13432 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__1_.mux_right_track_40.mux_l1_in_0__A0
timestamp 1679235063
transform 1 0 14076 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__1_.mux_right_track_40.mux_l1_in_0__A1
timestamp 1679235063
transform 1 0 15180 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__1_.mux_right_track_44.mux_l1_in_0__A0
timestamp 1679235063
transform 1 0 15180 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__1_.mux_right_track_44.mux_l1_in_0__A1
timestamp 1679235063
transform 1 0 16376 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__1_.mux_right_track_46.mux_l1_in_0__A0
timestamp 1679235063
transform 1 0 16468 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__1_.mux_right_track_46.mux_l1_in_0__A1
timestamp 1679235063
transform 1 0 17848 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__1_.mux_right_track_48.mux_l1_in_0__A0
timestamp 1679235063
transform 1 0 19228 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__1_.mux_right_track_48.mux_l1_in_0__A1
timestamp 1679235063
transform 1 0 20056 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__1_.mux_right_track_50.mux_l1_in_0__A0
timestamp 1679235063
transform 1 0 20700 0 1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__1_.mux_right_track_50.mux_l1_in_0__A1
timestamp 1679235063
transform 1 0 20884 0 1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__1_.mux_right_track_50.mux_l1_in_1__A1
timestamp 1679235063
transform 1 0 18768 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__1_.mux_right_track_52.mux_l1_in_0__A0
timestamp 1679235063
transform 1 0 18584 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__1_.mux_right_track_52.mux_l1_in_0__A1
timestamp 1679235063
transform 1 0 20240 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__1_.mux_right_track_54.mux_l1_in_0__A1
timestamp 1679235063
transform 1 0 18676 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__1_.mux_right_track_56.mux_l1_in_0__A0
timestamp 1679235063
transform 1 0 17756 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__1_.mux_right_track_56.mux_l1_in_0__A1
timestamp 1679235063
transform 1 0 18952 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__1_.mux_top_track_0.mux_l1_in_0__A0
timestamp 1679235063
transform 1 0 9108 0 1 42432
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__1_.mux_top_track_0.mux_l1_in_0__A1
timestamp 1679235063
transform 1 0 8924 0 1 42432
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__1_.mux_top_track_0.mux_l1_in_0__S
timestamp 1679235063
transform 1 0 10120 0 -1 43520
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__1_.mux_top_track_0.mux_l1_in_1__A1
timestamp 1679235063
transform 1 0 18124 0 -1 42432
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__1_.mux_top_track_0.mux_l1_in_1__S
timestamp 1679235063
transform 1 0 16744 0 -1 42432
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__1_.mux_top_track_0.mux_l1_in_2__A0
timestamp 1679235063
transform 1 0 14536 0 -1 38080
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__1_.mux_top_track_0.mux_l1_in_2__S
timestamp 1679235063
transform 1 0 13800 0 1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__1_.mux_top_track_0.mux_l1_in_3__A1
timestamp 1679235063
transform 1 0 10396 0 -1 38080
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__1_.mux_top_track_0.mux_l1_in_3__S
timestamp 1679235063
transform 1 0 9568 0 1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__1_.mux_top_track_2.mux_l1_in_0__A0
timestamp 1679235063
transform 1 0 18032 0 1 43520
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__1_.mux_top_track_2.mux_l1_in_0__A1
timestamp 1679235063
transform 1 0 16376 0 -1 43520
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__1_.mux_top_track_2.mux_l1_in_2__A0
timestamp 1679235063
transform 1 0 10764 0 1 35904
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__1_.mux_top_track_2.mux_l1_in_2__A1
timestamp 1679235063
transform 1 0 11132 0 1 35904
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__1_.mux_top_track_4.mux_l1_in_0__A0
timestamp 1679235063
transform 1 0 16008 0 -1 41344
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__1_.mux_top_track_4.mux_l1_in_0__A1
timestamp 1679235063
transform 1 0 14812 0 1 41344
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__1_.mux_top_track_4.mux_l1_in_0__S
timestamp 1679235063
transform 1 0 14628 0 1 41344
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__1_.mux_top_track_4.mux_l1_in_1__S
timestamp 1679235063
transform 1 0 18952 0 1 35904
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__1_.mux_top_track_4.mux_l1_in_2__A0
timestamp 1679235063
transform 1 0 10488 0 -1 33728
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__1_.mux_top_track_4.mux_l1_in_2__A1
timestamp 1679235063
transform 1 0 10488 0 1 32640
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__1_.mux_top_track_4.mux_l1_in_2__S
timestamp 1679235063
transform 1 0 11868 0 1 32640
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__1_.mux_top_track_6.mux_l1_in_0__A0
timestamp 1679235063
transform 1 0 8464 0 1 41344
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__1_.mux_top_track_6.mux_l1_in_0__A1
timestamp 1679235063
transform 1 0 8648 0 1 41344
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__1_.mux_top_track_6.mux_l1_in_0__S
timestamp 1679235063
transform 1 0 10764 0 -1 42432
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__1_.mux_top_track_6.mux_l1_in_1__A1
timestamp 1679235063
transform 1 0 18400 0 1 38080
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__1_.mux_top_track_6.mux_l1_in_1__S
timestamp 1679235063
transform 1 0 17480 0 -1 38080
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__1_.mux_top_track_6.mux_l1_in_2__A0
timestamp 1679235063
transform 1 0 13156 0 -1 32640
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__1_.mux_top_track_6.mux_l1_in_2__S
timestamp 1679235063
transform 1 0 13340 0 -1 32640
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__1_.mux_top_track_6.mux_l1_in_3__A1
timestamp 1679235063
transform 1 0 7360 0 1 30464
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__1_.mux_top_track_6.mux_l1_in_3__S
timestamp 1679235063
transform 1 0 8924 0 1 30464
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__1_.mux_top_track_10.mux_l1_in_0__A0
timestamp 1679235063
transform 1 0 11040 0 1 40256
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__1_.mux_top_track_10.mux_l1_in_0__A1
timestamp 1679235063
transform 1 0 11040 0 -1 40256
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__1_.mux_top_track_10.mux_l1_in_0__S
timestamp 1679235063
transform 1 0 11224 0 -1 40256
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__1_.mux_top_track_10.mux_l1_in_1__A1
timestamp 1679235063
transform 1 0 18952 0 1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__1_.mux_top_track_10.mux_l1_in_1__S
timestamp 1679235063
transform 1 0 17296 0 -1 38080
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__1_.mux_top_track_10.mux_l1_in_2__A0
timestamp 1679235063
transform 1 0 11960 0 1 30464
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__1_.mux_top_track_10.mux_l1_in_2__S
timestamp 1679235063
transform 1 0 12144 0 1 30464
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__1_.mux_top_track_10.mux_l1_in_3__A1
timestamp 1679235063
transform 1 0 6716 0 -1 31552
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__1_.mux_top_track_10.mux_l1_in_3__S
timestamp 1679235063
transform 1 0 6900 0 -1 31552
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__1_.mux_top_track_12.mux_l1_in_0__A0
timestamp 1679235063
transform 1 0 13524 0 -1 38080
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__1_.mux_top_track_12.mux_l1_in_0__A1
timestamp 1679235063
transform 1 0 13524 0 1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__1_.mux_top_track_12.mux_l1_in_0__S
timestamp 1679235063
transform 1 0 12144 0 -1 38080
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__1_.mux_top_track_12.mux_l1_in_1__S
timestamp 1679235063
transform 1 0 16652 0 -1 32640
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__1_.mux_top_track_12.mux_l1_in_2__A0
timestamp 1679235063
transform 1 0 6348 0 1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__1_.mux_top_track_12.mux_l1_in_2__A1
timestamp 1679235063
transform 1 0 7452 0 1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__1_.mux_top_track_12.mux_l1_in_2__S
timestamp 1679235063
transform 1 0 7636 0 1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__1_.mux_top_track_20.mux_l1_in_0__A0
timestamp 1679235063
transform 1 0 15456 0 -1 35904
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__1_.mux_top_track_20.mux_l1_in_0__A1
timestamp 1679235063
transform 1 0 14076 0 -1 35904
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__1_.mux_top_track_20.mux_l1_in_2__A0
timestamp 1679235063
transform 1 0 9200 0 -1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__1_.mux_top_track_20.mux_l1_in_2__A1
timestamp 1679235063
transform 1 0 9384 0 -1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__1_.mux_top_track_28.mux_l1_in_0__A0
timestamp 1679235063
transform 1 0 13708 0 -1 38080
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__1_.mux_top_track_28.mux_l1_in_0__A1
timestamp 1679235063
transform 1 0 11224 0 -1 38080
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__1_.mux_top_track_28.mux_l1_in_1__A0
timestamp 1679235063
transform 1 0 12420 0 -1 33728
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__1_.mux_top_track_28.mux_l2_in_1__A1
timestamp 1679235063
transform 1 0 4784 0 -1 32640
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__1_.mux_top_track_36.mux_l1_in_0__A0
timestamp 1679235063
transform 1 0 12880 0 -1 41344
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__1_.mux_top_track_36.mux_l1_in_0__A1
timestamp 1679235063
transform 1 0 10580 0 1 40256
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__1_.mux_top_track_36.mux_l2_in_0__A0
timestamp 1679235063
transform 1 0 13064 0 1 39168
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__1_.mux_top_track_36.mux_l2_in_1__A1
timestamp 1679235063
transform 1 0 8740 0 -1 39168
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__1_.mux_top_track_44.mux_l1_in_1__A1
timestamp 1679235063
transform 1 0 10580 0 -1 38080
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__1_.mux_top_track_52.mux_l2_in_1__A1
timestamp 1679235063
transform 1 0 14076 0 -1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__dfrtp_4  cby_0__1_.cby_0__1_.mem_right_ipin_0.sky130_fd_sc_hd__dfrtp_1_0_ pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1679235063
transform 1 0 3956 0 -1 8704
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_2  cby_0__1_.cby_0__1_.mem_right_ipin_0.sky130_fd_sc_hd__dfrtp_1_1_ pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1679235063
transform 1 0 9108 0 1 18496
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_1  cby_0__1_.cby_0__1_.mem_right_ipin_0.sky130_fd_sc_hd__dfrtp_1_2_ pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1679235063
transform 1 0 6256 0 1 22848
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  cby_0__1_.cby_0__1_.mem_right_ipin_0.sky130_fd_sc_hd__dfrtp_1_3_
timestamp 1679235063
transform 1 0 6532 0 -1 23936
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_4  cby_0__1_.cby_0__1_.mem_right_ipin_1.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1679235063
transform 1 0 7820 0 -1 21760
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_2  cby_0__1_.cby_0__1_.mem_right_ipin_1.sky130_fd_sc_hd__dfrtp_1_1_
timestamp 1679235063
transform 1 0 11776 0 -1 16320
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_1  cby_0__1_.cby_0__1_.mem_right_ipin_1.sky130_fd_sc_hd__dfrtp_1_2_
timestamp 1679235063
transform 1 0 8096 0 -1 14144
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  cby_0__1_.cby_0__1_.mem_right_ipin_1.sky130_fd_sc_hd__dfrtp_1_3_
timestamp 1679235063
transform 1 0 6716 0 1 15232
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_4  cby_0__1_.cby_0__1_.mem_right_ipin_2.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1679235063
transform 1 0 8096 0 -1 15232
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_2  cby_0__1_.cby_0__1_.mem_right_ipin_2.sky130_fd_sc_hd__dfrtp_1_1_
timestamp 1679235063
transform 1 0 10212 0 1 15232
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_1  cby_0__1_.cby_0__1_.mem_right_ipin_2.sky130_fd_sc_hd__dfrtp_1_2_
timestamp 1679235063
transform 1 0 5980 0 1 16320
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  cby_0__1_.cby_0__1_.mem_right_ipin_2.sky130_fd_sc_hd__dfrtp_1_3_
timestamp 1679235063
transform 1 0 4784 0 1 17408
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_4  cby_0__1_.cby_0__1_.mem_right_ipin_3.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1679235063
transform 1 0 6532 0 -1 18496
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_2  cby_0__1_.cby_0__1_.mem_right_ipin_3.sky130_fd_sc_hd__dfrtp_1_1_
timestamp 1679235063
transform 1 0 8096 0 -1 19584
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_1  cby_0__1_.cby_0__1_.mem_right_ipin_3.sky130_fd_sc_hd__dfrtp_1_2_
timestamp 1679235063
transform 1 0 5336 0 1 19584
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  cby_0__1_.cby_0__1_.mem_right_ipin_3.sky130_fd_sc_hd__dfrtp_1_3_
timestamp 1679235063
transform 1 0 4140 0 1 21760
box -38 -48 1878 592
use sky130_fd_sc_hd__mux2_1  cby_0__1_.cby_0__1_.mux_right_ipin_0.mux_l1_in_0_ pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1679235063
transform 1 0 12972 0 1 15232
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  cby_0__1_.cby_0__1_.mux_right_ipin_0.mux_l1_in_1_
timestamp 1679235063
transform 1 0 12972 0 1 18496
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  cby_0__1_.cby_0__1_.mux_right_ipin_0.mux_l1_in_2_
timestamp 1679235063
transform 1 0 14260 0 1 18496
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  cby_0__1_.cby_0__1_.mux_right_ipin_0.mux_l1_in_3_
timestamp 1679235063
transform 1 0 12144 0 -1 23936
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  cby_0__1_.cby_0__1_.mux_right_ipin_0.mux_l1_in_4_
timestamp 1679235063
transform 1 0 10396 0 -1 19584
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  cby_0__1_.cby_0__1_.mux_right_ipin_0.mux_l2_in_0_
timestamp 1679235063
transform 1 0 11224 0 1 19584
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  cby_0__1_.cby_0__1_.mux_right_ipin_0.mux_l2_in_1_
timestamp 1679235063
transform 1 0 11224 0 1 20672
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  cby_0__1_.cby_0__1_.mux_right_ipin_0.mux_l2_in_2_
timestamp 1679235063
transform 1 0 9108 0 1 21760
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  cby_0__1_.cby_0__1_.mux_right_ipin_0.mux_l2_in_3__248 pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1679235063
transform 1 0 10672 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  cby_0__1_.cby_0__1_.mux_right_ipin_0.mux_l2_in_3_
timestamp 1679235063
transform 1 0 9476 0 -1 25024
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  cby_0__1_.cby_0__1_.mux_right_ipin_0.mux_l3_in_0_
timestamp 1679235063
transform 1 0 9108 0 1 20672
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  cby_0__1_.cby_0__1_.mux_right_ipin_0.mux_l3_in_1_
timestamp 1679235063
transform 1 0 7544 0 1 21760
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  cby_0__1_.cby_0__1_.mux_right_ipin_0.mux_l4_in_0_
timestamp 1679235063
transform 1 0 6440 0 1 23936
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  cby_0__1_.cby_0__1_.mux_right_ipin_0.sky130_fd_sc_hd__buf_4_0_
timestamp 1679235063
transform 1 0 4048 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  cby_0__1_.cby_0__1_.mux_right_ipin_1.mux_l1_in_0_
timestamp 1679235063
transform 1 0 15180 0 1 11968
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  cby_0__1_.cby_0__1_.mux_right_ipin_1.mux_l1_in_1_
timestamp 1679235063
transform 1 0 15088 0 1 16320
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  cby_0__1_.cby_0__1_.mux_right_ipin_1.mux_l1_in_2_
timestamp 1679235063
transform 1 0 14720 0 1 21760
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  cby_0__1_.cby_0__1_.mux_right_ipin_1.mux_l1_in_3_
timestamp 1679235063
transform 1 0 13984 0 -1 18496
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  cby_0__1_.cby_0__1_.mux_right_ipin_1.mux_l1_in_4_
timestamp 1679235063
transform 1 0 11132 0 1 21760
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  cby_0__1_.cby_0__1_.mux_right_ipin_1.mux_l2_in_0_
timestamp 1679235063
transform 1 0 12972 0 1 14144
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  cby_0__1_.cby_0__1_.mux_right_ipin_1.mux_l2_in_1_
timestamp 1679235063
transform 1 0 11776 0 1 18496
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  cby_0__1_.cby_0__1_.mux_right_ipin_1.mux_l2_in_2_
timestamp 1679235063
transform 1 0 9568 0 -1 16320
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  cby_0__1_.cby_0__1_.mux_right_ipin_1.mux_l2_in_3_
timestamp 1679235063
transform 1 0 11684 0 -1 20672
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  cby_0__1_.cby_0__1_.mux_right_ipin_1.mux_l2_in_3__249
timestamp 1679235063
transform 1 0 10948 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  cby_0__1_.cby_0__1_.mux_right_ipin_1.mux_l3_in_0_
timestamp 1679235063
transform 1 0 10304 0 1 16320
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  cby_0__1_.cby_0__1_.mux_right_ipin_1.mux_l3_in_1_
timestamp 1679235063
transform 1 0 9108 0 1 16320
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  cby_0__1_.cby_0__1_.mux_right_ipin_1.mux_l4_in_0_
timestamp 1679235063
transform 1 0 6992 0 -1 16320
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  cby_0__1_.cby_0__1_.mux_right_ipin_1.sky130_fd_sc_hd__buf_4_0_
timestamp 1679235063
transform 1 0 4140 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  cby_0__1_.cby_0__1_.mux_right_ipin_2.mux_l1_in_0_
timestamp 1679235063
transform 1 0 16376 0 1 11968
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  cby_0__1_.cby_0__1_.mux_right_ipin_2.mux_l1_in_1_
timestamp 1679235063
transform 1 0 13340 0 -1 13056
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  cby_0__1_.cby_0__1_.mux_right_ipin_2.mux_l1_in_2_
timestamp 1679235063
transform 1 0 14260 0 -1 21760
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  cby_0__1_.cby_0__1_.mux_right_ipin_2.mux_l1_in_3_
timestamp 1679235063
transform 1 0 13064 0 -1 17408
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  cby_0__1_.cby_0__1_.mux_right_ipin_2.mux_l1_in_4_
timestamp 1679235063
transform 1 0 10396 0 -1 22848
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  cby_0__1_.cby_0__1_.mux_right_ipin_2.mux_l2_in_0_
timestamp 1679235063
transform 1 0 11776 0 -1 15232
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  cby_0__1_.cby_0__1_.mux_right_ipin_2.mux_l2_in_1_
timestamp 1679235063
transform 1 0 11684 0 -1 19584
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  cby_0__1_.cby_0__1_.mux_right_ipin_2.mux_l2_in_2_
timestamp 1679235063
transform 1 0 9108 0 1 19584
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  cby_0__1_.cby_0__1_.mux_right_ipin_2.mux_l2_in_3_
timestamp 1679235063
transform 1 0 9016 0 -1 18496
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  cby_0__1_.cby_0__1_.mux_right_ipin_2.mux_l2_in_3__250
timestamp 1679235063
transform 1 0 8372 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  cby_0__1_.cby_0__1_.mux_right_ipin_2.mux_l3_in_0_
timestamp 1679235063
transform 1 0 7452 0 -1 17408
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  cby_0__1_.cby_0__1_.mux_right_ipin_2.mux_l3_in_1_
timestamp 1679235063
transform 1 0 7084 0 1 17408
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  cby_0__1_.cby_0__1_.mux_right_ipin_2.mux_l4_in_0_
timestamp 1679235063
transform 1 0 5244 0 -1 18496
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  cby_0__1_.cby_0__1_.mux_right_ipin_2.sky130_fd_sc_hd__buf_4_0_
timestamp 1679235063
transform 1 0 3312 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  cby_0__1_.cby_0__1_.mux_right_ipin_3.mux_l1_in_0_
timestamp 1679235063
transform 1 0 12972 0 -1 15232
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  cby_0__1_.cby_0__1_.mux_right_ipin_3.mux_l1_in_1_
timestamp 1679235063
transform 1 0 12788 0 -1 18496
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  cby_0__1_.cby_0__1_.mux_right_ipin_3.mux_l1_in_2_
timestamp 1679235063
transform 1 0 13248 0 -1 19584
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  cby_0__1_.cby_0__1_.mux_right_ipin_3.mux_l1_in_3_
timestamp 1679235063
transform 1 0 11776 0 -1 25024
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  cby_0__1_.cby_0__1_.mux_right_ipin_3.mux_l1_in_4_
timestamp 1679235063
transform 1 0 9844 0 -1 17408
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  cby_0__1_.cby_0__1_.mux_right_ipin_3.mux_l2_in_0_
timestamp 1679235063
transform 1 0 10396 0 -1 18496
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  cby_0__1_.cby_0__1_.mux_right_ipin_3.mux_l2_in_1_
timestamp 1679235063
transform 1 0 10396 0 -1 21760
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  cby_0__1_.cby_0__1_.mux_right_ipin_3.mux_l2_in_2_
timestamp 1679235063
transform 1 0 8188 0 -1 20672
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  cby_0__1_.cby_0__1_.mux_right_ipin_3.mux_l2_in_3_
timestamp 1679235063
transform 1 0 9200 0 -1 23936
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  cby_0__1_.cby_0__1_.mux_right_ipin_3.mux_l2_in_3__251
timestamp 1679235063
transform 1 0 9568 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  cby_0__1_.cby_0__1_.mux_right_ipin_3.mux_l3_in_0_
timestamp 1679235063
transform 1 0 7820 0 1 19584
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  cby_0__1_.cby_0__1_.mux_right_ipin_3.mux_l3_in_1_
timestamp 1679235063
transform 1 0 6624 0 -1 21760
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  cby_0__1_.cby_0__1_.mux_right_ipin_3.mux_l4_in_0_
timestamp 1679235063
transform 1 0 5152 0 -1 21760
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  cby_0__1_.cby_0__1_.mux_right_ipin_3.sky130_fd_sc_hd__buf_4_0_
timestamp 1679235063
transform 1 0 3128 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_8  cby_0__1_.grid_io_left_left_0__1_.logical_tile_io_mode_io__0.logical_tile_io_mode_physical__iopad_0.io_0_.IN_PROTECT_GATE pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1679235063
transform 1 0 3588 0 -1 31552
box -38 -48 1970 592
use sky130_fd_sc_hd__inv_1  cby_0__1_.grid_io_left_left_0__1_.logical_tile_io_mode_io__0.logical_tile_io_mode_physical__iopad_0.io_0_.INV_SOC_DIR pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1679235063
transform 1 0 3220 0 -1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__or2b_2  cby_0__1_.grid_io_left_left_0__1_.logical_tile_io_mode_io__0.logical_tile_io_mode_physical__iopad_0.io_0_.ISOL_EN_GATE pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1679235063
transform 1 0 3956 0 1 26112
box -38 -48 682 592
use sky130_fd_sc_hd__ebufn_8  cby_0__1_.grid_io_left_left_0__1_.logical_tile_io_mode_io__0.logical_tile_io_mode_physical__iopad_0.io_0_.OUT_PROTECT_GATE
timestamp 1679235063
transform 1 0 2024 0 -1 28288
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_1  cby_0__1_.grid_io_left_left_0__1_.logical_tile_io_mode_io__0.logical_tile_io_mode_physical__iopad_0.io_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1679235063
transform 1 0 3956 0 1 23936
box -38 -48 1878 592
use sky130_fd_sc_hd__ebufn_8  cby_0__1_.grid_io_left_left_0__1_.logical_tile_io_mode_io__1.logical_tile_io_mode_physical__iopad_0.io_0_.IN_PROTECT_GATE
timestamp 1679235063
transform 1 0 3956 0 1 29376
box -38 -48 1970 592
use sky130_fd_sc_hd__inv_1  cby_0__1_.grid_io_left_left_0__1_.logical_tile_io_mode_io__1.logical_tile_io_mode_physical__iopad_0.io_0_.INV_SOC_DIR
timestamp 1679235063
transform 1 0 3956 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__or2b_2  cby_0__1_.grid_io_left_left_0__1_.logical_tile_io_mode_io__1.logical_tile_io_mode_physical__iopad_0.io_0_.ISOL_EN_GATE
timestamp 1679235063
transform 1 0 3956 0 -1 26112
box -38 -48 682 592
use sky130_fd_sc_hd__ebufn_8  cby_0__1_.grid_io_left_left_0__1_.logical_tile_io_mode_io__1.logical_tile_io_mode_physical__iopad_0.io_0_.OUT_PROTECT_GATE
timestamp 1679235063
transform 1 0 1656 0 -1 25024
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_1  cby_0__1_.grid_io_left_left_0__1_.logical_tile_io_mode_io__1.logical_tile_io_mode_physical__iopad_0.io_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1679235063
transform 1 0 3956 0 -1 25024
box -38 -48 1878 592
use sky130_fd_sc_hd__ebufn_8  cby_0__1_.grid_io_left_left_0__1_.logical_tile_io_mode_io__2.logical_tile_io_mode_physical__iopad_0.io_0_.IN_PROTECT_GATE
timestamp 1679235063
transform 1 0 3956 0 1 28288
box -38 -48 1970 592
use sky130_fd_sc_hd__inv_1  cby_0__1_.grid_io_left_left_0__1_.logical_tile_io_mode_io__2.logical_tile_io_mode_physical__iopad_0.io_0_.INV_SOC_DIR
timestamp 1679235063
transform 1 0 3312 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__or2b_2  cby_0__1_.grid_io_left_left_0__1_.logical_tile_io_mode_io__2.logical_tile_io_mode_physical__iopad_0.io_0_.ISOL_EN_GATE
timestamp 1679235063
transform 1 0 4324 0 -1 22848
box -38 -48 682 592
use sky130_fd_sc_hd__ebufn_8  cby_0__1_.grid_io_left_left_0__1_.logical_tile_io_mode_io__2.logical_tile_io_mode_physical__iopad_0.io_0_.OUT_PROTECT_GATE
timestamp 1679235063
transform 1 0 1564 0 1 22848
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_1  cby_0__1_.grid_io_left_left_0__1_.logical_tile_io_mode_io__2.logical_tile_io_mode_physical__iopad_0.io_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1679235063
transform 1 0 4140 0 1 20672
box -38 -48 1878 592
use sky130_fd_sc_hd__ebufn_8  cby_0__1_.grid_io_left_left_0__1_.logical_tile_io_mode_io__3.logical_tile_io_mode_physical__iopad_0.io_0_.IN_PROTECT_GATE
timestamp 1679235063
transform 1 0 3404 0 -1 27200
box -38 -48 1970 592
use sky130_fd_sc_hd__inv_1  cby_0__1_.grid_io_left_left_0__1_.logical_tile_io_mode_io__3.logical_tile_io_mode_physical__iopad_0.io_0_.INV_SOC_DIR
timestamp 1679235063
transform 1 0 3680 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__or2b_2  cby_0__1_.grid_io_left_left_0__1_.logical_tile_io_mode_io__3.logical_tile_io_mode_physical__iopad_0.io_0_.ISOL_EN_GATE
timestamp 1679235063
transform 1 0 6900 0 1 18496
box -38 -48 682 592
use sky130_fd_sc_hd__ebufn_8  cby_0__1_.grid_io_left_left_0__1_.logical_tile_io_mode_io__3.logical_tile_io_mode_physical__iopad_0.io_0_.OUT_PROTECT_GATE
timestamp 1679235063
transform 1 0 1840 0 -1 21760
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_2  cby_0__1_.grid_io_left_left_0__1_.logical_tile_io_mode_io__3.logical_tile_io_mode_physical__iopad_0.io_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1679235063
transform 1 0 10028 0 1 14144
box -38 -48 1970 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_0_prog_clk pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1679235063
transform 1 0 14628 0 1 29376
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_8  clkbuf_4_0_0_prog_clk pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1679235063
transform 1 0 9108 0 1 17408
box -38 -48 1050 592
use sky130_fd_sc_hd__clkbuf_8  clkbuf_4_1_0_prog_clk
timestamp 1679235063
transform 1 0 11684 0 -1 17408
box -38 -48 1050 592
use sky130_fd_sc_hd__clkbuf_8  clkbuf_4_2_0_prog_clk
timestamp 1679235063
transform 1 0 8188 0 -1 22848
box -38 -48 1050 592
use sky130_fd_sc_hd__clkbuf_8  clkbuf_4_3_0_prog_clk
timestamp 1679235063
transform 1 0 10212 0 1 22848
box -38 -48 1050 592
use sky130_fd_sc_hd__clkbuf_8  clkbuf_4_4_0_prog_clk
timestamp 1679235063
transform 1 0 17940 0 1 17408
box -38 -48 1050 592
use sky130_fd_sc_hd__clkbuf_8  clkbuf_4_5_0_prog_clk
timestamp 1679235063
transform 1 0 20424 0 -1 18496
box -38 -48 1050 592
use sky130_fd_sc_hd__clkbuf_8  clkbuf_4_6_0_prog_clk
timestamp 1679235063
transform 1 0 18032 0 -1 22848
box -38 -48 1050 592
use sky130_fd_sc_hd__clkbuf_8  clkbuf_4_7_0_prog_clk
timestamp 1679235063
transform 1 0 20516 0 -1 22848
box -38 -48 1050 592
use sky130_fd_sc_hd__clkbuf_8  clkbuf_4_8_0_prog_clk
timestamp 1679235063
transform 1 0 9108 0 -1 36992
box -38 -48 1050 592
use sky130_fd_sc_hd__clkbuf_8  clkbuf_4_9_0_prog_clk
timestamp 1679235063
transform 1 0 11500 0 1 35904
box -38 -48 1050 592
use sky130_fd_sc_hd__clkbuf_8  clkbuf_4_10_0_prog_clk
timestamp 1679235063
transform 1 0 9108 0 1 40256
box -38 -48 1050 592
use sky130_fd_sc_hd__clkbuf_8  clkbuf_4_11_0_prog_clk
timestamp 1679235063
transform 1 0 11684 0 -1 41344
box -38 -48 1050 592
use sky130_fd_sc_hd__clkbuf_8  clkbuf_4_12_0_prog_clk
timestamp 1679235063
transform 1 0 19412 0 1 38080
box -38 -48 1050 592
use sky130_fd_sc_hd__clkbuf_8  clkbuf_4_13_0_prog_clk
timestamp 1679235063
transform 1 0 21344 0 1 38080
box -38 -48 1050 592
use sky130_fd_sc_hd__clkbuf_8  clkbuf_4_14_0_prog_clk
timestamp 1679235063
transform 1 0 17940 0 1 42432
box -38 -48 1050 592
use sky130_fd_sc_hd__clkbuf_8  clkbuf_4_15_0_prog_clk
timestamp 1679235063
transform 1 0 20516 0 -1 43520
box -38 -48 1050 592
use sky130_fd_sc_hd__decap_3  FILLER_0_3 pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1679235063
transform 1 0 1380 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_10 pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1679235063
transform 1 0 2024 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_18
timestamp 1679235063
transform 1 0 2760 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_26 pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1679235063
transform 1 0 3496 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_29
timestamp 1679235063
transform 1 0 3772 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_35
timestamp 1679235063
transform 1 0 4324 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_49
timestamp 1679235063
transform 1 0 5612 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_53 pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1679235063
transform 1 0 5980 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_61
timestamp 1679235063
transform 1 0 6716 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_67
timestamp 1679235063
transform 1 0 7268 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_0_81
timestamp 1679235063
transform 1 0 8556 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_85
timestamp 1679235063
transform 1 0 8924 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_90
timestamp 1679235063
transform 1 0 9384 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_96
timestamp 1679235063
transform 1 0 9936 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_110
timestamp 1679235063
transform 1 0 11224 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_113
timestamp 1679235063
transform 1 0 11500 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_118
timestamp 1679235063
transform 1 0 11960 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_138
timestamp 1679235063
transform 1 0 13800 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_143
timestamp 1679235063
transform 1 0 14260 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_163
timestamp 1679235063
transform 1 0 16100 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_167
timestamp 1679235063
transform 1 0 16468 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_169
timestamp 1679235063
transform 1 0 16652 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_187
timestamp 1679235063
transform 1 0 18308 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_191
timestamp 1679235063
transform 1 0 18676 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_195
timestamp 1679235063
transform 1 0 19044 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_197
timestamp 1679235063
transform 1 0 19228 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_215 pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1679235063
transform 1 0 20884 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_223
timestamp 1679235063
transform 1 0 21620 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_225
timestamp 1679235063
transform 1 0 21804 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_243
timestamp 1679235063
transform 1 0 23460 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_251
timestamp 1679235063
transform 1 0 24196 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_253
timestamp 1679235063
transform 1 0 24380 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_264
timestamp 1679235063
transform 1 0 25392 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_1_5
timestamp 1679235063
transform 1 0 1564 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_1_11
timestamp 1679235063
transform 1 0 2116 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_19
timestamp 1679235063
transform 1 0 2852 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_1_33
timestamp 1679235063
transform 1 0 4140 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_1_37
timestamp 1679235063
transform 1 0 4508 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_1_40
timestamp 1679235063
transform 1 0 4784 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_1_46
timestamp 1679235063
transform 1 0 5336 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_1_54
timestamp 1679235063
transform 1 0 6072 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_1_59
timestamp 1679235063
transform 1 0 6532 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_1_66
timestamp 1679235063
transform 1 0 7176 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_74
timestamp 1679235063
transform 1 0 7912 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_82
timestamp 1679235063
transform 1 0 8648 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_96
timestamp 1679235063
transform 1 0 9936 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_1_110
timestamp 1679235063
transform 1 0 11224 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_1_113
timestamp 1679235063
transform 1 0 11500 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_1_119
timestamp 1679235063
transform 1 0 12052 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_139
timestamp 1679235063
transform 1 0 13892 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_1_159
timestamp 1679235063
transform 1 0 15732 0 -1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_1_167
timestamp 1679235063
transform 1 0 16468 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_1_169
timestamp 1679235063
transform 1 0 16652 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_1_187
timestamp 1679235063
transform 1 0 18308 0 -1 3264
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_1_207 pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1679235063
transform 1 0 20148 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_1_219
timestamp 1679235063
transform 1 0 21252 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_1_223
timestamp 1679235063
transform 1 0 21620 0 -1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_1_225
timestamp 1679235063
transform 1 0 21804 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_1_237 pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1679235063
transform 1 0 22908 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_1_243
timestamp 1679235063
transform 1 0 23460 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_1_264
timestamp 1679235063
transform 1 0 25392 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_2_3
timestamp 1679235063
transform 1 0 1380 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_2_10
timestamp 1679235063
transform 1 0 2024 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_2_16
timestamp 1679235063
transform 1 0 2576 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_2_25
timestamp 1679235063
transform 1 0 3404 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_2_29
timestamp 1679235063
transform 1 0 3772 0 1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_2_37
timestamp 1679235063
transform 1 0 4508 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_2_41
timestamp 1679235063
transform 1 0 4876 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_2_47
timestamp 1679235063
transform 1 0 5428 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_2_51
timestamp 1679235063
transform 1 0 5796 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_2_55
timestamp 1679235063
transform 1 0 6164 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_2_63
timestamp 1679235063
transform 1 0 6900 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_2_68
timestamp 1679235063
transform 1 0 7360 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_2_73
timestamp 1679235063
transform 1 0 7820 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_2_79
timestamp 1679235063
transform 1 0 8372 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_2_85
timestamp 1679235063
transform 1 0 8924 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_2_91
timestamp 1679235063
transform 1 0 9476 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_2_99
timestamp 1679235063
transform 1 0 10212 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_2_105
timestamp 1679235063
transform 1 0 10764 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_2_117
timestamp 1679235063
transform 1 0 11868 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_2_121
timestamp 1679235063
transform 1 0 12236 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_2_138
timestamp 1679235063
transform 1 0 13800 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_2_141
timestamp 1679235063
transform 1 0 14076 0 1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_2_149
timestamp 1679235063
transform 1 0 14812 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_2_167
timestamp 1679235063
transform 1 0 16468 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_2_187
timestamp 1679235063
transform 1 0 18308 0 1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_2_195
timestamp 1679235063
transform 1 0 19044 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_2_197
timestamp 1679235063
transform 1 0 19228 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_2_215
timestamp 1679235063
transform 1 0 20884 0 1 3264
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_2_235
timestamp 1679235063
transform 1 0 22724 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_2_247
timestamp 1679235063
transform 1 0 23828 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_2_251
timestamp 1679235063
transform 1 0 24196 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_2_253
timestamp 1679235063
transform 1 0 24380 0 1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_2_261
timestamp 1679235063
transform 1 0 25116 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_3_3
timestamp 1679235063
transform 1 0 1380 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_3_8
timestamp 1679235063
transform 1 0 1840 0 -1 4352
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_3_12
timestamp 1679235063
transform 1 0 2208 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_24
timestamp 1679235063
transform 1 0 3312 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_36
timestamp 1679235063
transform 1 0 4416 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_3_48
timestamp 1679235063
transform 1 0 5520 0 -1 4352
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_3_59
timestamp 1679235063
transform 1 0 6532 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_71
timestamp 1679235063
transform 1 0 7636 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_3_83
timestamp 1679235063
transform 1 0 8740 0 -1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_3_95
timestamp 1679235063
transform 1 0 9844 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_3_98
timestamp 1679235063
transform 1 0 10120 0 -1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_3_106
timestamp 1679235063
transform 1 0 10856 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_3_113
timestamp 1679235063
transform 1 0 11500 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_3_125
timestamp 1679235063
transform 1 0 12604 0 -1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_3_133
timestamp 1679235063
transform 1 0 13340 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_3_151
timestamp 1679235063
transform 1 0 14996 0 -1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_3_159
timestamp 1679235063
transform 1 0 15732 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_3_166
timestamp 1679235063
transform 1 0 16376 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_3_169
timestamp 1679235063
transform 1 0 16652 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_3_187
timestamp 1679235063
transform 1 0 18308 0 -1 4352
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_3_207
timestamp 1679235063
transform 1 0 20148 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_3_219
timestamp 1679235063
transform 1 0 21252 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_3_223
timestamp 1679235063
transform 1 0 21620 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_3_225
timestamp 1679235063
transform 1 0 21804 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_3_243
timestamp 1679235063
transform 1 0 23460 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_3_263
timestamp 1679235063
transform 1 0 25300 0 -1 4352
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_4_3
timestamp 1679235063
transform 1 0 1380 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_15
timestamp 1679235063
transform 1 0 2484 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_4_27
timestamp 1679235063
transform 1 0 3588 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_4_29
timestamp 1679235063
transform 1 0 3772 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_41
timestamp 1679235063
transform 1 0 4876 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_53
timestamp 1679235063
transform 1 0 5980 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_65
timestamp 1679235063
transform 1 0 7084 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_4_77
timestamp 1679235063
transform 1 0 8188 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_83
timestamp 1679235063
transform 1 0 8740 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_4_85
timestamp 1679235063
transform 1 0 8924 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_97
timestamp 1679235063
transform 1 0 10028 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_109
timestamp 1679235063
transform 1 0 11132 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_121
timestamp 1679235063
transform 1 0 12236 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_4_133
timestamp 1679235063
transform 1 0 13340 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_139
timestamp 1679235063
transform 1 0 13892 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_4_141
timestamp 1679235063
transform 1 0 14076 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_153
timestamp 1679235063
transform 1 0 15180 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_165
timestamp 1679235063
transform 1 0 16284 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_4_177
timestamp 1679235063
transform 1 0 17388 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_4_194
timestamp 1679235063
transform 1 0 18952 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_4_197
timestamp 1679235063
transform 1 0 19228 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_4_215
timestamp 1679235063
transform 1 0 20884 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_4_235
timestamp 1679235063
transform 1 0 22724 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_4_239
timestamp 1679235063
transform 1 0 23092 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_4_250
timestamp 1679235063
transform 1 0 24104 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_4_253
timestamp 1679235063
transform 1 0 24380 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_4_259
timestamp 1679235063
transform 1 0 24932 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_265
timestamp 1679235063
transform 1 0 25484 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_5_3
timestamp 1679235063
transform 1 0 1380 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_15
timestamp 1679235063
transform 1 0 2484 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_27
timestamp 1679235063
transform 1 0 3588 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_39
timestamp 1679235063
transform 1 0 4692 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_5_51
timestamp 1679235063
transform 1 0 5796 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_5_55
timestamp 1679235063
transform 1 0 6164 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_5_57
timestamp 1679235063
transform 1 0 6348 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_69
timestamp 1679235063
transform 1 0 7452 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_81
timestamp 1679235063
transform 1 0 8556 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_93
timestamp 1679235063
transform 1 0 9660 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_5_105
timestamp 1679235063
transform 1 0 10764 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_111
timestamp 1679235063
transform 1 0 11316 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_5_113
timestamp 1679235063
transform 1 0 11500 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_125
timestamp 1679235063
transform 1 0 12604 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_137
timestamp 1679235063
transform 1 0 13708 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_149
timestamp 1679235063
transform 1 0 14812 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_5_161
timestamp 1679235063
transform 1 0 15916 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_167
timestamp 1679235063
transform 1 0 16468 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_5_169
timestamp 1679235063
transform 1 0 16652 0 -1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_5_177
timestamp 1679235063
transform 1 0 17388 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_5_195
timestamp 1679235063
transform 1 0 19044 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_5_215
timestamp 1679235063
transform 1 0 20884 0 -1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_5_223
timestamp 1679235063
transform 1 0 21620 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_5_225
timestamp 1679235063
transform 1 0 21804 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_5_243
timestamp 1679235063
transform 1 0 23460 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_5_247
timestamp 1679235063
transform 1 0 23828 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_5_264
timestamp 1679235063
transform 1 0 25392 0 -1 5440
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_6_3
timestamp 1679235063
transform 1 0 1380 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_15
timestamp 1679235063
transform 1 0 2484 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_6_27
timestamp 1679235063
transform 1 0 3588 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_6_29
timestamp 1679235063
transform 1 0 3772 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_41
timestamp 1679235063
transform 1 0 4876 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_53
timestamp 1679235063
transform 1 0 5980 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_65
timestamp 1679235063
transform 1 0 7084 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_6_77
timestamp 1679235063
transform 1 0 8188 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_83
timestamp 1679235063
transform 1 0 8740 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_6_85
timestamp 1679235063
transform 1 0 8924 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_97
timestamp 1679235063
transform 1 0 10028 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_109
timestamp 1679235063
transform 1 0 11132 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_121
timestamp 1679235063
transform 1 0 12236 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_6_133
timestamp 1679235063
transform 1 0 13340 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_139
timestamp 1679235063
transform 1 0 13892 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_6_141
timestamp 1679235063
transform 1 0 14076 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_153
timestamp 1679235063
transform 1 0 15180 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_165
timestamp 1679235063
transform 1 0 16284 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_177
timestamp 1679235063
transform 1 0 17388 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_6_189
timestamp 1679235063
transform 1 0 18492 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_195
timestamp 1679235063
transform 1 0 19044 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_6_197
timestamp 1679235063
transform 1 0 19228 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_6_209
timestamp 1679235063
transform 1 0 20332 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_6_227
timestamp 1679235063
transform 1 0 21988 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_6_247
timestamp 1679235063
transform 1 0 23828 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_6_251
timestamp 1679235063
transform 1 0 24196 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_6_253
timestamp 1679235063
transform 1 0 24380 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_6_259
timestamp 1679235063
transform 1 0 24932 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_265
timestamp 1679235063
transform 1 0 25484 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_7_3
timestamp 1679235063
transform 1 0 1380 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_15
timestamp 1679235063
transform 1 0 2484 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_27
timestamp 1679235063
transform 1 0 3588 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_39
timestamp 1679235063
transform 1 0 4692 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_7_51
timestamp 1679235063
transform 1 0 5796 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_7_55
timestamp 1679235063
transform 1 0 6164 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_7_57
timestamp 1679235063
transform 1 0 6348 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_69
timestamp 1679235063
transform 1 0 7452 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_81
timestamp 1679235063
transform 1 0 8556 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_93
timestamp 1679235063
transform 1 0 9660 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_7_105
timestamp 1679235063
transform 1 0 10764 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_111
timestamp 1679235063
transform 1 0 11316 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_7_113
timestamp 1679235063
transform 1 0 11500 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_125
timestamp 1679235063
transform 1 0 12604 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_137
timestamp 1679235063
transform 1 0 13708 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_149
timestamp 1679235063
transform 1 0 14812 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_7_161
timestamp 1679235063
transform 1 0 15916 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_167
timestamp 1679235063
transform 1 0 16468 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_7_169
timestamp 1679235063
transform 1 0 16652 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_7_181
timestamp 1679235063
transform 1 0 17756 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_7_184
timestamp 1679235063
transform 1 0 18032 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_7_202
timestamp 1679235063
transform 1 0 19688 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_7_222
timestamp 1679235063
transform 1 0 21528 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_7_225
timestamp 1679235063
transform 1 0 21804 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_7_243
timestamp 1679235063
transform 1 0 23460 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_7_247
timestamp 1679235063
transform 1 0 23828 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_7_264
timestamp 1679235063
transform 1 0 25392 0 -1 6528
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_8_3
timestamp 1679235063
transform 1 0 1380 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_15
timestamp 1679235063
transform 1 0 2484 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_8_27
timestamp 1679235063
transform 1 0 3588 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_8_29
timestamp 1679235063
transform 1 0 3772 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_41
timestamp 1679235063
transform 1 0 4876 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_53
timestamp 1679235063
transform 1 0 5980 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_65
timestamp 1679235063
transform 1 0 7084 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_8_77
timestamp 1679235063
transform 1 0 8188 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_83
timestamp 1679235063
transform 1 0 8740 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_8_85
timestamp 1679235063
transform 1 0 8924 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_97
timestamp 1679235063
transform 1 0 10028 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_109
timestamp 1679235063
transform 1 0 11132 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_121
timestamp 1679235063
transform 1 0 12236 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_8_133
timestamp 1679235063
transform 1 0 13340 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_139
timestamp 1679235063
transform 1 0 13892 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_8_141
timestamp 1679235063
transform 1 0 14076 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_153
timestamp 1679235063
transform 1 0 15180 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_165
timestamp 1679235063
transform 1 0 16284 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_177
timestamp 1679235063
transform 1 0 17388 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_8_189
timestamp 1679235063
transform 1 0 18492 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_195
timestamp 1679235063
transform 1 0 19044 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_8_197
timestamp 1679235063
transform 1 0 19228 0 1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_8_205
timestamp 1679235063
transform 1 0 19964 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_8_209
timestamp 1679235063
transform 1 0 20332 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_8_213
timestamp 1679235063
transform 1 0 20700 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_8_230
timestamp 1679235063
transform 1 0 22264 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_8_250
timestamp 1679235063
transform 1 0 24104 0 1 6528
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_8_253
timestamp 1679235063
transform 1 0 24380 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_8_265
timestamp 1679235063
transform 1 0 25484 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_9_3
timestamp 1679235063
transform 1 0 1380 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_15
timestamp 1679235063
transform 1 0 2484 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_27
timestamp 1679235063
transform 1 0 3588 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_39
timestamp 1679235063
transform 1 0 4692 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_9_51
timestamp 1679235063
transform 1 0 5796 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_9_55
timestamp 1679235063
transform 1 0 6164 0 -1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_9_57
timestamp 1679235063
transform 1 0 6348 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_69
timestamp 1679235063
transform 1 0 7452 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_81
timestamp 1679235063
transform 1 0 8556 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_93
timestamp 1679235063
transform 1 0 9660 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_9_105
timestamp 1679235063
transform 1 0 10764 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_9_111
timestamp 1679235063
transform 1 0 11316 0 -1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_9_113
timestamp 1679235063
transform 1 0 11500 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_125
timestamp 1679235063
transform 1 0 12604 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_137
timestamp 1679235063
transform 1 0 13708 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_149
timestamp 1679235063
transform 1 0 14812 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_9_161
timestamp 1679235063
transform 1 0 15916 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_9_167
timestamp 1679235063
transform 1 0 16468 0 -1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_9_169
timestamp 1679235063
transform 1 0 16652 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_9_181
timestamp 1679235063
transform 1 0 17756 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_9_187
timestamp 1679235063
transform 1 0 18308 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_9_192
timestamp 1679235063
transform 1 0 18768 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_9_202
timestamp 1679235063
transform 1 0 19688 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_9_222
timestamp 1679235063
transform 1 0 21528 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_9_225
timestamp 1679235063
transform 1 0 21804 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_9_244
timestamp 1679235063
transform 1 0 23552 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_9_264
timestamp 1679235063
transform 1 0 25392 0 -1 7616
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_10_3
timestamp 1679235063
transform 1 0 1380 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_15
timestamp 1679235063
transform 1 0 2484 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_10_27
timestamp 1679235063
transform 1 0 3588 0 1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_10_29
timestamp 1679235063
transform 1 0 3772 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_41
timestamp 1679235063
transform 1 0 4876 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_53
timestamp 1679235063
transform 1 0 5980 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_65
timestamp 1679235063
transform 1 0 7084 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_10_77
timestamp 1679235063
transform 1 0 8188 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_10_83
timestamp 1679235063
transform 1 0 8740 0 1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_10_85
timestamp 1679235063
transform 1 0 8924 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_97
timestamp 1679235063
transform 1 0 10028 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_109
timestamp 1679235063
transform 1 0 11132 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_121
timestamp 1679235063
transform 1 0 12236 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_10_133
timestamp 1679235063
transform 1 0 13340 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_10_139
timestamp 1679235063
transform 1 0 13892 0 1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_10_141
timestamp 1679235063
transform 1 0 14076 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_153
timestamp 1679235063
transform 1 0 15180 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_165
timestamp 1679235063
transform 1 0 16284 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_177
timestamp 1679235063
transform 1 0 17388 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_10_189
timestamp 1679235063
transform 1 0 18492 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_10_195
timestamp 1679235063
transform 1 0 19044 0 1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_10_197
timestamp 1679235063
transform 1 0 19228 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_10_209
timestamp 1679235063
transform 1 0 20332 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_10_213
timestamp 1679235063
transform 1 0 20700 0 1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_10_224
timestamp 1679235063
transform 1 0 21712 0 1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_10_232
timestamp 1679235063
transform 1 0 22448 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_10_250
timestamp 1679235063
transform 1 0 24104 0 1 7616
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_10_253
timestamp 1679235063
transform 1 0 24380 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_10_265
timestamp 1679235063
transform 1 0 25484 0 1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_11_3
timestamp 1679235063
transform 1 0 1380 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_15
timestamp 1679235063
transform 1 0 2484 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_11_27
timestamp 1679235063
transform 1 0 3588 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_11_54
timestamp 1679235063
transform 1 0 6072 0 -1 8704
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_11_59
timestamp 1679235063
transform 1 0 6532 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_71
timestamp 1679235063
transform 1 0 7636 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_83
timestamp 1679235063
transform 1 0 8740 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_95
timestamp 1679235063
transform 1 0 9844 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_11_107
timestamp 1679235063
transform 1 0 10948 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_11_111
timestamp 1679235063
transform 1 0 11316 0 -1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_11_113
timestamp 1679235063
transform 1 0 11500 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_125
timestamp 1679235063
transform 1 0 12604 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_137
timestamp 1679235063
transform 1 0 13708 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_149
timestamp 1679235063
transform 1 0 14812 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_11_161
timestamp 1679235063
transform 1 0 15916 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_11_167
timestamp 1679235063
transform 1 0 16468 0 -1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_11_169
timestamp 1679235063
transform 1 0 16652 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_11_181
timestamp 1679235063
transform 1 0 17756 0 -1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_11_189
timestamp 1679235063
transform 1 0 18492 0 -1 8704
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_11_196
timestamp 1679235063
transform 1 0 19136 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_11_208
timestamp 1679235063
transform 1 0 20240 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_11_212
timestamp 1679235063
transform 1 0 20608 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_11_217
timestamp 1679235063
transform 1 0 21068 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_11_223
timestamp 1679235063
transform 1 0 21620 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_11_225
timestamp 1679235063
transform 1 0 21804 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_11_244
timestamp 1679235063
transform 1 0 23552 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_11_264
timestamp 1679235063
transform 1 0 25392 0 -1 8704
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_12_3
timestamp 1679235063
transform 1 0 1380 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_15
timestamp 1679235063
transform 1 0 2484 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_12_27
timestamp 1679235063
transform 1 0 3588 0 1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_12_29
timestamp 1679235063
transform 1 0 3772 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_41
timestamp 1679235063
transform 1 0 4876 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_53
timestamp 1679235063
transform 1 0 5980 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_12_74
timestamp 1679235063
transform 1 0 7912 0 1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_12_82
timestamp 1679235063
transform 1 0 8648 0 1 8704
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_12_85
timestamp 1679235063
transform 1 0 8924 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_97
timestamp 1679235063
transform 1 0 10028 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_109
timestamp 1679235063
transform 1 0 11132 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_121
timestamp 1679235063
transform 1 0 12236 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_12_133
timestamp 1679235063
transform 1 0 13340 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_12_139
timestamp 1679235063
transform 1 0 13892 0 1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_12_141
timestamp 1679235063
transform 1 0 14076 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_153
timestamp 1679235063
transform 1 0 15180 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_165
timestamp 1679235063
transform 1 0 16284 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_177
timestamp 1679235063
transform 1 0 17388 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_12_189
timestamp 1679235063
transform 1 0 18492 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_12_195
timestamp 1679235063
transform 1 0 19044 0 1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_12_197
timestamp 1679235063
transform 1 0 19228 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_209
timestamp 1679235063
transform 1 0 20332 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_221
timestamp 1679235063
transform 1 0 21436 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_233
timestamp 1679235063
transform 1 0 22540 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_12_245
timestamp 1679235063
transform 1 0 23644 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_12_250
timestamp 1679235063
transform 1 0 24104 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_12_253
timestamp 1679235063
transform 1 0 24380 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_12_259
timestamp 1679235063
transform 1 0 24932 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_12_265
timestamp 1679235063
transform 1 0 25484 0 1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_13_3
timestamp 1679235063
transform 1 0 1380 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_15
timestamp 1679235063
transform 1 0 2484 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_27
timestamp 1679235063
transform 1 0 3588 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_39
timestamp 1679235063
transform 1 0 4692 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_13_51
timestamp 1679235063
transform 1 0 5796 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_13_55
timestamp 1679235063
transform 1 0 6164 0 -1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_13_57
timestamp 1679235063
transform 1 0 6348 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_13_69
timestamp 1679235063
transform 1 0 7452 0 -1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_13_73
timestamp 1679235063
transform 1 0 7820 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_85
timestamp 1679235063
transform 1 0 8924 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_97
timestamp 1679235063
transform 1 0 10028 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_13_109
timestamp 1679235063
transform 1 0 11132 0 -1 9792
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_13_113
timestamp 1679235063
transform 1 0 11500 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_125
timestamp 1679235063
transform 1 0 12604 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_137
timestamp 1679235063
transform 1 0 13708 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_149
timestamp 1679235063
transform 1 0 14812 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_13_161
timestamp 1679235063
transform 1 0 15916 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_13_167
timestamp 1679235063
transform 1 0 16468 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_13_169
timestamp 1679235063
transform 1 0 16652 0 -1 9792
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_13_175
timestamp 1679235063
transform 1 0 17204 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_13_187
timestamp 1679235063
transform 1 0 18308 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_13_191
timestamp 1679235063
transform 1 0 18676 0 -1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_13_196
timestamp 1679235063
transform 1 0 19136 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_208
timestamp 1679235063
transform 1 0 20240 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_13_220
timestamp 1679235063
transform 1 0 21344 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_13_225
timestamp 1679235063
transform 1 0 21804 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_13_231
timestamp 1679235063
transform 1 0 22356 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_13_235
timestamp 1679235063
transform 1 0 22724 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_13_239
timestamp 1679235063
transform 1 0 23092 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_13_243
timestamp 1679235063
transform 1 0 23460 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_13_247
timestamp 1679235063
transform 1 0 23828 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_13_264
timestamp 1679235063
transform 1 0 25392 0 -1 9792
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_14_3
timestamp 1679235063
transform 1 0 1380 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_15
timestamp 1679235063
transform 1 0 2484 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_14_27
timestamp 1679235063
transform 1 0 3588 0 1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_14_29
timestamp 1679235063
transform 1 0 3772 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_41
timestamp 1679235063
transform 1 0 4876 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_53
timestamp 1679235063
transform 1 0 5980 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_65
timestamp 1679235063
transform 1 0 7084 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_14_77
timestamp 1679235063
transform 1 0 8188 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_14_83
timestamp 1679235063
transform 1 0 8740 0 1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_14_85
timestamp 1679235063
transform 1 0 8924 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_97
timestamp 1679235063
transform 1 0 10028 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_109
timestamp 1679235063
transform 1 0 11132 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_121
timestamp 1679235063
transform 1 0 12236 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_14_133
timestamp 1679235063
transform 1 0 13340 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_14_139
timestamp 1679235063
transform 1 0 13892 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_14_141
timestamp 1679235063
transform 1 0 14076 0 1 9792
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_14_149
timestamp 1679235063
transform 1 0 14812 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_14_161
timestamp 1679235063
transform 1 0 15916 0 1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_14_169
timestamp 1679235063
transform 1 0 16652 0 1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_14_174
timestamp 1679235063
transform 1 0 17112 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_14_186
timestamp 1679235063
transform 1 0 18216 0 1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_14_194
timestamp 1679235063
transform 1 0 18952 0 1 9792
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_14_197
timestamp 1679235063
transform 1 0 19228 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_209
timestamp 1679235063
transform 1 0 20332 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_14_221
timestamp 1679235063
transform 1 0 21436 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_14_230
timestamp 1679235063
transform 1 0 22264 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_14_250
timestamp 1679235063
transform 1 0 24104 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_14_253
timestamp 1679235063
transform 1 0 24380 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_14_259
timestamp 1679235063
transform 1 0 24932 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_14_265
timestamp 1679235063
transform 1 0 25484 0 1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_15_3
timestamp 1679235063
transform 1 0 1380 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_15
timestamp 1679235063
transform 1 0 2484 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_27
timestamp 1679235063
transform 1 0 3588 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_39
timestamp 1679235063
transform 1 0 4692 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_15_51
timestamp 1679235063
transform 1 0 5796 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_15_55
timestamp 1679235063
transform 1 0 6164 0 -1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_15_57
timestamp 1679235063
transform 1 0 6348 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_69
timestamp 1679235063
transform 1 0 7452 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_81
timestamp 1679235063
transform 1 0 8556 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_93
timestamp 1679235063
transform 1 0 9660 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_15_105
timestamp 1679235063
transform 1 0 10764 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_15_111
timestamp 1679235063
transform 1 0 11316 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_15_113
timestamp 1679235063
transform 1 0 11500 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_15_121
timestamp 1679235063
transform 1 0 12236 0 -1 10880
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_15_125
timestamp 1679235063
transform 1 0 12604 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_137
timestamp 1679235063
transform 1 0 13708 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_149
timestamp 1679235063
transform 1 0 14812 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_15_161
timestamp 1679235063
transform 1 0 15916 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_15_167
timestamp 1679235063
transform 1 0 16468 0 -1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_15_169
timestamp 1679235063
transform 1 0 16652 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_15_181
timestamp 1679235063
transform 1 0 17756 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_15_190
timestamp 1679235063
transform 1 0 18584 0 -1 10880
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_15_205
timestamp 1679235063
transform 1 0 19964 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_15_217
timestamp 1679235063
transform 1 0 21068 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_15_221
timestamp 1679235063
transform 1 0 21436 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_15_225
timestamp 1679235063
transform 1 0 21804 0 -1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_15_233
timestamp 1679235063
transform 1 0 22540 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_15_238
timestamp 1679235063
transform 1 0 23000 0 -1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_15_246
timestamp 1679235063
transform 1 0 23736 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_15_264
timestamp 1679235063
transform 1 0 25392 0 -1 10880
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_16_3
timestamp 1679235063
transform 1 0 1380 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_15
timestamp 1679235063
transform 1 0 2484 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_16_27
timestamp 1679235063
transform 1 0 3588 0 1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_16_29
timestamp 1679235063
transform 1 0 3772 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_41
timestamp 1679235063
transform 1 0 4876 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_53
timestamp 1679235063
transform 1 0 5980 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_65
timestamp 1679235063
transform 1 0 7084 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_16_77
timestamp 1679235063
transform 1 0 8188 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_16_83
timestamp 1679235063
transform 1 0 8740 0 1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_16_85
timestamp 1679235063
transform 1 0 8924 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_97
timestamp 1679235063
transform 1 0 10028 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_109
timestamp 1679235063
transform 1 0 11132 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_121
timestamp 1679235063
transform 1 0 12236 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_16_133
timestamp 1679235063
transform 1 0 13340 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_16_139
timestamp 1679235063
transform 1 0 13892 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_16_141
timestamp 1679235063
transform 1 0 14076 0 1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_16_157
timestamp 1679235063
transform 1 0 15548 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_16_165
timestamp 1679235063
transform 1 0 16284 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_16_172
timestamp 1679235063
transform 1 0 16928 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_16_176
timestamp 1679235063
transform 1 0 17296 0 1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_16_184
timestamp 1679235063
transform 1 0 18032 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_16_191
timestamp 1679235063
transform 1 0 18676 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_16_195
timestamp 1679235063
transform 1 0 19044 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_16_197
timestamp 1679235063
transform 1 0 19228 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_16_203
timestamp 1679235063
transform 1 0 19780 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_16_210
timestamp 1679235063
transform 1 0 20424 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_16_214
timestamp 1679235063
transform 1 0 20792 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_16_219
timestamp 1679235063
transform 1 0 21252 0 1 10880
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_16_227
timestamp 1679235063
transform 1 0 21988 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_16_239
timestamp 1679235063
transform 1 0 23092 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_16_243
timestamp 1679235063
transform 1 0 23460 0 1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_16_251
timestamp 1679235063
transform 1 0 24196 0 1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_16_253
timestamp 1679235063
transform 1 0 24380 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_16_265
timestamp 1679235063
transform 1 0 25484 0 1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_17_3
timestamp 1679235063
transform 1 0 1380 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_15
timestamp 1679235063
transform 1 0 2484 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_27
timestamp 1679235063
transform 1 0 3588 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_39
timestamp 1679235063
transform 1 0 4692 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_17_51
timestamp 1679235063
transform 1 0 5796 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_17_55
timestamp 1679235063
transform 1 0 6164 0 -1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_17_57
timestamp 1679235063
transform 1 0 6348 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_69
timestamp 1679235063
transform 1 0 7452 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_81
timestamp 1679235063
transform 1 0 8556 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_17_93
timestamp 1679235063
transform 1 0 9660 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_17_107
timestamp 1679235063
transform 1 0 10948 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_17_111
timestamp 1679235063
transform 1 0 11316 0 -1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_17_115
timestamp 1679235063
transform 1 0 11684 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_17_127
timestamp 1679235063
transform 1 0 12788 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_17_149
timestamp 1679235063
transform 1 0 14812 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_17_162
timestamp 1679235063
transform 1 0 16008 0 -1 11968
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_17_169
timestamp 1679235063
transform 1 0 16652 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_17_181
timestamp 1679235063
transform 1 0 17756 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_17_203
timestamp 1679235063
transform 1 0 19780 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_17_215
timestamp 1679235063
transform 1 0 20884 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_17_219
timestamp 1679235063
transform 1 0 21252 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_17_223
timestamp 1679235063
transform 1 0 21620 0 -1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_17_225
timestamp 1679235063
transform 1 0 21804 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_17_237
timestamp 1679235063
transform 1 0 22908 0 -1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_17_245
timestamp 1679235063
transform 1 0 23644 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_17_264
timestamp 1679235063
transform 1 0 25392 0 -1 11968
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_18_3
timestamp 1679235063
transform 1 0 1380 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_15
timestamp 1679235063
transform 1 0 2484 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_18_27
timestamp 1679235063
transform 1 0 3588 0 1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_18_29
timestamp 1679235063
transform 1 0 3772 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_41
timestamp 1679235063
transform 1 0 4876 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_53
timestamp 1679235063
transform 1 0 5980 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_65
timestamp 1679235063
transform 1 0 7084 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_18_77
timestamp 1679235063
transform 1 0 8188 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_18_83
timestamp 1679235063
transform 1 0 8740 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_18_85
timestamp 1679235063
transform 1 0 8924 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_18_91
timestamp 1679235063
transform 1 0 9476 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_18_112
timestamp 1679235063
transform 1 0 11408 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_18_136
timestamp 1679235063
transform 1 0 13616 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_18_141
timestamp 1679235063
transform 1 0 14076 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_18_147
timestamp 1679235063
transform 1 0 14628 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_18_151
timestamp 1679235063
transform 1 0 14996 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_18_162
timestamp 1679235063
transform 1 0 16008 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_18_175
timestamp 1679235063
transform 1 0 17204 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_18_182
timestamp 1679235063
transform 1 0 17848 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_18_194
timestamp 1679235063
transform 1 0 18952 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_18_197
timestamp 1679235063
transform 1 0 19228 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_18_221
timestamp 1679235063
transform 1 0 21436 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_18_228
timestamp 1679235063
transform 1 0 22080 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_18_232
timestamp 1679235063
transform 1 0 22448 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_18_237
timestamp 1679235063
transform 1 0 22908 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_18_244
timestamp 1679235063
transform 1 0 23552 0 1 11968
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_18_253
timestamp 1679235063
transform 1 0 24380 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_18_265
timestamp 1679235063
transform 1 0 25484 0 1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_19_3
timestamp 1679235063
transform 1 0 1380 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_15
timestamp 1679235063
transform 1 0 2484 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_27
timestamp 1679235063
transform 1 0 3588 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_39
timestamp 1679235063
transform 1 0 4692 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_19_51
timestamp 1679235063
transform 1 0 5796 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_19_55
timestamp 1679235063
transform 1 0 6164 0 -1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_19_57
timestamp 1679235063
transform 1 0 6348 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_69
timestamp 1679235063
transform 1 0 7452 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_19_81
timestamp 1679235063
transform 1 0 8556 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_19_104
timestamp 1679235063
transform 1 0 10672 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_19_108
timestamp 1679235063
transform 1 0 11040 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_19_113
timestamp 1679235063
transform 1 0 11500 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_19_123
timestamp 1679235063
transform 1 0 12420 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_19_131
timestamp 1679235063
transform 1 0 13156 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_19_142
timestamp 1679235063
transform 1 0 14168 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_19_166
timestamp 1679235063
transform 1 0 16376 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_19_169
timestamp 1679235063
transform 1 0 16652 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_19_175
timestamp 1679235063
transform 1 0 17204 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_19_179
timestamp 1679235063
transform 1 0 17572 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_19_202
timestamp 1679235063
transform 1 0 19688 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_19_208
timestamp 1679235063
transform 1 0 20240 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_19_212
timestamp 1679235063
transform 1 0 20608 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_19_222
timestamp 1679235063
transform 1 0 21528 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_19_225
timestamp 1679235063
transform 1 0 21804 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_19_231
timestamp 1679235063
transform 1 0 22356 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_19_238
timestamp 1679235063
transform 1 0 23000 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_19_242
timestamp 1679235063
transform 1 0 23368 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_19_264
timestamp 1679235063
transform 1 0 25392 0 -1 13056
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_20_3
timestamp 1679235063
transform 1 0 1380 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_15
timestamp 1679235063
transform 1 0 2484 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_20_27
timestamp 1679235063
transform 1 0 3588 0 1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_20_29
timestamp 1679235063
transform 1 0 3772 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_41
timestamp 1679235063
transform 1 0 4876 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_53
timestamp 1679235063
transform 1 0 5980 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_65
timestamp 1679235063
transform 1 0 7084 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_20_77
timestamp 1679235063
transform 1 0 8188 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_20_83
timestamp 1679235063
transform 1 0 8740 0 1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_20_85
timestamp 1679235063
transform 1 0 8924 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_20_97
timestamp 1679235063
transform 1 0 10028 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_20_109
timestamp 1679235063
transform 1 0 11132 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_20_113
timestamp 1679235063
transform 1 0 11500 0 1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_20_122
timestamp 1679235063
transform 1 0 12328 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_20_138
timestamp 1679235063
transform 1 0 13800 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_20_141
timestamp 1679235063
transform 1 0 14076 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_20_151
timestamp 1679235063
transform 1 0 14996 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_20_159
timestamp 1679235063
transform 1 0 15732 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_20_163
timestamp 1679235063
transform 1 0 16100 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_20_176
timestamp 1679235063
transform 1 0 17296 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_20_189
timestamp 1679235063
transform 1 0 18492 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_20_193
timestamp 1679235063
transform 1 0 18860 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_20_197
timestamp 1679235063
transform 1 0 19228 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_20_203
timestamp 1679235063
transform 1 0 19780 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_20_211
timestamp 1679235063
transform 1 0 20516 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_20_215
timestamp 1679235063
transform 1 0 20884 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_20_225
timestamp 1679235063
transform 1 0 21804 0 1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_20_233
timestamp 1679235063
transform 1 0 22540 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_20_250
timestamp 1679235063
transform 1 0 24104 0 1 13056
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_20_253
timestamp 1679235063
transform 1 0 24380 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_20_265
timestamp 1679235063
transform 1 0 25484 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_21_3
timestamp 1679235063
transform 1 0 1380 0 -1 14144
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_21_21
timestamp 1679235063
transform 1 0 3036 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_33
timestamp 1679235063
transform 1 0 4140 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_21_45
timestamp 1679235063
transform 1 0 5244 0 -1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_21_53
timestamp 1679235063
transform 1 0 5980 0 -1 14144
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_21_57
timestamp 1679235063
transform 1 0 6348 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_21_69
timestamp 1679235063
transform 1 0 7452 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_21_75
timestamp 1679235063
transform 1 0 8004 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_21_96
timestamp 1679235063
transform 1 0 9936 0 -1 14144
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_21_100
timestamp 1679235063
transform 1 0 10304 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_21_113
timestamp 1679235063
transform 1 0 11500 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_21_121
timestamp 1679235063
transform 1 0 12236 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_21_132
timestamp 1679235063
transform 1 0 13248 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_21_136
timestamp 1679235063
transform 1 0 13616 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_21_140
timestamp 1679235063
transform 1 0 13984 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_21_147
timestamp 1679235063
transform 1 0 14628 0 -1 14144
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_21_151
timestamp 1679235063
transform 1 0 14996 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_21_166
timestamp 1679235063
transform 1 0 16376 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_21_169
timestamp 1679235063
transform 1 0 16652 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_21_179
timestamp 1679235063
transform 1 0 17572 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_21_185
timestamp 1679235063
transform 1 0 18124 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_21_197
timestamp 1679235063
transform 1 0 19228 0 -1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_21_205
timestamp 1679235063
transform 1 0 19964 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_21_215
timestamp 1679235063
transform 1 0 20884 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_21_222
timestamp 1679235063
transform 1 0 21528 0 -1 14144
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_21_225
timestamp 1679235063
transform 1 0 21804 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_21_237
timestamp 1679235063
transform 1 0 22908 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_21_241
timestamp 1679235063
transform 1 0 23276 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_21_247
timestamp 1679235063
transform 1 0 23828 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_21_264
timestamp 1679235063
transform 1 0 25392 0 -1 14144
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_22_3
timestamp 1679235063
transform 1 0 1380 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_15
timestamp 1679235063
transform 1 0 2484 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_22_27
timestamp 1679235063
transform 1 0 3588 0 1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_22_29
timestamp 1679235063
transform 1 0 3772 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_41
timestamp 1679235063
transform 1 0 4876 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_53
timestamp 1679235063
transform 1 0 5980 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_22_65
timestamp 1679235063
transform 1 0 7084 0 1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_22_73
timestamp 1679235063
transform 1 0 7820 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_22_82
timestamp 1679235063
transform 1 0 8648 0 1 14144
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_22_85
timestamp 1679235063
transform 1 0 8924 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_22_118
timestamp 1679235063
transform 1 0 11960 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_22_124
timestamp 1679235063
transform 1 0 12512 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_22_127
timestamp 1679235063
transform 1 0 12788 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_22_138
timestamp 1679235063
transform 1 0 13800 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_22_141
timestamp 1679235063
transform 1 0 14076 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_22_147
timestamp 1679235063
transform 1 0 14628 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_22_151
timestamp 1679235063
transform 1 0 14996 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_22_174
timestamp 1679235063
transform 1 0 17112 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_22_182
timestamp 1679235063
transform 1 0 17848 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_22_186
timestamp 1679235063
transform 1 0 18216 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_22_191
timestamp 1679235063
transform 1 0 18676 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_22_195
timestamp 1679235063
transform 1 0 19044 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_22_197
timestamp 1679235063
transform 1 0 19228 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_22_202
timestamp 1679235063
transform 1 0 19688 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_22_210
timestamp 1679235063
transform 1 0 20424 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_22_236
timestamp 1679235063
transform 1 0 22816 0 1 14144
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_22_240
timestamp 1679235063
transform 1 0 23184 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_253
timestamp 1679235063
transform 1 0 24380 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_22_265
timestamp 1679235063
transform 1 0 25484 0 1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_23_3
timestamp 1679235063
transform 1 0 1380 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_15
timestamp 1679235063
transform 1 0 2484 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_27
timestamp 1679235063
transform 1 0 3588 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_39
timestamp 1679235063
transform 1 0 4692 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_23_51
timestamp 1679235063
transform 1 0 5796 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_23_55
timestamp 1679235063
transform 1 0 6164 0 -1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_23_57
timestamp 1679235063
transform 1 0 6348 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_23_69
timestamp 1679235063
transform 1 0 7452 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_23_74
timestamp 1679235063
transform 1 0 7912 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_23_99
timestamp 1679235063
transform 1 0 10212 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_23_103
timestamp 1679235063
transform 1 0 10580 0 -1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_23_111
timestamp 1679235063
transform 1 0 11316 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_23_113
timestamp 1679235063
transform 1 0 11500 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_23_125
timestamp 1679235063
transform 1 0 12604 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_23_138
timestamp 1679235063
transform 1 0 13800 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_23_151
timestamp 1679235063
transform 1 0 14996 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_23_155
timestamp 1679235063
transform 1 0 15364 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_23_166
timestamp 1679235063
transform 1 0 16376 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_23_169
timestamp 1679235063
transform 1 0 16652 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_23_175
timestamp 1679235063
transform 1 0 17204 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_23_188
timestamp 1679235063
transform 1 0 18400 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_23_212
timestamp 1679235063
transform 1 0 20608 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_23_219
timestamp 1679235063
transform 1 0 21252 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_23_223
timestamp 1679235063
transform 1 0 21620 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_23_225
timestamp 1679235063
transform 1 0 21804 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_23_231
timestamp 1679235063
transform 1 0 22356 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_23_236
timestamp 1679235063
transform 1 0 22816 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_23_244
timestamp 1679235063
transform 1 0 23552 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_23_264
timestamp 1679235063
transform 1 0 25392 0 -1 15232
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_24_3
timestamp 1679235063
transform 1 0 1380 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_15
timestamp 1679235063
transform 1 0 2484 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_24_27
timestamp 1679235063
transform 1 0 3588 0 1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_24_29
timestamp 1679235063
transform 1 0 3772 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_41
timestamp 1679235063
transform 1 0 4876 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_24_53
timestamp 1679235063
transform 1 0 5980 0 1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_24_81
timestamp 1679235063
transform 1 0 8556 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_24_85
timestamp 1679235063
transform 1 0 8924 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_24_95
timestamp 1679235063
transform 1 0 9844 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_24_120
timestamp 1679235063
transform 1 0 12144 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_24_127
timestamp 1679235063
transform 1 0 12788 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_24_138
timestamp 1679235063
transform 1 0 13800 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_24_143
timestamp 1679235063
transform 1 0 14260 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_24_149
timestamp 1679235063
transform 1 0 14812 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_24_153
timestamp 1679235063
transform 1 0 15180 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_24_157
timestamp 1679235063
transform 1 0 15548 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_24_178
timestamp 1679235063
transform 1 0 17480 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_24_182
timestamp 1679235063
transform 1 0 17848 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_24_192
timestamp 1679235063
transform 1 0 18768 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_24_197
timestamp 1679235063
transform 1 0 19228 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_24_208
timestamp 1679235063
transform 1 0 20240 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_24_215
timestamp 1679235063
transform 1 0 20884 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_24_222
timestamp 1679235063
transform 1 0 21528 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_24_229
timestamp 1679235063
transform 1 0 22172 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_24_233
timestamp 1679235063
transform 1 0 22540 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_24_250
timestamp 1679235063
transform 1 0 24104 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_24_253
timestamp 1679235063
transform 1 0 24380 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_24_263
timestamp 1679235063
transform 1 0 25300 0 1 15232
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_25_3
timestamp 1679235063
transform 1 0 1380 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_15
timestamp 1679235063
transform 1 0 2484 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_27
timestamp 1679235063
transform 1 0 3588 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_39
timestamp 1679235063
transform 1 0 4692 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_25_51
timestamp 1679235063
transform 1 0 5796 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_25_55
timestamp 1679235063
transform 1 0 6164 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_25_57
timestamp 1679235063
transform 1 0 6348 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_25_63
timestamp 1679235063
transform 1 0 6900 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_25_73
timestamp 1679235063
transform 1 0 7820 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_25_85
timestamp 1679235063
transform 1 0 8924 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_25_90
timestamp 1679235063
transform 1 0 9384 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_25_101
timestamp 1679235063
transform 1 0 10396 0 -1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_25_109
timestamp 1679235063
transform 1 0 11132 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_25_113
timestamp 1679235063
transform 1 0 11500 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_25_137
timestamp 1679235063
transform 1 0 13708 0 -1 16320
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_25_141
timestamp 1679235063
transform 1 0 14076 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_25_153
timestamp 1679235063
transform 1 0 15180 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_25_161
timestamp 1679235063
transform 1 0 15916 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_25_165
timestamp 1679235063
transform 1 0 16284 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_25_169
timestamp 1679235063
transform 1 0 16652 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_25_177
timestamp 1679235063
transform 1 0 17388 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_25_180
timestamp 1679235063
transform 1 0 17664 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_25_183
timestamp 1679235063
transform 1 0 17940 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_25_189
timestamp 1679235063
transform 1 0 18492 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_25_194
timestamp 1679235063
transform 1 0 18952 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_25_205
timestamp 1679235063
transform 1 0 19964 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_25_218
timestamp 1679235063
transform 1 0 21160 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_25_225
timestamp 1679235063
transform 1 0 21804 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_25_236
timestamp 1679235063
transform 1 0 22816 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_25_243
timestamp 1679235063
transform 1 0 23460 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_25_247
timestamp 1679235063
transform 1 0 23828 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_25_264
timestamp 1679235063
transform 1 0 25392 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_26_3
timestamp 1679235063
transform 1 0 1380 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_26_21
timestamp 1679235063
transform 1 0 3036 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_26_27
timestamp 1679235063
transform 1 0 3588 0 1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_26_29
timestamp 1679235063
transform 1 0 3772 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_41
timestamp 1679235063
transform 1 0 4876 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_26_73
timestamp 1679235063
transform 1 0 7820 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_26_77
timestamp 1679235063
transform 1 0 8188 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_26_85
timestamp 1679235063
transform 1 0 8924 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_26_96
timestamp 1679235063
transform 1 0 9936 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_26_109
timestamp 1679235063
transform 1 0 11132 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_26_121
timestamp 1679235063
transform 1 0 12236 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_26_125
timestamp 1679235063
transform 1 0 12604 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_26_130
timestamp 1679235063
transform 1 0 13064 0 1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_26_138
timestamp 1679235063
transform 1 0 13800 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_26_141
timestamp 1679235063
transform 1 0 14076 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_26_147
timestamp 1679235063
transform 1 0 14628 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_26_150
timestamp 1679235063
transform 1 0 14904 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_26_161
timestamp 1679235063
transform 1 0 15916 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_26_165
timestamp 1679235063
transform 1 0 16284 0 1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_26_168
timestamp 1679235063
transform 1 0 16560 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_26_180
timestamp 1679235063
transform 1 0 17664 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_26_191
timestamp 1679235063
transform 1 0 18676 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_26_195
timestamp 1679235063
transform 1 0 19044 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_26_199
timestamp 1679235063
transform 1 0 19412 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_26_204
timestamp 1679235063
transform 1 0 19872 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_26_212
timestamp 1679235063
transform 1 0 20608 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_26_220
timestamp 1679235063
transform 1 0 21344 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_26_244
timestamp 1679235063
transform 1 0 23552 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_26_248
timestamp 1679235063
transform 1 0 23920 0 1 16320
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_26_253
timestamp 1679235063
transform 1 0 24380 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_26_265
timestamp 1679235063
transform 1 0 25484 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_27_3
timestamp 1679235063
transform 1 0 1380 0 -1 17408
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_27_15
timestamp 1679235063
transform 1 0 2484 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_27
timestamp 1679235063
transform 1 0 3588 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_27_39
timestamp 1679235063
transform 1 0 4692 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_27_45
timestamp 1679235063
transform 1 0 5244 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_27_54
timestamp 1679235063
transform 1 0 6072 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_27_57
timestamp 1679235063
transform 1 0 6348 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_27_62
timestamp 1679235063
transform 1 0 6808 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_27_68
timestamp 1679235063
transform 1 0 7360 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_27_78
timestamp 1679235063
transform 1 0 8280 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_27_91
timestamp 1679235063
transform 1 0 9476 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_27_104
timestamp 1679235063
transform 1 0 10672 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_27_108
timestamp 1679235063
transform 1 0 11040 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_27_113
timestamp 1679235063
transform 1 0 11500 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_27_126
timestamp 1679235063
transform 1 0 12696 0 -1 17408
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_27_139
timestamp 1679235063
transform 1 0 13892 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_27_151
timestamp 1679235063
transform 1 0 14996 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_27_155
timestamp 1679235063
transform 1 0 15364 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_27_166
timestamp 1679235063
transform 1 0 16376 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_27_169
timestamp 1679235063
transform 1 0 16652 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_27_191
timestamp 1679235063
transform 1 0 18676 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_27_204
timestamp 1679235063
transform 1 0 19872 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_27_208
timestamp 1679235063
transform 1 0 20240 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_27_220
timestamp 1679235063
transform 1 0 21344 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_27_225
timestamp 1679235063
transform 1 0 21804 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_27_235
timestamp 1679235063
transform 1 0 22724 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_27_243
timestamp 1679235063
transform 1 0 23460 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_27_247
timestamp 1679235063
transform 1 0 23828 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_27_264
timestamp 1679235063
transform 1 0 25392 0 -1 17408
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_28_3
timestamp 1679235063
transform 1 0 1380 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_15
timestamp 1679235063
transform 1 0 2484 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_28_27
timestamp 1679235063
transform 1 0 3588 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_28_29
timestamp 1679235063
transform 1 0 3772 0 1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_28_37
timestamp 1679235063
transform 1 0 4508 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_28_60
timestamp 1679235063
transform 1 0 6624 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_28_64
timestamp 1679235063
transform 1 0 6992 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_28_74
timestamp 1679235063
transform 1 0 7912 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_28_78
timestamp 1679235063
transform 1 0 8280 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_28_82
timestamp 1679235063
transform 1 0 8648 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_28_85
timestamp 1679235063
transform 1 0 8924 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_28_98
timestamp 1679235063
transform 1 0 10120 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_28_104
timestamp 1679235063
transform 1 0 10672 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_28_128
timestamp 1679235063
transform 1 0 12880 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_28_132
timestamp 1679235063
transform 1 0 13248 0 1 17408
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_28_141
timestamp 1679235063
transform 1 0 14076 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_28_153
timestamp 1679235063
transform 1 0 15180 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_28_158
timestamp 1679235063
transform 1 0 15640 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_28_162
timestamp 1679235063
transform 1 0 16008 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_28_167
timestamp 1679235063
transform 1 0 16468 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_28_179
timestamp 1679235063
transform 1 0 17572 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_28_194
timestamp 1679235063
transform 1 0 18952 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_28_199
timestamp 1679235063
transform 1 0 19412 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_28_222
timestamp 1679235063
transform 1 0 21528 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_28_246
timestamp 1679235063
transform 1 0 23736 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_28_250
timestamp 1679235063
transform 1 0 24104 0 1 17408
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_28_253
timestamp 1679235063
transform 1 0 24380 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_28_265
timestamp 1679235063
transform 1 0 25484 0 1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_29_3
timestamp 1679235063
transform 1 0 1380 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_15
timestamp 1679235063
transform 1 0 2484 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_27
timestamp 1679235063
transform 1 0 3588 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_29_39
timestamp 1679235063
transform 1 0 4692 0 -1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_29_54
timestamp 1679235063
transform 1 0 6072 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_29_57
timestamp 1679235063
transform 1 0 6348 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_29_82
timestamp 1679235063
transform 1 0 8648 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_29_95
timestamp 1679235063
transform 1 0 9844 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_29_99
timestamp 1679235063
transform 1 0 10212 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_29_110
timestamp 1679235063
transform 1 0 11224 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_29_113
timestamp 1679235063
transform 1 0 11500 0 -1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_29_125
timestamp 1679235063
transform 1 0 12604 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_29_136
timestamp 1679235063
transform 1 0 13616 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_29_149
timestamp 1679235063
transform 1 0 14812 0 -1 18496
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_29_153
timestamp 1679235063
transform 1 0 15180 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_29_165
timestamp 1679235063
transform 1 0 16284 0 -1 18496
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_29_169
timestamp 1679235063
transform 1 0 16652 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_29_181
timestamp 1679235063
transform 1 0 17756 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_29_202
timestamp 1679235063
transform 1 0 19688 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_29_208
timestamp 1679235063
transform 1 0 20240 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_29_221
timestamp 1679235063
transform 1 0 21436 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_29_225
timestamp 1679235063
transform 1 0 21804 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_29_244
timestamp 1679235063
transform 1 0 23552 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_29_264
timestamp 1679235063
transform 1 0 25392 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_30_3
timestamp 1679235063
transform 1 0 1380 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_30_21
timestamp 1679235063
transform 1 0 3036 0 1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_30_27
timestamp 1679235063
transform 1 0 3588 0 1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_30_29
timestamp 1679235063
transform 1 0 3772 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_30_41
timestamp 1679235063
transform 1 0 4876 0 1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_30_49
timestamp 1679235063
transform 1 0 5612 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_30_59
timestamp 1679235063
transform 1 0 6532 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_30_70
timestamp 1679235063
transform 1 0 7544 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_30_82
timestamp 1679235063
transform 1 0 8648 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_30_85
timestamp 1679235063
transform 1 0 8924 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_30_108
timestamp 1679235063
transform 1 0 11040 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_30_114
timestamp 1679235063
transform 1 0 11592 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_30_125
timestamp 1679235063
transform 1 0 12604 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_30_138
timestamp 1679235063
transform 1 0 13800 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_30_141
timestamp 1679235063
transform 1 0 14076 0 1 18496
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_30_152
timestamp 1679235063
transform 1 0 15088 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_30_164
timestamp 1679235063
transform 1 0 16192 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_30_169
timestamp 1679235063
transform 1 0 16652 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_30_180
timestamp 1679235063
transform 1 0 17664 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_30_184
timestamp 1679235063
transform 1 0 18032 0 1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_30_194
timestamp 1679235063
transform 1 0 18952 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_30_199
timestamp 1679235063
transform 1 0 19412 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_30_211
timestamp 1679235063
transform 1 0 20516 0 1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_30_226
timestamp 1679235063
transform 1 0 21896 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_30_250
timestamp 1679235063
transform 1 0 24104 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_30_253
timestamp 1679235063
transform 1 0 24380 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_30_263
timestamp 1679235063
transform 1 0 25300 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_31_3
timestamp 1679235063
transform 1 0 1380 0 -1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_31_9
timestamp 1679235063
transform 1 0 1932 0 -1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_31_14
timestamp 1679235063
transform 1 0 2392 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_26
timestamp 1679235063
transform 1 0 3496 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_38
timestamp 1679235063
transform 1 0 4600 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_31_50
timestamp 1679235063
transform 1 0 5704 0 -1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_31_57
timestamp 1679235063
transform 1 0 6348 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_31_63
timestamp 1679235063
transform 1 0 6900 0 -1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_31_69
timestamp 1679235063
transform 1 0 7452 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_31_72
timestamp 1679235063
transform 1 0 7728 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_31_97
timestamp 1679235063
transform 1 0 10028 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_31_110
timestamp 1679235063
transform 1 0 11224 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_31_113
timestamp 1679235063
transform 1 0 11500 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_31_124
timestamp 1679235063
transform 1 0 12512 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_31_130
timestamp 1679235063
transform 1 0 13064 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_31_141
timestamp 1679235063
transform 1 0 14076 0 -1 19584
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_31_149
timestamp 1679235063
transform 1 0 14812 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_31_161
timestamp 1679235063
transform 1 0 15916 0 -1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_31_167
timestamp 1679235063
transform 1 0 16468 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_31_169
timestamp 1679235063
transform 1 0 16652 0 -1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_31_177
timestamp 1679235063
transform 1 0 17388 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_31_181
timestamp 1679235063
transform 1 0 17756 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_31_188
timestamp 1679235063
transform 1 0 18400 0 -1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_31_215
timestamp 1679235063
transform 1 0 20884 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_31_219
timestamp 1679235063
transform 1 0 21252 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_31_223
timestamp 1679235063
transform 1 0 21620 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_31_225
timestamp 1679235063
transform 1 0 21804 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_31_247
timestamp 1679235063
transform 1 0 23828 0 -1 19584
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_31_253
timestamp 1679235063
transform 1 0 24380 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_31_265
timestamp 1679235063
transform 1 0 25484 0 -1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_32_3
timestamp 1679235063
transform 1 0 1380 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_15
timestamp 1679235063
transform 1 0 2484 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_32_27
timestamp 1679235063
transform 1 0 3588 0 1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_32_29
timestamp 1679235063
transform 1 0 3772 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_32_41
timestamp 1679235063
transform 1 0 4876 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_32_45
timestamp 1679235063
transform 1 0 5244 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_32_66
timestamp 1679235063
transform 1 0 7176 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_32_70
timestamp 1679235063
transform 1 0 7544 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_32_82
timestamp 1679235063
transform 1 0 8648 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_32_85
timestamp 1679235063
transform 1 0 8924 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_32_96
timestamp 1679235063
transform 1 0 9936 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_32_105
timestamp 1679235063
transform 1 0 10764 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_32_109
timestamp 1679235063
transform 1 0 11132 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_32_119
timestamp 1679235063
transform 1 0 12052 0 1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_32_127
timestamp 1679235063
transform 1 0 12788 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_32_137
timestamp 1679235063
transform 1 0 13708 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_32_141
timestamp 1679235063
transform 1 0 14076 0 1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_32_149
timestamp 1679235063
transform 1 0 14812 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_32_154
timestamp 1679235063
transform 1 0 15272 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_32_158
timestamp 1679235063
transform 1 0 15640 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_32_163
timestamp 1679235063
transform 1 0 16100 0 1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_32_174
timestamp 1679235063
transform 1 0 17112 0 1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_32_184
timestamp 1679235063
transform 1 0 18032 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_32_191
timestamp 1679235063
transform 1 0 18676 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_32_195
timestamp 1679235063
transform 1 0 19044 0 1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_32_197
timestamp 1679235063
transform 1 0 19228 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_32_213
timestamp 1679235063
transform 1 0 20700 0 1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_32_221
timestamp 1679235063
transform 1 0 21436 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_32_230
timestamp 1679235063
transform 1 0 22264 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_32_250
timestamp 1679235063
transform 1 0 24104 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_32_253
timestamp 1679235063
transform 1 0 24380 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_32_259
timestamp 1679235063
transform 1 0 24932 0 1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_32_265
timestamp 1679235063
transform 1 0 25484 0 1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_33_3
timestamp 1679235063
transform 1 0 1380 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_33_15
timestamp 1679235063
transform 1 0 2484 0 -1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_33_23
timestamp 1679235063
transform 1 0 3220 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_33_27
timestamp 1679235063
transform 1 0 3588 0 -1 20672
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_33_36
timestamp 1679235063
transform 1 0 4416 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_33_48
timestamp 1679235063
transform 1 0 5520 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_33_52
timestamp 1679235063
transform 1 0 5888 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_33_55
timestamp 1679235063
transform 1 0 6164 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_33_57
timestamp 1679235063
transform 1 0 6348 0 -1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_33_73
timestamp 1679235063
transform 1 0 7820 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_33_86
timestamp 1679235063
transform 1 0 9016 0 -1 20672
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_33_92
timestamp 1679235063
transform 1 0 9568 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_33_104
timestamp 1679235063
transform 1 0 10672 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_33_110
timestamp 1679235063
transform 1 0 11224 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_33_113
timestamp 1679235063
transform 1 0 11500 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_33_124
timestamp 1679235063
transform 1 0 12512 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_33_128
timestamp 1679235063
transform 1 0 12880 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_33_152
timestamp 1679235063
transform 1 0 15088 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_33_164
timestamp 1679235063
transform 1 0 16192 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_33_169
timestamp 1679235063
transform 1 0 16652 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_33_174
timestamp 1679235063
transform 1 0 17112 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_33_178
timestamp 1679235063
transform 1 0 17480 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_33_183
timestamp 1679235063
transform 1 0 17940 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_33_187
timestamp 1679235063
transform 1 0 18308 0 -1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_33_202
timestamp 1679235063
transform 1 0 19688 0 -1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_33_210
timestamp 1679235063
transform 1 0 20424 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_33_220
timestamp 1679235063
transform 1 0 21344 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_33_225
timestamp 1679235063
transform 1 0 21804 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_33_244
timestamp 1679235063
transform 1 0 23552 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_33_264
timestamp 1679235063
transform 1 0 25392 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_34_3
timestamp 1679235063
transform 1 0 1380 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_34_21
timestamp 1679235063
transform 1 0 3036 0 1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_34_27
timestamp 1679235063
transform 1 0 3588 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_34_29
timestamp 1679235063
transform 1 0 3772 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_34_53
timestamp 1679235063
transform 1 0 5980 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_34_65
timestamp 1679235063
transform 1 0 7084 0 1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_34_73
timestamp 1679235063
transform 1 0 7820 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_34_82
timestamp 1679235063
transform 1 0 8648 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_34_85
timestamp 1679235063
transform 1 0 8924 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_34_96
timestamp 1679235063
transform 1 0 9936 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_34_100
timestamp 1679235063
transform 1 0 10304 0 1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_34_108
timestamp 1679235063
transform 1 0 11040 0 1 20672
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_34_119
timestamp 1679235063
transform 1 0 12052 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_34_131
timestamp 1679235063
transform 1 0 13156 0 1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_34_139
timestamp 1679235063
transform 1 0 13892 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_34_141
timestamp 1679235063
transform 1 0 14076 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_34_163
timestamp 1679235063
transform 1 0 16100 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_34_170
timestamp 1679235063
transform 1 0 16744 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_34_174
timestamp 1679235063
transform 1 0 17112 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_34_185
timestamp 1679235063
transform 1 0 18124 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_34_192
timestamp 1679235063
transform 1 0 18768 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_34_197
timestamp 1679235063
transform 1 0 19228 0 1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_34_203
timestamp 1679235063
transform 1 0 19780 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_34_224
timestamp 1679235063
transform 1 0 21712 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_34_228
timestamp 1679235063
transform 1 0 22080 0 1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_34_250
timestamp 1679235063
transform 1 0 24104 0 1 20672
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_34_253
timestamp 1679235063
transform 1 0 24380 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_34_265
timestamp 1679235063
transform 1 0 25484 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_35_3
timestamp 1679235063
transform 1 0 1380 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_35_7
timestamp 1679235063
transform 1 0 1748 0 -1 21760
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_35_29
timestamp 1679235063
transform 1 0 3772 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_35_41
timestamp 1679235063
transform 1 0 4876 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_35_53
timestamp 1679235063
transform 1 0 5980 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_35_57
timestamp 1679235063
transform 1 0 6348 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_35_69
timestamp 1679235063
transform 1 0 7452 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_35_96
timestamp 1679235063
transform 1 0 9936 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_35_100
timestamp 1679235063
transform 1 0 10304 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_35_110
timestamp 1679235063
transform 1 0 11224 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_35_113
timestamp 1679235063
transform 1 0 11500 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_35_117
timestamp 1679235063
transform 1 0 11868 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_35_120
timestamp 1679235063
transform 1 0 12144 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_35_123
timestamp 1679235063
transform 1 0 12420 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_35_127
timestamp 1679235063
transform 1 0 12788 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_35_131
timestamp 1679235063
transform 1 0 13156 0 -1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_35_141
timestamp 1679235063
transform 1 0 14076 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_35_152
timestamp 1679235063
transform 1 0 15088 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_35_156
timestamp 1679235063
transform 1 0 15456 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_35_159
timestamp 1679235063
transform 1 0 15732 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_35_166
timestamp 1679235063
transform 1 0 16376 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_35_169
timestamp 1679235063
transform 1 0 16652 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_35_172
timestamp 1679235063
transform 1 0 16928 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_35_183
timestamp 1679235063
transform 1 0 17940 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_35_207
timestamp 1679235063
transform 1 0 20148 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_35_219
timestamp 1679235063
transform 1 0 21252 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_35_223
timestamp 1679235063
transform 1 0 21620 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_35_225
timestamp 1679235063
transform 1 0 21804 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_35_236
timestamp 1679235063
transform 1 0 22816 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_35_260
timestamp 1679235063
transform 1 0 25024 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_35_264
timestamp 1679235063
transform 1 0 25392 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_36_3
timestamp 1679235063
transform 1 0 1380 0 1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_36_9
timestamp 1679235063
transform 1 0 1932 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_36_13
timestamp 1679235063
transform 1 0 2300 0 1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_36_21
timestamp 1679235063
transform 1 0 3036 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_36_25
timestamp 1679235063
transform 1 0 3404 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_36_29
timestamp 1679235063
transform 1 0 3772 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_36_53
timestamp 1679235063
transform 1 0 5980 0 1 21760
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_36_57
timestamp 1679235063
transform 1 0 6348 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_36_69
timestamp 1679235063
transform 1 0 7452 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_36_79
timestamp 1679235063
transform 1 0 8372 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_36_85
timestamp 1679235063
transform 1 0 8924 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_36_96
timestamp 1679235063
transform 1 0 9936 0 1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_36_104
timestamp 1679235063
transform 1 0 10672 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_36_107
timestamp 1679235063
transform 1 0 10948 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_36_118
timestamp 1679235063
transform 1 0 11960 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_36_122
timestamp 1679235063
transform 1 0 12328 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_36_132
timestamp 1679235063
transform 1 0 13248 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_36_136
timestamp 1679235063
transform 1 0 13616 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_36_145
timestamp 1679235063
transform 1 0 14444 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_36_157
timestamp 1679235063
transform 1 0 15548 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_36_170
timestamp 1679235063
transform 1 0 16744 0 1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_36_176
timestamp 1679235063
transform 1 0 17296 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_36_186
timestamp 1679235063
transform 1 0 18216 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_36_193
timestamp 1679235063
transform 1 0 18860 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_36_197
timestamp 1679235063
transform 1 0 19228 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_36_207
timestamp 1679235063
transform 1 0 20148 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_36_215
timestamp 1679235063
transform 1 0 20884 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_36_238
timestamp 1679235063
transform 1 0 23000 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_36_250
timestamp 1679235063
transform 1 0 24104 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_36_253
timestamp 1679235063
transform 1 0 24380 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_36_259
timestamp 1679235063
transform 1 0 24932 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_36_263
timestamp 1679235063
transform 1 0 25300 0 1 21760
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_37_3
timestamp 1679235063
transform 1 0 1380 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_15
timestamp 1679235063
transform 1 0 2484 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_37_27
timestamp 1679235063
transform 1 0 3588 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_37_33
timestamp 1679235063
transform 1 0 4140 0 -1 22848
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_37_42
timestamp 1679235063
transform 1 0 4968 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_37_54
timestamp 1679235063
transform 1 0 6072 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_37_57
timestamp 1679235063
transform 1 0 6348 0 -1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_37_73
timestamp 1679235063
transform 1 0 7820 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_37_88
timestamp 1679235063
transform 1 0 9200 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_37_92
timestamp 1679235063
transform 1 0 9568 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_37_96
timestamp 1679235063
transform 1 0 9936 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_37_99
timestamp 1679235063
transform 1 0 10212 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_37_110
timestamp 1679235063
transform 1 0 11224 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_37_113
timestamp 1679235063
transform 1 0 11500 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_37_118
timestamp 1679235063
transform 1 0 11960 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_37_122
timestamp 1679235063
transform 1 0 12328 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_37_125
timestamp 1679235063
transform 1 0 12604 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_37_130
timestamp 1679235063
transform 1 0 13064 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_37_143
timestamp 1679235063
transform 1 0 14260 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_37_155
timestamp 1679235063
transform 1 0 15364 0 -1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_37_166
timestamp 1679235063
transform 1 0 16376 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_37_169
timestamp 1679235063
transform 1 0 16652 0 -1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_37_177
timestamp 1679235063
transform 1 0 17388 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_37_182
timestamp 1679235063
transform 1 0 17848 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_37_195
timestamp 1679235063
transform 1 0 19044 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_37_207
timestamp 1679235063
transform 1 0 20148 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_37_222
timestamp 1679235063
transform 1 0 21528 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_37_225
timestamp 1679235063
transform 1 0 21804 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_37_251
timestamp 1679235063
transform 1 0 24196 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_37_258
timestamp 1679235063
transform 1 0 24840 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_37_262
timestamp 1679235063
transform 1 0 25208 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_38_3
timestamp 1679235063
transform 1 0 1380 0 1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_38_26
timestamp 1679235063
transform 1 0 3496 0 1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_38_29
timestamp 1679235063
transform 1 0 3772 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_38_33
timestamp 1679235063
transform 1 0 4140 0 1 22848
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_38_42
timestamp 1679235063
transform 1 0 4968 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_38_54
timestamp 1679235063
transform 1 0 6072 0 1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_38_76
timestamp 1679235063
transform 1 0 8096 0 1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_38_80
timestamp 1679235063
transform 1 0 8464 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_38_85
timestamp 1679235063
transform 1 0 8924 0 1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_38_91
timestamp 1679235063
transform 1 0 9476 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_38_95
timestamp 1679235063
transform 1 0 9844 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_38_110
timestamp 1679235063
transform 1 0 11224 0 1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_38_116
timestamp 1679235063
transform 1 0 11776 0 1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_38_138
timestamp 1679235063
transform 1 0 13800 0 1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_38_141
timestamp 1679235063
transform 1 0 14076 0 1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_38_152
timestamp 1679235063
transform 1 0 15088 0 1 22848
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_38_156
timestamp 1679235063
transform 1 0 15456 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_38_168
timestamp 1679235063
transform 1 0 16560 0 1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_38_194
timestamp 1679235063
transform 1 0 18952 0 1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_38_197
timestamp 1679235063
transform 1 0 19228 0 1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_38_219
timestamp 1679235063
transform 1 0 21252 0 1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_38_223
timestamp 1679235063
transform 1 0 21620 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_38_230
timestamp 1679235063
transform 1 0 22264 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_38_250
timestamp 1679235063
transform 1 0 24104 0 1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_38_253
timestamp 1679235063
transform 1 0 24380 0 1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_38_264
timestamp 1679235063
transform 1 0 25392 0 1 22848
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_39_3
timestamp 1679235063
transform 1 0 1380 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_15
timestamp 1679235063
transform 1 0 2484 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_39_27
timestamp 1679235063
transform 1 0 3588 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_39_31
timestamp 1679235063
transform 1 0 3956 0 -1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_39_39
timestamp 1679235063
transform 1 0 4692 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_39_49
timestamp 1679235063
transform 1 0 5612 0 -1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_39_55
timestamp 1679235063
transform 1 0 6164 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_39_57
timestamp 1679235063
transform 1 0 6348 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_39_79
timestamp 1679235063
transform 1 0 8372 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_39_83
timestamp 1679235063
transform 1 0 8740 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_39_87
timestamp 1679235063
transform 1 0 9108 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_39_97
timestamp 1679235063
transform 1 0 10028 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_39_110
timestamp 1679235063
transform 1 0 11224 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_39_113
timestamp 1679235063
transform 1 0 11500 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_39_118
timestamp 1679235063
transform 1 0 11960 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_39_129
timestamp 1679235063
transform 1 0 12972 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_39_142
timestamp 1679235063
transform 1 0 14168 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_39_148
timestamp 1679235063
transform 1 0 14720 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_39_153
timestamp 1679235063
transform 1 0 15180 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_39_164
timestamp 1679235063
transform 1 0 16192 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_39_169
timestamp 1679235063
transform 1 0 16652 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_39_180
timestamp 1679235063
transform 1 0 17664 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_39_187
timestamp 1679235063
transform 1 0 18308 0 -1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_39_193
timestamp 1679235063
transform 1 0 18860 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_39_196
timestamp 1679235063
transform 1 0 19136 0 -1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_39_222
timestamp 1679235063
transform 1 0 21528 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_39_227
timestamp 1679235063
transform 1 0 21988 0 -1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_39_235
timestamp 1679235063
transform 1 0 22724 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_39_256
timestamp 1679235063
transform 1 0 24656 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_39_264
timestamp 1679235063
transform 1 0 25392 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_40_3
timestamp 1679235063
transform 1 0 1380 0 1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_40_9
timestamp 1679235063
transform 1 0 1932 0 1 23936
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_40_13
timestamp 1679235063
transform 1 0 2300 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_40_25
timestamp 1679235063
transform 1 0 3404 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_40_29
timestamp 1679235063
transform 1 0 3772 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_40_51
timestamp 1679235063
transform 1 0 5796 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_40_55
timestamp 1679235063
transform 1 0 6164 0 1 23936
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_40_67
timestamp 1679235063
transform 1 0 7268 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_40_79
timestamp 1679235063
transform 1 0 8372 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_40_83
timestamp 1679235063
transform 1 0 8740 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_40_85
timestamp 1679235063
transform 1 0 8924 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_40_90
timestamp 1679235063
transform 1 0 9384 0 1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_40_96
timestamp 1679235063
transform 1 0 9936 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_40_99
timestamp 1679235063
transform 1 0 10212 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_40_104
timestamp 1679235063
transform 1 0 10672 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_40_127
timestamp 1679235063
transform 1 0 12788 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_40_135
timestamp 1679235063
transform 1 0 13524 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_40_139
timestamp 1679235063
transform 1 0 13892 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_40_141
timestamp 1679235063
transform 1 0 14076 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_40_151
timestamp 1679235063
transform 1 0 14996 0 1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_40_157
timestamp 1679235063
transform 1 0 15548 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_40_178
timestamp 1679235063
transform 1 0 17480 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_40_190
timestamp 1679235063
transform 1 0 18584 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_40_194
timestamp 1679235063
transform 1 0 18952 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_40_199
timestamp 1679235063
transform 1 0 19412 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_40_203
timestamp 1679235063
transform 1 0 19780 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_40_214
timestamp 1679235063
transform 1 0 20792 0 1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_40_220
timestamp 1679235063
transform 1 0 21344 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_40_230
timestamp 1679235063
transform 1 0 22264 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_40_250
timestamp 1679235063
transform 1 0 24104 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_40_253
timestamp 1679235063
transform 1 0 24380 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_40_259
timestamp 1679235063
transform 1 0 24932 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_40_263
timestamp 1679235063
transform 1 0 25300 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_41_3
timestamp 1679235063
transform 1 0 1380 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_41_27
timestamp 1679235063
transform 1 0 3588 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_41_51
timestamp 1679235063
transform 1 0 5796 0 -1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_41_55
timestamp 1679235063
transform 1 0 6164 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_41_57
timestamp 1679235063
transform 1 0 6348 0 -1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_41_67
timestamp 1679235063
transform 1 0 7268 0 -1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_41_73
timestamp 1679235063
transform 1 0 7820 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_41_76
timestamp 1679235063
transform 1 0 8096 0 -1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_41_87
timestamp 1679235063
transform 1 0 9108 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_41_100
timestamp 1679235063
transform 1 0 10304 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_41_107
timestamp 1679235063
transform 1 0 10948 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_41_113
timestamp 1679235063
transform 1 0 11500 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_41_125
timestamp 1679235063
transform 1 0 12604 0 -1 25024
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_41_138
timestamp 1679235063
transform 1 0 13800 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_41_153
timestamp 1679235063
transform 1 0 15180 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_41_166
timestamp 1679235063
transform 1 0 16376 0 -1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_41_169
timestamp 1679235063
transform 1 0 16652 0 -1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_41_175
timestamp 1679235063
transform 1 0 17204 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_41_196
timestamp 1679235063
transform 1 0 19136 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_41_200
timestamp 1679235063
transform 1 0 19504 0 -1 25024
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_41_210
timestamp 1679235063
transform 1 0 20424 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_41_222
timestamp 1679235063
transform 1 0 21528 0 -1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_41_229
timestamp 1679235063
transform 1 0 22172 0 -1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_41_234
timestamp 1679235063
transform 1 0 22632 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_41_258
timestamp 1679235063
transform 1 0 24840 0 -1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_41_262
timestamp 1679235063
transform 1 0 25208 0 -1 25024
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_42_3
timestamp 1679235063
transform 1 0 1380 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_15
timestamp 1679235063
transform 1 0 2484 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_42_27
timestamp 1679235063
transform 1 0 3588 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_42_29
timestamp 1679235063
transform 1 0 3772 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_42_35
timestamp 1679235063
transform 1 0 4324 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_42_39
timestamp 1679235063
transform 1 0 4692 0 1 25024
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_42_48
timestamp 1679235063
transform 1 0 5520 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_42_60
timestamp 1679235063
transform 1 0 6624 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_42_64
timestamp 1679235063
transform 1 0 6992 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_42_67
timestamp 1679235063
transform 1 0 7268 0 1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_42_78
timestamp 1679235063
transform 1 0 8280 0 1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  FILLER_42_85
timestamp 1679235063
transform 1 0 8924 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_42_108
timestamp 1679235063
transform 1 0 11040 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_42_112
timestamp 1679235063
transform 1 0 11408 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_42_116
timestamp 1679235063
transform 1 0 11776 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_42_129
timestamp 1679235063
transform 1 0 12972 0 1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_42_137
timestamp 1679235063
transform 1 0 13708 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_42_141
timestamp 1679235063
transform 1 0 14076 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_42_145
timestamp 1679235063
transform 1 0 14444 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_42_155
timestamp 1679235063
transform 1 0 15364 0 1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_42_163
timestamp 1679235063
transform 1 0 16100 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_42_168
timestamp 1679235063
transform 1 0 16560 0 1 25024
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_42_179
timestamp 1679235063
transform 1 0 17572 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_42_191
timestamp 1679235063
transform 1 0 18676 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_42_195
timestamp 1679235063
transform 1 0 19044 0 1 25024
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_42_197
timestamp 1679235063
transform 1 0 19228 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_42_229
timestamp 1679235063
transform 1 0 22172 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_42_241
timestamp 1679235063
transform 1 0 23276 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_42_245
timestamp 1679235063
transform 1 0 23644 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_42_250
timestamp 1679235063
transform 1 0 24104 0 1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_42_253
timestamp 1679235063
transform 1 0 24380 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_42_259
timestamp 1679235063
transform 1 0 24932 0 1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_42_265
timestamp 1679235063
transform 1 0 25484 0 1 25024
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_43_3
timestamp 1679235063
transform 1 0 1380 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_43_15
timestamp 1679235063
transform 1 0 2484 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_43_19
timestamp 1679235063
transform 1 0 2852 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_43_22
timestamp 1679235063
transform 1 0 3128 0 -1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_43_27
timestamp 1679235063
transform 1 0 3588 0 -1 26112
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_43_38
timestamp 1679235063
transform 1 0 4600 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_43_50
timestamp 1679235063
transform 1 0 5704 0 -1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_43_57
timestamp 1679235063
transform 1 0 6348 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_43_61
timestamp 1679235063
transform 1 0 6716 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_43_65
timestamp 1679235063
transform 1 0 7084 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_43_89
timestamp 1679235063
transform 1 0 9292 0 -1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_43_93
timestamp 1679235063
transform 1 0 9660 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_43_97
timestamp 1679235063
transform 1 0 10028 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_43_107
timestamp 1679235063
transform 1 0 10948 0 -1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_43_111
timestamp 1679235063
transform 1 0 11316 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_43_113
timestamp 1679235063
transform 1 0 11500 0 -1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_43_118
timestamp 1679235063
transform 1 0 11960 0 -1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_43_122
timestamp 1679235063
transform 1 0 12328 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_43_134
timestamp 1679235063
transform 1 0 13432 0 -1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_43_142
timestamp 1679235063
transform 1 0 14168 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_43_166
timestamp 1679235063
transform 1 0 16376 0 -1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_43_171
timestamp 1679235063
transform 1 0 16836 0 -1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_43_179
timestamp 1679235063
transform 1 0 17572 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_43_191
timestamp 1679235063
transform 1 0 18676 0 -1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_43_206
timestamp 1679235063
transform 1 0 20056 0 -1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_43_214
timestamp 1679235063
transform 1 0 20792 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_43_217
timestamp 1679235063
transform 1 0 21068 0 -1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_43_222
timestamp 1679235063
transform 1 0 21528 0 -1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_43_225
timestamp 1679235063
transform 1 0 21804 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_43_237
timestamp 1679235063
transform 1 0 22908 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_43_244
timestamp 1679235063
transform 1 0 23552 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_43_264
timestamp 1679235063
transform 1 0 25392 0 -1 26112
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_44_3
timestamp 1679235063
transform 1 0 1380 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_44_15
timestamp 1679235063
transform 1 0 2484 0 1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_44_23
timestamp 1679235063
transform 1 0 3220 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_44_29
timestamp 1679235063
transform 1 0 3772 0 1 26112
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_44_38
timestamp 1679235063
transform 1 0 4600 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_44_50
timestamp 1679235063
transform 1 0 5704 0 1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_44_78
timestamp 1679235063
transform 1 0 8280 0 1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_44_82
timestamp 1679235063
transform 1 0 8648 0 1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_44_85
timestamp 1679235063
transform 1 0 8924 0 1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_44_89
timestamp 1679235063
transform 1 0 9292 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_44_98
timestamp 1679235063
transform 1 0 10120 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_44_103
timestamp 1679235063
transform 1 0 10580 0 1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_44_114
timestamp 1679235063
transform 1 0 11592 0 1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_44_125
timestamp 1679235063
transform 1 0 12604 0 1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_44_138
timestamp 1679235063
transform 1 0 13800 0 1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_44_143
timestamp 1679235063
transform 1 0 14260 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_44_148
timestamp 1679235063
transform 1 0 14720 0 1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_44_159
timestamp 1679235063
transform 1 0 15732 0 1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_44_171
timestamp 1679235063
transform 1 0 16836 0 1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_44_179
timestamp 1679235063
transform 1 0 17572 0 1 26112
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_44_184
timestamp 1679235063
transform 1 0 18032 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_44_197
timestamp 1679235063
transform 1 0 19228 0 1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_44_208
timestamp 1679235063
transform 1 0 20240 0 1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_44_212
timestamp 1679235063
transform 1 0 20608 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_44_217
timestamp 1679235063
transform 1 0 21068 0 1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_44_228
timestamp 1679235063
transform 1 0 22080 0 1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_44_241
timestamp 1679235063
transform 1 0 23276 0 1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_44_245
timestamp 1679235063
transform 1 0 23644 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_44_250
timestamp 1679235063
transform 1 0 24104 0 1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_44_253
timestamp 1679235063
transform 1 0 24380 0 1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_44_263
timestamp 1679235063
transform 1 0 25300 0 1 26112
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_45_3
timestamp 1679235063
transform 1 0 1380 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_45_15
timestamp 1679235063
transform 1 0 2484 0 -1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_45_23
timestamp 1679235063
transform 1 0 3220 0 -1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_45_46
timestamp 1679235063
transform 1 0 5336 0 -1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_45_54
timestamp 1679235063
transform 1 0 6072 0 -1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_45_57
timestamp 1679235063
transform 1 0 6348 0 -1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_45_79
timestamp 1679235063
transform 1 0 8372 0 -1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_45_85
timestamp 1679235063
transform 1 0 8924 0 -1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_45_96
timestamp 1679235063
transform 1 0 9936 0 -1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_45_102
timestamp 1679235063
transform 1 0 10488 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_45_107
timestamp 1679235063
transform 1 0 10948 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_45_111
timestamp 1679235063
transform 1 0 11316 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_45_113
timestamp 1679235063
transform 1 0 11500 0 -1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_45_123
timestamp 1679235063
transform 1 0 12420 0 -1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_45_131
timestamp 1679235063
transform 1 0 13156 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_45_152
timestamp 1679235063
transform 1 0 15088 0 -1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_45_156
timestamp 1679235063
transform 1 0 15456 0 -1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_45_164
timestamp 1679235063
transform 1 0 16192 0 -1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_45_169
timestamp 1679235063
transform 1 0 16652 0 -1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_45_180
timestamp 1679235063
transform 1 0 17664 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_45_193
timestamp 1679235063
transform 1 0 18860 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_45_200
timestamp 1679235063
transform 1 0 19504 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_45_207
timestamp 1679235063
transform 1 0 20148 0 -1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_45_211
timestamp 1679235063
transform 1 0 20516 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_45_222
timestamp 1679235063
transform 1 0 21528 0 -1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_45_225
timestamp 1679235063
transform 1 0 21804 0 -1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_45_248
timestamp 1679235063
transform 1 0 23920 0 -1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_45_252
timestamp 1679235063
transform 1 0 24288 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_45_259
timestamp 1679235063
transform 1 0 24932 0 -1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_45_263
timestamp 1679235063
transform 1 0 25300 0 -1 27200
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_46_3
timestamp 1679235063
transform 1 0 1380 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_15
timestamp 1679235063
transform 1 0 2484 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_46_27
timestamp 1679235063
transform 1 0 3588 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_46_29
timestamp 1679235063
transform 1 0 3772 0 1 27200
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_46_34
timestamp 1679235063
transform 1 0 4232 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_46
timestamp 1679235063
transform 1 0 5336 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_46_58
timestamp 1679235063
transform 1 0 6440 0 1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_46_68
timestamp 1679235063
transform 1 0 7360 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_46_73
timestamp 1679235063
transform 1 0 7820 0 1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_46_81
timestamp 1679235063
transform 1 0 8556 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_46_85
timestamp 1679235063
transform 1 0 8924 0 1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_46_91
timestamp 1679235063
transform 1 0 9476 0 1 27200
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_46_95
timestamp 1679235063
transform 1 0 9844 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_46_107
timestamp 1679235063
transform 1 0 10948 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_46_110
timestamp 1679235063
transform 1 0 11224 0 1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_46_121
timestamp 1679235063
transform 1 0 12236 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_46_127
timestamp 1679235063
transform 1 0 12788 0 1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_46_138
timestamp 1679235063
transform 1 0 13800 0 1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_46_141
timestamp 1679235063
transform 1 0 14076 0 1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_46_151
timestamp 1679235063
transform 1 0 14996 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_46_176
timestamp 1679235063
transform 1 0 17296 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_46_189
timestamp 1679235063
transform 1 0 18492 0 1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_46_193
timestamp 1679235063
transform 1 0 18860 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_46_197
timestamp 1679235063
transform 1 0 19228 0 1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_46_208
timestamp 1679235063
transform 1 0 20240 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_46_221
timestamp 1679235063
transform 1 0 21436 0 1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_46_229
timestamp 1679235063
transform 1 0 22172 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_46_250
timestamp 1679235063
transform 1 0 24104 0 1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_46_253
timestamp 1679235063
transform 1 0 24380 0 1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_46_259
timestamp 1679235063
transform 1 0 24932 0 1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_46_265
timestamp 1679235063
transform 1 0 25484 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_47_3
timestamp 1679235063
transform 1 0 1380 0 -1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_47_9
timestamp 1679235063
transform 1 0 1932 0 -1 28288
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_47_31
timestamp 1679235063
transform 1 0 3956 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_43
timestamp 1679235063
transform 1 0 5060 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_47_55
timestamp 1679235063
transform 1 0 6164 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_47_57
timestamp 1679235063
transform 1 0 6348 0 -1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_47_79
timestamp 1679235063
transform 1 0 8372 0 -1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_47_83
timestamp 1679235063
transform 1 0 8740 0 -1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_47_87
timestamp 1679235063
transform 1 0 9108 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_47_108
timestamp 1679235063
transform 1 0 11040 0 -1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_47_113
timestamp 1679235063
transform 1 0 11500 0 -1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_47_123
timestamp 1679235063
transform 1 0 12420 0 -1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_47_149
timestamp 1679235063
transform 1 0 14812 0 -1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_47_153
timestamp 1679235063
transform 1 0 15180 0 -1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_47_163
timestamp 1679235063
transform 1 0 16100 0 -1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_47_167
timestamp 1679235063
transform 1 0 16468 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_47_169
timestamp 1679235063
transform 1 0 16652 0 -1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_47_175
timestamp 1679235063
transform 1 0 17204 0 -1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_47_186
timestamp 1679235063
transform 1 0 18216 0 -1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_47_192
timestamp 1679235063
transform 1 0 18768 0 -1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_47_216
timestamp 1679235063
transform 1 0 20976 0 -1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_47_220
timestamp 1679235063
transform 1 0 21344 0 -1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_47_225
timestamp 1679235063
transform 1 0 21804 0 -1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_47_248
timestamp 1679235063
transform 1 0 23920 0 -1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_47_252
timestamp 1679235063
transform 1 0 24288 0 -1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_47_259
timestamp 1679235063
transform 1 0 24932 0 -1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_47_263
timestamp 1679235063
transform 1 0 25300 0 -1 28288
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_48_3
timestamp 1679235063
transform 1 0 1380 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_15
timestamp 1679235063
transform 1 0 2484 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_48_27
timestamp 1679235063
transform 1 0 3588 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_48_29
timestamp 1679235063
transform 1 0 3772 0 1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_48_52
timestamp 1679235063
transform 1 0 5888 0 1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_48_56
timestamp 1679235063
transform 1 0 6256 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_48_59
timestamp 1679235063
transform 1 0 6532 0 1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_48_69
timestamp 1679235063
transform 1 0 7452 0 1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_48_82
timestamp 1679235063
transform 1 0 8648 0 1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_48_85
timestamp 1679235063
transform 1 0 8924 0 1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_48_107
timestamp 1679235063
transform 1 0 10948 0 1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_48_111
timestamp 1679235063
transform 1 0 11316 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_48_121
timestamp 1679235063
transform 1 0 12236 0 1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_48_134
timestamp 1679235063
transform 1 0 13432 0 1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_48_141
timestamp 1679235063
transform 1 0 14076 0 1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_48_152
timestamp 1679235063
transform 1 0 15088 0 1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_48_158
timestamp 1679235063
transform 1 0 15640 0 1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_48_173
timestamp 1679235063
transform 1 0 17020 0 1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_48_177
timestamp 1679235063
transform 1 0 17388 0 1 28288
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_48_184
timestamp 1679235063
transform 1 0 18032 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_197
timestamp 1679235063
transform 1 0 19228 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_48_209
timestamp 1679235063
transform 1 0 20332 0 1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_48_215
timestamp 1679235063
transform 1 0 20884 0 1 28288
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_48_226
timestamp 1679235063
transform 1 0 21896 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_48_238
timestamp 1679235063
transform 1 0 23000 0 1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_48_246
timestamp 1679235063
transform 1 0 23736 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_48_250
timestamp 1679235063
transform 1 0 24104 0 1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_48_253
timestamp 1679235063
transform 1 0 24380 0 1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_48_258
timestamp 1679235063
transform 1 0 24840 0 1 28288
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_49_3
timestamp 1679235063
transform 1 0 1380 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_49_15
timestamp 1679235063
transform 1 0 2484 0 -1 29376
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_49_26
timestamp 1679235063
transform 1 0 3496 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_38
timestamp 1679235063
transform 1 0 4600 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_49_50
timestamp 1679235063
transform 1 0 5704 0 -1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_49_57
timestamp 1679235063
transform 1 0 6348 0 -1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_49_63
timestamp 1679235063
transform 1 0 6900 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_49_84
timestamp 1679235063
transform 1 0 8832 0 -1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_49_92
timestamp 1679235063
transform 1 0 9568 0 -1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_49_103
timestamp 1679235063
transform 1 0 10580 0 -1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_49_109
timestamp 1679235063
transform 1 0 11132 0 -1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_49_115
timestamp 1679235063
transform 1 0 11684 0 -1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_49_127
timestamp 1679235063
transform 1 0 12788 0 -1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_49_131
timestamp 1679235063
transform 1 0 13156 0 -1 29376
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_49_143
timestamp 1679235063
transform 1 0 14260 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_49_155
timestamp 1679235063
transform 1 0 15364 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_49_165
timestamp 1679235063
transform 1 0 16284 0 -1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_49_169
timestamp 1679235063
transform 1 0 16652 0 -1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_49_180
timestamp 1679235063
transform 1 0 17664 0 -1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_49_193
timestamp 1679235063
transform 1 0 18860 0 -1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_49_201
timestamp 1679235063
transform 1 0 19596 0 -1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_49_212
timestamp 1679235063
transform 1 0 20608 0 -1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_49_216
timestamp 1679235063
transform 1 0 20976 0 -1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_49_222
timestamp 1679235063
transform 1 0 21528 0 -1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_49_225
timestamp 1679235063
transform 1 0 21804 0 -1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_49_236
timestamp 1679235063
transform 1 0 22816 0 -1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_49_246
timestamp 1679235063
transform 1 0 23736 0 -1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_49_251
timestamp 1679235063
transform 1 0 24196 0 -1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_49_259
timestamp 1679235063
transform 1 0 24932 0 -1 29376
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_50_3
timestamp 1679235063
transform 1 0 1380 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_15
timestamp 1679235063
transform 1 0 2484 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_50_27
timestamp 1679235063
transform 1 0 3588 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_50_29
timestamp 1679235063
transform 1 0 3772 0 1 29376
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_50_52
timestamp 1679235063
transform 1 0 5888 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_50_64
timestamp 1679235063
transform 1 0 6992 0 1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_50_68
timestamp 1679235063
transform 1 0 7360 0 1 29376
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_50_71
timestamp 1679235063
transform 1 0 7636 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_50_83
timestamp 1679235063
transform 1 0 8740 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_50_85
timestamp 1679235063
transform 1 0 8924 0 1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_50_113
timestamp 1679235063
transform 1 0 11500 0 1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_50_125
timestamp 1679235063
transform 1 0 12604 0 1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_50_129
timestamp 1679235063
transform 1 0 12972 0 1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_50_137
timestamp 1679235063
transform 1 0 13708 0 1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_50_141
timestamp 1679235063
transform 1 0 14076 0 1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_50_167
timestamp 1679235063
transform 1 0 16468 0 1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_50_171
timestamp 1679235063
transform 1 0 16836 0 1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_50_182
timestamp 1679235063
transform 1 0 17848 0 1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_50_189
timestamp 1679235063
transform 1 0 18492 0 1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_50_195
timestamp 1679235063
transform 1 0 19044 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_50_197
timestamp 1679235063
transform 1 0 19228 0 1 29376
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_50_209
timestamp 1679235063
transform 1 0 20332 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_221
timestamp 1679235063
transform 1 0 21436 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_50_233
timestamp 1679235063
transform 1 0 22540 0 1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_50_245
timestamp 1679235063
transform 1 0 23644 0 1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_50_251
timestamp 1679235063
transform 1 0 24196 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_50_253
timestamp 1679235063
transform 1 0 24380 0 1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_50_264
timestamp 1679235063
transform 1 0 25392 0 1 29376
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_51_3
timestamp 1679235063
transform 1 0 1380 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_15
timestamp 1679235063
transform 1 0 2484 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_27
timestamp 1679235063
transform 1 0 3588 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_39
timestamp 1679235063
transform 1 0 4692 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_51_51
timestamp 1679235063
transform 1 0 5796 0 -1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_51_55
timestamp 1679235063
transform 1 0 6164 0 -1 30464
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_51_57
timestamp 1679235063
transform 1 0 6348 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_69
timestamp 1679235063
transform 1 0 7452 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_51_81
timestamp 1679235063
transform 1 0 8556 0 -1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_51_92
timestamp 1679235063
transform 1 0 9568 0 -1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_51_96
timestamp 1679235063
transform 1 0 9936 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_51_99
timestamp 1679235063
transform 1 0 10212 0 -1 30464
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_51_110
timestamp 1679235063
transform 1 0 11224 0 -1 30464
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_51_113
timestamp 1679235063
transform 1 0 11500 0 -1 30464
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_51_118
timestamp 1679235063
transform 1 0 11960 0 -1 30464
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_51_133
timestamp 1679235063
transform 1 0 13340 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_51_145
timestamp 1679235063
transform 1 0 14444 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_51_166
timestamp 1679235063
transform 1 0 16376 0 -1 30464
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_51_171
timestamp 1679235063
transform 1 0 16836 0 -1 30464
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_51_175
timestamp 1679235063
transform 1 0 17204 0 -1 30464
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_51_186
timestamp 1679235063
transform 1 0 18216 0 -1 30464
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_51_190
timestamp 1679235063
transform 1 0 18584 0 -1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_51_196
timestamp 1679235063
transform 1 0 19136 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_51_199
timestamp 1679235063
transform 1 0 19412 0 -1 30464
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_51_204
timestamp 1679235063
transform 1 0 19872 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_51_216
timestamp 1679235063
transform 1 0 20976 0 -1 30464
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_51_225
timestamp 1679235063
transform 1 0 21804 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_51_237
timestamp 1679235063
transform 1 0 22908 0 -1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_51_241
timestamp 1679235063
transform 1 0 23276 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_51_262
timestamp 1679235063
transform 1 0 25208 0 -1 30464
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_52_3
timestamp 1679235063
transform 1 0 1380 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_15
timestamp 1679235063
transform 1 0 2484 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_52_27
timestamp 1679235063
transform 1 0 3588 0 1 30464
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_52_29
timestamp 1679235063
transform 1 0 3772 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_41
timestamp 1679235063
transform 1 0 4876 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_53
timestamp 1679235063
transform 1 0 5980 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_52_65
timestamp 1679235063
transform 1 0 7084 0 1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_52_70
timestamp 1679235063
transform 1 0 7544 0 1 30464
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_52_81
timestamp 1679235063
transform 1 0 8556 0 1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_52_87
timestamp 1679235063
transform 1 0 9108 0 1 30464
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_52_101
timestamp 1679235063
transform 1 0 10396 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_52_113
timestamp 1679235063
transform 1 0 11500 0 1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_52_117
timestamp 1679235063
transform 1 0 11868 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_52_122
timestamp 1679235063
transform 1 0 12328 0 1 30464
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_52_133
timestamp 1679235063
transform 1 0 13340 0 1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_52_139
timestamp 1679235063
transform 1 0 13892 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_52_141
timestamp 1679235063
transform 1 0 14076 0 1 30464
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_52_152
timestamp 1679235063
transform 1 0 15088 0 1 30464
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_52_158
timestamp 1679235063
transform 1 0 15640 0 1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_52_170
timestamp 1679235063
transform 1 0 16744 0 1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_52_194
timestamp 1679235063
transform 1 0 18952 0 1 30464
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_52_197
timestamp 1679235063
transform 1 0 19228 0 1 30464
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_52_208
timestamp 1679235063
transform 1 0 20240 0 1 30464
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_52_212
timestamp 1679235063
transform 1 0 20608 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_52_224
timestamp 1679235063
transform 1 0 21712 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_52_234
timestamp 1679235063
transform 1 0 22632 0 1 30464
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_52_238
timestamp 1679235063
transform 1 0 23000 0 1 30464
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_52_249
timestamp 1679235063
transform 1 0 24012 0 1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_52_253
timestamp 1679235063
transform 1 0 24380 0 1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_52_259
timestamp 1679235063
transform 1 0 24932 0 1 30464
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_52_264
timestamp 1679235063
transform 1 0 25392 0 1 30464
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_53_3
timestamp 1679235063
transform 1 0 1380 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_15
timestamp 1679235063
transform 1 0 2484 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_53_48
timestamp 1679235063
transform 1 0 5520 0 -1 31552
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_53_57
timestamp 1679235063
transform 1 0 6348 0 -1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_53_65
timestamp 1679235063
transform 1 0 7084 0 -1 31552
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_53_76
timestamp 1679235063
transform 1 0 8096 0 -1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_53_83
timestamp 1679235063
transform 1 0 8740 0 -1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_53_89
timestamp 1679235063
transform 1 0 9292 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_53_110
timestamp 1679235063
transform 1 0 11224 0 -1 31552
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_53_115
timestamp 1679235063
transform 1 0 11684 0 -1 31552
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_53_123
timestamp 1679235063
transform 1 0 12420 0 -1 31552
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_53_145
timestamp 1679235063
transform 1 0 14444 0 -1 31552
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_53_149
timestamp 1679235063
transform 1 0 14812 0 -1 31552
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_53_157
timestamp 1679235063
transform 1 0 15548 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_53_166
timestamp 1679235063
transform 1 0 16376 0 -1 31552
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_53_169
timestamp 1679235063
transform 1 0 16652 0 -1 31552
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_53_180
timestamp 1679235063
transform 1 0 17664 0 -1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_53_184
timestamp 1679235063
transform 1 0 18032 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_53_194
timestamp 1679235063
transform 1 0 18952 0 -1 31552
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_53_209
timestamp 1679235063
transform 1 0 20332 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_53_221
timestamp 1679235063
transform 1 0 21436 0 -1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_53_225
timestamp 1679235063
transform 1 0 21804 0 -1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_53_248
timestamp 1679235063
transform 1 0 23920 0 -1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_53_255
timestamp 1679235063
transform 1 0 24564 0 -1 31552
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_53_259
timestamp 1679235063
transform 1 0 24932 0 -1 31552
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_53_264
timestamp 1679235063
transform 1 0 25392 0 -1 31552
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_54_3
timestamp 1679235063
transform 1 0 1380 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_15
timestamp 1679235063
transform 1 0 2484 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_54_27
timestamp 1679235063
transform 1 0 3588 0 1 31552
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_54_29
timestamp 1679235063
transform 1 0 3772 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_41
timestamp 1679235063
transform 1 0 4876 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_54_53
timestamp 1679235063
transform 1 0 5980 0 1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_54_76
timestamp 1679235063
transform 1 0 8096 0 1 31552
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_54_82
timestamp 1679235063
transform 1 0 8648 0 1 31552
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_54_85
timestamp 1679235063
transform 1 0 8924 0 1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_54_111
timestamp 1679235063
transform 1 0 11316 0 1 31552
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_54_117
timestamp 1679235063
transform 1 0 11868 0 1 31552
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_54_128
timestamp 1679235063
transform 1 0 12880 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_141
timestamp 1679235063
transform 1 0 14076 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_54_153
timestamp 1679235063
transform 1 0 15180 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_54_174
timestamp 1679235063
transform 1 0 17112 0 1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_54_187
timestamp 1679235063
transform 1 0 18308 0 1 31552
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_54_195
timestamp 1679235063
transform 1 0 19044 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_54_201
timestamp 1679235063
transform 1 0 19596 0 1 31552
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_54_212
timestamp 1679235063
transform 1 0 20608 0 1 31552
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_54_218
timestamp 1679235063
transform 1 0 21160 0 1 31552
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_54_226
timestamp 1679235063
transform 1 0 21896 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_54_236
timestamp 1679235063
transform 1 0 22816 0 1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_54_250
timestamp 1679235063
transform 1 0 24104 0 1 31552
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_54_253
timestamp 1679235063
transform 1 0 24380 0 1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_54_259
timestamp 1679235063
transform 1 0 24932 0 1 31552
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_54_264
timestamp 1679235063
transform 1 0 25392 0 1 31552
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_55_3
timestamp 1679235063
transform 1 0 1380 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_15
timestamp 1679235063
transform 1 0 2484 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_27
timestamp 1679235063
transform 1 0 3588 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_55_39
timestamp 1679235063
transform 1 0 4692 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_55_42
timestamp 1679235063
transform 1 0 4968 0 -1 32640
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_55_53
timestamp 1679235063
transform 1 0 5980 0 -1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_55_57
timestamp 1679235063
transform 1 0 6348 0 -1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_55_63
timestamp 1679235063
transform 1 0 6900 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_55_67
timestamp 1679235063
transform 1 0 7268 0 -1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_55_92
timestamp 1679235063
transform 1 0 9568 0 -1 32640
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_55_96
timestamp 1679235063
transform 1 0 9936 0 -1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_55_107
timestamp 1679235063
transform 1 0 10948 0 -1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_55_111
timestamp 1679235063
transform 1 0 11316 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_55_113
timestamp 1679235063
transform 1 0 11500 0 -1 32640
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_55_118
timestamp 1679235063
transform 1 0 11960 0 -1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_55_127
timestamp 1679235063
transform 1 0 12788 0 -1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_55_135
timestamp 1679235063
transform 1 0 13524 0 -1 32640
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_55_146
timestamp 1679235063
transform 1 0 14536 0 -1 32640
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_55_154
timestamp 1679235063
transform 1 0 15272 0 -1 32640
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_55_164
timestamp 1679235063
transform 1 0 16192 0 -1 32640
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_55_171
timestamp 1679235063
transform 1 0 16836 0 -1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_55_186
timestamp 1679235063
transform 1 0 18216 0 -1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_55_199
timestamp 1679235063
transform 1 0 19412 0 -1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_55_212
timestamp 1679235063
transform 1 0 20608 0 -1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_55_219
timestamp 1679235063
transform 1 0 21252 0 -1 32640
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_55_223
timestamp 1679235063
transform 1 0 21620 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_55_225
timestamp 1679235063
transform 1 0 21804 0 -1 32640
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_55_230
timestamp 1679235063
transform 1 0 22264 0 -1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_55_237
timestamp 1679235063
transform 1 0 22908 0 -1 32640
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_55_244
timestamp 1679235063
transform 1 0 23552 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_55_256
timestamp 1679235063
transform 1 0 24656 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_55_259
timestamp 1679235063
transform 1 0 24932 0 -1 32640
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_55_264
timestamp 1679235063
transform 1 0 25392 0 -1 32640
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_56_3
timestamp 1679235063
transform 1 0 1380 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_15
timestamp 1679235063
transform 1 0 2484 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_56_27
timestamp 1679235063
transform 1 0 3588 0 1 32640
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_56_29
timestamp 1679235063
transform 1 0 3772 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_56_41
timestamp 1679235063
transform 1 0 4876 0 1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_56_45
timestamp 1679235063
transform 1 0 5244 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_56_66
timestamp 1679235063
transform 1 0 7176 0 1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_56_79
timestamp 1679235063
transform 1 0 8372 0 1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_56_83
timestamp 1679235063
transform 1 0 8740 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_56_85
timestamp 1679235063
transform 1 0 8924 0 1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_56_89
timestamp 1679235063
transform 1 0 9292 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_56_99
timestamp 1679235063
transform 1 0 10212 0 1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_56_104
timestamp 1679235063
transform 1 0 10672 0 1 32640
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_56_115
timestamp 1679235063
transform 1 0 11684 0 1 32640
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_56_119
timestamp 1679235063
transform 1 0 12052 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_56_131
timestamp 1679235063
transform 1 0 13156 0 1 32640
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_56_139
timestamp 1679235063
transform 1 0 13892 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_56_141
timestamp 1679235063
transform 1 0 14076 0 1 32640
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_56_152
timestamp 1679235063
transform 1 0 15088 0 1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_56_164
timestamp 1679235063
transform 1 0 16192 0 1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_56_177
timestamp 1679235063
transform 1 0 17388 0 1 32640
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_56_181
timestamp 1679235063
transform 1 0 17756 0 1 32640
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_56_189
timestamp 1679235063
transform 1 0 18492 0 1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_56_197
timestamp 1679235063
transform 1 0 19228 0 1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_56_209
timestamp 1679235063
transform 1 0 20332 0 1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_56_213
timestamp 1679235063
transform 1 0 20700 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_56_223
timestamp 1679235063
transform 1 0 21620 0 1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_56_236
timestamp 1679235063
transform 1 0 22816 0 1 32640
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_56_246
timestamp 1679235063
transform 1 0 23736 0 1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_56_253
timestamp 1679235063
transform 1 0 24380 0 1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_56_259
timestamp 1679235063
transform 1 0 24932 0 1 32640
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_56_264
timestamp 1679235063
transform 1 0 25392 0 1 32640
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_57_3
timestamp 1679235063
transform 1 0 1380 0 -1 33728
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_57_8
timestamp 1679235063
transform 1 0 1840 0 -1 33728
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_57_12
timestamp 1679235063
transform 1 0 2208 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_24
timestamp 1679235063
transform 1 0 3312 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_36
timestamp 1679235063
transform 1 0 4416 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_57_48
timestamp 1679235063
transform 1 0 5520 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_57_52
timestamp 1679235063
transform 1 0 5888 0 -1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_57_57
timestamp 1679235063
transform 1 0 6348 0 -1 33728
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_57_65
timestamp 1679235063
transform 1 0 7084 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_57_68
timestamp 1679235063
transform 1 0 7360 0 -1 33728
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_57_78
timestamp 1679235063
transform 1 0 8280 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_57_90
timestamp 1679235063
transform 1 0 9384 0 -1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_57_97
timestamp 1679235063
transform 1 0 10028 0 -1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_57_101
timestamp 1679235063
transform 1 0 10396 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_57_104
timestamp 1679235063
transform 1 0 10672 0 -1 33728
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_57_113
timestamp 1679235063
transform 1 0 11500 0 -1 33728
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_57_121
timestamp 1679235063
transform 1 0 12236 0 -1 33728
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_57_136
timestamp 1679235063
transform 1 0 13616 0 -1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_57_160
timestamp 1679235063
transform 1 0 15824 0 -1 33728
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_57_164
timestamp 1679235063
transform 1 0 16192 0 -1 33728
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_57_169
timestamp 1679235063
transform 1 0 16652 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_57_181
timestamp 1679235063
transform 1 0 17756 0 -1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_57_207
timestamp 1679235063
transform 1 0 20148 0 -1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_57_220
timestamp 1679235063
transform 1 0 21344 0 -1 33728
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_57_225
timestamp 1679235063
transform 1 0 21804 0 -1 33728
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_57_236
timestamp 1679235063
transform 1 0 22816 0 -1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_57_242
timestamp 1679235063
transform 1 0 23368 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_57_264
timestamp 1679235063
transform 1 0 25392 0 -1 33728
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_58_3
timestamp 1679235063
transform 1 0 1380 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_15
timestamp 1679235063
transform 1 0 2484 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_58_27
timestamp 1679235063
transform 1 0 3588 0 1 33728
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_58_29
timestamp 1679235063
transform 1 0 3772 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_58_41
timestamp 1679235063
transform 1 0 4876 0 1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_58_47
timestamp 1679235063
transform 1 0 5428 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_58_69
timestamp 1679235063
transform 1 0 7452 0 1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_58_82
timestamp 1679235063
transform 1 0 8648 0 1 33728
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_58_85
timestamp 1679235063
transform 1 0 8924 0 1 33728
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_58_95
timestamp 1679235063
transform 1 0 9844 0 1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_58_108
timestamp 1679235063
transform 1 0 11040 0 1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_58_132
timestamp 1679235063
transform 1 0 13248 0 1 33728
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_58_136
timestamp 1679235063
transform 1 0 13616 0 1 33728
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_58_141
timestamp 1679235063
transform 1 0 14076 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_58_153
timestamp 1679235063
transform 1 0 15180 0 1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_58_157
timestamp 1679235063
transform 1 0 15548 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_58_178
timestamp 1679235063
transform 1 0 17480 0 1 33728
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_58_182
timestamp 1679235063
transform 1 0 17848 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_58_194
timestamp 1679235063
transform 1 0 18952 0 1 33728
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_58_197
timestamp 1679235063
transform 1 0 19228 0 1 33728
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_58_201
timestamp 1679235063
transform 1 0 19596 0 1 33728
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_58_211
timestamp 1679235063
transform 1 0 20516 0 1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_58_223
timestamp 1679235063
transform 1 0 21620 0 1 33728
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_58_227
timestamp 1679235063
transform 1 0 21988 0 1 33728
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_58_240
timestamp 1679235063
transform 1 0 23184 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_58_253
timestamp 1679235063
transform 1 0 24380 0 1 33728
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_58_258
timestamp 1679235063
transform 1 0 24840 0 1 33728
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_59_3
timestamp 1679235063
transform 1 0 1380 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_15
timestamp 1679235063
transform 1 0 2484 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_27
timestamp 1679235063
transform 1 0 3588 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_39
timestamp 1679235063
transform 1 0 4692 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_59_51
timestamp 1679235063
transform 1 0 5796 0 -1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_59_55
timestamp 1679235063
transform 1 0 6164 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_59_57
timestamp 1679235063
transform 1 0 6348 0 -1 34816
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_59_65
timestamp 1679235063
transform 1 0 7084 0 -1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_59_70
timestamp 1679235063
transform 1 0 7544 0 -1 34816
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_59_92
timestamp 1679235063
transform 1 0 9568 0 -1 34816
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_59_96
timestamp 1679235063
transform 1 0 9936 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_59_108
timestamp 1679235063
transform 1 0 11040 0 -1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_59_113
timestamp 1679235063
transform 1 0 11500 0 -1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_59_124
timestamp 1679235063
transform 1 0 12512 0 -1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_59_139
timestamp 1679235063
transform 1 0 13892 0 -1 34816
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_59_143
timestamp 1679235063
transform 1 0 14260 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_59_155
timestamp 1679235063
transform 1 0 15364 0 -1 34816
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_59_166
timestamp 1679235063
transform 1 0 16376 0 -1 34816
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_59_169
timestamp 1679235063
transform 1 0 16652 0 -1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_59_175
timestamp 1679235063
transform 1 0 17204 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_59_184
timestamp 1679235063
transform 1 0 18032 0 -1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_59_197
timestamp 1679235063
transform 1 0 19228 0 -1 34816
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_59_201
timestamp 1679235063
transform 1 0 19596 0 -1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_59_208
timestamp 1679235063
transform 1 0 20240 0 -1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_59_221
timestamp 1679235063
transform 1 0 21436 0 -1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_59_225
timestamp 1679235063
transform 1 0 21804 0 -1 34816
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_59_236
timestamp 1679235063
transform 1 0 22816 0 -1 34816
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_59_240
timestamp 1679235063
transform 1 0 23184 0 -1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_59_249
timestamp 1679235063
transform 1 0 24012 0 -1 34816
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_59_253
timestamp 1679235063
transform 1 0 24380 0 -1 34816
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_59_264
timestamp 1679235063
transform 1 0 25392 0 -1 34816
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_60_3
timestamp 1679235063
transform 1 0 1380 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_15
timestamp 1679235063
transform 1 0 2484 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_60_27
timestamp 1679235063
transform 1 0 3588 0 1 34816
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_60_29
timestamp 1679235063
transform 1 0 3772 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_60_41
timestamp 1679235063
transform 1 0 4876 0 1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_60_52
timestamp 1679235063
transform 1 0 5888 0 1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_60_76
timestamp 1679235063
transform 1 0 8096 0 1 34816
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_60_80
timestamp 1679235063
transform 1 0 8464 0 1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_60_85
timestamp 1679235063
transform 1 0 8924 0 1 34816
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_60_96
timestamp 1679235063
transform 1 0 9936 0 1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_60_120
timestamp 1679235063
transform 1 0 12144 0 1 34816
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_60_124
timestamp 1679235063
transform 1 0 12512 0 1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_60_136
timestamp 1679235063
transform 1 0 13616 0 1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_60_141
timestamp 1679235063
transform 1 0 14076 0 1 34816
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_60_151
timestamp 1679235063
transform 1 0 14996 0 1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_60_155
timestamp 1679235063
transform 1 0 15364 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_60_176
timestamp 1679235063
transform 1 0 17296 0 1 34816
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_60_180
timestamp 1679235063
transform 1 0 17664 0 1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_60_194
timestamp 1679235063
transform 1 0 18952 0 1 34816
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_60_197
timestamp 1679235063
transform 1 0 19228 0 1 34816
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_60_219
timestamp 1679235063
transform 1 0 21252 0 1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_60_226
timestamp 1679235063
transform 1 0 21896 0 1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_60_250
timestamp 1679235063
transform 1 0 24104 0 1 34816
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_60_253
timestamp 1679235063
transform 1 0 24380 0 1 34816
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_60_263
timestamp 1679235063
transform 1 0 25300 0 1 34816
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_61_3
timestamp 1679235063
transform 1 0 1380 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_15
timestamp 1679235063
transform 1 0 2484 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_61_27
timestamp 1679235063
transform 1 0 3588 0 -1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_61_33
timestamp 1679235063
transform 1 0 4140 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_61_54
timestamp 1679235063
transform 1 0 6072 0 -1 35904
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_61_59
timestamp 1679235063
transform 1 0 6532 0 -1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_61_63
timestamp 1679235063
transform 1 0 6900 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_61_72
timestamp 1679235063
transform 1 0 7728 0 -1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_61_96
timestamp 1679235063
transform 1 0 9936 0 -1 35904
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_61_100
timestamp 1679235063
transform 1 0 10304 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_61_113
timestamp 1679235063
transform 1 0 11500 0 -1 35904
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_61_135
timestamp 1679235063
transform 1 0 13524 0 -1 35904
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_61_139
timestamp 1679235063
transform 1 0 13892 0 -1 35904
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_61_143
timestamp 1679235063
transform 1 0 14260 0 -1 35904
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_61_154
timestamp 1679235063
transform 1 0 15272 0 -1 35904
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_61_158
timestamp 1679235063
transform 1 0 15640 0 -1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_61_164
timestamp 1679235063
transform 1 0 16192 0 -1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_61_169
timestamp 1679235063
transform 1 0 16652 0 -1 35904
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_61_177
timestamp 1679235063
transform 1 0 17388 0 -1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_61_200
timestamp 1679235063
transform 1 0 19504 0 -1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_61_213
timestamp 1679235063
transform 1 0 20700 0 -1 35904
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_61_217
timestamp 1679235063
transform 1 0 21068 0 -1 35904
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_61_221
timestamp 1679235063
transform 1 0 21436 0 -1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_61_225
timestamp 1679235063
transform 1 0 21804 0 -1 35904
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_61_236
timestamp 1679235063
transform 1 0 22816 0 -1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_61_261
timestamp 1679235063
transform 1 0 25116 0 -1 35904
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_61_265
timestamp 1679235063
transform 1 0 25484 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_62_3
timestamp 1679235063
transform 1 0 1380 0 1 35904
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_62_8
timestamp 1679235063
transform 1 0 1840 0 1 35904
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_62_12
timestamp 1679235063
transform 1 0 2208 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_62_24
timestamp 1679235063
transform 1 0 3312 0 1 35904
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_62_29
timestamp 1679235063
transform 1 0 3772 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_62_41
timestamp 1679235063
transform 1 0 4876 0 1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_62_65
timestamp 1679235063
transform 1 0 7084 0 1 35904
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_62_69
timestamp 1679235063
transform 1 0 7452 0 1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_62_81
timestamp 1679235063
transform 1 0 8556 0 1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_62_85
timestamp 1679235063
transform 1 0 8924 0 1 35904
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_62_96
timestamp 1679235063
transform 1 0 9936 0 1 35904
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_62_104
timestamp 1679235063
transform 1 0 10672 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_62_111
timestamp 1679235063
transform 1 0 11316 0 1 35904
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_62_124
timestamp 1679235063
transform 1 0 12512 0 1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_62_137
timestamp 1679235063
transform 1 0 13708 0 1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_62_141
timestamp 1679235063
transform 1 0 14076 0 1 35904
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_62_152
timestamp 1679235063
transform 1 0 15088 0 1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_62_159
timestamp 1679235063
transform 1 0 15732 0 1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_62_163
timestamp 1679235063
transform 1 0 16100 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_62_173
timestamp 1679235063
transform 1 0 17020 0 1 35904
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_62_180
timestamp 1679235063
transform 1 0 17664 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_62_192
timestamp 1679235063
transform 1 0 18768 0 1 35904
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_62_197
timestamp 1679235063
transform 1 0 19228 0 1 35904
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_62_208
timestamp 1679235063
transform 1 0 20240 0 1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_62_214
timestamp 1679235063
transform 1 0 20792 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_62_224
timestamp 1679235063
transform 1 0 21712 0 1 35904
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_62_232
timestamp 1679235063
transform 1 0 22448 0 1 35904
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_62_237
timestamp 1679235063
transform 1 0 22908 0 1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_62_250
timestamp 1679235063
transform 1 0 24104 0 1 35904
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_62_259
timestamp 1679235063
transform 1 0 24932 0 1 35904
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_62_264
timestamp 1679235063
transform 1 0 25392 0 1 35904
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_63_3
timestamp 1679235063
transform 1 0 1380 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_63_15
timestamp 1679235063
transform 1 0 2484 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_63_27
timestamp 1679235063
transform 1 0 3588 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_63_39
timestamp 1679235063
transform 1 0 4692 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_63_51
timestamp 1679235063
transform 1 0 5796 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_63_55
timestamp 1679235063
transform 1 0 6164 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_63_57
timestamp 1679235063
transform 1 0 6348 0 -1 36992
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_63_69
timestamp 1679235063
transform 1 0 7452 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_63_81
timestamp 1679235063
transform 1 0 8556 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_63_84
timestamp 1679235063
transform 1 0 8832 0 -1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_63_98
timestamp 1679235063
transform 1 0 10120 0 -1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_63_102
timestamp 1679235063
transform 1 0 10488 0 -1 36992
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_63_110
timestamp 1679235063
transform 1 0 11224 0 -1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_63_115
timestamp 1679235063
transform 1 0 11684 0 -1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_63_125
timestamp 1679235063
transform 1 0 12604 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_63_138
timestamp 1679235063
transform 1 0 13800 0 -1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_63_143
timestamp 1679235063
transform 1 0 14260 0 -1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_63_154
timestamp 1679235063
transform 1 0 15272 0 -1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_63_158
timestamp 1679235063
transform 1 0 15640 0 -1 36992
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_63_166
timestamp 1679235063
transform 1 0 16376 0 -1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_63_171
timestamp 1679235063
transform 1 0 16836 0 -1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_63_182
timestamp 1679235063
transform 1 0 17848 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_63_194
timestamp 1679235063
transform 1 0 18952 0 -1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_63_200
timestamp 1679235063
transform 1 0 19504 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_63_203
timestamp 1679235063
transform 1 0 19780 0 -1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_63_214
timestamp 1679235063
transform 1 0 20792 0 -1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_63_218
timestamp 1679235063
transform 1 0 21160 0 -1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_63_227
timestamp 1679235063
transform 1 0 21988 0 -1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_63_232
timestamp 1679235063
transform 1 0 22448 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_63_256
timestamp 1679235063
transform 1 0 24656 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_63_260
timestamp 1679235063
transform 1 0 25024 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_63_264
timestamp 1679235063
transform 1 0 25392 0 -1 36992
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_64_3
timestamp 1679235063
transform 1 0 1380 0 1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_64_15
timestamp 1679235063
transform 1 0 2484 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_64_27
timestamp 1679235063
transform 1 0 3588 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_64_29
timestamp 1679235063
transform 1 0 3772 0 1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_64_52
timestamp 1679235063
transform 1 0 5888 0 1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_64_56
timestamp 1679235063
transform 1 0 6256 0 1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_64_82
timestamp 1679235063
transform 1 0 8648 0 1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_64_85
timestamp 1679235063
transform 1 0 8924 0 1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_64_90
timestamp 1679235063
transform 1 0 9384 0 1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_64_94
timestamp 1679235063
transform 1 0 9752 0 1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_64_105
timestamp 1679235063
transform 1 0 10764 0 1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_64_109
timestamp 1679235063
transform 1 0 11132 0 1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_64_120
timestamp 1679235063
transform 1 0 12144 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_64_133
timestamp 1679235063
transform 1 0 13340 0 1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_64_137
timestamp 1679235063
transform 1 0 13708 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_64_141
timestamp 1679235063
transform 1 0 14076 0 1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_64_146
timestamp 1679235063
transform 1 0 14536 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_64_159
timestamp 1679235063
transform 1 0 15732 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_64_172
timestamp 1679235063
transform 1 0 16928 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_64_185
timestamp 1679235063
transform 1 0 18124 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_64_192
timestamp 1679235063
transform 1 0 18768 0 1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_64_199
timestamp 1679235063
transform 1 0 19412 0 1 36992
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_64_216
timestamp 1679235063
transform 1 0 20976 0 1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_64_220
timestamp 1679235063
transform 1 0 21344 0 1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_64_231
timestamp 1679235063
transform 1 0 22356 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_64_238
timestamp 1679235063
transform 1 0 23000 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_64_250
timestamp 1679235063
transform 1 0 24104 0 1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_64_253
timestamp 1679235063
transform 1 0 24380 0 1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_64_263
timestamp 1679235063
transform 1 0 25300 0 1 36992
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_65_3
timestamp 1679235063
transform 1 0 1380 0 -1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_65_15
timestamp 1679235063
transform 1 0 2484 0 -1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_65_27
timestamp 1679235063
transform 1 0 3588 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_65_39
timestamp 1679235063
transform 1 0 4692 0 -1 38080
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_65_45
timestamp 1679235063
transform 1 0 5244 0 -1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_65_54
timestamp 1679235063
transform 1 0 6072 0 -1 38080
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_65_57
timestamp 1679235063
transform 1 0 6348 0 -1 38080
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_65_82
timestamp 1679235063
transform 1 0 8648 0 -1 38080
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_65_88
timestamp 1679235063
transform 1 0 9200 0 -1 38080
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_65_99
timestamp 1679235063
transform 1 0 10212 0 -1 38080
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_65_105
timestamp 1679235063
transform 1 0 10764 0 -1 38080
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_65_109
timestamp 1679235063
transform 1 0 11132 0 -1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_65_113
timestamp 1679235063
transform 1 0 11500 0 -1 38080
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_65_118
timestamp 1679235063
transform 1 0 11960 0 -1 38080
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_65_122
timestamp 1679235063
transform 1 0 12328 0 -1 38080
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_65_133
timestamp 1679235063
transform 1 0 13340 0 -1 38080
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_65_141
timestamp 1679235063
transform 1 0 14076 0 -1 38080
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_65_145
timestamp 1679235063
transform 1 0 14444 0 -1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_65_148
timestamp 1679235063
transform 1 0 14720 0 -1 38080
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_65_160
timestamp 1679235063
transform 1 0 15824 0 -1 38080
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_65_169
timestamp 1679235063
transform 1 0 16652 0 -1 38080
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_65_174
timestamp 1679235063
transform 1 0 17112 0 -1 38080
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_65_180
timestamp 1679235063
transform 1 0 17664 0 -1 38080
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_65_192
timestamp 1679235063
transform 1 0 18768 0 -1 38080
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_65_205
timestamp 1679235063
transform 1 0 19964 0 -1 38080
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_65_209
timestamp 1679235063
transform 1 0 20332 0 -1 38080
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_65_221
timestamp 1679235063
transform 1 0 21436 0 -1 38080
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_65_225
timestamp 1679235063
transform 1 0 21804 0 -1 38080
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_65_236
timestamp 1679235063
transform 1 0 22816 0 -1 38080
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_65_242
timestamp 1679235063
transform 1 0 23368 0 -1 38080
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_65_264
timestamp 1679235063
transform 1 0 25392 0 -1 38080
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_66_3
timestamp 1679235063
transform 1 0 1380 0 1 38080
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_66_8
timestamp 1679235063
transform 1 0 1840 0 1 38080
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_66_12
timestamp 1679235063
transform 1 0 2208 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_66_24
timestamp 1679235063
transform 1 0 3312 0 1 38080
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_66_29
timestamp 1679235063
transform 1 0 3772 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_66_41
timestamp 1679235063
transform 1 0 4876 0 1 38080
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_66_67
timestamp 1679235063
transform 1 0 7268 0 1 38080
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_66_80
timestamp 1679235063
transform 1 0 8464 0 1 38080
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_66_85
timestamp 1679235063
transform 1 0 8924 0 1 38080
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_66_97
timestamp 1679235063
transform 1 0 10028 0 1 38080
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_66_110
timestamp 1679235063
transform 1 0 11224 0 1 38080
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_66_138
timestamp 1679235063
transform 1 0 13800 0 1 38080
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_66_141
timestamp 1679235063
transform 1 0 14076 0 1 38080
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_66_146
timestamp 1679235063
transform 1 0 14536 0 1 38080
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_66_154
timestamp 1679235063
transform 1 0 15272 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_66_158
timestamp 1679235063
transform 1 0 15640 0 1 38080
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_66_162
timestamp 1679235063
transform 1 0 16008 0 1 38080
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_66_173
timestamp 1679235063
transform 1 0 17020 0 1 38080
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_66_186
timestamp 1679235063
transform 1 0 18216 0 1 38080
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_66_197
timestamp 1679235063
transform 1 0 19228 0 1 38080
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_66_210
timestamp 1679235063
transform 1 0 20424 0 1 38080
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_66_218
timestamp 1679235063
transform 1 0 21160 0 1 38080
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_66_231
timestamp 1679235063
transform 1 0 22356 0 1 38080
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_66_244
timestamp 1679235063
transform 1 0 23552 0 1 38080
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_66_253
timestamp 1679235063
transform 1 0 24380 0 1 38080
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_66_264
timestamp 1679235063
transform 1 0 25392 0 1 38080
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_67_3
timestamp 1679235063
transform 1 0 1380 0 -1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_67_15
timestamp 1679235063
transform 1 0 2484 0 -1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_67_27
timestamp 1679235063
transform 1 0 3588 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_67_39
timestamp 1679235063
transform 1 0 4692 0 -1 39168
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_67_45
timestamp 1679235063
transform 1 0 5244 0 -1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_67_54
timestamp 1679235063
transform 1 0 6072 0 -1 39168
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_67_57
timestamp 1679235063
transform 1 0 6348 0 -1 39168
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_67_68
timestamp 1679235063
transform 1 0 7360 0 -1 39168
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_67_80
timestamp 1679235063
transform 1 0 8464 0 -1 39168
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_67_85
timestamp 1679235063
transform 1 0 8924 0 -1 39168
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_67_96
timestamp 1679235063
transform 1 0 9936 0 -1 39168
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_67_100
timestamp 1679235063
transform 1 0 10304 0 -1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_67_110
timestamp 1679235063
transform 1 0 11224 0 -1 39168
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_67_113
timestamp 1679235063
transform 1 0 11500 0 -1 39168
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_67_130
timestamp 1679235063
transform 1 0 13064 0 -1 39168
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_67_142
timestamp 1679235063
transform 1 0 14168 0 -1 39168
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_67_159
timestamp 1679235063
transform 1 0 15732 0 -1 39168
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_67_163
timestamp 1679235063
transform 1 0 16100 0 -1 39168
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_67_167
timestamp 1679235063
transform 1 0 16468 0 -1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_67_169
timestamp 1679235063
transform 1 0 16652 0 -1 39168
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_67_191
timestamp 1679235063
transform 1 0 18676 0 -1 39168
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_67_195
timestamp 1679235063
transform 1 0 19044 0 -1 39168
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_67_208
timestamp 1679235063
transform 1 0 20240 0 -1 39168
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_67_221
timestamp 1679235063
transform 1 0 21436 0 -1 39168
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_67_229
timestamp 1679235063
transform 1 0 22172 0 -1 39168
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_67_251
timestamp 1679235063
transform 1 0 24196 0 -1 39168
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_67_263
timestamp 1679235063
transform 1 0 25300 0 -1 39168
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_68_3
timestamp 1679235063
transform 1 0 1380 0 1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_68_15
timestamp 1679235063
transform 1 0 2484 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_68_27
timestamp 1679235063
transform 1 0 3588 0 1 39168
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_68_29
timestamp 1679235063
transform 1 0 3772 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_68_41
timestamp 1679235063
transform 1 0 4876 0 1 39168
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_68_64
timestamp 1679235063
transform 1 0 6992 0 1 39168
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_68_68
timestamp 1679235063
transform 1 0 7360 0 1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_68_77
timestamp 1679235063
transform 1 0 8188 0 1 39168
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_68_83
timestamp 1679235063
transform 1 0 8740 0 1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_68_85
timestamp 1679235063
transform 1 0 8924 0 1 39168
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_68_90
timestamp 1679235063
transform 1 0 9384 0 1 39168
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_68_103
timestamp 1679235063
transform 1 0 10580 0 1 39168
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_68_127
timestamp 1679235063
transform 1 0 12788 0 1 39168
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_68_136
timestamp 1679235063
transform 1 0 13616 0 1 39168
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_68_143
timestamp 1679235063
transform 1 0 14260 0 1 39168
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_68_154
timestamp 1679235063
transform 1 0 15272 0 1 39168
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_68_167
timestamp 1679235063
transform 1 0 16468 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_68_179
timestamp 1679235063
transform 1 0 17572 0 1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_68_188
timestamp 1679235063
transform 1 0 18400 0 1 39168
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_68_197
timestamp 1679235063
transform 1 0 19228 0 1 39168
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_68_208
timestamp 1679235063
transform 1 0 20240 0 1 39168
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_68_212
timestamp 1679235063
transform 1 0 20608 0 1 39168
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_68_229
timestamp 1679235063
transform 1 0 22172 0 1 39168
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_68_242
timestamp 1679235063
transform 1 0 23368 0 1 39168
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_68_249
timestamp 1679235063
transform 1 0 24012 0 1 39168
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_68_253
timestamp 1679235063
transform 1 0 24380 0 1 39168
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_68_264
timestamp 1679235063
transform 1 0 25392 0 1 39168
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_69_3
timestamp 1679235063
transform 1 0 1380 0 -1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_69_15
timestamp 1679235063
transform 1 0 2484 0 -1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_69_27
timestamp 1679235063
transform 1 0 3588 0 -1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_69_39
timestamp 1679235063
transform 1 0 4692 0 -1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_69_51
timestamp 1679235063
transform 1 0 5796 0 -1 40256
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_69_55
timestamp 1679235063
transform 1 0 6164 0 -1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_69_57
timestamp 1679235063
transform 1 0 6348 0 -1 40256
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_69_61
timestamp 1679235063
transform 1 0 6716 0 -1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_69_65
timestamp 1679235063
transform 1 0 7084 0 -1 40256
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_69_78
timestamp 1679235063
transform 1 0 8280 0 -1 40256
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_69_105
timestamp 1679235063
transform 1 0 10764 0 -1 40256
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_69_113
timestamp 1679235063
transform 1 0 11500 0 -1 40256
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_69_124
timestamp 1679235063
transform 1 0 12512 0 -1 40256
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_69_128
timestamp 1679235063
transform 1 0 12880 0 -1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_69_149
timestamp 1679235063
transform 1 0 14812 0 -1 40256
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_69_153
timestamp 1679235063
transform 1 0 15180 0 -1 40256
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_69_166
timestamp 1679235063
transform 1 0 16376 0 -1 40256
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_69_169
timestamp 1679235063
transform 1 0 16652 0 -1 40256
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_69_179
timestamp 1679235063
transform 1 0 17572 0 -1 40256
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_69_185
timestamp 1679235063
transform 1 0 18124 0 -1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_69_195
timestamp 1679235063
transform 1 0 19044 0 -1 40256
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_69_208
timestamp 1679235063
transform 1 0 20240 0 -1 40256
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_69_221
timestamp 1679235063
transform 1 0 21436 0 -1 40256
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_69_233
timestamp 1679235063
transform 1 0 22540 0 -1 40256
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_69_240
timestamp 1679235063
transform 1 0 23184 0 -1 40256
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_69_263
timestamp 1679235063
transform 1 0 25300 0 -1 40256
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_70_3
timestamp 1679235063
transform 1 0 1380 0 1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_70_15
timestamp 1679235063
transform 1 0 2484 0 1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_70_27
timestamp 1679235063
transform 1 0 3588 0 1 40256
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_70_29
timestamp 1679235063
transform 1 0 3772 0 1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_70_41
timestamp 1679235063
transform 1 0 4876 0 1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_70_53
timestamp 1679235063
transform 1 0 5980 0 1 40256
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_70_57
timestamp 1679235063
transform 1 0 6348 0 1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_70_78
timestamp 1679235063
transform 1 0 8280 0 1 40256
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_70_85
timestamp 1679235063
transform 1 0 8924 0 1 40256
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_70_98
timestamp 1679235063
transform 1 0 10120 0 1 40256
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_70_102
timestamp 1679235063
transform 1 0 10488 0 1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_70_107
timestamp 1679235063
transform 1 0 10948 0 1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_70_110
timestamp 1679235063
transform 1 0 11224 0 1 40256
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_70_121
timestamp 1679235063
transform 1 0 12236 0 1 40256
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_70_134
timestamp 1679235063
transform 1 0 13432 0 1 40256
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_70_138
timestamp 1679235063
transform 1 0 13800 0 1 40256
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_70_141
timestamp 1679235063
transform 1 0 14076 0 1 40256
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_70_152
timestamp 1679235063
transform 1 0 15088 0 1 40256
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_70_164
timestamp 1679235063
transform 1 0 16192 0 1 40256
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_70_179
timestamp 1679235063
transform 1 0 17572 0 1 40256
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_70_191
timestamp 1679235063
transform 1 0 18676 0 1 40256
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_70_195
timestamp 1679235063
transform 1 0 19044 0 1 40256
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_70_197
timestamp 1679235063
transform 1 0 19228 0 1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_70_209
timestamp 1679235063
transform 1 0 20332 0 1 40256
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_70_224
timestamp 1679235063
transform 1 0 21712 0 1 40256
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_70_230
timestamp 1679235063
transform 1 0 22264 0 1 40256
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_70_241
timestamp 1679235063
transform 1 0 23276 0 1 40256
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_70_245
timestamp 1679235063
transform 1 0 23644 0 1 40256
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_70_250
timestamp 1679235063
transform 1 0 24104 0 1 40256
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_70_253
timestamp 1679235063
transform 1 0 24380 0 1 40256
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_70_263
timestamp 1679235063
transform 1 0 25300 0 1 40256
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_71_3
timestamp 1679235063
transform 1 0 1380 0 -1 41344
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_71_8
timestamp 1679235063
transform 1 0 1840 0 -1 41344
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_71_12
timestamp 1679235063
transform 1 0 2208 0 -1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_71_24
timestamp 1679235063
transform 1 0 3312 0 -1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_71_29
timestamp 1679235063
transform 1 0 3772 0 -1 41344
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_71_33
timestamp 1679235063
transform 1 0 4140 0 -1 41344
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_71_41
timestamp 1679235063
transform 1 0 4876 0 -1 41344
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_71_45
timestamp 1679235063
transform 1 0 5244 0 -1 41344
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_71_53
timestamp 1679235063
transform 1 0 5980 0 -1 41344
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_71_57
timestamp 1679235063
transform 1 0 6348 0 -1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_71_69
timestamp 1679235063
transform 1 0 7452 0 -1 41344
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_71_73
timestamp 1679235063
transform 1 0 7820 0 -1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_71_82
timestamp 1679235063
transform 1 0 8648 0 -1 41344
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_71_106
timestamp 1679235063
transform 1 0 10856 0 -1 41344
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_71_113
timestamp 1679235063
transform 1 0 11500 0 -1 41344
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_71_126
timestamp 1679235063
transform 1 0 12696 0 -1 41344
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_71_132
timestamp 1679235063
transform 1 0 13248 0 -1 41344
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_71_158
timestamp 1679235063
transform 1 0 15640 0 -1 41344
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_71_164
timestamp 1679235063
transform 1 0 16192 0 -1 41344
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_71_169
timestamp 1679235063
transform 1 0 16652 0 -1 41344
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_71_192
timestamp 1679235063
transform 1 0 18768 0 -1 41344
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_71_196
timestamp 1679235063
transform 1 0 19136 0 -1 41344
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_71_207
timestamp 1679235063
transform 1 0 20148 0 -1 41344
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_71_211
timestamp 1679235063
transform 1 0 20516 0 -1 41344
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_71_222
timestamp 1679235063
transform 1 0 21528 0 -1 41344
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_71_225
timestamp 1679235063
transform 1 0 21804 0 -1 41344
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_71_230
timestamp 1679235063
transform 1 0 22264 0 -1 41344
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_71_234
timestamp 1679235063
transform 1 0 22632 0 -1 41344
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_71_256
timestamp 1679235063
transform 1 0 24656 0 -1 41344
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_71_260
timestamp 1679235063
transform 1 0 25024 0 -1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_71_264
timestamp 1679235063
transform 1 0 25392 0 -1 41344
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_72_3
timestamp 1679235063
transform 1 0 1380 0 1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_72_15
timestamp 1679235063
transform 1 0 2484 0 1 41344
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_72_23
timestamp 1679235063
transform 1 0 3220 0 1 41344
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_72_29
timestamp 1679235063
transform 1 0 3772 0 1 41344
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_72_35
timestamp 1679235063
transform 1 0 4324 0 1 41344
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_72_43
timestamp 1679235063
transform 1 0 5060 0 1 41344
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_72_47
timestamp 1679235063
transform 1 0 5428 0 1 41344
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_72_73
timestamp 1679235063
transform 1 0 7820 0 1 41344
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_72_79
timestamp 1679235063
transform 1 0 8372 0 1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_72_85
timestamp 1679235063
transform 1 0 8924 0 1 41344
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_72_96
timestamp 1679235063
transform 1 0 9936 0 1 41344
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_72_109
timestamp 1679235063
transform 1 0 11132 0 1 41344
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_72_122
timestamp 1679235063
transform 1 0 12328 0 1 41344
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_72_134
timestamp 1679235063
transform 1 0 13432 0 1 41344
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_72_141
timestamp 1679235063
transform 1 0 14076 0 1 41344
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_72_151
timestamp 1679235063
transform 1 0 14996 0 1 41344
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_72_162
timestamp 1679235063
transform 1 0 16008 0 1 41344
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_72_175
timestamp 1679235063
transform 1 0 17204 0 1 41344
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_72_179
timestamp 1679235063
transform 1 0 17572 0 1 41344
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_72_194
timestamp 1679235063
transform 1 0 18952 0 1 41344
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_72_199
timestamp 1679235063
transform 1 0 19412 0 1 41344
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_72_210
timestamp 1679235063
transform 1 0 20424 0 1 41344
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_72_218
timestamp 1679235063
transform 1 0 21160 0 1 41344
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_72_229
timestamp 1679235063
transform 1 0 22172 0 1 41344
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_72_233
timestamp 1679235063
transform 1 0 22540 0 1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_72_243
timestamp 1679235063
transform 1 0 23460 0 1 41344
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_72_250
timestamp 1679235063
transform 1 0 24104 0 1 41344
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_72_253
timestamp 1679235063
transform 1 0 24380 0 1 41344
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_72_263
timestamp 1679235063
transform 1 0 25300 0 1 41344
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_73_3
timestamp 1679235063
transform 1 0 1380 0 -1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_73_15
timestamp 1679235063
transform 1 0 2484 0 -1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_73_27
timestamp 1679235063
transform 1 0 3588 0 -1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_73_39
timestamp 1679235063
transform 1 0 4692 0 -1 42432
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_73_47
timestamp 1679235063
transform 1 0 5428 0 -1 42432
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_73_53
timestamp 1679235063
transform 1 0 5980 0 -1 42432
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_73_57
timestamp 1679235063
transform 1 0 6348 0 -1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_73_69
timestamp 1679235063
transform 1 0 7452 0 -1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_73_90
timestamp 1679235063
transform 1 0 9384 0 -1 42432
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_73_103
timestamp 1679235063
transform 1 0 10580 0 -1 42432
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_73_109
timestamp 1679235063
transform 1 0 11132 0 -1 42432
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_73_113
timestamp 1679235063
transform 1 0 11500 0 -1 42432
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_73_124
timestamp 1679235063
transform 1 0 12512 0 -1 42432
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_73_137
timestamp 1679235063
transform 1 0 13708 0 -1 42432
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_73_144
timestamp 1679235063
transform 1 0 14352 0 -1 42432
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_73_152
timestamp 1679235063
transform 1 0 15088 0 -1 42432
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_73_163
timestamp 1679235063
transform 1 0 16100 0 -1 42432
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_73_167
timestamp 1679235063
transform 1 0 16468 0 -1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_73_169
timestamp 1679235063
transform 1 0 16652 0 -1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_73_172
timestamp 1679235063
transform 1 0 16928 0 -1 42432
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_73_183
timestamp 1679235063
transform 1 0 17940 0 -1 42432
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_73_187
timestamp 1679235063
transform 1 0 18308 0 -1 42432
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_73_191
timestamp 1679235063
transform 1 0 18676 0 -1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_73_212
timestamp 1679235063
transform 1 0 20608 0 -1 42432
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_73_216
timestamp 1679235063
transform 1 0 20976 0 -1 42432
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_73_222
timestamp 1679235063
transform 1 0 21528 0 -1 42432
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_73_229
timestamp 1679235063
transform 1 0 22172 0 -1 42432
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_73_239
timestamp 1679235063
transform 1 0 23092 0 -1 42432
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_73_263
timestamp 1679235063
transform 1 0 25300 0 -1 42432
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_74_3
timestamp 1679235063
transform 1 0 1380 0 1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_74_15
timestamp 1679235063
transform 1 0 2484 0 1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_74_27
timestamp 1679235063
transform 1 0 3588 0 1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_74_29
timestamp 1679235063
transform 1 0 3772 0 1 42432
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_74_37
timestamp 1679235063
transform 1 0 4508 0 1 42432
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_74_43
timestamp 1679235063
transform 1 0 5060 0 1 42432
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_74_47
timestamp 1679235063
transform 1 0 5428 0 1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_74_59
timestamp 1679235063
transform 1 0 6532 0 1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_74_71
timestamp 1679235063
transform 1 0 7636 0 1 42432
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_74_81
timestamp 1679235063
transform 1 0 8556 0 1 42432
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_74_89
timestamp 1679235063
transform 1 0 9292 0 1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_74_92
timestamp 1679235063
transform 1 0 9568 0 1 42432
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_74_102
timestamp 1679235063
transform 1 0 10488 0 1 42432
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_74_126
timestamp 1679235063
transform 1 0 12696 0 1 42432
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_74_130
timestamp 1679235063
transform 1 0 13064 0 1 42432
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_74_138
timestamp 1679235063
transform 1 0 13800 0 1 42432
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_74_141
timestamp 1679235063
transform 1 0 14076 0 1 42432
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_74_147
timestamp 1679235063
transform 1 0 14628 0 1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_74_168
timestamp 1679235063
transform 1 0 16560 0 1 42432
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_74_172
timestamp 1679235063
transform 1 0 16928 0 1 42432
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_74_178
timestamp 1679235063
transform 1 0 17480 0 1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_74_181
timestamp 1679235063
transform 1 0 17756 0 1 42432
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_74_194
timestamp 1679235063
transform 1 0 18952 0 1 42432
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_74_197
timestamp 1679235063
transform 1 0 19228 0 1 42432
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_74_221
timestamp 1679235063
transform 1 0 21436 0 1 42432
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_74_234
timestamp 1679235063
transform 1 0 22632 0 1 42432
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_74_238
timestamp 1679235063
transform 1 0 23000 0 1 42432
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_74_250
timestamp 1679235063
transform 1 0 24104 0 1 42432
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_74_253
timestamp 1679235063
transform 1 0 24380 0 1 42432
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_74_264
timestamp 1679235063
transform 1 0 25392 0 1 42432
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_75_3
timestamp 1679235063
transform 1 0 1380 0 -1 43520
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_75_9
timestamp 1679235063
transform 1 0 1932 0 -1 43520
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_75_13
timestamp 1679235063
transform 1 0 2300 0 -1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_75_25
timestamp 1679235063
transform 1 0 3404 0 -1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_75_37
timestamp 1679235063
transform 1 0 4508 0 -1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_75_49
timestamp 1679235063
transform 1 0 5612 0 -1 43520
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_75_55
timestamp 1679235063
transform 1 0 6164 0 -1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_75_57
timestamp 1679235063
transform 1 0 6348 0 -1 43520
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_75_65
timestamp 1679235063
transform 1 0 7084 0 -1 43520
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_75_70
timestamp 1679235063
transform 1 0 7544 0 -1 43520
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_75_75
timestamp 1679235063
transform 1 0 8004 0 -1 43520
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_75_83
timestamp 1679235063
transform 1 0 8740 0 -1 43520
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_75_96
timestamp 1679235063
transform 1 0 9936 0 -1 43520
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_75_100
timestamp 1679235063
transform 1 0 10304 0 -1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_75_113
timestamp 1679235063
transform 1 0 11500 0 -1 43520
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_75_121
timestamp 1679235063
transform 1 0 12236 0 -1 43520
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_75_145
timestamp 1679235063
transform 1 0 14444 0 -1 43520
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_75_158
timestamp 1679235063
transform 1 0 15640 0 -1 43520
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_75_164
timestamp 1679235063
transform 1 0 16192 0 -1 43520
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_75_169
timestamp 1679235063
transform 1 0 16652 0 -1 43520
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_75_181
timestamp 1679235063
transform 1 0 17756 0 -1 43520
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_75_185
timestamp 1679235063
transform 1 0 18124 0 -1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_75_206
timestamp 1679235063
transform 1 0 20056 0 -1 43520
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_75_210
timestamp 1679235063
transform 1 0 20424 0 -1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_75_222
timestamp 1679235063
transform 1 0 21528 0 -1 43520
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_75_225
timestamp 1679235063
transform 1 0 21804 0 -1 43520
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_75_236
timestamp 1679235063
transform 1 0 22816 0 -1 43520
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_75_242
timestamp 1679235063
transform 1 0 23368 0 -1 43520
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_75_264
timestamp 1679235063
transform 1 0 25392 0 -1 43520
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_76_3
timestamp 1679235063
transform 1 0 1380 0 1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_76_15
timestamp 1679235063
transform 1 0 2484 0 1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_76_27
timestamp 1679235063
transform 1 0 3588 0 1 43520
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_76_29
timestamp 1679235063
transform 1 0 3772 0 1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_76_41
timestamp 1679235063
transform 1 0 4876 0 1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_76_53
timestamp 1679235063
transform 1 0 5980 0 1 43520
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_76_63
timestamp 1679235063
transform 1 0 6900 0 1 43520
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_76_67
timestamp 1679235063
transform 1 0 7268 0 1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_76_82
timestamp 1679235063
transform 1 0 8648 0 1 43520
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_76_85
timestamp 1679235063
transform 1 0 8924 0 1 43520
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_76_108
timestamp 1679235063
transform 1 0 11040 0 1 43520
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_76_112
timestamp 1679235063
transform 1 0 11408 0 1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_76_124
timestamp 1679235063
transform 1 0 12512 0 1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_76_136
timestamp 1679235063
transform 1 0 13616 0 1 43520
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_76_141
timestamp 1679235063
transform 1 0 14076 0 1 43520
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_76_151
timestamp 1679235063
transform 1 0 14996 0 1 43520
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_76_163
timestamp 1679235063
transform 1 0 16100 0 1 43520
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_76_171
timestamp 1679235063
transform 1 0 16836 0 1 43520
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_76_182
timestamp 1679235063
transform 1 0 17848 0 1 43520
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_76_188
timestamp 1679235063
transform 1 0 18400 0 1 43520
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_76_193
timestamp 1679235063
transform 1 0 18860 0 1 43520
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_76_197
timestamp 1679235063
transform 1 0 19228 0 1 43520
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_76_207
timestamp 1679235063
transform 1 0 20148 0 1 43520
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_76_213
timestamp 1679235063
transform 1 0 20700 0 1 43520
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_76_223
timestamp 1679235063
transform 1 0 21620 0 1 43520
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_76_227
timestamp 1679235063
transform 1 0 21988 0 1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_76_237
timestamp 1679235063
transform 1 0 22908 0 1 43520
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_76_249
timestamp 1679235063
transform 1 0 24012 0 1 43520
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_76_253
timestamp 1679235063
transform 1 0 24380 0 1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_76_258
timestamp 1679235063
transform 1 0 24840 0 1 43520
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_76_264
timestamp 1679235063
transform 1 0 25392 0 1 43520
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_77_3
timestamp 1679235063
transform 1 0 1380 0 -1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_77_15
timestamp 1679235063
transform 1 0 2484 0 -1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_77_27
timestamp 1679235063
transform 1 0 3588 0 -1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_77_39
timestamp 1679235063
transform 1 0 4692 0 -1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_77_54
timestamp 1679235063
transform 1 0 6072 0 -1 44608
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_77_57
timestamp 1679235063
transform 1 0 6348 0 -1 44608
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_77_63
timestamp 1679235063
transform 1 0 6900 0 -1 44608
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_77_71
timestamp 1679235063
transform 1 0 7636 0 -1 44608
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_77_75
timestamp 1679235063
transform 1 0 8004 0 -1 44608
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_77_83
timestamp 1679235063
transform 1 0 8740 0 -1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_77_88
timestamp 1679235063
transform 1 0 9200 0 -1 44608
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_77_92
timestamp 1679235063
transform 1 0 9568 0 -1 44608
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_77_96
timestamp 1679235063
transform 1 0 9936 0 -1 44608
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_77_102
timestamp 1679235063
transform 1 0 10488 0 -1 44608
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_77_110
timestamp 1679235063
transform 1 0 11224 0 -1 44608
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_77_115
timestamp 1679235063
transform 1 0 11684 0 -1 44608
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_77_126
timestamp 1679235063
transform 1 0 12696 0 -1 44608
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_77_150
timestamp 1679235063
transform 1 0 14904 0 -1 44608
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_77_154
timestamp 1679235063
transform 1 0 15272 0 -1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_77_166
timestamp 1679235063
transform 1 0 16376 0 -1 44608
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_77_169
timestamp 1679235063
transform 1 0 16652 0 -1 44608
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_77_191
timestamp 1679235063
transform 1 0 18676 0 -1 44608
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_77_203
timestamp 1679235063
transform 1 0 19780 0 -1 44608
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_77_215
timestamp 1679235063
transform 1 0 20884 0 -1 44608
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_77_223
timestamp 1679235063
transform 1 0 21620 0 -1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_77_225
timestamp 1679235063
transform 1 0 21804 0 -1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_77_228
timestamp 1679235063
transform 1 0 22080 0 -1 44608
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_77_250
timestamp 1679235063
transform 1 0 24104 0 -1 44608
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_77_264
timestamp 1679235063
transform 1 0 25392 0 -1 44608
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_78_3
timestamp 1679235063
transform 1 0 1380 0 1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_78_15
timestamp 1679235063
transform 1 0 2484 0 1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_78_27
timestamp 1679235063
transform 1 0 3588 0 1 44608
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_78_29
timestamp 1679235063
transform 1 0 3772 0 1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_78_41
timestamp 1679235063
transform 1 0 4876 0 1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_78_53
timestamp 1679235063
transform 1 0 5980 0 1 44608
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_78_59
timestamp 1679235063
transform 1 0 6532 0 1 44608
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_78_69
timestamp 1679235063
transform 1 0 7452 0 1 44608
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_78_75
timestamp 1679235063
transform 1 0 8004 0 1 44608
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_78_82
timestamp 1679235063
transform 1 0 8648 0 1 44608
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_78_85
timestamp 1679235063
transform 1 0 8924 0 1 44608
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_78_91
timestamp 1679235063
transform 1 0 9476 0 1 44608
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_78_95
timestamp 1679235063
transform 1 0 9844 0 1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_78_107
timestamp 1679235063
transform 1 0 10948 0 1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_78_112
timestamp 1679235063
transform 1 0 11408 0 1 44608
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_78_118
timestamp 1679235063
transform 1 0 11960 0 1 44608
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_78_124
timestamp 1679235063
transform 1 0 12512 0 1 44608
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_78_128
timestamp 1679235063
transform 1 0 12880 0 1 44608
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_78_138
timestamp 1679235063
transform 1 0 13800 0 1 44608
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_78_141
timestamp 1679235063
transform 1 0 14076 0 1 44608
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_78_149
timestamp 1679235063
transform 1 0 14812 0 1 44608
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_78_172
timestamp 1679235063
transform 1 0 16928 0 1 44608
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_78_176
timestamp 1679235063
transform 1 0 17296 0 1 44608
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_78_184
timestamp 1679235063
transform 1 0 18032 0 1 44608
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_78_194
timestamp 1679235063
transform 1 0 18952 0 1 44608
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_78_197
timestamp 1679235063
transform 1 0 19228 0 1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_78_200
timestamp 1679235063
transform 1 0 19504 0 1 44608
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_78_222
timestamp 1679235063
transform 1 0 21528 0 1 44608
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_78_226
timestamp 1679235063
transform 1 0 21896 0 1 44608
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_78_250
timestamp 1679235063
transform 1 0 24104 0 1 44608
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_78_253
timestamp 1679235063
transform 1 0 24380 0 1 44608
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_78_263
timestamp 1679235063
transform 1 0 25300 0 1 44608
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_79_3
timestamp 1679235063
transform 1 0 1380 0 -1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_79_15
timestamp 1679235063
transform 1 0 2484 0 -1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_79_27
timestamp 1679235063
transform 1 0 3588 0 -1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_79_39
timestamp 1679235063
transform 1 0 4692 0 -1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_79_51
timestamp 1679235063
transform 1 0 5796 0 -1 45696
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_79_55
timestamp 1679235063
transform 1 0 6164 0 -1 45696
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_79_57
timestamp 1679235063
transform 1 0 6348 0 -1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_79_69
timestamp 1679235063
transform 1 0 7452 0 -1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_79_81
timestamp 1679235063
transform 1 0 8556 0 -1 45696
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_79_85
timestamp 1679235063
transform 1 0 8924 0 -1 45696
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_79_107
timestamp 1679235063
transform 1 0 10948 0 -1 45696
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_79_111
timestamp 1679235063
transform 1 0 11316 0 -1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_79_113
timestamp 1679235063
transform 1 0 11500 0 -1 45696
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_79_119
timestamp 1679235063
transform 1 0 12052 0 -1 45696
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_79_123
timestamp 1679235063
transform 1 0 12420 0 -1 45696
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_79_140
timestamp 1679235063
transform 1 0 13984 0 -1 45696
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_79_164
timestamp 1679235063
transform 1 0 16192 0 -1 45696
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_79_169
timestamp 1679235063
transform 1 0 16652 0 -1 45696
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_79_179
timestamp 1679235063
transform 1 0 17572 0 -1 45696
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_79_185
timestamp 1679235063
transform 1 0 18124 0 -1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_79_206
timestamp 1679235063
transform 1 0 20056 0 -1 45696
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_79_219
timestamp 1679235063
transform 1 0 21252 0 -1 45696
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_79_223
timestamp 1679235063
transform 1 0 21620 0 -1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_79_225
timestamp 1679235063
transform 1 0 21804 0 -1 45696
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_79_248
timestamp 1679235063
transform 1 0 23920 0 -1 45696
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_79_252
timestamp 1679235063
transform 1 0 24288 0 -1 45696
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_79_264
timestamp 1679235063
transform 1 0 25392 0 -1 45696
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_80_3
timestamp 1679235063
transform 1 0 1380 0 1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_80_15
timestamp 1679235063
transform 1 0 2484 0 1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_80_27
timestamp 1679235063
transform 1 0 3588 0 1 45696
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_80_29
timestamp 1679235063
transform 1 0 3772 0 1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_80_41
timestamp 1679235063
transform 1 0 4876 0 1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_80_53
timestamp 1679235063
transform 1 0 5980 0 1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_80_65
timestamp 1679235063
transform 1 0 7084 0 1 45696
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_80_73
timestamp 1679235063
transform 1 0 7820 0 1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_80_78
timestamp 1679235063
transform 1 0 8280 0 1 45696
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_80_82
timestamp 1679235063
transform 1 0 8648 0 1 45696
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_80_85
timestamp 1679235063
transform 1 0 8924 0 1 45696
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_80_90
timestamp 1679235063
transform 1 0 9384 0 1 45696
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_80_96
timestamp 1679235063
transform 1 0 9936 0 1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_80_100
timestamp 1679235063
transform 1 0 10304 0 1 45696
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_80_113
timestamp 1679235063
transform 1 0 11500 0 1 45696
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_80_138
timestamp 1679235063
transform 1 0 13800 0 1 45696
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_80_143
timestamp 1679235063
transform 1 0 14260 0 1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_80_155
timestamp 1679235063
transform 1 0 15364 0 1 45696
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_80_159
timestamp 1679235063
transform 1 0 15732 0 1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_80_168
timestamp 1679235063
transform 1 0 16560 0 1 45696
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_80_172
timestamp 1679235063
transform 1 0 16928 0 1 45696
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_80_194
timestamp 1679235063
transform 1 0 18952 0 1 45696
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_80_197
timestamp 1679235063
transform 1 0 19228 0 1 45696
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_80_220
timestamp 1679235063
transform 1 0 21344 0 1 45696
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_80_224
timestamp 1679235063
transform 1 0 21712 0 1 45696
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_80_228
timestamp 1679235063
transform 1 0 22080 0 1 45696
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_80_239
timestamp 1679235063
transform 1 0 23092 0 1 45696
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_80_245
timestamp 1679235063
transform 1 0 23644 0 1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_80_253
timestamp 1679235063
transform 1 0 24380 0 1 45696
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_80_263
timestamp 1679235063
transform 1 0 25300 0 1 45696
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_81_3
timestamp 1679235063
transform 1 0 1380 0 -1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_81_15
timestamp 1679235063
transform 1 0 2484 0 -1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_81_27
timestamp 1679235063
transform 1 0 3588 0 -1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_81_39
timestamp 1679235063
transform 1 0 4692 0 -1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_81_51
timestamp 1679235063
transform 1 0 5796 0 -1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_81_55
timestamp 1679235063
transform 1 0 6164 0 -1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_81_57
timestamp 1679235063
transform 1 0 6348 0 -1 46784
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_81_65
timestamp 1679235063
transform 1 0 7084 0 -1 46784
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_81_70
timestamp 1679235063
transform 1 0 7544 0 -1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_81_82
timestamp 1679235063
transform 1 0 8648 0 -1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_81_94
timestamp 1679235063
transform 1 0 9752 0 -1 46784
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_81_110
timestamp 1679235063
transform 1 0 11224 0 -1 46784
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_81_113
timestamp 1679235063
transform 1 0 11500 0 -1 46784
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_81_118
timestamp 1679235063
transform 1 0 11960 0 -1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_81_142
timestamp 1679235063
transform 1 0 14168 0 -1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_81_166
timestamp 1679235063
transform 1 0 16376 0 -1 46784
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_81_169
timestamp 1679235063
transform 1 0 16652 0 -1 46784
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_81_191
timestamp 1679235063
transform 1 0 18676 0 -1 46784
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_81_200
timestamp 1679235063
transform 1 0 19504 0 -1 46784
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_81_211
timestamp 1679235063
transform 1 0 20516 0 -1 46784
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_81_219
timestamp 1679235063
transform 1 0 21252 0 -1 46784
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_81_225
timestamp 1679235063
transform 1 0 21804 0 -1 46784
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_81_236
timestamp 1679235063
transform 1 0 22816 0 -1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_81_248
timestamp 1679235063
transform 1 0 23920 0 -1 46784
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_81_252
timestamp 1679235063
transform 1 0 24288 0 -1 46784
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_81_264
timestamp 1679235063
transform 1 0 25392 0 -1 46784
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_82_3
timestamp 1679235063
transform 1 0 1380 0 1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_82_15
timestamp 1679235063
transform 1 0 2484 0 1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_82_27
timestamp 1679235063
transform 1 0 3588 0 1 46784
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_82_29
timestamp 1679235063
transform 1 0 3772 0 1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_82_41
timestamp 1679235063
transform 1 0 4876 0 1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_82_53
timestamp 1679235063
transform 1 0 5980 0 1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_82_65
timestamp 1679235063
transform 1 0 7084 0 1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_82_77
timestamp 1679235063
transform 1 0 8188 0 1 46784
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_82_83
timestamp 1679235063
transform 1 0 8740 0 1 46784
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_82_85
timestamp 1679235063
transform 1 0 8924 0 1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_82_97
timestamp 1679235063
transform 1 0 10028 0 1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_82_118
timestamp 1679235063
transform 1 0 11960 0 1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_82_130
timestamp 1679235063
transform 1 0 13064 0 1 46784
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_82_138
timestamp 1679235063
transform 1 0 13800 0 1 46784
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_82_141
timestamp 1679235063
transform 1 0 14076 0 1 46784
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_82_144
timestamp 1679235063
transform 1 0 14352 0 1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_82_156
timestamp 1679235063
transform 1 0 15456 0 1 46784
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_82_179
timestamp 1679235063
transform 1 0 17572 0 1 46784
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_82_183
timestamp 1679235063
transform 1 0 17940 0 1 46784
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_82_194
timestamp 1679235063
transform 1 0 18952 0 1 46784
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_82_197
timestamp 1679235063
transform 1 0 19228 0 1 46784
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_82_207
timestamp 1679235063
transform 1 0 20148 0 1 46784
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_82_219
timestamp 1679235063
transform 1 0 21252 0 1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_82_231
timestamp 1679235063
transform 1 0 22356 0 1 46784
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_82_239
timestamp 1679235063
transform 1 0 23092 0 1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_82_250
timestamp 1679235063
transform 1 0 24104 0 1 46784
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_82_255
timestamp 1679235063
transform 1 0 24564 0 1 46784
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_82_261
timestamp 1679235063
transform 1 0 25116 0 1 46784
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_83_3
timestamp 1679235063
transform 1 0 1380 0 -1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_83_15
timestamp 1679235063
transform 1 0 2484 0 -1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_83_27
timestamp 1679235063
transform 1 0 3588 0 -1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_83_39
timestamp 1679235063
transform 1 0 4692 0 -1 47872
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_83_51
timestamp 1679235063
transform 1 0 5796 0 -1 47872
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_83_55
timestamp 1679235063
transform 1 0 6164 0 -1 47872
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_83_57
timestamp 1679235063
transform 1 0 6348 0 -1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_83_69
timestamp 1679235063
transform 1 0 7452 0 -1 47872
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_83_81
timestamp 1679235063
transform 1 0 8556 0 -1 47872
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_83_87
timestamp 1679235063
transform 1 0 9108 0 -1 47872
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_83_91
timestamp 1679235063
transform 1 0 9476 0 -1 47872
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_83_103
timestamp 1679235063
transform 1 0 10580 0 -1 47872
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_83_111
timestamp 1679235063
transform 1 0 11316 0 -1 47872
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_83_113
timestamp 1679235063
transform 1 0 11500 0 -1 47872
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_83_117
timestamp 1679235063
transform 1 0 11868 0 -1 47872
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_83_120
timestamp 1679235063
transform 1 0 12144 0 -1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_83_132
timestamp 1679235063
transform 1 0 13248 0 -1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_83_144
timestamp 1679235063
transform 1 0 14352 0 -1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_83_156
timestamp 1679235063
transform 1 0 15456 0 -1 47872
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_83_169
timestamp 1679235063
transform 1 0 16652 0 -1 47872
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_83_180
timestamp 1679235063
transform 1 0 17664 0 -1 47872
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_83_193
timestamp 1679235063
transform 1 0 18860 0 -1 47872
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_83_199
timestamp 1679235063
transform 1 0 19412 0 -1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_83_211
timestamp 1679235063
transform 1 0 20516 0 -1 47872
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_83_223
timestamp 1679235063
transform 1 0 21620 0 -1 47872
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_83_225
timestamp 1679235063
transform 1 0 21804 0 -1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_83_237
timestamp 1679235063
transform 1 0 22908 0 -1 47872
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_83_249
timestamp 1679235063
transform 1 0 24012 0 -1 47872
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_83_253
timestamp 1679235063
transform 1 0 24380 0 -1 47872
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_83_264
timestamp 1679235063
transform 1 0 25392 0 -1 47872
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_84_3
timestamp 1679235063
transform 1 0 1380 0 1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_84_15
timestamp 1679235063
transform 1 0 2484 0 1 47872
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_84_27
timestamp 1679235063
transform 1 0 3588 0 1 47872
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_84_29
timestamp 1679235063
transform 1 0 3772 0 1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_84_41
timestamp 1679235063
transform 1 0 4876 0 1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_84_53
timestamp 1679235063
transform 1 0 5980 0 1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_84_65
timestamp 1679235063
transform 1 0 7084 0 1 47872
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_84_77
timestamp 1679235063
transform 1 0 8188 0 1 47872
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_84_83
timestamp 1679235063
transform 1 0 8740 0 1 47872
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_84_85
timestamp 1679235063
transform 1 0 8924 0 1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_84_97
timestamp 1679235063
transform 1 0 10028 0 1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_84_109
timestamp 1679235063
transform 1 0 11132 0 1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_84_121
timestamp 1679235063
transform 1 0 12236 0 1 47872
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_84_133
timestamp 1679235063
transform 1 0 13340 0 1 47872
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_84_139
timestamp 1679235063
transform 1 0 13892 0 1 47872
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_84_141
timestamp 1679235063
transform 1 0 14076 0 1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_84_153
timestamp 1679235063
transform 1 0 15180 0 1 47872
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_84_165
timestamp 1679235063
transform 1 0 16284 0 1 47872
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_84_173
timestamp 1679235063
transform 1 0 17020 0 1 47872
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_84_182
timestamp 1679235063
transform 1 0 17848 0 1 47872
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_84_186
timestamp 1679235063
transform 1 0 18216 0 1 47872
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_84_194
timestamp 1679235063
transform 1 0 18952 0 1 47872
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_84_197
timestamp 1679235063
transform 1 0 19228 0 1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_84_209
timestamp 1679235063
transform 1 0 20332 0 1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_84_221
timestamp 1679235063
transform 1 0 21436 0 1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_84_233
timestamp 1679235063
transform 1 0 22540 0 1 47872
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_84_245
timestamp 1679235063
transform 1 0 23644 0 1 47872
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_84_251
timestamp 1679235063
transform 1 0 24196 0 1 47872
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_84_253
timestamp 1679235063
transform 1 0 24380 0 1 47872
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_84_261
timestamp 1679235063
transform 1 0 25116 0 1 47872
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_85_3
timestamp 1679235063
transform 1 0 1380 0 -1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_85_15
timestamp 1679235063
transform 1 0 2484 0 -1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_85_27
timestamp 1679235063
transform 1 0 3588 0 -1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_85_39
timestamp 1679235063
transform 1 0 4692 0 -1 48960
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_85_51
timestamp 1679235063
transform 1 0 5796 0 -1 48960
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_85_55
timestamp 1679235063
transform 1 0 6164 0 -1 48960
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_85_57
timestamp 1679235063
transform 1 0 6348 0 -1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_85_69
timestamp 1679235063
transform 1 0 7452 0 -1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_85_81
timestamp 1679235063
transform 1 0 8556 0 -1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_85_93
timestamp 1679235063
transform 1 0 9660 0 -1 48960
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_85_105
timestamp 1679235063
transform 1 0 10764 0 -1 48960
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_85_111
timestamp 1679235063
transform 1 0 11316 0 -1 48960
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_85_113
timestamp 1679235063
transform 1 0 11500 0 -1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_85_125
timestamp 1679235063
transform 1 0 12604 0 -1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_85_137
timestamp 1679235063
transform 1 0 13708 0 -1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_85_149
timestamp 1679235063
transform 1 0 14812 0 -1 48960
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_85_161
timestamp 1679235063
transform 1 0 15916 0 -1 48960
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_85_167
timestamp 1679235063
transform 1 0 16468 0 -1 48960
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_85_169
timestamp 1679235063
transform 1 0 16652 0 -1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_85_181
timestamp 1679235063
transform 1 0 17756 0 -1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_85_193
timestamp 1679235063
transform 1 0 18860 0 -1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_85_205
timestamp 1679235063
transform 1 0 19964 0 -1 48960
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_85_217
timestamp 1679235063
transform 1 0 21068 0 -1 48960
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_85_223
timestamp 1679235063
transform 1 0 21620 0 -1 48960
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_85_225
timestamp 1679235063
transform 1 0 21804 0 -1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_85_237
timestamp 1679235063
transform 1 0 22908 0 -1 48960
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_85_249
timestamp 1679235063
transform 1 0 24012 0 -1 48960
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_85_253
timestamp 1679235063
transform 1 0 24380 0 -1 48960
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_85_264
timestamp 1679235063
transform 1 0 25392 0 -1 48960
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_86_3
timestamp 1679235063
transform 1 0 1380 0 1 48960
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_86_21
timestamp 1679235063
transform 1 0 3036 0 1 48960
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_86_25
timestamp 1679235063
transform 1 0 3404 0 1 48960
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_86_29
timestamp 1679235063
transform 1 0 3772 0 1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_86_41
timestamp 1679235063
transform 1 0 4876 0 1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_86_53
timestamp 1679235063
transform 1 0 5980 0 1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_86_65
timestamp 1679235063
transform 1 0 7084 0 1 48960
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_86_77
timestamp 1679235063
transform 1 0 8188 0 1 48960
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_86_83
timestamp 1679235063
transform 1 0 8740 0 1 48960
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_86_85
timestamp 1679235063
transform 1 0 8924 0 1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_86_97
timestamp 1679235063
transform 1 0 10028 0 1 48960
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_86_109
timestamp 1679235063
transform 1 0 11132 0 1 48960
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_86_113
timestamp 1679235063
transform 1 0 11500 0 1 48960
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_86_117
timestamp 1679235063
transform 1 0 11868 0 1 48960
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_86_125
timestamp 1679235063
transform 1 0 12604 0 1 48960
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_86_129
timestamp 1679235063
transform 1 0 12972 0 1 48960
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_86_137
timestamp 1679235063
transform 1 0 13708 0 1 48960
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_86_141
timestamp 1679235063
transform 1 0 14076 0 1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_86_153
timestamp 1679235063
transform 1 0 15180 0 1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_86_165
timestamp 1679235063
transform 1 0 16284 0 1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_86_177
timestamp 1679235063
transform 1 0 17388 0 1 48960
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_86_189
timestamp 1679235063
transform 1 0 18492 0 1 48960
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_86_195
timestamp 1679235063
transform 1 0 19044 0 1 48960
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_86_197
timestamp 1679235063
transform 1 0 19228 0 1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_86_209
timestamp 1679235063
transform 1 0 20332 0 1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_86_221
timestamp 1679235063
transform 1 0 21436 0 1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_86_233
timestamp 1679235063
transform 1 0 22540 0 1 48960
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_86_245
timestamp 1679235063
transform 1 0 23644 0 1 48960
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_86_251
timestamp 1679235063
transform 1 0 24196 0 1 48960
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_86_253
timestamp 1679235063
transform 1 0 24380 0 1 48960
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_86_259
timestamp 1679235063
transform 1 0 24932 0 1 48960
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_86_264
timestamp 1679235063
transform 1 0 25392 0 1 48960
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_87_3
timestamp 1679235063
transform 1 0 1380 0 -1 50048
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_87_25
timestamp 1679235063
transform 1 0 3404 0 -1 50048
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_87_54
timestamp 1679235063
transform 1 0 6072 0 -1 50048
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_87_61
timestamp 1679235063
transform 1 0 6716 0 -1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_87_73
timestamp 1679235063
transform 1 0 7820 0 -1 50048
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_87_85
timestamp 1679235063
transform 1 0 8924 0 -1 50048
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_87_91
timestamp 1679235063
transform 1 0 9476 0 -1 50048
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_87_103
timestamp 1679235063
transform 1 0 10580 0 -1 50048
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_87_111
timestamp 1679235063
transform 1 0 11316 0 -1 50048
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_87_113
timestamp 1679235063
transform 1 0 11500 0 -1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_87_125
timestamp 1679235063
transform 1 0 12604 0 -1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_87_137
timestamp 1679235063
transform 1 0 13708 0 -1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_87_149
timestamp 1679235063
transform 1 0 14812 0 -1 50048
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_87_161
timestamp 1679235063
transform 1 0 15916 0 -1 50048
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_87_167
timestamp 1679235063
transform 1 0 16468 0 -1 50048
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_87_169
timestamp 1679235063
transform 1 0 16652 0 -1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_87_181
timestamp 1679235063
transform 1 0 17756 0 -1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_87_193
timestamp 1679235063
transform 1 0 18860 0 -1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_87_205
timestamp 1679235063
transform 1 0 19964 0 -1 50048
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_87_217
timestamp 1679235063
transform 1 0 21068 0 -1 50048
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_87_223
timestamp 1679235063
transform 1 0 21620 0 -1 50048
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_87_225
timestamp 1679235063
transform 1 0 21804 0 -1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_87_237
timestamp 1679235063
transform 1 0 22908 0 -1 50048
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_87_249
timestamp 1679235063
transform 1 0 24012 0 -1 50048
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_87_253
timestamp 1679235063
transform 1 0 24380 0 -1 50048
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_87_264
timestamp 1679235063
transform 1 0 25392 0 -1 50048
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_88_3
timestamp 1679235063
transform 1 0 1380 0 1 50048
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_88_9
timestamp 1679235063
transform 1 0 1932 0 1 50048
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_88_26
timestamp 1679235063
transform 1 0 3496 0 1 50048
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_88_29
timestamp 1679235063
transform 1 0 3772 0 1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_88_41
timestamp 1679235063
transform 1 0 4876 0 1 50048
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_88_53
timestamp 1679235063
transform 1 0 5980 0 1 50048
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_88_61
timestamp 1679235063
transform 1 0 6716 0 1 50048
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_88_65
timestamp 1679235063
transform 1 0 7084 0 1 50048
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_88_77
timestamp 1679235063
transform 1 0 8188 0 1 50048
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_88_83
timestamp 1679235063
transform 1 0 8740 0 1 50048
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_88_85
timestamp 1679235063
transform 1 0 8924 0 1 50048
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_88_91
timestamp 1679235063
transform 1 0 9476 0 1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_88_103
timestamp 1679235063
transform 1 0 10580 0 1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_88_115
timestamp 1679235063
transform 1 0 11684 0 1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_88_127
timestamp 1679235063
transform 1 0 12788 0 1 50048
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_88_139
timestamp 1679235063
transform 1 0 13892 0 1 50048
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_88_141
timestamp 1679235063
transform 1 0 14076 0 1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_88_153
timestamp 1679235063
transform 1 0 15180 0 1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_88_165
timestamp 1679235063
transform 1 0 16284 0 1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_88_177
timestamp 1679235063
transform 1 0 17388 0 1 50048
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_88_189
timestamp 1679235063
transform 1 0 18492 0 1 50048
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_88_195
timestamp 1679235063
transform 1 0 19044 0 1 50048
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_88_197
timestamp 1679235063
transform 1 0 19228 0 1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_88_209
timestamp 1679235063
transform 1 0 20332 0 1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_88_221
timestamp 1679235063
transform 1 0 21436 0 1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_88_233
timestamp 1679235063
transform 1 0 22540 0 1 50048
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_88_245
timestamp 1679235063
transform 1 0 23644 0 1 50048
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_88_251
timestamp 1679235063
transform 1 0 24196 0 1 50048
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_88_253
timestamp 1679235063
transform 1 0 24380 0 1 50048
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_88_259
timestamp 1679235063
transform 1 0 24932 0 1 50048
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_88_264
timestamp 1679235063
transform 1 0 25392 0 1 50048
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_89_3
timestamp 1679235063
transform 1 0 1380 0 -1 51136
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_89_11
timestamp 1679235063
transform 1 0 2116 0 -1 51136
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_89_29
timestamp 1679235063
transform 1 0 3772 0 -1 51136
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_89_49
timestamp 1679235063
transform 1 0 5612 0 -1 51136
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_89_55
timestamp 1679235063
transform 1 0 6164 0 -1 51136
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_89_57
timestamp 1679235063
transform 1 0 6348 0 -1 51136
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_89_65
timestamp 1679235063
transform 1 0 7084 0 -1 51136
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_89_79
timestamp 1679235063
transform 1 0 8372 0 -1 51136
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_89_87
timestamp 1679235063
transform 1 0 9108 0 -1 51136
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_89_93
timestamp 1679235063
transform 1 0 9660 0 -1 51136
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_89_105
timestamp 1679235063
transform 1 0 10764 0 -1 51136
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_89_111
timestamp 1679235063
transform 1 0 11316 0 -1 51136
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_89_113
timestamp 1679235063
transform 1 0 11500 0 -1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_89_125
timestamp 1679235063
transform 1 0 12604 0 -1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_89_137
timestamp 1679235063
transform 1 0 13708 0 -1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_89_149
timestamp 1679235063
transform 1 0 14812 0 -1 51136
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_89_161
timestamp 1679235063
transform 1 0 15916 0 -1 51136
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_89_167
timestamp 1679235063
transform 1 0 16468 0 -1 51136
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_89_169
timestamp 1679235063
transform 1 0 16652 0 -1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_89_181
timestamp 1679235063
transform 1 0 17756 0 -1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_89_193
timestamp 1679235063
transform 1 0 18860 0 -1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_89_205
timestamp 1679235063
transform 1 0 19964 0 -1 51136
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_89_217
timestamp 1679235063
transform 1 0 21068 0 -1 51136
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_89_223
timestamp 1679235063
transform 1 0 21620 0 -1 51136
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_89_225
timestamp 1679235063
transform 1 0 21804 0 -1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_89_237
timestamp 1679235063
transform 1 0 22908 0 -1 51136
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_89_249
timestamp 1679235063
transform 1 0 24012 0 -1 51136
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_89_255
timestamp 1679235063
transform 1 0 24564 0 -1 51136
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_89_258
timestamp 1679235063
transform 1 0 24840 0 -1 51136
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_89_264
timestamp 1679235063
transform 1 0 25392 0 -1 51136
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_90_3
timestamp 1679235063
transform 1 0 1380 0 1 51136
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_90_9
timestamp 1679235063
transform 1 0 1932 0 1 51136
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_90_26
timestamp 1679235063
transform 1 0 3496 0 1 51136
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_90_29
timestamp 1679235063
transform 1 0 3772 0 1 51136
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_90_41
timestamp 1679235063
transform 1 0 4876 0 1 51136
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_90_61
timestamp 1679235063
transform 1 0 6716 0 1 51136
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_90_81
timestamp 1679235063
transform 1 0 8556 0 1 51136
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_90_85
timestamp 1679235063
transform 1 0 8924 0 1 51136
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_90_97
timestamp 1679235063
transform 1 0 10028 0 1 51136
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_90_102
timestamp 1679235063
transform 1 0 10488 0 1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_90_114
timestamp 1679235063
transform 1 0 11592 0 1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_90_126
timestamp 1679235063
transform 1 0 12696 0 1 51136
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_90_138
timestamp 1679235063
transform 1 0 13800 0 1 51136
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_90_141
timestamp 1679235063
transform 1 0 14076 0 1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_90_153
timestamp 1679235063
transform 1 0 15180 0 1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_90_165
timestamp 1679235063
transform 1 0 16284 0 1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_90_177
timestamp 1679235063
transform 1 0 17388 0 1 51136
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_90_189
timestamp 1679235063
transform 1 0 18492 0 1 51136
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_90_195
timestamp 1679235063
transform 1 0 19044 0 1 51136
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_90_197
timestamp 1679235063
transform 1 0 19228 0 1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_90_209
timestamp 1679235063
transform 1 0 20332 0 1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_90_221
timestamp 1679235063
transform 1 0 21436 0 1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_90_233
timestamp 1679235063
transform 1 0 22540 0 1 51136
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_90_245
timestamp 1679235063
transform 1 0 23644 0 1 51136
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_90_251
timestamp 1679235063
transform 1 0 24196 0 1 51136
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_90_253
timestamp 1679235063
transform 1 0 24380 0 1 51136
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_90_259
timestamp 1679235063
transform 1 0 24932 0 1 51136
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_90_264
timestamp 1679235063
transform 1 0 25392 0 1 51136
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_91_3
timestamp 1679235063
transform 1 0 1380 0 -1 52224
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_91_15
timestamp 1679235063
transform 1 0 2484 0 -1 52224
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_91_34
timestamp 1679235063
transform 1 0 4232 0 -1 52224
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_91_54
timestamp 1679235063
transform 1 0 6072 0 -1 52224
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_91_57
timestamp 1679235063
transform 1 0 6348 0 -1 52224
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_91_61
timestamp 1679235063
transform 1 0 6716 0 -1 52224
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_91_66
timestamp 1679235063
transform 1 0 7176 0 -1 52224
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_91_72
timestamp 1679235063
transform 1 0 7728 0 -1 52224
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_91_89
timestamp 1679235063
transform 1 0 9292 0 -1 52224
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_91_109
timestamp 1679235063
transform 1 0 11132 0 -1 52224
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_91_113
timestamp 1679235063
transform 1 0 11500 0 -1 52224
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_91_118
timestamp 1679235063
transform 1 0 11960 0 -1 52224
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_91_125
timestamp 1679235063
transform 1 0 12604 0 -1 52224
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_91_133
timestamp 1679235063
transform 1 0 13340 0 -1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_91_145
timestamp 1679235063
transform 1 0 14444 0 -1 52224
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_91_157
timestamp 1679235063
transform 1 0 15548 0 -1 52224
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_91_165
timestamp 1679235063
transform 1 0 16284 0 -1 52224
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_91_169
timestamp 1679235063
transform 1 0 16652 0 -1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_91_181
timestamp 1679235063
transform 1 0 17756 0 -1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_91_193
timestamp 1679235063
transform 1 0 18860 0 -1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_91_205
timestamp 1679235063
transform 1 0 19964 0 -1 52224
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_91_217
timestamp 1679235063
transform 1 0 21068 0 -1 52224
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_91_223
timestamp 1679235063
transform 1 0 21620 0 -1 52224
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_91_225
timestamp 1679235063
transform 1 0 21804 0 -1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_91_237
timestamp 1679235063
transform 1 0 22908 0 -1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_91_249
timestamp 1679235063
transform 1 0 24012 0 -1 52224
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_91_261
timestamp 1679235063
transform 1 0 25116 0 -1 52224
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_92_3
timestamp 1679235063
transform 1 0 1380 0 1 52224
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_92_9
timestamp 1679235063
transform 1 0 1932 0 1 52224
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_92_26
timestamp 1679235063
transform 1 0 3496 0 1 52224
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_92_29
timestamp 1679235063
transform 1 0 3772 0 1 52224
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_92_41
timestamp 1679235063
transform 1 0 4876 0 1 52224
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_92_45
timestamp 1679235063
transform 1 0 5244 0 1 52224
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_92_62
timestamp 1679235063
transform 1 0 6808 0 1 52224
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_92_82
timestamp 1679235063
transform 1 0 8648 0 1 52224
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_92_85
timestamp 1679235063
transform 1 0 8924 0 1 52224
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_92_97
timestamp 1679235063
transform 1 0 10028 0 1 52224
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_92_121
timestamp 1679235063
transform 1 0 12236 0 1 52224
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_92_128
timestamp 1679235063
transform 1 0 12880 0 1 52224
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_92_132
timestamp 1679235063
transform 1 0 13248 0 1 52224
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_92_137
timestamp 1679235063
transform 1 0 13708 0 1 52224
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_92_143
timestamp 1679235063
transform 1 0 14260 0 1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_92_155
timestamp 1679235063
transform 1 0 15364 0 1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_92_167
timestamp 1679235063
transform 1 0 16468 0 1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_92_179
timestamp 1679235063
transform 1 0 17572 0 1 52224
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_92_191
timestamp 1679235063
transform 1 0 18676 0 1 52224
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_92_195
timestamp 1679235063
transform 1 0 19044 0 1 52224
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_92_197
timestamp 1679235063
transform 1 0 19228 0 1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_92_209
timestamp 1679235063
transform 1 0 20332 0 1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_92_221
timestamp 1679235063
transform 1 0 21436 0 1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_92_233
timestamp 1679235063
transform 1 0 22540 0 1 52224
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_92_245
timestamp 1679235063
transform 1 0 23644 0 1 52224
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_92_251
timestamp 1679235063
transform 1 0 24196 0 1 52224
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_92_253
timestamp 1679235063
transform 1 0 24380 0 1 52224
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_92_258
timestamp 1679235063
transform 1 0 24840 0 1 52224
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_92_264
timestamp 1679235063
transform 1 0 25392 0 1 52224
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_93_3
timestamp 1679235063
transform 1 0 1380 0 -1 53312
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_93_8
timestamp 1679235063
transform 1 0 1840 0 -1 53312
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_93_12
timestamp 1679235063
transform 1 0 2208 0 -1 53312
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_93_34
timestamp 1679235063
transform 1 0 4232 0 -1 53312
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_93_54
timestamp 1679235063
transform 1 0 6072 0 -1 53312
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_93_57
timestamp 1679235063
transform 1 0 6348 0 -1 53312
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_93_69
timestamp 1679235063
transform 1 0 7452 0 -1 53312
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_93_73
timestamp 1679235063
transform 1 0 7820 0 -1 53312
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_93_90
timestamp 1679235063
transform 1 0 9384 0 -1 53312
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_93_110
timestamp 1679235063
transform 1 0 11224 0 -1 53312
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_93_113
timestamp 1679235063
transform 1 0 11500 0 -1 53312
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_93_133
timestamp 1679235063
transform 1 0 13340 0 -1 53312
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_93_141
timestamp 1679235063
transform 1 0 14076 0 -1 53312
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_93_148
timestamp 1679235063
transform 1 0 14720 0 -1 53312
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_93_152
timestamp 1679235063
transform 1 0 15088 0 -1 53312
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_93_160
timestamp 1679235063
transform 1 0 15824 0 -1 53312
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_93_164
timestamp 1679235063
transform 1 0 16192 0 -1 53312
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_93_169
timestamp 1679235063
transform 1 0 16652 0 -1 53312
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_93_177
timestamp 1679235063
transform 1 0 17388 0 -1 53312
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_93_189
timestamp 1679235063
transform 1 0 18492 0 -1 53312
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_93_196
timestamp 1679235063
transform 1 0 19136 0 -1 53312
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_93_204
timestamp 1679235063
transform 1 0 19872 0 -1 53312
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_93_208
timestamp 1679235063
transform 1 0 20240 0 -1 53312
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_93_212
timestamp 1679235063
transform 1 0 20608 0 -1 53312
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_93_220
timestamp 1679235063
transform 1 0 21344 0 -1 53312
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_93_227
timestamp 1679235063
transform 1 0 21988 0 -1 53312
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_93_232
timestamp 1679235063
transform 1 0 22448 0 -1 53312
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_93_235
timestamp 1679235063
transform 1 0 22724 0 -1 53312
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_93_239
timestamp 1679235063
transform 1 0 23092 0 -1 53312
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_93_244
timestamp 1679235063
transform 1 0 23552 0 -1 53312
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_93_251
timestamp 1679235063
transform 1 0 24196 0 -1 53312
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_93_255
timestamp 1679235063
transform 1 0 24564 0 -1 53312
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_93_258
timestamp 1679235063
transform 1 0 24840 0 -1 53312
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_93_264
timestamp 1679235063
transform 1 0 25392 0 -1 53312
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_94_3
timestamp 1679235063
transform 1 0 1380 0 1 53312
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_94_9
timestamp 1679235063
transform 1 0 1932 0 1 53312
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_94_26
timestamp 1679235063
transform 1 0 3496 0 1 53312
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_94_29
timestamp 1679235063
transform 1 0 3772 0 1 53312
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_94_41
timestamp 1679235063
transform 1 0 4876 0 1 53312
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_94_45
timestamp 1679235063
transform 1 0 5244 0 1 53312
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_94_62
timestamp 1679235063
transform 1 0 6808 0 1 53312
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_94_82
timestamp 1679235063
transform 1 0 8648 0 1 53312
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_94_85
timestamp 1679235063
transform 1 0 8924 0 1 53312
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_94_97
timestamp 1679235063
transform 1 0 10028 0 1 53312
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_94_117
timestamp 1679235063
transform 1 0 11868 0 1 53312
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_94_137
timestamp 1679235063
transform 1 0 13708 0 1 53312
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_94_141
timestamp 1679235063
transform 1 0 14076 0 1 53312
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_94_147
timestamp 1679235063
transform 1 0 14628 0 1 53312
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_94_151
timestamp 1679235063
transform 1 0 14996 0 1 53312
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_94_161
timestamp 1679235063
transform 1 0 15916 0 1 53312
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_94_167
timestamp 1679235063
transform 1 0 16468 0 1 53312
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_94_173
timestamp 1679235063
transform 1 0 17020 0 1 53312
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_94_180
timestamp 1679235063
transform 1 0 17664 0 1 53312
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_94_184
timestamp 1679235063
transform 1 0 18032 0 1 53312
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_94_189
timestamp 1679235063
transform 1 0 18492 0 1 53312
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_94_195
timestamp 1679235063
transform 1 0 19044 0 1 53312
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_94_197
timestamp 1679235063
transform 1 0 19228 0 1 53312
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_94_203
timestamp 1679235063
transform 1 0 19780 0 1 53312
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_94_211
timestamp 1679235063
transform 1 0 20516 0 1 53312
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_94_215
timestamp 1679235063
transform 1 0 20884 0 1 53312
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_94_221
timestamp 1679235063
transform 1 0 21436 0 1 53312
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_94_228
timestamp 1679235063
transform 1 0 22080 0 1 53312
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_94_235
timestamp 1679235063
transform 1 0 22724 0 1 53312
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_94_242
timestamp 1679235063
transform 1 0 23368 0 1 53312
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_94_250
timestamp 1679235063
transform 1 0 24104 0 1 53312
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_94_255
timestamp 1679235063
transform 1 0 24564 0 1 53312
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_94_264
timestamp 1679235063
transform 1 0 25392 0 1 53312
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_95_3
timestamp 1679235063
transform 1 0 1380 0 -1 54400
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_95_9
timestamp 1679235063
transform 1 0 1932 0 -1 54400
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_95_26
timestamp 1679235063
transform 1 0 3496 0 -1 54400
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_95_29
timestamp 1679235063
transform 1 0 3772 0 -1 54400
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_95_37
timestamp 1679235063
transform 1 0 4508 0 -1 54400
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_95_54
timestamp 1679235063
transform 1 0 6072 0 -1 54400
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_95_57
timestamp 1679235063
transform 1 0 6348 0 -1 54400
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_95_65
timestamp 1679235063
transform 1 0 7084 0 -1 54400
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_95_82
timestamp 1679235063
transform 1 0 8648 0 -1 54400
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_95_85
timestamp 1679235063
transform 1 0 8924 0 -1 54400
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_95_93
timestamp 1679235063
transform 1 0 9660 0 -1 54400
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_95_110
timestamp 1679235063
transform 1 0 11224 0 -1 54400
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_95_113
timestamp 1679235063
transform 1 0 11500 0 -1 54400
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_95_118
timestamp 1679235063
transform 1 0 11960 0 -1 54400
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_95_138
timestamp 1679235063
transform 1 0 13800 0 -1 54400
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_95_143
timestamp 1679235063
transform 1 0 14260 0 -1 54400
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_95_147
timestamp 1679235063
transform 1 0 14628 0 -1 54400
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_95_153
timestamp 1679235063
transform 1 0 15180 0 -1 54400
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_95_161
timestamp 1679235063
transform 1 0 15916 0 -1 54400
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_95_165
timestamp 1679235063
transform 1 0 16284 0 -1 54400
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_95_169
timestamp 1679235063
transform 1 0 16652 0 -1 54400
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_95_175
timestamp 1679235063
transform 1 0 17204 0 -1 54400
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_95_183
timestamp 1679235063
transform 1 0 17940 0 -1 54400
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_95_191
timestamp 1679235063
transform 1 0 18676 0 -1 54400
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_95_195
timestamp 1679235063
transform 1 0 19044 0 -1 54400
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_95_197
timestamp 1679235063
transform 1 0 19228 0 -1 54400
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_95_203
timestamp 1679235063
transform 1 0 19780 0 -1 54400
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_95_211
timestamp 1679235063
transform 1 0 20516 0 -1 54400
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_95_219
timestamp 1679235063
transform 1 0 21252 0 -1 54400
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_95_223
timestamp 1679235063
transform 1 0 21620 0 -1 54400
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_95_225
timestamp 1679235063
transform 1 0 21804 0 -1 54400
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_95_231
timestamp 1679235063
transform 1 0 22356 0 -1 54400
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_95_239
timestamp 1679235063
transform 1 0 23092 0 -1 54400
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_95_243
timestamp 1679235063
transform 1 0 23460 0 -1 54400
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_95_250
timestamp 1679235063
transform 1 0 24104 0 -1 54400
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_95_257
timestamp 1679235063
transform 1 0 24748 0 -1 54400
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_95_264
timestamp 1679235063
transform 1 0 25392 0 -1 54400
box -38 -48 222 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold1 pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1679235063
transform 1 0 19412 0 1 46784
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold2
timestamp 1679235063
transform 1 0 7728 0 -1 39168
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold3
timestamp 1679235063
transform 1 0 15364 0 -1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold4
timestamp 1679235063
transform 1 0 17940 0 1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold5
timestamp 1679235063
transform 1 0 19780 0 1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold6
timestamp 1679235063
transform 1 0 7912 0 -1 41344
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold7
timestamp 1679235063
transform 1 0 14260 0 1 43520
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold8
timestamp 1679235063
transform 1 0 13064 0 1 44608
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold9
timestamp 1679235063
transform 1 0 20516 0 -1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold10
timestamp 1679235063
transform 1 0 20608 0 -1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold11
timestamp 1679235063
transform 1 0 14812 0 1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold12
timestamp 1679235063
transform 1 0 9660 0 1 30464
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold13
timestamp 1679235063
transform 1 0 16836 0 1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold14
timestamp 1679235063
transform 1 0 18216 0 1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold15
timestamp 1679235063
transform 1 0 11684 0 -1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold16
timestamp 1679235063
transform 1 0 13432 0 -1 39168
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold17
timestamp 1679235063
transform 1 0 15640 0 -1 31552
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold18
timestamp 1679235063
transform 1 0 5336 0 -1 39168
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold19
timestamp 1679235063
transform 1 0 16836 0 -1 40256
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold20
timestamp 1679235063
transform 1 0 20148 0 -1 44608
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold21
timestamp 1679235063
transform 1 0 4784 0 1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold22
timestamp 1679235063
transform 1 0 12972 0 1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold23
timestamp 1679235063
transform 1 0 6532 0 -1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold24
timestamp 1679235063
transform 1 0 4232 0 1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold25
timestamp 1679235063
transform 1 0 16836 0 -1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold26
timestamp 1679235063
transform 1 0 21068 0 1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold27
timestamp 1679235063
transform 1 0 20884 0 1 43520
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold28
timestamp 1679235063
transform 1 0 9384 0 1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold29
timestamp 1679235063
transform 1 0 12328 0 1 46784
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold30
timestamp 1679235063
transform 1 0 10212 0 -1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold31
timestamp 1679235063
transform 1 0 20148 0 -1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold32
timestamp 1679235063
transform 1 0 14260 0 1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold33
timestamp 1679235063
transform 1 0 5796 0 1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold34
timestamp 1679235063
transform 1 0 18216 0 1 34816
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold35
timestamp 1679235063
transform 1 0 24564 0 1 34816
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold36
timestamp 1679235063
transform 1 0 8188 0 -1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold37
timestamp 1679235063
transform 1 0 15640 0 -1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold38
timestamp 1679235063
transform 1 0 7820 0 1 42432
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold39
timestamp 1679235063
transform 1 0 20516 0 1 46784
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold40
timestamp 1679235063
transform 1 0 17112 0 1 47872
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold41
timestamp 1679235063
transform 1 0 21988 0 -1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold42
timestamp 1679235063
transform 1 0 14260 0 1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold43
timestamp 1679235063
transform 1 0 20792 0 -1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold44
timestamp 1679235063
transform 1 0 21528 0 1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold45
timestamp 1679235063
transform 1 0 23368 0 1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold46
timestamp 1679235063
transform 1 0 15456 0 -1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold47
timestamp 1679235063
transform 1 0 18492 0 -1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold48
timestamp 1679235063
transform 1 0 16008 0 1 30464
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold49
timestamp 1679235063
transform 1 0 16100 0 1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold50
timestamp 1679235063
transform 1 0 24564 0 1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold51
timestamp 1679235063
transform 1 0 16836 0 -1 45696
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold52
timestamp 1679235063
transform 1 0 23368 0 1 31552
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold53
timestamp 1679235063
transform 1 0 24656 0 1 42432
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold54
timestamp 1679235063
transform 1 0 14260 0 1 34816
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold55
timestamp 1679235063
transform 1 0 20608 0 -1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold56
timestamp 1679235063
transform 1 0 4876 0 -1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold57
timestamp 1679235063
transform 1 0 11684 0 -1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold58
timestamp 1679235063
transform 1 0 24564 0 -1 39168
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold59
timestamp 1679235063
transform 1 0 7084 0 -1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold60
timestamp 1679235063
transform 1 0 22540 0 1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold61
timestamp 1679235063
transform 1 0 8832 0 -1 30464
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold62
timestamp 1679235063
transform 1 0 7544 0 -1 33728
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold63
timestamp 1679235063
transform 1 0 9108 0 1 33728
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold64
timestamp 1679235063
transform 1 0 24564 0 1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold65
timestamp 1679235063
transform 1 0 18216 0 -1 36992
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold66
timestamp 1679235063
transform 1 0 6624 0 1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold67
timestamp 1679235063
transform 1 0 24564 0 1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold68
timestamp 1679235063
transform 1 0 24564 0 1 45696
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold69
timestamp 1679235063
transform 1 0 7912 0 1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold70
timestamp 1679235063
transform 1 0 7452 0 1 39168
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold71
timestamp 1679235063
transform 1 0 10488 0 -1 46784
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold72
timestamp 1679235063
transform 1 0 20884 0 1 33728
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold73
timestamp 1679235063
transform 1 0 17296 0 -1 34816
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold74
timestamp 1679235063
transform 1 0 17940 0 1 40256
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold75
timestamp 1679235063
transform 1 0 5152 0 1 34816
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold76
timestamp 1679235063
transform 1 0 11776 0 -1 34816
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold77
timestamp 1679235063
transform 1 0 6716 0 1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold78
timestamp 1679235063
transform 1 0 18216 0 1 44608
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold79
timestamp 1679235063
transform 1 0 19412 0 1 43520
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold80
timestamp 1679235063
transform 1 0 15456 0 1 32640
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold81
timestamp 1679235063
transform 1 0 15456 0 -1 32640
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold82
timestamp 1679235063
transform 1 0 11868 0 -1 36992
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold83
timestamp 1679235063
transform 1 0 14628 0 -1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold84
timestamp 1679235063
transform 1 0 15824 0 1 45696
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold85
timestamp 1679235063
transform 1 0 12696 0 1 41344
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold86
timestamp 1679235063
transform 1 0 9108 0 1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold87
timestamp 1679235063
transform 1 0 24564 0 1 40256
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold88
timestamp 1679235063
transform 1 0 6992 0 -1 35904
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold89
timestamp 1679235063
transform 1 0 19044 0 -1 44608
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold90
timestamp 1679235063
transform 1 0 7084 0 -1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold91
timestamp 1679235063
transform 1 0 9752 0 1 42432
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold92
timestamp 1679235063
transform 1 0 22356 0 -1 42432
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s50_1  hold93 pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1679235063
transform 1 0 15456 0 1 40256
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold94
timestamp 1679235063
transform 1 0 5336 0 -1 38080
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold95
timestamp 1679235063
transform 1 0 5336 0 -1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold96
timestamp 1679235063
transform 1 0 24564 0 1 44608
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold97
timestamp 1679235063
transform 1 0 11868 0 1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold98
timestamp 1679235063
transform 1 0 11592 0 1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold99
timestamp 1679235063
transform 1 0 14260 0 1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold100
timestamp 1679235063
transform 1 0 11500 0 1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold101
timestamp 1679235063
transform 1 0 17848 0 1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold102
timestamp 1679235063
transform 1 0 19780 0 1 33728
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold103
timestamp 1679235063
transform 1 0 24564 0 1 36992
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold104
timestamp 1679235063
transform 1 0 7912 0 1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold105
timestamp 1679235063
transform 1 0 23368 0 1 36992
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold106
timestamp 1679235063
transform 1 0 17664 0 1 39168
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold107
timestamp 1679235063
transform 1 0 19412 0 1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold108
timestamp 1679235063
transform 1 0 10212 0 -1 32640
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold109
timestamp 1679235063
transform 1 0 24564 0 1 41344
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold110
timestamp 1679235063
transform 1 0 15364 0 1 43520
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold111
timestamp 1679235063
transform 1 0 19412 0 -1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold112
timestamp 1679235063
transform 1 0 11684 0 -1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold113
timestamp 1679235063
transform 1 0 7912 0 1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold114
timestamp 1679235063
transform 1 0 23276 0 1 43520
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold115
timestamp 1679235063
transform 1 0 6348 0 1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__clkbuf_1  input1
timestamp 1679235063
transform 1 0 1564 0 -1 53312
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input2
timestamp 1679235063
transform 1 0 1564 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input3
timestamp 1679235063
transform 1 0 22356 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input4
timestamp 1679235063
transform 1 0 25116 0 -1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input5
timestamp 1679235063
transform 1 0 25116 0 1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input6
timestamp 1679235063
transform 1 0 25116 0 -1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input7
timestamp 1679235063
transform 1 0 22724 0 1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input8
timestamp 1679235063
transform 1 0 22172 0 -1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input9
timestamp 1679235063
transform 1 0 25116 0 -1 41344
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input10
timestamp 1679235063
transform 1 0 23828 0 1 40256
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input11
timestamp 1679235063
transform 1 0 23828 0 1 41344
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input12
timestamp 1679235063
transform 1 0 25116 0 1 43520
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input13
timestamp 1679235063
transform 1 0 21252 0 -1 42432
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input14
timestamp 1679235063
transform 1 0 21252 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input15
timestamp 1679235063
transform 1 0 23184 0 1 42432
box -38 -48 958 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input16
timestamp 1679235063
transform 1 0 24472 0 -1 44608
box -38 -48 958 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input17
timestamp 1679235063
transform 1 0 24472 0 -1 45696
box -38 -48 958 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input18
timestamp 1679235063
transform 1 0 24472 0 -1 46784
box -38 -48 958 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input19
timestamp 1679235063
transform 1 0 23184 0 1 46784
box -38 -48 958 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input20
timestamp 1679235063
transform 1 0 24472 0 -1 48960
box -38 -48 958 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input21
timestamp 1679235063
transform 1 0 24472 0 -1 47872
box -38 -48 958 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input22
timestamp 1679235063
transform 1 0 24472 0 -1 50048
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_1  input23
timestamp 1679235063
transform 1 0 25116 0 1 48960
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input24
timestamp 1679235063
transform 1 0 25116 0 1 50048
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input25
timestamp 1679235063
transform 1 0 23920 0 -1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input26
timestamp 1679235063
transform 1 0 23828 0 1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input27
timestamp 1679235063
transform 1 0 25116 0 1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input28
timestamp 1679235063
transform 1 0 25116 0 1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input29
timestamp 1679235063
transform 1 0 25116 0 -1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input30
timestamp 1679235063
transform 1 0 25116 0 1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input31
timestamp 1679235063
transform 1 0 25116 0 1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input32
timestamp 1679235063
transform 1 0 25116 0 -1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input33
timestamp 1679235063
transform 1 0 1748 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  input34 pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1679235063
transform 1 0 4968 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  input35
timestamp 1679235063
transform 1 0 5704 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  input36
timestamp 1679235063
transform 1 0 5888 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  input37
timestamp 1679235063
transform 1 0 6532 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  input38
timestamp 1679235063
transform 1 0 6808 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  input39
timestamp 1679235063
transform 1 0 6900 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input40
timestamp 1679235063
transform 1 0 7636 0 1 2176
box -38 -48 958 592
use sky130_fd_sc_hd__buf_2  input41
timestamp 1679235063
transform 1 0 8004 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  input42
timestamp 1679235063
transform 1 0 7544 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  input43
timestamp 1679235063
transform 1 0 8280 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input44
timestamp 1679235063
transform 1 0 1748 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input45
timestamp 1679235063
transform 1 0 9016 0 -1 3264
box -38 -48 958 592
use sky130_fd_sc_hd__buf_2  input46
timestamp 1679235063
transform 1 0 9108 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  input47
timestamp 1679235063
transform 1 0 9844 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  input48
timestamp 1679235063
transform 1 0 9568 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input49
timestamp 1679235063
transform 1 0 10304 0 -1 3264
box -38 -48 958 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input50
timestamp 1679235063
transform 1 0 10948 0 1 3264
box -38 -48 958 592
use sky130_fd_sc_hd__buf_2  input51
timestamp 1679235063
transform 1 0 11684 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input52
timestamp 1679235063
transform 1 0 11684 0 -1 4352
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_1  input53
timestamp 1679235063
transform 1 0 11684 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input54
timestamp 1679235063
transform 1 0 10304 0 1 2176
box -38 -48 958 592
use sky130_fd_sc_hd__buf_2  input55
timestamp 1679235063
transform 1 0 1656 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  input56
timestamp 1679235063
transform 1 0 2484 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input57
timestamp 1679235063
transform 1 0 3220 0 -1 3264
box -38 -48 958 592
use sky130_fd_sc_hd__buf_2  input58
timestamp 1679235063
transform 1 0 2392 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input59
timestamp 1679235063
transform 1 0 3128 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  input60
timestamp 1679235063
transform 1 0 3956 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input61
timestamp 1679235063
transform 1 0 4692 0 1 2176
box -38 -48 958 592
use sky130_fd_sc_hd__buf_2  input62
timestamp 1679235063
transform 1 0 5060 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  input63
timestamp 1679235063
transform 1 0 11684 0 -1 54400
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  input64
timestamp 1679235063
transform 1 0 16652 0 1 53312
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  input65
timestamp 1679235063
transform 1 0 17572 0 -1 54400
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  input66
timestamp 1679235063
transform 1 0 17388 0 1 53312
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  input67
timestamp 1679235063
transform 1 0 18308 0 -1 54400
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input68
timestamp 1679235063
transform 1 0 18124 0 1 53312
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  input69
timestamp 1679235063
transform 1 0 19412 0 -1 54400
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  input70
timestamp 1679235063
transform 1 0 18860 0 -1 53312
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  input71
timestamp 1679235063
transform 1 0 19412 0 1 53312
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  input72
timestamp 1679235063
transform 1 0 20148 0 -1 54400
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input73
timestamp 1679235063
transform 1 0 20148 0 1 53312
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input74
timestamp 1679235063
transform 1 0 13340 0 1 52224
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  input75
timestamp 1679235063
transform 1 0 20332 0 -1 53312
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  input76
timestamp 1679235063
transform 1 0 20884 0 -1 54400
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  input77
timestamp 1679235063
transform 1 0 21068 0 1 53312
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  input78
timestamp 1679235063
transform 1 0 21988 0 -1 54400
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  input79
timestamp 1679235063
transform 1 0 21804 0 1 53312
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input80
timestamp 1679235063
transform 1 0 22448 0 1 53312
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  input81
timestamp 1679235063
transform 1 0 22724 0 -1 54400
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  input82
timestamp 1679235063
transform 1 0 23092 0 1 53312
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input83
timestamp 1679235063
transform 1 0 23276 0 -1 53312
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input84
timestamp 1679235063
transform 1 0 23920 0 -1 53312
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  input85
timestamp 1679235063
transform 1 0 13708 0 -1 53312
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  input86
timestamp 1679235063
transform 1 0 14260 0 1 53312
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  input87
timestamp 1679235063
transform 1 0 14444 0 -1 53312
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  input88
timestamp 1679235063
transform 1 0 14812 0 -1 54400
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  input89
timestamp 1679235063
transform 1 0 15548 0 -1 54400
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input90
timestamp 1679235063
transform 1 0 15548 0 1 53312
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  input91
timestamp 1679235063
transform 1 0 15916 0 -1 53312
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  input92
timestamp 1679235063
transform 1 0 16836 0 -1 54400
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  input93
timestamp 1679235063
transform 1 0 1564 0 -1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input94
timestamp 1679235063
transform 1 0 1564 0 1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input95
timestamp 1679235063
transform 1 0 1564 0 1 38080
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input96
timestamp 1679235063
transform 1 0 1564 0 -1 41344
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  input97
timestamp 1679235063
transform 1 0 1564 0 -1 43520
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_16  input98
timestamp 1679235063
transform 1 0 23552 0 -1 3264
box -38 -48 1878 592
use sky130_fd_sc_hd__buf_2  input99
timestamp 1679235063
transform 1 0 25024 0 -1 51136
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  input100
timestamp 1679235063
transform 1 0 25024 0 1 51136
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  input101
timestamp 1679235063
transform 1 0 25024 0 1 52224
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  input102
timestamp 1679235063
transform 1 0 25024 0 -1 53312
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  input103
timestamp 1679235063
transform 1 0 25024 0 -1 54400
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  input104 pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1679235063
transform 1 0 24840 0 1 53312
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  input105
timestamp 1679235063
transform 1 0 23736 0 -1 54400
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input106
timestamp 1679235063
transform 1 0 23736 0 1 53312
box -38 -48 406 592
use sky130_fd_sc_hd__conb_1  left_tile_202
timestamp 1679235063
transform 1 0 25116 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__buf_12  output107 pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1679235063
transform 1 0 18216 0 -1 6528
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output108
timestamp 1679235063
transform 1 0 1564 0 1 48960
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output109
timestamp 1679235063
transform 1 0 22632 0 1 9792
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output110
timestamp 1679235063
transform 1 0 23920 0 -1 9792
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output111
timestamp 1679235063
transform 1 0 23920 0 -1 10880
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output112
timestamp 1679235063
transform 1 0 23920 0 -1 11968
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output113
timestamp 1679235063
transform 1 0 22632 0 1 13056
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output114
timestamp 1679235063
transform 1 0 23920 0 -1 13056
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output115
timestamp 1679235063
transform 1 0 23920 0 -1 14144
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output116
timestamp 1679235063
transform 1 0 22632 0 1 15232
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output117
timestamp 1679235063
transform 1 0 23920 0 -1 15232
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output118
timestamp 1679235063
transform 1 0 23920 0 -1 16320
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output119
timestamp 1679235063
transform 1 0 20056 0 -1 7616
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output120
timestamp 1679235063
transform 1 0 22080 0 -1 18496
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output121
timestamp 1679235063
transform 1 0 23920 0 -1 17408
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output122
timestamp 1679235063
transform 1 0 23920 0 -1 18496
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output123
timestamp 1679235063
transform 1 0 22632 0 1 19584
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output124
timestamp 1679235063
transform 1 0 22080 0 -1 20672
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output125
timestamp 1679235063
transform 1 0 22632 0 1 20672
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output126
timestamp 1679235063
transform 1 0 23920 0 -1 20672
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output127
timestamp 1679235063
transform 1 0 22632 0 1 22848
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output128
timestamp 1679235063
transform 1 0 22632 0 1 23936
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output129
timestamp 1679235063
transform 1 0 23920 0 -1 26112
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output130
timestamp 1679235063
transform 1 0 22080 0 -1 8704
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output131
timestamp 1679235063
transform 1 0 17572 0 -1 5440
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output132
timestamp 1679235063
transform 1 0 22632 0 1 7616
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output133
timestamp 1679235063
transform 1 0 23920 0 -1 5440
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output134
timestamp 1679235063
transform 1 0 22632 0 1 6528
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output135
timestamp 1679235063
transform 1 0 23920 0 -1 6528
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output136
timestamp 1679235063
transform 1 0 23920 0 -1 7616
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output137
timestamp 1679235063
transform 1 0 23920 0 -1 8704
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output138
timestamp 1679235063
transform 1 0 12328 0 1 3264
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output139
timestamp 1679235063
transform 1 0 16836 0 -1 4352
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output140
timestamp 1679235063
transform 1 0 19412 0 1 2176
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output141
timestamp 1679235063
transform 1 0 18676 0 -1 3264
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output142
timestamp 1679235063
transform 1 0 18676 0 -1 4352
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output143
timestamp 1679235063
transform 1 0 19412 0 1 3264
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output144
timestamp 1679235063
transform 1 0 21988 0 1 2176
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output145
timestamp 1679235063
transform 1 0 19412 0 1 4352
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output146
timestamp 1679235063
transform 1 0 21252 0 1 3264
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output147
timestamp 1679235063
transform 1 0 19412 0 -1 5440
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output148
timestamp 1679235063
transform 1 0 21252 0 1 4352
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output149
timestamp 1679235063
transform 1 0 12420 0 -1 3264
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output150
timestamp 1679235063
transform 1 0 21988 0 -1 4352
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output151
timestamp 1679235063
transform 1 0 20516 0 1 5440
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output152
timestamp 1679235063
transform 1 0 21988 0 -1 5440
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output153
timestamp 1679235063
transform 1 0 23828 0 -1 4352
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output154
timestamp 1679235063
transform 1 0 22356 0 1 5440
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output155
timestamp 1679235063
transform 1 0 21988 0 -1 6528
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output156
timestamp 1679235063
transform 1 0 22080 0 -1 7616
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output157
timestamp 1679235063
transform 1 0 20056 0 -1 6528
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output158
timestamp 1679235063
transform 1 0 20792 0 1 6528
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output159
timestamp 1679235063
transform 1 0 17480 0 1 4352
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output160
timestamp 1679235063
transform 1 0 13524 0 -1 4352
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output161
timestamp 1679235063
transform 1 0 12328 0 1 2176
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output162
timestamp 1679235063
transform 1 0 14260 0 -1 3264
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output163
timestamp 1679235063
transform 1 0 14628 0 1 2176
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output164
timestamp 1679235063
transform 1 0 14996 0 1 3264
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output165
timestamp 1679235063
transform 1 0 16836 0 1 2176
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output166
timestamp 1679235063
transform 1 0 16836 0 -1 3264
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output167
timestamp 1679235063
transform 1 0 16836 0 1 3264
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output168
timestamp 1679235063
transform 1 0 1932 0 -1 50048
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output169
timestamp 1679235063
transform 1 0 2024 0 1 53312
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output170
timestamp 1679235063
transform 1 0 2024 0 -1 54400
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output171
timestamp 1679235063
transform 1 0 4600 0 -1 53312
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output172
timestamp 1679235063
transform 1 0 5336 0 1 52224
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output173
timestamp 1679235063
transform 1 0 7084 0 1 51136
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output174
timestamp 1679235063
transform 1 0 5336 0 1 53312
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output175
timestamp 1679235063
transform 1 0 7176 0 1 52224
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output176
timestamp 1679235063
transform 1 0 4600 0 -1 54400
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output177
timestamp 1679235063
transform 1 0 7820 0 -1 52224
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output178
timestamp 1679235063
transform 1 0 7176 0 1 53312
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output179
timestamp 1679235063
transform 1 0 2024 0 1 50048
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output180
timestamp 1679235063
transform 1 0 7912 0 -1 53312
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output181
timestamp 1679235063
transform 1 0 9660 0 -1 52224
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output182
timestamp 1679235063
transform 1 0 7176 0 -1 54400
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output183
timestamp 1679235063
transform 1 0 9752 0 -1 53312
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output184
timestamp 1679235063
transform 1 0 10764 0 1 52224
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output185
timestamp 1679235063
transform 1 0 10396 0 1 53312
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output186
timestamp 1679235063
transform 1 0 9752 0 -1 54400
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output187
timestamp 1679235063
transform 1 0 11868 0 -1 53312
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output188
timestamp 1679235063
transform 1 0 12236 0 1 53312
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output189
timestamp 1679235063
transform 1 0 12328 0 -1 54400
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output190
timestamp 1679235063
transform 1 0 2300 0 -1 51136
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output191
timestamp 1679235063
transform 1 0 2024 0 1 51136
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output192
timestamp 1679235063
transform 1 0 2760 0 -1 52224
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output193
timestamp 1679235063
transform 1 0 2024 0 1 52224
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output194
timestamp 1679235063
transform 1 0 4140 0 -1 51136
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output195
timestamp 1679235063
transform 1 0 2760 0 -1 53312
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output196
timestamp 1679235063
transform 1 0 4600 0 -1 52224
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output197
timestamp 1679235063
transform 1 0 5244 0 1 51136
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output198
timestamp 1679235063
transform 1 0 1564 0 -1 14144
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output199
timestamp 1679235063
transform 1 0 1564 0 1 16320
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output200
timestamp 1679235063
transform 1 0 1564 0 1 18496
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output201
timestamp 1679235063
transform 1 0 1564 0 1 20672
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_3  PHY_0
timestamp 1679235063
transform 1 0 1104 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_1
timestamp 1679235063
transform -1 0 25852 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_2
timestamp 1679235063
transform 1 0 1104 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_3
timestamp 1679235063
transform -1 0 25852 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_4
timestamp 1679235063
transform 1 0 1104 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_5
timestamp 1679235063
transform -1 0 25852 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_6
timestamp 1679235063
transform 1 0 1104 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_7
timestamp 1679235063
transform -1 0 25852 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_8
timestamp 1679235063
transform 1 0 1104 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_9
timestamp 1679235063
transform -1 0 25852 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_10
timestamp 1679235063
transform 1 0 1104 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_11
timestamp 1679235063
transform -1 0 25852 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_12
timestamp 1679235063
transform 1 0 1104 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_13
timestamp 1679235063
transform -1 0 25852 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_14
timestamp 1679235063
transform 1 0 1104 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_15
timestamp 1679235063
transform -1 0 25852 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_16
timestamp 1679235063
transform 1 0 1104 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_17
timestamp 1679235063
transform -1 0 25852 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_18
timestamp 1679235063
transform 1 0 1104 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_19
timestamp 1679235063
transform -1 0 25852 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_20
timestamp 1679235063
transform 1 0 1104 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_21
timestamp 1679235063
transform -1 0 25852 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_22
timestamp 1679235063
transform 1 0 1104 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_23
timestamp 1679235063
transform -1 0 25852 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_24
timestamp 1679235063
transform 1 0 1104 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_25
timestamp 1679235063
transform -1 0 25852 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_26
timestamp 1679235063
transform 1 0 1104 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_27
timestamp 1679235063
transform -1 0 25852 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_28
timestamp 1679235063
transform 1 0 1104 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_29
timestamp 1679235063
transform -1 0 25852 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_30
timestamp 1679235063
transform 1 0 1104 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_31
timestamp 1679235063
transform -1 0 25852 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_32
timestamp 1679235063
transform 1 0 1104 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_33
timestamp 1679235063
transform -1 0 25852 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_34
timestamp 1679235063
transform 1 0 1104 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_35
timestamp 1679235063
transform -1 0 25852 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_36
timestamp 1679235063
transform 1 0 1104 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_37
timestamp 1679235063
transform -1 0 25852 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_38
timestamp 1679235063
transform 1 0 1104 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_39
timestamp 1679235063
transform -1 0 25852 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_40
timestamp 1679235063
transform 1 0 1104 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_41
timestamp 1679235063
transform -1 0 25852 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_42
timestamp 1679235063
transform 1 0 1104 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_43
timestamp 1679235063
transform -1 0 25852 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_44
timestamp 1679235063
transform 1 0 1104 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_45
timestamp 1679235063
transform -1 0 25852 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_46
timestamp 1679235063
transform 1 0 1104 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_47
timestamp 1679235063
transform -1 0 25852 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_48
timestamp 1679235063
transform 1 0 1104 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_49
timestamp 1679235063
transform -1 0 25852 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_50
timestamp 1679235063
transform 1 0 1104 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_51
timestamp 1679235063
transform -1 0 25852 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_52
timestamp 1679235063
transform 1 0 1104 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_53
timestamp 1679235063
transform -1 0 25852 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_54
timestamp 1679235063
transform 1 0 1104 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_55
timestamp 1679235063
transform -1 0 25852 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_56
timestamp 1679235063
transform 1 0 1104 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_57
timestamp 1679235063
transform -1 0 25852 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_58
timestamp 1679235063
transform 1 0 1104 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_59
timestamp 1679235063
transform -1 0 25852 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_60
timestamp 1679235063
transform 1 0 1104 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_61
timestamp 1679235063
transform -1 0 25852 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_62
timestamp 1679235063
transform 1 0 1104 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_63
timestamp 1679235063
transform -1 0 25852 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_64
timestamp 1679235063
transform 1 0 1104 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_65
timestamp 1679235063
transform -1 0 25852 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_66
timestamp 1679235063
transform 1 0 1104 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_67
timestamp 1679235063
transform -1 0 25852 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_68
timestamp 1679235063
transform 1 0 1104 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_69
timestamp 1679235063
transform -1 0 25852 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_70
timestamp 1679235063
transform 1 0 1104 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_71
timestamp 1679235063
transform -1 0 25852 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_72
timestamp 1679235063
transform 1 0 1104 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_73
timestamp 1679235063
transform -1 0 25852 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_74
timestamp 1679235063
transform 1 0 1104 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_75
timestamp 1679235063
transform -1 0 25852 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_76
timestamp 1679235063
transform 1 0 1104 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_77
timestamp 1679235063
transform -1 0 25852 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_78
timestamp 1679235063
transform 1 0 1104 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_79
timestamp 1679235063
transform -1 0 25852 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_80
timestamp 1679235063
transform 1 0 1104 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_81
timestamp 1679235063
transform -1 0 25852 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_82
timestamp 1679235063
transform 1 0 1104 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_83
timestamp 1679235063
transform -1 0 25852 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_84
timestamp 1679235063
transform 1 0 1104 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_85
timestamp 1679235063
transform -1 0 25852 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_86
timestamp 1679235063
transform 1 0 1104 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_87
timestamp 1679235063
transform -1 0 25852 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_88
timestamp 1679235063
transform 1 0 1104 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_89
timestamp 1679235063
transform -1 0 25852 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_90
timestamp 1679235063
transform 1 0 1104 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_91
timestamp 1679235063
transform -1 0 25852 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_92
timestamp 1679235063
transform 1 0 1104 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_93
timestamp 1679235063
transform -1 0 25852 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_94
timestamp 1679235063
transform 1 0 1104 0 -1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_95
timestamp 1679235063
transform -1 0 25852 0 -1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_96
timestamp 1679235063
transform 1 0 1104 0 1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_97
timestamp 1679235063
transform -1 0 25852 0 1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_98
timestamp 1679235063
transform 1 0 1104 0 -1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_99
timestamp 1679235063
transform -1 0 25852 0 -1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_100
timestamp 1679235063
transform 1 0 1104 0 1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_101
timestamp 1679235063
transform -1 0 25852 0 1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_102
timestamp 1679235063
transform 1 0 1104 0 -1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_103
timestamp 1679235063
transform -1 0 25852 0 -1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_104
timestamp 1679235063
transform 1 0 1104 0 1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_105
timestamp 1679235063
transform -1 0 25852 0 1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_106
timestamp 1679235063
transform 1 0 1104 0 -1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_107
timestamp 1679235063
transform -1 0 25852 0 -1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_108
timestamp 1679235063
transform 1 0 1104 0 1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_109
timestamp 1679235063
transform -1 0 25852 0 1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_110
timestamp 1679235063
transform 1 0 1104 0 -1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_111
timestamp 1679235063
transform -1 0 25852 0 -1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_112
timestamp 1679235063
transform 1 0 1104 0 1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_113
timestamp 1679235063
transform -1 0 25852 0 1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_114
timestamp 1679235063
transform 1 0 1104 0 -1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_115
timestamp 1679235063
transform -1 0 25852 0 -1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_116
timestamp 1679235063
transform 1 0 1104 0 1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_117
timestamp 1679235063
transform -1 0 25852 0 1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_118
timestamp 1679235063
transform 1 0 1104 0 -1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_119
timestamp 1679235063
transform -1 0 25852 0 -1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_120
timestamp 1679235063
transform 1 0 1104 0 1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_121
timestamp 1679235063
transform -1 0 25852 0 1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_122
timestamp 1679235063
transform 1 0 1104 0 -1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_123
timestamp 1679235063
transform -1 0 25852 0 -1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_124
timestamp 1679235063
transform 1 0 1104 0 1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_125
timestamp 1679235063
transform -1 0 25852 0 1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_126
timestamp 1679235063
transform 1 0 1104 0 -1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_127
timestamp 1679235063
transform -1 0 25852 0 -1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_128
timestamp 1679235063
transform 1 0 1104 0 1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_129
timestamp 1679235063
transform -1 0 25852 0 1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_130
timestamp 1679235063
transform 1 0 1104 0 -1 38080
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_131
timestamp 1679235063
transform -1 0 25852 0 -1 38080
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_132
timestamp 1679235063
transform 1 0 1104 0 1 38080
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_133
timestamp 1679235063
transform -1 0 25852 0 1 38080
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_134
timestamp 1679235063
transform 1 0 1104 0 -1 39168
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_135
timestamp 1679235063
transform -1 0 25852 0 -1 39168
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_136
timestamp 1679235063
transform 1 0 1104 0 1 39168
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_137
timestamp 1679235063
transform -1 0 25852 0 1 39168
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_138
timestamp 1679235063
transform 1 0 1104 0 -1 40256
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_139
timestamp 1679235063
transform -1 0 25852 0 -1 40256
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_140
timestamp 1679235063
transform 1 0 1104 0 1 40256
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_141
timestamp 1679235063
transform -1 0 25852 0 1 40256
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_142
timestamp 1679235063
transform 1 0 1104 0 -1 41344
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_143
timestamp 1679235063
transform -1 0 25852 0 -1 41344
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_144
timestamp 1679235063
transform 1 0 1104 0 1 41344
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_145
timestamp 1679235063
transform -1 0 25852 0 1 41344
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_146
timestamp 1679235063
transform 1 0 1104 0 -1 42432
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_147
timestamp 1679235063
transform -1 0 25852 0 -1 42432
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_148
timestamp 1679235063
transform 1 0 1104 0 1 42432
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_149
timestamp 1679235063
transform -1 0 25852 0 1 42432
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_150
timestamp 1679235063
transform 1 0 1104 0 -1 43520
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_151
timestamp 1679235063
transform -1 0 25852 0 -1 43520
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_152
timestamp 1679235063
transform 1 0 1104 0 1 43520
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_153
timestamp 1679235063
transform -1 0 25852 0 1 43520
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_154
timestamp 1679235063
transform 1 0 1104 0 -1 44608
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_155
timestamp 1679235063
transform -1 0 25852 0 -1 44608
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_156
timestamp 1679235063
transform 1 0 1104 0 1 44608
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_157
timestamp 1679235063
transform -1 0 25852 0 1 44608
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_158
timestamp 1679235063
transform 1 0 1104 0 -1 45696
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_159
timestamp 1679235063
transform -1 0 25852 0 -1 45696
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_160
timestamp 1679235063
transform 1 0 1104 0 1 45696
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_161
timestamp 1679235063
transform -1 0 25852 0 1 45696
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_162
timestamp 1679235063
transform 1 0 1104 0 -1 46784
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_163
timestamp 1679235063
transform -1 0 25852 0 -1 46784
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_164
timestamp 1679235063
transform 1 0 1104 0 1 46784
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_165
timestamp 1679235063
transform -1 0 25852 0 1 46784
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_166
timestamp 1679235063
transform 1 0 1104 0 -1 47872
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_167
timestamp 1679235063
transform -1 0 25852 0 -1 47872
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_168
timestamp 1679235063
transform 1 0 1104 0 1 47872
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_169
timestamp 1679235063
transform -1 0 25852 0 1 47872
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_170
timestamp 1679235063
transform 1 0 1104 0 -1 48960
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_171
timestamp 1679235063
transform -1 0 25852 0 -1 48960
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_172
timestamp 1679235063
transform 1 0 1104 0 1 48960
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_173
timestamp 1679235063
transform -1 0 25852 0 1 48960
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_174
timestamp 1679235063
transform 1 0 1104 0 -1 50048
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_175
timestamp 1679235063
transform -1 0 25852 0 -1 50048
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_176
timestamp 1679235063
transform 1 0 1104 0 1 50048
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_177
timestamp 1679235063
transform -1 0 25852 0 1 50048
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_178
timestamp 1679235063
transform 1 0 1104 0 -1 51136
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_179
timestamp 1679235063
transform -1 0 25852 0 -1 51136
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_180
timestamp 1679235063
transform 1 0 1104 0 1 51136
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_181
timestamp 1679235063
transform -1 0 25852 0 1 51136
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_182
timestamp 1679235063
transform 1 0 1104 0 -1 52224
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_183
timestamp 1679235063
transform -1 0 25852 0 -1 52224
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_184
timestamp 1679235063
transform 1 0 1104 0 1 52224
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_185
timestamp 1679235063
transform -1 0 25852 0 1 52224
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_186
timestamp 1679235063
transform 1 0 1104 0 -1 53312
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_187
timestamp 1679235063
transform -1 0 25852 0 -1 53312
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_188
timestamp 1679235063
transform 1 0 1104 0 1 53312
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_189
timestamp 1679235063
transform -1 0 25852 0 1 53312
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_190
timestamp 1679235063
transform 1 0 1104 0 -1 54400
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_191
timestamp 1679235063
transform -1 0 25852 0 -1 54400
box -38 -48 314 592
use sky130_fd_sc_hd__dfrtp_2  sb_0__1_.mem_bottom_track_1.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1679235063
transform 1 0 18952 0 -1 19584
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__1_.mem_bottom_track_1.sky130_fd_sc_hd__dfrtp_1_1_
timestamp 1679235063
transform 1 0 17112 0 1 22848
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__1_.mem_bottom_track_1.sky130_fd_sc_hd__dfrtp_1_2_
timestamp 1679235063
transform 1 0 18308 0 -1 21760
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__1_.mem_bottom_track_3.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1679235063
transform 1 0 19412 0 1 22848
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__1_.mem_bottom_track_3.sky130_fd_sc_hd__dfrtp_1_1_
timestamp 1679235063
transform 1 0 19688 0 -1 23936
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__1_.mem_bottom_track_3.sky130_fd_sc_hd__dfrtp_1_2_
timestamp 1679235063
transform 1 0 19872 0 1 20672
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_2  sb_0__1_.mem_bottom_track_5.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1679235063
transform 1 0 21068 0 1 21760
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__1_.mem_bottom_track_5.sky130_fd_sc_hd__dfrtp_1_1_
timestamp 1679235063
transform 1 0 22816 0 -1 23936
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__1_.mem_bottom_track_5.sky130_fd_sc_hd__dfrtp_1_2_
timestamp 1679235063
transform 1 0 23184 0 -1 21760
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_4  sb_0__1_.mem_bottom_track_7.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1679235063
transform 1 0 22080 0 -1 22848
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__1_.mem_bottom_track_7.sky130_fd_sc_hd__dfrtp_1_1_
timestamp 1679235063
transform 1 0 17296 0 -1 25024
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__1_.mem_bottom_track_7.sky130_fd_sc_hd__dfrtp_1_2_
timestamp 1679235063
transform 1 0 15640 0 1 23936
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_4  sb_0__1_.mem_bottom_track_11.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1679235063
transform 1 0 14260 0 -1 26112
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__1_.mem_bottom_track_11.sky130_fd_sc_hd__dfrtp_1_1_
timestamp 1679235063
transform 1 0 12972 0 -1 28288
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__1_.mem_bottom_track_11.sky130_fd_sc_hd__dfrtp_1_2_
timestamp 1679235063
transform 1 0 13248 0 -1 27200
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_2  sb_0__1_.mem_bottom_track_13.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1679235063
transform 1 0 15364 0 1 27200
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__1_.mem_bottom_track_13.sky130_fd_sc_hd__dfrtp_1_1_
timestamp 1679235063
transform 1 0 19136 0 -1 28288
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__1_.mem_bottom_track_13.sky130_fd_sc_hd__dfrtp_1_2_
timestamp 1679235063
transform 1 0 20332 0 1 25024
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_2  sb_0__1_.mem_bottom_track_21.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1679235063
transform 1 0 21988 0 -1 27200
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__1_.mem_bottom_track_21.sky130_fd_sc_hd__dfrtp_1_1_
timestamp 1679235063
transform 1 0 22264 0 1 27200
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__1_.mem_bottom_track_21.sky130_fd_sc_hd__dfrtp_1_2_
timestamp 1679235063
transform 1 0 23000 0 -1 25024
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_2  sb_0__1_.mem_bottom_track_29.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1679235063
transform 1 0 21988 0 -1 28288
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__1_.mem_bottom_track_29.sky130_fd_sc_hd__dfrtp_1_1_
timestamp 1679235063
transform 1 0 17112 0 1 30464
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__1_.mem_bottom_track_29.sky130_fd_sc_hd__dfrtp_1_2_
timestamp 1679235063
transform 1 0 14536 0 -1 30464
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__1_.mem_bottom_track_37.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1679235063
transform 1 0 15272 0 1 31552
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__1_.mem_bottom_track_37.sky130_fd_sc_hd__dfrtp_1_1_
timestamp 1679235063
transform 1 0 13984 0 -1 33728
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__1_.mem_bottom_track_37.sky130_fd_sc_hd__dfrtp_1_2_
timestamp 1679235063
transform 1 0 12604 0 -1 31552
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__1_.mem_bottom_track_45.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1679235063
transform 1 0 15640 0 1 33728
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__1_.mem_bottom_track_45.sky130_fd_sc_hd__dfrtp_1_1_
timestamp 1679235063
transform 1 0 19412 0 1 34816
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__1_.mem_bottom_track_45.sky130_fd_sc_hd__dfrtp_1_2_
timestamp 1679235063
transform 1 0 18308 0 -1 33728
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__1_.mem_bottom_track_53.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1679235063
transform 1 0 15456 0 1 34816
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_2  sb_0__1_.mem_bottom_track_53.sky130_fd_sc_hd__dfrtp_1_1_
timestamp 1679235063
transform 1 0 9108 0 1 43520
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__1_.mem_right_track_0.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1679235063
transform 1 0 17664 0 -1 35904
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__1_.mem_right_track_0.sky130_fd_sc_hd__dfrtp_1_1_
timestamp 1679235063
transform 1 0 22080 0 -1 31552
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__1_.mem_right_track_0.sky130_fd_sc_hd__dfrtp_1_2_
timestamp 1679235063
transform 1 0 23368 0 -1 30464
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_2  sb_0__1_.mem_right_track_2.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1679235063
transform 1 0 23460 0 -1 33728
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__1_.mem_right_track_2.sky130_fd_sc_hd__dfrtp_1_1_
timestamp 1679235063
transform 1 0 22816 0 -1 41344
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__1_.mem_right_track_2.sky130_fd_sc_hd__dfrtp_1_2_
timestamp 1679235063
transform 1 0 23552 0 -1 43520
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__1_.mem_right_track_4.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1679235063
transform 1 0 23460 0 -1 42432
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__1_.mem_right_track_4.sky130_fd_sc_hd__dfrtp_1_1_
timestamp 1679235063
transform 1 0 22356 0 -1 39168
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__1_.mem_right_track_4.sky130_fd_sc_hd__dfrtp_1_2_
timestamp 1679235063
transform 1 0 22264 0 1 34816
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_2  sb_0__1_.mem_right_track_6.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1679235063
transform 1 0 23184 0 -1 35904
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__1_.mem_right_track_6.sky130_fd_sc_hd__dfrtp_1_1_
timestamp 1679235063
transform 1 0 22816 0 -1 36992
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__1_.mem_right_track_6.sky130_fd_sc_hd__dfrtp_1_2_
timestamp 1679235063
transform 1 0 23552 0 -1 38080
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_2  sb_0__1_.mem_right_track_8.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1679235063
transform 1 0 23368 0 -1 40256
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__1_.mem_right_track_8.sky130_fd_sc_hd__dfrtp_1_1_
timestamp 1679235063
transform 1 0 22264 0 -1 44608
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__1_.mem_right_track_8.sky130_fd_sc_hd__dfrtp_1_2_
timestamp 1679235063
transform 1 0 22264 0 1 44608
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__1_.mem_right_track_10.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1679235063
transform 1 0 22080 0 -1 45696
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__1_.mem_right_track_10.sky130_fd_sc_hd__dfrtp_1_1_
timestamp 1679235063
transform 1 0 19596 0 1 42432
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__1_.mem_right_track_10.sky130_fd_sc_hd__dfrtp_1_2_
timestamp 1679235063
transform 1 0 18768 0 -1 42432
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__1_.mem_right_track_12.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1679235063
transform 1 0 19688 0 1 44608
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__1_.mem_right_track_12.sky130_fd_sc_hd__dfrtp_1_1_
timestamp 1679235063
transform 1 0 19504 0 1 45696
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__1_.mem_right_track_12.sky130_fd_sc_hd__dfrtp_1_2_
timestamp 1679235063
transform 1 0 18216 0 -1 43520
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__1_.mem_right_track_14.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1679235063
transform 1 0 18216 0 -1 45696
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__1_.mem_right_track_14.sky130_fd_sc_hd__dfrtp_1_1_
timestamp 1679235063
transform 1 0 17112 0 1 45696
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__1_.mem_right_track_14.sky130_fd_sc_hd__dfrtp_1_2_
timestamp 1679235063
transform 1 0 16836 0 -1 44608
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__1_.mem_right_track_16.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1679235063
transform 1 0 16836 0 -1 46784
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__1_.mem_right_track_16.sky130_fd_sc_hd__dfrtp_1_1_
timestamp 1679235063
transform 1 0 15732 0 1 46784
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__1_.mem_right_track_16.sky130_fd_sc_hd__dfrtp_1_2_
timestamp 1679235063
transform 1 0 15088 0 1 44608
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__1_.mem_right_track_18.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1679235063
transform 1 0 14536 0 -1 46784
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__1_.mem_right_track_18.sky130_fd_sc_hd__dfrtp_1_1_
timestamp 1679235063
transform 1 0 14352 0 -1 45696
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__1_.mem_right_track_18.sky130_fd_sc_hd__dfrtp_1_2_
timestamp 1679235063
transform 1 0 13800 0 -1 41344
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__1_.mem_right_track_20.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1679235063
transform 1 0 12972 0 -1 40256
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__1_.mem_right_track_20.sky130_fd_sc_hd__dfrtp_1_1_
timestamp 1679235063
transform 1 0 11960 0 1 38080
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__1_.mem_right_track_20.sky130_fd_sc_hd__dfrtp_1_2_
timestamp 1679235063
transform 1 0 11408 0 1 33728
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__1_.mem_right_track_22.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1679235063
transform 1 0 11684 0 -1 35904
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__1_.mem_right_track_22.sky130_fd_sc_hd__dfrtp_1_1_
timestamp 1679235063
transform 1 0 10304 0 1 34816
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__1_.mem_right_track_22.sky130_fd_sc_hd__dfrtp_1_2_
timestamp 1679235063
transform 1 0 9384 0 -1 31552
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__1_.mem_right_track_24.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1679235063
transform 1 0 9660 0 1 29376
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__1_.mem_right_track_24.sky130_fd_sc_hd__dfrtp_1_1_
timestamp 1679235063
transform 1 0 9200 0 -1 28288
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__1_.mem_right_track_26.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1679235063
transform 1 0 9108 0 1 28288
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__1_.mem_right_track_26.sky130_fd_sc_hd__dfrtp_1_1_
timestamp 1679235063
transform 1 0 6992 0 -1 29376
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__1_.mem_right_track_28.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1679235063
transform 1 0 6532 0 -1 28288
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__1_.mem_right_track_28.sky130_fd_sc_hd__dfrtp_1_1_
timestamp 1679235063
transform 1 0 6532 0 -1 27200
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__1_.mem_right_track_30.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1679235063
transform 1 0 6440 0 1 26112
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__1_.mem_right_track_30.sky130_fd_sc_hd__dfrtp_1_1_
timestamp 1679235063
transform 1 0 7452 0 -1 26112
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__1_.mem_right_track_32.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1679235063
transform 1 0 9200 0 1 25024
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__1_.mem_right_track_32.sky130_fd_sc_hd__dfrtp_1_1_
timestamp 1679235063
transform 1 0 10948 0 1 23936
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__1_.mem_right_track_34.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1679235063
transform 1 0 11960 0 1 22848
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__1_.mem_right_track_34.sky130_fd_sc_hd__dfrtp_1_1_
timestamp 1679235063
transform 1 0 14260 0 1 20672
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__1_.mem_right_track_36.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1679235063
transform 1 0 13248 0 -1 20672
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__1_.mem_right_track_36.sky130_fd_sc_hd__dfrtp_1_1_
timestamp 1679235063
transform 1 0 11040 0 1 17408
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__1_.mem_right_track_36.sky130_fd_sc_hd__dfrtp_1_2_
timestamp 1679235063
transform 1 0 8832 0 -1 13056
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__1_.mem_right_track_38.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1679235063
transform 1 0 9568 0 1 11968
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__1_.mem_right_track_38.sky130_fd_sc_hd__dfrtp_1_1_
timestamp 1679235063
transform 1 0 11776 0 1 11968
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__1_.mem_right_track_40.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1679235063
transform 1 0 12972 0 -1 11968
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__1_.mem_right_track_40.sky130_fd_sc_hd__dfrtp_1_1_
timestamp 1679235063
transform 1 0 14536 0 -1 13056
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__1_.mem_right_track_44.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1679235063
transform 1 0 15272 0 1 14144
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__1_.mem_right_track_44.sky130_fd_sc_hd__dfrtp_1_1_
timestamp 1679235063
transform 1 0 15640 0 1 15232
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__1_.mem_right_track_46.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1679235063
transform 1 0 16836 0 -1 17408
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__1_.mem_right_track_46.sky130_fd_sc_hd__dfrtp_1_1_
timestamp 1679235063
transform 1 0 17848 0 -1 18496
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__1_.mem_right_track_48.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1679235063
transform 1 0 19688 0 1 17408
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__1_.mem_right_track_48.sky130_fd_sc_hd__dfrtp_1_1_
timestamp 1679235063
transform 1 0 21896 0 1 17408
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__1_.mem_right_track_50.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1679235063
transform 1 0 22264 0 1 18496
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__1_.mem_right_track_50.sky130_fd_sc_hd__dfrtp_1_1_
timestamp 1679235063
transform 1 0 21988 0 -1 19584
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__1_.mem_right_track_52.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1679235063
transform 1 0 21712 0 1 16320
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__1_.mem_right_track_52.sky130_fd_sc_hd__dfrtp_1_1_
timestamp 1679235063
transform 1 0 20976 0 1 14144
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__1_.mem_right_track_54.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1679235063
transform 1 0 19596 0 1 11968
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__1_.mem_right_track_54.sky130_fd_sc_hd__dfrtp_1_1_
timestamp 1679235063
transform 1 0 17940 0 -1 11968
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__1_.mem_right_track_56.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1679235063
transform 1 0 17848 0 -1 13056
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__1_.mem_right_track_56.sky130_fd_sc_hd__dfrtp_1_1_
timestamp 1679235063
transform 1 0 18768 0 -1 15232
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_4  sb_0__1_.mem_top_track_0.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1679235063
transform 1 0 3956 0 -1 50048
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__1_.mem_top_track_0.sky130_fd_sc_hd__dfrtp_1_1_
timestamp 1679235063
transform 1 0 9108 0 -1 45696
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__1_.mem_top_track_0.sky130_fd_sc_hd__dfrtp_1_2_
timestamp 1679235063
transform 1 0 10120 0 1 46784
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_2  sb_0__1_.mem_top_track_2.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1679235063
transform 1 0 11868 0 1 45696
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__1_.mem_top_track_2.sky130_fd_sc_hd__dfrtp_1_1_
timestamp 1679235063
transform 1 0 13064 0 -1 44608
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__1_.mem_top_track_2.sky130_fd_sc_hd__dfrtp_1_2_
timestamp 1679235063
transform 1 0 12328 0 -1 46784
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_2  sb_0__1_.mem_top_track_4.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1679235063
transform 1 0 12512 0 -1 43520
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__1_.mem_top_track_4.sky130_fd_sc_hd__dfrtp_1_1_
timestamp 1679235063
transform 1 0 10948 0 1 39168
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__1_.mem_top_track_4.sky130_fd_sc_hd__dfrtp_1_2_
timestamp 1679235063
transform 1 0 9016 0 -1 41344
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_4  sb_0__1_.mem_top_track_6.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1679235063
transform 1 0 8648 0 -1 40256
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__1_.mem_top_track_6.sky130_fd_sc_hd__dfrtp_1_1_
timestamp 1679235063
transform 1 0 6808 0 1 36992
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__1_.mem_top_track_6.sky130_fd_sc_hd__dfrtp_1_2_
timestamp 1679235063
transform 1 0 5428 0 1 38080
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_4  sb_0__1_.mem_top_track_10.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1679235063
transform 1 0 6532 0 -1 38080
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__1_.mem_top_track_10.sky130_fd_sc_hd__dfrtp_1_1_
timestamp 1679235063
transform 1 0 5244 0 1 35904
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__1_.mem_top_track_10.sky130_fd_sc_hd__dfrtp_1_2_
timestamp 1679235063
transform 1 0 4232 0 -1 35904
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_2  sb_0__1_.mem_top_track_12.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1679235063
transform 1 0 5520 0 1 33728
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__1_.mem_top_track_12.sky130_fd_sc_hd__dfrtp_1_1_
timestamp 1679235063
transform 1 0 6256 0 1 31552
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__1_.mem_top_track_12.sky130_fd_sc_hd__dfrtp_1_2_
timestamp 1679235063
transform 1 0 5336 0 1 32640
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_2  sb_0__1_.mem_top_track_20.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1679235063
transform 1 0 7636 0 -1 32640
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__1_.mem_top_track_20.sky130_fd_sc_hd__dfrtp_1_1_
timestamp 1679235063
transform 1 0 9476 0 1 31552
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__1_.mem_top_track_20.sky130_fd_sc_hd__dfrtp_1_2_
timestamp 1679235063
transform 1 0 7728 0 -1 34816
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__1_.mem_top_track_28.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1679235063
transform 1 0 8096 0 -1 35904
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__1_.mem_top_track_28.sky130_fd_sc_hd__dfrtp_1_1_
timestamp 1679235063
transform 1 0 6256 0 1 34816
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__1_.mem_top_track_28.sky130_fd_sc_hd__dfrtp_1_2_
timestamp 1679235063
transform 1 0 4048 0 1 36992
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__1_.mem_top_track_36.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1679235063
transform 1 0 5152 0 1 39168
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__1_.mem_top_track_36.sky130_fd_sc_hd__dfrtp_1_1_
timestamp 1679235063
transform 1 0 6440 0 1 40256
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__1_.mem_top_track_36.sky130_fd_sc_hd__dfrtp_1_2_
timestamp 1679235063
transform 1 0 5980 0 1 41344
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__1_.mem_top_track_44.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1679235063
transform 1 0 7544 0 -1 42432
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__1_.mem_top_track_44.sky130_fd_sc_hd__dfrtp_1_1_
timestamp 1679235063
transform 1 0 10856 0 1 42432
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__1_.mem_top_track_52.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1679235063
transform 1 0 14720 0 1 42432
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__1_.mem_top_track_52.sky130_fd_sc_hd__dfrtp_1_1_
timestamp 1679235063
transform 1 0 16928 0 -1 41344
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__1_.mem_top_track_52.sky130_fd_sc_hd__dfrtp_1_2_
timestamp 1679235063
transform 1 0 16836 0 -1 39168
box -38 -48 1878 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_bottom_track_1.mux_l1_in_0_
timestamp 1679235063
transform 1 0 17388 0 -1 28288
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_bottom_track_1.mux_l1_in_1_
timestamp 1679235063
transform 1 0 18584 0 -1 32640
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_bottom_track_1.mux_l1_in_2_
timestamp 1679235063
transform 1 0 13432 0 -1 22848
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_bottom_track_1.mux_l2_in_0_
timestamp 1679235063
transform 1 0 17848 0 -1 26112
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_bottom_track_1.mux_l2_in_1_
timestamp 1679235063
transform 1 0 17112 0 -1 21760
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  sb_0__1_.mux_bottom_track_1.mux_l2_in_1__252
timestamp 1679235063
transform 1 0 16100 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_bottom_track_1.mux_l3_in_0_
timestamp 1679235063
transform 1 0 17388 0 1 21760
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_2  sb_0__1_.mux_bottom_track_1.sky130_fd_sc_hd__buf_4_0_
timestamp 1679235063
transform 1 0 16100 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_bottom_track_3.mux_l1_in_0_
timestamp 1679235063
transform 1 0 19412 0 1 27200
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_bottom_track_3.mux_l1_in_1_
timestamp 1679235063
transform 1 0 19780 0 1 31552
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_bottom_track_3.mux_l2_in_0_
timestamp 1679235063
transform 1 0 19228 0 -1 26112
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  sb_0__1_.mux_bottom_track_3.mux_l2_in_1__203
timestamp 1679235063
transform 1 0 18584 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_bottom_track_3.mux_l2_in_1_
timestamp 1679235063
transform 1 0 17296 0 1 20672
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_bottom_track_3.mux_l3_in_0_
timestamp 1679235063
transform 1 0 18860 0 -1 20672
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  sb_0__1_.mux_bottom_track_3.sky130_fd_sc_hd__buf_4_0_
timestamp 1679235063
transform 1 0 16100 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_bottom_track_5.mux_l1_in_0_
timestamp 1679235063
transform 1 0 19780 0 -1 29376
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_bottom_track_5.mux_l1_in_1_
timestamp 1679235063
transform 1 0 21804 0 1 30464
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_bottom_track_5.mux_l1_in_2_
timestamp 1679235063
transform 1 0 19964 0 1 23936
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_bottom_track_5.mux_l2_in_0_
timestamp 1679235063
transform 1 0 22448 0 1 26112
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_bottom_track_5.mux_l2_in_1_
timestamp 1679235063
transform 1 0 24564 0 1 22848
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  sb_0__1_.mux_bottom_track_5.mux_l2_in_1__206
timestamp 1679235063
transform 1 0 21988 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_bottom_track_5.mux_l3_in_0_
timestamp 1679235063
transform 1 0 21988 0 -1 21760
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  sb_0__1_.mux_bottom_track_5.sky130_fd_sc_hd__buf_4_0_
timestamp 1679235063
transform 1 0 20976 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_bottom_track_7.mux_l1_in_0_
timestamp 1679235063
transform 1 0 16836 0 -1 29376
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_bottom_track_7.mux_l1_in_1_
timestamp 1679235063
transform 1 0 19780 0 -1 32640
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_bottom_track_7.mux_l1_in_2_
timestamp 1679235063
transform 1 0 16744 0 1 25024
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  sb_0__1_.mux_bottom_track_7.mux_l1_in_3__208
timestamp 1679235063
transform 1 0 14904 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_bottom_track_7.mux_l1_in_3_
timestamp 1679235063
transform 1 0 15364 0 -1 23936
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_bottom_track_7.mux_l2_in_0_
timestamp 1679235063
transform 1 0 17664 0 1 27200
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_bottom_track_7.mux_l2_in_1_
timestamp 1679235063
transform 1 0 15548 0 -1 25024
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_bottom_track_7.mux_l3_in_0_
timestamp 1679235063
transform 1 0 16836 0 -1 23936
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_2  sb_0__1_.mux_bottom_track_7.sky130_fd_sc_hd__buf_4_0_
timestamp 1679235063
transform 1 0 15732 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_bottom_track_11.mux_l1_in_0_
timestamp 1679235063
transform 1 0 17480 0 1 31552
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_bottom_track_11.mux_l1_in_1_
timestamp 1679235063
transform 1 0 18400 0 -1 34816
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_bottom_track_11.mux_l1_in_2_
timestamp 1679235063
transform 1 0 14904 0 1 26112
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_bottom_track_11.mux_l1_in_3_
timestamp 1679235063
transform 1 0 12144 0 1 25024
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  sb_0__1_.mux_bottom_track_11.mux_l1_in_3__253
timestamp 1679235063
transform 1 0 11500 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_bottom_track_11.mux_l2_in_0_
timestamp 1679235063
transform 1 0 15456 0 -1 29376
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_bottom_track_11.mux_l2_in_1_
timestamp 1679235063
transform 1 0 12972 0 1 26112
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_bottom_track_11.mux_l3_in_0_
timestamp 1679235063
transform 1 0 14536 0 1 25024
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  sb_0__1_.mux_bottom_track_11.sky130_fd_sc_hd__buf_4_0_
timestamp 1679235063
transform 1 0 15364 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_bottom_track_13.mux_l1_in_0_
timestamp 1679235063
transform 1 0 17388 0 -1 30464
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_bottom_track_13.mux_l1_in_1_
timestamp 1679235063
transform 1 0 20608 0 -1 34816
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_bottom_track_13.mux_l1_in_2_
timestamp 1679235063
transform 1 0 18032 0 -1 27200
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_bottom_track_13.mux_l2_in_0_
timestamp 1679235063
transform 1 0 19504 0 1 29376
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  sb_0__1_.mux_bottom_track_13.mux_l2_in_1__254
timestamp 1679235063
transform 1 0 19872 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_bottom_track_13.mux_l2_in_1_
timestamp 1679235063
transform 1 0 19412 0 1 26112
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_bottom_track_13.mux_l3_in_0_
timestamp 1679235063
transform 1 0 19596 0 -1 25024
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  sb_0__1_.mux_bottom_track_13.sky130_fd_sc_hd__buf_4_0_
timestamp 1679235063
transform 1 0 18124 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_bottom_track_21.mux_l1_in_0_
timestamp 1679235063
transform 1 0 19412 0 1 30464
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_bottom_track_21.mux_l1_in_1_
timestamp 1679235063
transform 1 0 21988 0 -1 34816
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_bottom_track_21.mux_l1_in_2_
timestamp 1679235063
transform 1 0 20608 0 1 27200
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_bottom_track_21.mux_l2_in_0_
timestamp 1679235063
transform 1 0 21988 0 -1 29376
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  sb_0__1_.mux_bottom_track_21.mux_l2_in_1__255
timestamp 1679235063
transform 1 0 23276 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_bottom_track_21.mux_l2_in_1_
timestamp 1679235063
transform 1 0 22080 0 -1 26112
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_bottom_track_21.mux_l3_in_0_
timestamp 1679235063
transform 1 0 21436 0 1 23936
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  sb_0__1_.mux_bottom_track_21.sky130_fd_sc_hd__buf_4_0_
timestamp 1679235063
transform 1 0 21896 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_bottom_track_29.mux_l1_in_0_
timestamp 1679235063
transform 1 0 16560 0 1 32640
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_bottom_track_29.mux_l1_in_1_
timestamp 1679235063
transform 1 0 20148 0 1 36992
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_bottom_track_29.mux_l1_in_2_
timestamp 1679235063
transform 1 0 18032 0 -1 29376
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_bottom_track_29.mux_l2_in_0_
timestamp 1679235063
transform 1 0 17388 0 -1 32640
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  sb_0__1_.mux_bottom_track_29.mux_l2_in_1__256
timestamp 1679235063
transform 1 0 18216 0 1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_bottom_track_29.mux_l2_in_1_
timestamp 1679235063
transform 1 0 17020 0 1 29376
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_bottom_track_29.mux_l3_in_0_
timestamp 1679235063
transform 1 0 16192 0 1 28288
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  sb_0__1_.mux_bottom_track_29.sky130_fd_sc_hd__buf_4_0_
timestamp 1679235063
transform 1 0 16468 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_bottom_track_37.mux_l1_in_0_
timestamp 1679235063
transform 1 0 17940 0 -1 38080
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_bottom_track_37.mux_l1_in_1_
timestamp 1679235063
transform 1 0 19872 0 -1 35904
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_bottom_track_37.mux_l2_in_0_
timestamp 1679235063
transform 1 0 15548 0 -1 34816
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_bottom_track_37.mux_l2_in_1_
timestamp 1679235063
transform 1 0 11408 0 1 28288
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  sb_0__1_.mux_bottom_track_37.mux_l2_in_1__204
timestamp 1679235063
transform 1 0 12328 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_bottom_track_37.mux_l3_in_0_
timestamp 1679235063
transform 1 0 13432 0 -1 29376
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  sb_0__1_.mux_bottom_track_37.sky130_fd_sc_hd__buf_4_0_
timestamp 1679235063
transform 1 0 12788 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_bottom_track_45.mux_l1_in_0_
timestamp 1679235063
transform 1 0 20608 0 -1 39168
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_bottom_track_45.mux_l2_in_0_
timestamp 1679235063
transform 1 0 20884 0 1 35904
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  sb_0__1_.mux_bottom_track_45.mux_l2_in_1__205
timestamp 1679235063
transform 1 0 21620 0 1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_bottom_track_45.mux_l2_in_1_
timestamp 1679235063
transform 1 0 21988 0 -1 33728
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_bottom_track_45.mux_l3_in_0_
timestamp 1679235063
transform 1 0 19504 0 -1 31552
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  sb_0__1_.mux_bottom_track_45.sky130_fd_sc_hd__buf_4_0_
timestamp 1679235063
transform 1 0 18400 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_bottom_track_53.mux_l1_in_0_
timestamp 1679235063
transform 1 0 14904 0 -1 39168
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  sb_0__1_.mux_bottom_track_53.mux_l1_in_1__207
timestamp 1679235063
transform 1 0 15364 0 1 38080
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_bottom_track_53.mux_l1_in_1_
timestamp 1679235063
transform 1 0 14996 0 -1 38080
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_bottom_track_53.mux_l2_in_0_
timestamp 1679235063
transform 1 0 11316 0 1 36992
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_2  sb_0__1_.mux_bottom_track_53.sky130_fd_sc_hd__buf_4_0_
timestamp 1679235063
transform 1 0 10580 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_right_track_0.mux_l1_in_0_
timestamp 1679235063
transform 1 0 20792 0 1 32640
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_right_track_0.mux_l1_in_1_
timestamp 1679235063
transform 1 0 21988 0 1 32640
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_right_track_0.mux_l2_in_0_
timestamp 1679235063
transform 1 0 21988 0 1 31552
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  sb_0__1_.mux_right_track_0.mux_l2_in_1__209
timestamp 1679235063
transform 1 0 21252 0 -1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_right_track_0.mux_l2_in_1_
timestamp 1679235063
transform 1 0 21068 0 1 28288
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_right_track_0.mux_l3_in_0_
timestamp 1679235063
transform 1 0 22816 0 1 29376
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  sb_0__1_.mux_right_track_0.sky130_fd_sc_hd__buf_4_0_
timestamp 1679235063
transform 1 0 24564 0 1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_right_track_2.mux_l1_in_0_
timestamp 1679235063
transform 1 0 22264 0 1 45696
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_right_track_2.mux_l1_in_1_
timestamp 1679235063
transform 1 0 21344 0 1 39168
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_right_track_2.mux_l1_in_2_
timestamp 1679235063
transform 1 0 19964 0 -1 36992
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_right_track_2.mux_l2_in_0_
timestamp 1679235063
transform 1 0 22632 0 1 41344
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  sb_0__1_.mux_right_track_2.mux_l2_in_1__215
timestamp 1679235063
transform 1 0 23736 0 1 39168
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_right_track_2.mux_l2_in_1_
timestamp 1679235063
transform 1 0 22540 0 1 39168
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_right_track_2.mux_l3_in_0_
timestamp 1679235063
transform 1 0 24564 0 1 39168
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  sb_0__1_.mux_right_track_2.sky130_fd_sc_hd__buf_4_0_
timestamp 1679235063
transform 1 0 24564 0 1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_right_track_4.mux_l1_in_0_
timestamp 1679235063
transform 1 0 22080 0 1 43520
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_right_track_4.mux_l1_in_1_
timestamp 1679235063
transform 1 0 21988 0 -1 38080
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_right_track_4.mux_l2_in_0_
timestamp 1679235063
transform 1 0 22724 0 1 38080
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  sb_0__1_.mux_right_track_4.mux_l2_in_1__226
timestamp 1679235063
transform 1 0 19964 0 -1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_right_track_4.mux_l2_in_1_
timestamp 1679235063
transform 1 0 20516 0 -1 33728
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_right_track_4.mux_l3_in_0_
timestamp 1679235063
transform 1 0 22356 0 1 33728
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  sb_0__1_.mux_right_track_4.sky130_fd_sc_hd__buf_4_0_
timestamp 1679235063
transform 1 0 23736 0 1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_right_track_6.mux_l1_in_0_
timestamp 1679235063
transform 1 0 21988 0 -1 43520
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_right_track_6.mux_l1_in_1_
timestamp 1679235063
transform 1 0 21528 0 1 36992
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_right_track_6.mux_l1_in_2_
timestamp 1679235063
transform 1 0 19504 0 1 32640
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_right_track_6.mux_l2_in_0_
timestamp 1679235063
transform 1 0 24564 0 1 38080
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  sb_0__1_.mux_right_track_6.mux_l2_in_1__235
timestamp 1679235063
transform 1 0 22632 0 1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_right_track_6.mux_l2_in_1_
timestamp 1679235063
transform 1 0 21988 0 -1 35904
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_right_track_6.mux_l3_in_0_
timestamp 1679235063
transform 1 0 23276 0 1 35904
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  sb_0__1_.mux_right_track_6.sky130_fd_sc_hd__buf_4_0_
timestamp 1679235063
transform 1 0 24288 0 -1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_right_track_8.mux_l1_in_0_
timestamp 1679235063
transform 1 0 21988 0 -1 46784
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_right_track_8.mux_l1_in_1_
timestamp 1679235063
transform 1 0 20884 0 1 40256
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_right_track_8.mux_l1_in_2_
timestamp 1679235063
transform 1 0 19136 0 -1 38080
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_right_track_8.mux_l2_in_0_
timestamp 1679235063
transform 1 0 21804 0 1 42432
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_right_track_8.mux_l2_in_1_
timestamp 1679235063
transform 1 0 21344 0 1 41344
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  sb_0__1_.mux_right_track_8.mux_l2_in_1__236
timestamp 1679235063
transform 1 0 21988 0 -1 41344
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_right_track_8.mux_l3_in_0_
timestamp 1679235063
transform 1 0 22448 0 1 40256
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  sb_0__1_.mux_right_track_8.sky130_fd_sc_hd__buf_4_0_
timestamp 1679235063
transform 1 0 23736 0 -1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_right_track_10.mux_l1_in_0_
timestamp 1679235063
transform 1 0 20424 0 -1 45696
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_right_track_10.mux_l1_in_1_
timestamp 1679235063
transform 1 0 20608 0 -1 40256
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_right_track_10.mux_l2_in_0_
timestamp 1679235063
transform 1 0 19596 0 1 41344
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  sb_0__1_.mux_right_track_10.mux_l2_in_1__210
timestamp 1679235063
transform 1 0 17388 0 1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_right_track_10.mux_l2_in_1_
timestamp 1679235063
transform 1 0 16192 0 1 35904
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_right_track_10.mux_l3_in_0_
timestamp 1679235063
transform 1 0 20608 0 -1 38080
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  sb_0__1_.mux_right_track_10.sky130_fd_sc_hd__buf_4_0_
timestamp 1679235063
transform 1 0 23276 0 -1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_right_track_12.mux_l1_in_0_
timestamp 1679235063
transform 1 0 19688 0 -1 46784
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_right_track_12.mux_l2_in_0_
timestamp 1679235063
transform 1 0 19320 0 -1 41344
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  sb_0__1_.mux_right_track_12.mux_l2_in_1__211
timestamp 1679235063
transform 1 0 18492 0 1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_right_track_12.mux_l2_in_1_
timestamp 1679235063
transform 1 0 17020 0 -1 36992
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_right_track_12.mux_l3_in_0_
timestamp 1679235063
transform 1 0 19412 0 -1 40256
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  sb_0__1_.mux_right_track_12.sky130_fd_sc_hd__buf_4_0_
timestamp 1679235063
transform 1 0 22632 0 -1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_right_track_14.mux_l1_in_0_
timestamp 1679235063
transform 1 0 18124 0 1 46784
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_right_track_14.mux_l2_in_0_
timestamp 1679235063
transform 1 0 18124 0 1 41344
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_right_track_14.mux_l2_in_1_
timestamp 1679235063
transform 1 0 16192 0 1 38080
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  sb_0__1_.mux_right_track_14.mux_l2_in_1__212
timestamp 1679235063
transform 1 0 16836 0 -1 38080
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_right_track_14.mux_l3_in_0_
timestamp 1679235063
transform 1 0 18216 0 -1 40256
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  sb_0__1_.mux_right_track_14.sky130_fd_sc_hd__buf_4_0_
timestamp 1679235063
transform 1 0 21988 0 -1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_right_track_16.mux_l1_in_0_
timestamp 1679235063
transform 1 0 18032 0 -1 47872
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_right_track_16.mux_l2_in_0_
timestamp 1679235063
transform 1 0 17020 0 1 43520
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_right_track_16.mux_l2_in_1_
timestamp 1679235063
transform 1 0 14444 0 1 39168
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  sb_0__1_.mux_right_track_16.mux_l2_in_1__213
timestamp 1679235063
transform 1 0 14260 0 1 38080
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_right_track_16.mux_l3_in_0_
timestamp 1679235063
transform 1 0 16744 0 1 40256
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  sb_0__1_.mux_right_track_16.sky130_fd_sc_hd__buf_4_0_
timestamp 1679235063
transform 1 0 20976 0 -1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_right_track_18.mux_l1_in_0_
timestamp 1679235063
transform 1 0 16836 0 -1 47872
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_right_track_18.mux_l2_in_0_
timestamp 1679235063
transform 1 0 16376 0 1 41344
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  sb_0__1_.mux_right_track_18.mux_l2_in_1__214
timestamp 1679235063
transform 1 0 14260 0 1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_right_track_18.mux_l2_in_1_
timestamp 1679235063
transform 1 0 12972 0 -1 36992
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_right_track_18.mux_l3_in_0_
timestamp 1679235063
transform 1 0 16100 0 1 36992
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  sb_0__1_.mux_right_track_18.sky130_fd_sc_hd__buf_4_0_
timestamp 1679235063
transform 1 0 19596 0 -1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_right_track_20.mux_l1_in_0_
timestamp 1679235063
transform 1 0 14812 0 -1 43520
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_right_track_20.mux_l2_in_0_
timestamp 1679235063
transform 1 0 14444 0 -1 36992
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  sb_0__1_.mux_right_track_20.mux_l2_in_1__216
timestamp 1679235063
transform 1 0 12512 0 -1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_right_track_20.mux_l2_in_1_
timestamp 1679235063
transform 1 0 12052 0 1 31552
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_right_track_20.mux_l3_in_0_
timestamp 1679235063
transform 1 0 14260 0 1 32640
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  sb_0__1_.mux_right_track_20.sky130_fd_sc_hd__buf_4_0_
timestamp 1679235063
transform 1 0 19228 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_right_track_22.mux_l1_in_0_
timestamp 1679235063
transform 1 0 12604 0 1 40256
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_right_track_22.mux_l2_in_0_
timestamp 1679235063
transform 1 0 13064 0 -1 34816
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  sb_0__1_.mux_right_track_22.mux_l2_in_1__217
timestamp 1679235063
transform 1 0 11684 0 -1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_right_track_22.mux_l2_in_1_
timestamp 1679235063
transform 1 0 10396 0 -1 30464
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_right_track_22.mux_l3_in_0_
timestamp 1679235063
transform 1 0 12512 0 -1 30464
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  sb_0__1_.mux_right_track_22.sky130_fd_sc_hd__buf_4_0_
timestamp 1679235063
transform 1 0 18032 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_right_track_24.mux_l1_in_0_
timestamp 1679235063
transform 1 0 14260 0 1 28288
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_right_track_24.mux_l1_in_1_
timestamp 1679235063
transform 1 0 10764 0 1 26112
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  sb_0__1_.mux_right_track_24.mux_l1_in_1__218
timestamp 1679235063
transform 1 0 11684 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_right_track_24.mux_l2_in_0_
timestamp 1679235063
transform 1 0 12604 0 -1 26112
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  sb_0__1_.mux_right_track_24.sky130_fd_sc_hd__buf_4_0_
timestamp 1679235063
transform 1 0 18492 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_right_track_26.mux_l1_in_0_
timestamp 1679235063
transform 1 0 14260 0 1 30464
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  sb_0__1_.mux_right_track_26.mux_l1_in_1__219
timestamp 1679235063
transform 1 0 9568 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_right_track_26.mux_l1_in_1_
timestamp 1679235063
transform 1 0 9108 0 -1 27200
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_right_track_26.mux_l2_in_0_
timestamp 1679235063
transform 1 0 11408 0 1 27200
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  sb_0__1_.mux_right_track_26.sky130_fd_sc_hd__buf_4_0_
timestamp 1679235063
transform 1 0 16100 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_right_track_28.mux_l1_in_0_
timestamp 1679235063
transform 1 0 11960 0 -1 29376
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  sb_0__1_.mux_right_track_28.mux_l1_in_1__220
timestamp 1679235063
transform 1 0 6808 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_right_track_28.mux_l1_in_1_
timestamp 1679235063
transform 1 0 7452 0 1 25024
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_right_track_28.mux_l2_in_0_
timestamp 1679235063
transform 1 0 10120 0 -1 26112
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  sb_0__1_.mux_right_track_28.sky130_fd_sc_hd__buf_4_0_
timestamp 1679235063
transform 1 0 16836 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_right_track_30.mux_l1_in_0_
timestamp 1679235063
transform 1 0 12604 0 1 28288
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_right_track_30.mux_l1_in_1_
timestamp 1679235063
transform 1 0 8280 0 -1 25024
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  sb_0__1_.mux_right_track_30.mux_l1_in_1__221
timestamp 1679235063
transform 1 0 9108 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_right_track_30.mux_l2_in_0_
timestamp 1679235063
transform 1 0 12972 0 -1 25024
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  sb_0__1_.mux_right_track_30.sky130_fd_sc_hd__buf_4_0_
timestamp 1679235063
transform 1 0 16836 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_right_track_32.mux_l1_in_0_
timestamp 1679235063
transform 1 0 12972 0 1 27200
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_right_track_32.mux_l1_in_1_
timestamp 1679235063
transform 1 0 10396 0 -1 23936
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  sb_0__1_.mux_right_track_32.mux_l1_in_1__222
timestamp 1679235063
transform 1 0 11684 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_right_track_32.mux_l2_in_0_
timestamp 1679235063
transform 1 0 14260 0 1 22848
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  sb_0__1_.mux_right_track_32.sky130_fd_sc_hd__buf_4_0_
timestamp 1679235063
transform 1 0 17480 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_right_track_34.mux_l1_in_0_
timestamp 1679235063
transform 1 0 16836 0 -1 27200
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_right_track_34.mux_l1_in_1_
timestamp 1679235063
transform 1 0 12420 0 1 21760
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  sb_0__1_.mux_right_track_34.mux_l1_in_1__223
timestamp 1679235063
transform 1 0 12880 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_right_track_34.mux_l2_in_0_
timestamp 1679235063
transform 1 0 15916 0 1 21760
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  sb_0__1_.mux_right_track_34.sky130_fd_sc_hd__buf_4_0_
timestamp 1679235063
transform 1 0 20608 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_right_track_36.mux_l1_in_0_
timestamp 1679235063
transform 1 0 13340 0 -1 23936
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_right_track_36.mux_l2_in_0_
timestamp 1679235063
transform 1 0 8648 0 -1 17408
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  sb_0__1_.mux_right_track_36.mux_l2_in_1__224
timestamp 1679235063
transform 1 0 7544 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_right_track_36.mux_l2_in_1_
timestamp 1679235063
transform 1 0 7084 0 1 8704
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_right_track_36.mux_l3_in_0_
timestamp 1679235063
transform 1 0 10304 0 1 13056
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  sb_0__1_.mux_right_track_36.sky130_fd_sc_hd__buf_4_0_
timestamp 1679235063
transform 1 0 16652 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_right_track_38.mux_l1_in_0_
timestamp 1679235063
transform 1 0 12420 0 -1 14144
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  sb_0__1_.mux_right_track_38.mux_l2_in_0__225
timestamp 1679235063
transform 1 0 17572 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_right_track_38.mux_l2_in_0_
timestamp 1679235063
transform 1 0 15180 0 -1 11968
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  sb_0__1_.mux_right_track_38.sky130_fd_sc_hd__buf_4_0_
timestamp 1679235063
transform 1 0 18308 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_right_track_40.mux_l1_in_0_
timestamp 1679235063
transform 1 0 14168 0 -1 15232
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_right_track_40.mux_l2_in_0_
timestamp 1679235063
transform 1 0 16468 0 1 13056
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  sb_0__1_.mux_right_track_40.mux_l2_in_0__227
timestamp 1679235063
transform 1 0 16928 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  sb_0__1_.mux_right_track_40.sky130_fd_sc_hd__buf_4_0_
timestamp 1679235063
transform 1 0 20148 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_right_track_44.mux_l1_in_0_
timestamp 1679235063
transform 1 0 15548 0 -1 17408
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_right_track_44.mux_l2_in_0_
timestamp 1679235063
transform 1 0 17572 0 -1 15232
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  sb_0__1_.mux_right_track_44.mux_l2_in_0__228
timestamp 1679235063
transform 1 0 19412 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  sb_0__1_.mux_right_track_44.sky130_fd_sc_hd__buf_4_0_
timestamp 1679235063
transform 1 0 21804 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_right_track_46.mux_l1_in_0_
timestamp 1679235063
transform 1 0 16836 0 1 18496
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_right_track_46.mux_l2_in_0_
timestamp 1679235063
transform 1 0 20332 0 -1 16320
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  sb_0__1_.mux_right_track_46.mux_l2_in_0__229
timestamp 1679235063
transform 1 0 21252 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  sb_0__1_.mux_right_track_46.sky130_fd_sc_hd__buf_4_0_
timestamp 1679235063
transform 1 0 22632 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_right_track_48.mux_l1_in_0_
timestamp 1679235063
transform 1 0 19044 0 -1 17408
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  sb_0__1_.mux_right_track_48.mux_l2_in_0__230
timestamp 1679235063
transform 1 0 23184 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_right_track_48.mux_l2_in_0_
timestamp 1679235063
transform 1 0 21988 0 -1 16320
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  sb_0__1_.mux_right_track_48.sky130_fd_sc_hd__buf_4_0_
timestamp 1679235063
transform 1 0 23276 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_right_track_50.mux_l1_in_0_
timestamp 1679235063
transform 1 0 21252 0 1 26112
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  sb_0__1_.mux_right_track_50.mux_l1_in_1__231
timestamp 1679235063
transform 1 0 19596 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_right_track_50.mux_l1_in_1_
timestamp 1679235063
transform 1 0 19136 0 -1 16320
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_right_track_50.mux_l2_in_0_
timestamp 1679235063
transform 1 0 21068 0 1 18496
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  sb_0__1_.mux_right_track_50.sky130_fd_sc_hd__buf_4_0_
timestamp 1679235063
transform 1 0 23000 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_right_track_52.mux_l1_in_0_
timestamp 1679235063
transform 1 0 19412 0 1 15232
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  sb_0__1_.mux_right_track_52.mux_l2_in_0__232
timestamp 1679235063
transform 1 0 22724 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_right_track_52.mux_l2_in_0_
timestamp 1679235063
transform 1 0 20700 0 -1 13056
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  sb_0__1_.mux_right_track_52.sky130_fd_sc_hd__buf_4_0_
timestamp 1679235063
transform 1 0 22724 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_right_track_54.mux_l1_in_0_
timestamp 1679235063
transform 1 0 17664 0 1 13056
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  sb_0__1_.mux_right_track_54.mux_l2_in_0__233
timestamp 1679235063
transform 1 0 19504 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_right_track_54.mux_l2_in_0_
timestamp 1679235063
transform 1 0 19136 0 -1 10880
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  sb_0__1_.mux_right_track_54.sky130_fd_sc_hd__buf_4_0_
timestamp 1679235063
transform 1 0 21436 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_right_track_56.mux_l1_in_0_
timestamp 1679235063
transform 1 0 17940 0 1 15232
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  sb_0__1_.mux_right_track_56.mux_l2_in_0__234
timestamp 1679235063
transform 1 0 21252 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_right_track_56.mux_l2_in_0_
timestamp 1679235063
transform 1 0 20056 0 -1 14144
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  sb_0__1_.mux_right_track_56.sky130_fd_sc_hd__buf_4_0_
timestamp 1679235063
transform 1 0 21988 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_top_track_0.mux_l1_in_0_
timestamp 1679235063
transform 1 0 9108 0 -1 43520
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_top_track_0.mux_l1_in_1_
timestamp 1679235063
transform 1 0 17112 0 -1 42432
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_top_track_0.mux_l1_in_2_
timestamp 1679235063
transform 1 0 14904 0 1 36992
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_top_track_0.mux_l1_in_3_
timestamp 1679235063
transform 1 0 9936 0 1 36992
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  sb_0__1_.mux_top_track_0.mux_l1_in_3__237
timestamp 1679235063
transform 1 0 9108 0 1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_top_track_0.mux_l2_in_0_
timestamp 1679235063
transform 1 0 11868 0 -1 44608
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_top_track_0.mux_l2_in_1_
timestamp 1679235063
transform 1 0 11500 0 1 41344
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_top_track_0.mux_l3_in_0_
timestamp 1679235063
transform 1 0 10672 0 1 45696
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  sb_0__1_.mux_top_track_0.sky130_fd_sc_hd__buf_4_0_
timestamp 1679235063
transform 1 0 11592 0 1 48960
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_top_track_2.mux_l1_in_0_
timestamp 1679235063
transform 1 0 16928 0 -1 43520
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_top_track_2.mux_l1_in_1_
timestamp 1679235063
transform 1 0 19412 0 -1 39168
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_top_track_2.mux_l1_in_2_
timestamp 1679235063
transform 1 0 12880 0 1 35904
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_top_track_2.mux_l2_in_0_
timestamp 1679235063
transform 1 0 15272 0 -1 42432
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  sb_0__1_.mux_top_track_2.mux_l2_in_1__240
timestamp 1679235063
transform 1 0 14076 0 -1 42432
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_top_track_2.mux_l2_in_1_
timestamp 1679235063
transform 1 0 12880 0 -1 42432
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_top_track_2.mux_l3_in_0_
timestamp 1679235063
transform 1 0 13156 0 -1 45696
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  sb_0__1_.mux_top_track_2.sky130_fd_sc_hd__buf_4_0_
timestamp 1679235063
transform 1 0 12696 0 1 48960
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_top_track_4.mux_l1_in_0_
timestamp 1679235063
transform 1 0 15180 0 1 41344
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_top_track_4.mux_l1_in_1_
timestamp 1679235063
transform 1 0 19412 0 1 35904
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_top_track_4.mux_l1_in_2_
timestamp 1679235063
transform 1 0 10856 0 1 32640
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_top_track_4.mux_l2_in_0_
timestamp 1679235063
transform 1 0 14260 0 1 40256
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_top_track_4.mux_l2_in_1_
timestamp 1679235063
transform 1 0 10396 0 -1 39168
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  sb_0__1_.mux_top_track_4.mux_l2_in_1__244
timestamp 1679235063
transform 1 0 11684 0 -1 38080
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_top_track_4.mux_l3_in_0_
timestamp 1679235063
transform 1 0 10304 0 1 41344
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  sb_0__1_.mux_top_track_4.sky130_fd_sc_hd__buf_4_0_
timestamp 1679235063
transform 1 0 11684 0 -1 46784
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_top_track_6.mux_l1_in_0_
timestamp 1679235063
transform 1 0 9108 0 1 41344
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_top_track_6.mux_l1_in_1_
timestamp 1679235063
transform 1 0 17388 0 1 38080
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_top_track_6.mux_l1_in_2_
timestamp 1679235063
transform 1 0 13708 0 -1 32640
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  sb_0__1_.mux_top_track_6.mux_l1_in_3__247
timestamp 1679235063
transform 1 0 11684 0 -1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_top_track_6.mux_l1_in_3_
timestamp 1679235063
transform 1 0 7728 0 1 30464
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_top_track_6.mux_l2_in_0_
timestamp 1679235063
transform 1 0 9752 0 1 39168
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_top_track_6.mux_l2_in_1_
timestamp 1679235063
transform 1 0 9108 0 1 34816
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_top_track_6.mux_l3_in_0_
timestamp 1679235063
transform 1 0 7452 0 -1 40256
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  sb_0__1_.mux_top_track_6.sky130_fd_sc_hd__buf_4_0_
timestamp 1679235063
transform 1 0 9108 0 1 45696
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_top_track_10.mux_l1_in_0_
timestamp 1679235063
transform 1 0 11684 0 -1 40256
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_top_track_10.mux_l1_in_1_
timestamp 1679235063
transform 1 0 17296 0 1 36992
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_top_track_10.mux_l1_in_2_
timestamp 1679235063
transform 1 0 12512 0 1 30464
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  sb_0__1_.mux_top_track_10.mux_l1_in_3__238
timestamp 1679235063
transform 1 0 8464 0 -1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_top_track_10.mux_l1_in_3_
timestamp 1679235063
transform 1 0 7268 0 -1 31552
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_top_track_10.mux_l2_in_0_
timestamp 1679235063
transform 1 0 9200 0 1 38080
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_top_track_10.mux_l2_in_1_
timestamp 1679235063
transform 1 0 7820 0 1 33728
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_top_track_10.mux_l3_in_0_
timestamp 1679235063
transform 1 0 7636 0 1 38080
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  sb_0__1_.mux_top_track_10.sky130_fd_sc_hd__buf_4_0_
timestamp 1679235063
transform 1 0 8372 0 1 44608
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_top_track_12.mux_l1_in_0_
timestamp 1679235063
transform 1 0 12512 0 1 36992
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_top_track_12.mux_l1_in_1_
timestamp 1679235063
transform 1 0 16836 0 -1 31552
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_top_track_12.mux_l1_in_2_
timestamp 1679235063
transform 1 0 7820 0 1 28288
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_top_track_12.mux_l2_in_0_
timestamp 1679235063
transform 1 0 10212 0 1 33728
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_top_track_12.mux_l2_in_1_
timestamp 1679235063
transform 1 0 7544 0 1 32640
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  sb_0__1_.mux_top_track_12.mux_l2_in_1__239
timestamp 1679235063
transform 1 0 6992 0 -1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_top_track_12.mux_l3_in_0_
timestamp 1679235063
transform 1 0 7728 0 1 35904
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  sb_0__1_.mux_top_track_12.sky130_fd_sc_hd__buf_4_0_
timestamp 1679235063
transform 1 0 7728 0 -1 43520
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_top_track_20.mux_l1_in_0_
timestamp 1679235063
transform 1 0 14444 0 -1 35904
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_top_track_20.mux_l1_in_1_
timestamp 1679235063
transform 1 0 18124 0 -1 31552
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_top_track_20.mux_l1_in_2_
timestamp 1679235063
transform 1 0 9752 0 -1 29376
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_top_track_20.mux_l2_in_0_
timestamp 1679235063
transform 1 0 12788 0 1 34816
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  sb_0__1_.mux_top_track_20.mux_l2_in_1__241
timestamp 1679235063
transform 1 0 9752 0 -1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_top_track_20.mux_l2_in_1_
timestamp 1679235063
transform 1 0 9384 0 1 32640
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_top_track_20.mux_l3_in_0_
timestamp 1679235063
transform 1 0 9384 0 -1 38080
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  sb_0__1_.mux_top_track_20.sky130_fd_sc_hd__buf_4_0_
timestamp 1679235063
transform 1 0 8372 0 1 43520
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_top_track_28.mux_l1_in_0_
timestamp 1679235063
transform 1 0 12512 0 -1 38080
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_top_track_28.mux_l1_in_1_
timestamp 1679235063
transform 1 0 12788 0 -1 33728
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_top_track_28.mux_l2_in_0_
timestamp 1679235063
transform 1 0 9108 0 1 35904
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  sb_0__1_.mux_top_track_28.mux_l2_in_1__242
timestamp 1679235063
transform 1 0 5612 0 -1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_top_track_28.mux_l2_in_1_
timestamp 1679235063
transform 1 0 5152 0 -1 32640
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_top_track_28.mux_l3_in_0_
timestamp 1679235063
transform 1 0 6532 0 -1 39168
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  sb_0__1_.mux_top_track_28.sky130_fd_sc_hd__buf_4_0_
timestamp 1679235063
transform 1 0 5796 0 -1 44608
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_top_track_36.mux_l1_in_0_
timestamp 1679235063
transform 1 0 11408 0 1 40256
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_top_track_36.mux_l2_in_0_
timestamp 1679235063
transform 1 0 12236 0 -1 39168
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  sb_0__1_.mux_top_track_36.mux_l2_in_1__243
timestamp 1679235063
transform 1 0 6808 0 -1 40256
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_top_track_36.mux_l2_in_1_
timestamp 1679235063
transform 1 0 9108 0 -1 39168
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_top_track_36.mux_l3_in_0_
timestamp 1679235063
transform 1 0 9752 0 -1 42432
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  sb_0__1_.mux_top_track_36.sky130_fd_sc_hd__buf_4_0_
timestamp 1679235063
transform 1 0 7268 0 -1 46784
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_top_track_44.mux_l1_in_0_
timestamp 1679235063
transform 1 0 15548 0 -1 40256
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  sb_0__1_.mux_top_track_44.mux_l1_in_1__245
timestamp 1679235063
transform 1 0 9108 0 1 39168
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_top_track_44.mux_l1_in_1_
timestamp 1679235063
transform 1 0 10396 0 1 38080
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_top_track_44.mux_l2_in_0_
timestamp 1679235063
transform 1 0 11684 0 -1 42432
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  sb_0__1_.mux_top_track_44.sky130_fd_sc_hd__buf_4_0_
timestamp 1679235063
transform 1 0 9200 0 -1 47872
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_top_track_52.mux_l1_in_0_
timestamp 1679235063
transform 1 0 20700 0 -1 41344
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_top_track_52.mux_l2_in_0_
timestamp 1679235063
transform 1 0 19412 0 1 39168
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  sb_0__1_.mux_top_track_52.mux_l2_in_1__246
timestamp 1679235063
transform 1 0 15456 0 1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_top_track_52.mux_l2_in_1_
timestamp 1679235063
transform 1 0 14260 0 1 35904
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_top_track_52.mux_l3_in_0_
timestamp 1679235063
transform 1 0 15640 0 1 39168
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  sb_0__1_.mux_top_track_52.sky130_fd_sc_hd__buf_4_0_
timestamp 1679235063
transform 1 0 10028 0 1 45696
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_192 pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1679235063
transform 1 0 3680 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_193
timestamp 1679235063
transform 1 0 6256 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_194
timestamp 1679235063
transform 1 0 8832 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_195
timestamp 1679235063
transform 1 0 11408 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_196
timestamp 1679235063
transform 1 0 13984 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_197
timestamp 1679235063
transform 1 0 16560 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_198
timestamp 1679235063
transform 1 0 19136 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_199
timestamp 1679235063
transform 1 0 21712 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_200
timestamp 1679235063
transform 1 0 24288 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_201
timestamp 1679235063
transform 1 0 6256 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_202
timestamp 1679235063
transform 1 0 11408 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_203
timestamp 1679235063
transform 1 0 16560 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_204
timestamp 1679235063
transform 1 0 21712 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_205
timestamp 1679235063
transform 1 0 3680 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_206
timestamp 1679235063
transform 1 0 8832 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_207
timestamp 1679235063
transform 1 0 13984 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_208
timestamp 1679235063
transform 1 0 19136 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_209
timestamp 1679235063
transform 1 0 24288 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_210
timestamp 1679235063
transform 1 0 6256 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_211
timestamp 1679235063
transform 1 0 11408 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_212
timestamp 1679235063
transform 1 0 16560 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_213
timestamp 1679235063
transform 1 0 21712 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_214
timestamp 1679235063
transform 1 0 3680 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_215
timestamp 1679235063
transform 1 0 8832 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_216
timestamp 1679235063
transform 1 0 13984 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_217
timestamp 1679235063
transform 1 0 19136 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_218
timestamp 1679235063
transform 1 0 24288 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_219
timestamp 1679235063
transform 1 0 6256 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_220
timestamp 1679235063
transform 1 0 11408 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_221
timestamp 1679235063
transform 1 0 16560 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_222
timestamp 1679235063
transform 1 0 21712 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_223
timestamp 1679235063
transform 1 0 3680 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_224
timestamp 1679235063
transform 1 0 8832 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_225
timestamp 1679235063
transform 1 0 13984 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_226
timestamp 1679235063
transform 1 0 19136 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_227
timestamp 1679235063
transform 1 0 24288 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_228
timestamp 1679235063
transform 1 0 6256 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_229
timestamp 1679235063
transform 1 0 11408 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_230
timestamp 1679235063
transform 1 0 16560 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_231
timestamp 1679235063
transform 1 0 21712 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_232
timestamp 1679235063
transform 1 0 3680 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_233
timestamp 1679235063
transform 1 0 8832 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_234
timestamp 1679235063
transform 1 0 13984 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_235
timestamp 1679235063
transform 1 0 19136 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_236
timestamp 1679235063
transform 1 0 24288 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_237
timestamp 1679235063
transform 1 0 6256 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_238
timestamp 1679235063
transform 1 0 11408 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_239
timestamp 1679235063
transform 1 0 16560 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_240
timestamp 1679235063
transform 1 0 21712 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_241
timestamp 1679235063
transform 1 0 3680 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_242
timestamp 1679235063
transform 1 0 8832 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_243
timestamp 1679235063
transform 1 0 13984 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_244
timestamp 1679235063
transform 1 0 19136 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_245
timestamp 1679235063
transform 1 0 24288 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_246
timestamp 1679235063
transform 1 0 6256 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_247
timestamp 1679235063
transform 1 0 11408 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_248
timestamp 1679235063
transform 1 0 16560 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_249
timestamp 1679235063
transform 1 0 21712 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_250
timestamp 1679235063
transform 1 0 3680 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_251
timestamp 1679235063
transform 1 0 8832 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_252
timestamp 1679235063
transform 1 0 13984 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_253
timestamp 1679235063
transform 1 0 19136 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_254
timestamp 1679235063
transform 1 0 24288 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_255
timestamp 1679235063
transform 1 0 6256 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_256
timestamp 1679235063
transform 1 0 11408 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_257
timestamp 1679235063
transform 1 0 16560 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_258
timestamp 1679235063
transform 1 0 21712 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_259
timestamp 1679235063
transform 1 0 3680 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_260
timestamp 1679235063
transform 1 0 8832 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_261
timestamp 1679235063
transform 1 0 13984 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_262
timestamp 1679235063
transform 1 0 19136 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_263
timestamp 1679235063
transform 1 0 24288 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_264
timestamp 1679235063
transform 1 0 6256 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_265
timestamp 1679235063
transform 1 0 11408 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_266
timestamp 1679235063
transform 1 0 16560 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_267
timestamp 1679235063
transform 1 0 21712 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_268
timestamp 1679235063
transform 1 0 3680 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_269
timestamp 1679235063
transform 1 0 8832 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_270
timestamp 1679235063
transform 1 0 13984 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_271
timestamp 1679235063
transform 1 0 19136 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_272
timestamp 1679235063
transform 1 0 24288 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_273
timestamp 1679235063
transform 1 0 6256 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_274
timestamp 1679235063
transform 1 0 11408 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_275
timestamp 1679235063
transform 1 0 16560 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_276
timestamp 1679235063
transform 1 0 21712 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_277
timestamp 1679235063
transform 1 0 3680 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_278
timestamp 1679235063
transform 1 0 8832 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_279
timestamp 1679235063
transform 1 0 13984 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_280
timestamp 1679235063
transform 1 0 19136 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_281
timestamp 1679235063
transform 1 0 24288 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_282
timestamp 1679235063
transform 1 0 6256 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_283
timestamp 1679235063
transform 1 0 11408 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_284
timestamp 1679235063
transform 1 0 16560 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_285
timestamp 1679235063
transform 1 0 21712 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_286
timestamp 1679235063
transform 1 0 3680 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_287
timestamp 1679235063
transform 1 0 8832 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_288
timestamp 1679235063
transform 1 0 13984 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_289
timestamp 1679235063
transform 1 0 19136 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_290
timestamp 1679235063
transform 1 0 24288 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_291
timestamp 1679235063
transform 1 0 6256 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_292
timestamp 1679235063
transform 1 0 11408 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_293
timestamp 1679235063
transform 1 0 16560 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_294
timestamp 1679235063
transform 1 0 21712 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_295
timestamp 1679235063
transform 1 0 3680 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_296
timestamp 1679235063
transform 1 0 8832 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_297
timestamp 1679235063
transform 1 0 13984 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_298
timestamp 1679235063
transform 1 0 19136 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_299
timestamp 1679235063
transform 1 0 24288 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_300
timestamp 1679235063
transform 1 0 6256 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_301
timestamp 1679235063
transform 1 0 11408 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_302
timestamp 1679235063
transform 1 0 16560 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_303
timestamp 1679235063
transform 1 0 21712 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_304
timestamp 1679235063
transform 1 0 3680 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_305
timestamp 1679235063
transform 1 0 8832 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_306
timestamp 1679235063
transform 1 0 13984 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_307
timestamp 1679235063
transform 1 0 19136 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_308
timestamp 1679235063
transform 1 0 24288 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_309
timestamp 1679235063
transform 1 0 6256 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_310
timestamp 1679235063
transform 1 0 11408 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_311
timestamp 1679235063
transform 1 0 16560 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_312
timestamp 1679235063
transform 1 0 21712 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_313
timestamp 1679235063
transform 1 0 3680 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_314
timestamp 1679235063
transform 1 0 8832 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_315
timestamp 1679235063
transform 1 0 13984 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_316
timestamp 1679235063
transform 1 0 19136 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_317
timestamp 1679235063
transform 1 0 24288 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_318
timestamp 1679235063
transform 1 0 6256 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_319
timestamp 1679235063
transform 1 0 11408 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_320
timestamp 1679235063
transform 1 0 16560 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_321
timestamp 1679235063
transform 1 0 21712 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_322
timestamp 1679235063
transform 1 0 3680 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_323
timestamp 1679235063
transform 1 0 8832 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_324
timestamp 1679235063
transform 1 0 13984 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_325
timestamp 1679235063
transform 1 0 19136 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_326
timestamp 1679235063
transform 1 0 24288 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_327
timestamp 1679235063
transform 1 0 6256 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_328
timestamp 1679235063
transform 1 0 11408 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_329
timestamp 1679235063
transform 1 0 16560 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_330
timestamp 1679235063
transform 1 0 21712 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_331
timestamp 1679235063
transform 1 0 3680 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_332
timestamp 1679235063
transform 1 0 8832 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_333
timestamp 1679235063
transform 1 0 13984 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_334
timestamp 1679235063
transform 1 0 19136 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_335
timestamp 1679235063
transform 1 0 24288 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_336
timestamp 1679235063
transform 1 0 6256 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_337
timestamp 1679235063
transform 1 0 11408 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_338
timestamp 1679235063
transform 1 0 16560 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_339
timestamp 1679235063
transform 1 0 21712 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_340
timestamp 1679235063
transform 1 0 3680 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_341
timestamp 1679235063
transform 1 0 8832 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_342
timestamp 1679235063
transform 1 0 13984 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_343
timestamp 1679235063
transform 1 0 19136 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_344
timestamp 1679235063
transform 1 0 24288 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_345
timestamp 1679235063
transform 1 0 6256 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_346
timestamp 1679235063
transform 1 0 11408 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_347
timestamp 1679235063
transform 1 0 16560 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_348
timestamp 1679235063
transform 1 0 21712 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_349
timestamp 1679235063
transform 1 0 3680 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_350
timestamp 1679235063
transform 1 0 8832 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_351
timestamp 1679235063
transform 1 0 13984 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_352
timestamp 1679235063
transform 1 0 19136 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_353
timestamp 1679235063
transform 1 0 24288 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_354
timestamp 1679235063
transform 1 0 6256 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_355
timestamp 1679235063
transform 1 0 11408 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_356
timestamp 1679235063
transform 1 0 16560 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_357
timestamp 1679235063
transform 1 0 21712 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_358
timestamp 1679235063
transform 1 0 3680 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_359
timestamp 1679235063
transform 1 0 8832 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_360
timestamp 1679235063
transform 1 0 13984 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_361
timestamp 1679235063
transform 1 0 19136 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_362
timestamp 1679235063
transform 1 0 24288 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_363
timestamp 1679235063
transform 1 0 6256 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_364
timestamp 1679235063
transform 1 0 11408 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_365
timestamp 1679235063
transform 1 0 16560 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_366
timestamp 1679235063
transform 1 0 21712 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_367
timestamp 1679235063
transform 1 0 3680 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_368
timestamp 1679235063
transform 1 0 8832 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_369
timestamp 1679235063
transform 1 0 13984 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_370
timestamp 1679235063
transform 1 0 19136 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_371
timestamp 1679235063
transform 1 0 24288 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_372
timestamp 1679235063
transform 1 0 6256 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_373
timestamp 1679235063
transform 1 0 11408 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_374
timestamp 1679235063
transform 1 0 16560 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_375
timestamp 1679235063
transform 1 0 21712 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_376
timestamp 1679235063
transform 1 0 3680 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_377
timestamp 1679235063
transform 1 0 8832 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_378
timestamp 1679235063
transform 1 0 13984 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_379
timestamp 1679235063
transform 1 0 19136 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_380
timestamp 1679235063
transform 1 0 24288 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_381
timestamp 1679235063
transform 1 0 6256 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_382
timestamp 1679235063
transform 1 0 11408 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_383
timestamp 1679235063
transform 1 0 16560 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_384
timestamp 1679235063
transform 1 0 21712 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_385
timestamp 1679235063
transform 1 0 3680 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_386
timestamp 1679235063
transform 1 0 8832 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_387
timestamp 1679235063
transform 1 0 13984 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_388
timestamp 1679235063
transform 1 0 19136 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_389
timestamp 1679235063
transform 1 0 24288 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_390
timestamp 1679235063
transform 1 0 6256 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_391
timestamp 1679235063
transform 1 0 11408 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_392
timestamp 1679235063
transform 1 0 16560 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_393
timestamp 1679235063
transform 1 0 21712 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_394
timestamp 1679235063
transform 1 0 3680 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_395
timestamp 1679235063
transform 1 0 8832 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_396
timestamp 1679235063
transform 1 0 13984 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_397
timestamp 1679235063
transform 1 0 19136 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_398
timestamp 1679235063
transform 1 0 24288 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_399
timestamp 1679235063
transform 1 0 6256 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_400
timestamp 1679235063
transform 1 0 11408 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_401
timestamp 1679235063
transform 1 0 16560 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_402
timestamp 1679235063
transform 1 0 21712 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_403
timestamp 1679235063
transform 1 0 3680 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_404
timestamp 1679235063
transform 1 0 8832 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_405
timestamp 1679235063
transform 1 0 13984 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_406
timestamp 1679235063
transform 1 0 19136 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_407
timestamp 1679235063
transform 1 0 24288 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_408
timestamp 1679235063
transform 1 0 6256 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_409
timestamp 1679235063
transform 1 0 11408 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_410
timestamp 1679235063
transform 1 0 16560 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_411
timestamp 1679235063
transform 1 0 21712 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_412
timestamp 1679235063
transform 1 0 3680 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_413
timestamp 1679235063
transform 1 0 8832 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_414
timestamp 1679235063
transform 1 0 13984 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_415
timestamp 1679235063
transform 1 0 19136 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_416
timestamp 1679235063
transform 1 0 24288 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_417
timestamp 1679235063
transform 1 0 6256 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_418
timestamp 1679235063
transform 1 0 11408 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_419
timestamp 1679235063
transform 1 0 16560 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_420
timestamp 1679235063
transform 1 0 21712 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_421
timestamp 1679235063
transform 1 0 3680 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_422
timestamp 1679235063
transform 1 0 8832 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_423
timestamp 1679235063
transform 1 0 13984 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_424
timestamp 1679235063
transform 1 0 19136 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_425
timestamp 1679235063
transform 1 0 24288 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_426
timestamp 1679235063
transform 1 0 6256 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_427
timestamp 1679235063
transform 1 0 11408 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_428
timestamp 1679235063
transform 1 0 16560 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_429
timestamp 1679235063
transform 1 0 21712 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_430
timestamp 1679235063
transform 1 0 3680 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_431
timestamp 1679235063
transform 1 0 8832 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_432
timestamp 1679235063
transform 1 0 13984 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_433
timestamp 1679235063
transform 1 0 19136 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_434
timestamp 1679235063
transform 1 0 24288 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_435
timestamp 1679235063
transform 1 0 6256 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_436
timestamp 1679235063
transform 1 0 11408 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_437
timestamp 1679235063
transform 1 0 16560 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_438
timestamp 1679235063
transform 1 0 21712 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_439
timestamp 1679235063
transform 1 0 3680 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_440
timestamp 1679235063
transform 1 0 8832 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_441
timestamp 1679235063
transform 1 0 13984 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_442
timestamp 1679235063
transform 1 0 19136 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_443
timestamp 1679235063
transform 1 0 24288 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_444
timestamp 1679235063
transform 1 0 6256 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_445
timestamp 1679235063
transform 1 0 11408 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_446
timestamp 1679235063
transform 1 0 16560 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_447
timestamp 1679235063
transform 1 0 21712 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_448
timestamp 1679235063
transform 1 0 3680 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_449
timestamp 1679235063
transform 1 0 8832 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_450
timestamp 1679235063
transform 1 0 13984 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_451
timestamp 1679235063
transform 1 0 19136 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_452
timestamp 1679235063
transform 1 0 24288 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_453
timestamp 1679235063
transform 1 0 6256 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_454
timestamp 1679235063
transform 1 0 11408 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_455
timestamp 1679235063
transform 1 0 16560 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_456
timestamp 1679235063
transform 1 0 21712 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_457
timestamp 1679235063
transform 1 0 3680 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_458
timestamp 1679235063
transform 1 0 8832 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_459
timestamp 1679235063
transform 1 0 13984 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_460
timestamp 1679235063
transform 1 0 19136 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_461
timestamp 1679235063
transform 1 0 24288 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_462
timestamp 1679235063
transform 1 0 6256 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_463
timestamp 1679235063
transform 1 0 11408 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_464
timestamp 1679235063
transform 1 0 16560 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_465
timestamp 1679235063
transform 1 0 21712 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_466
timestamp 1679235063
transform 1 0 3680 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_467
timestamp 1679235063
transform 1 0 8832 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_468
timestamp 1679235063
transform 1 0 13984 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_469
timestamp 1679235063
transform 1 0 19136 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_470
timestamp 1679235063
transform 1 0 24288 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_471
timestamp 1679235063
transform 1 0 6256 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_472
timestamp 1679235063
transform 1 0 11408 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_473
timestamp 1679235063
transform 1 0 16560 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_474
timestamp 1679235063
transform 1 0 21712 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_475
timestamp 1679235063
transform 1 0 3680 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_476
timestamp 1679235063
transform 1 0 8832 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_477
timestamp 1679235063
transform 1 0 13984 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_478
timestamp 1679235063
transform 1 0 19136 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_479
timestamp 1679235063
transform 1 0 24288 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_480
timestamp 1679235063
transform 1 0 6256 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_481
timestamp 1679235063
transform 1 0 11408 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_482
timestamp 1679235063
transform 1 0 16560 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_483
timestamp 1679235063
transform 1 0 21712 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_484
timestamp 1679235063
transform 1 0 3680 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_485
timestamp 1679235063
transform 1 0 8832 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_486
timestamp 1679235063
transform 1 0 13984 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_487
timestamp 1679235063
transform 1 0 19136 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_488
timestamp 1679235063
transform 1 0 24288 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_489
timestamp 1679235063
transform 1 0 6256 0 -1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_490
timestamp 1679235063
transform 1 0 11408 0 -1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_491
timestamp 1679235063
transform 1 0 16560 0 -1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_492
timestamp 1679235063
transform 1 0 21712 0 -1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_493
timestamp 1679235063
transform 1 0 3680 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_494
timestamp 1679235063
transform 1 0 8832 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_495
timestamp 1679235063
transform 1 0 13984 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_496
timestamp 1679235063
transform 1 0 19136 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_497
timestamp 1679235063
transform 1 0 24288 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_498
timestamp 1679235063
transform 1 0 6256 0 -1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_499
timestamp 1679235063
transform 1 0 11408 0 -1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_500
timestamp 1679235063
transform 1 0 16560 0 -1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_501
timestamp 1679235063
transform 1 0 21712 0 -1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_502
timestamp 1679235063
transform 1 0 3680 0 1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_503
timestamp 1679235063
transform 1 0 8832 0 1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_504
timestamp 1679235063
transform 1 0 13984 0 1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_505
timestamp 1679235063
transform 1 0 19136 0 1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_506
timestamp 1679235063
transform 1 0 24288 0 1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_507
timestamp 1679235063
transform 1 0 6256 0 -1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_508
timestamp 1679235063
transform 1 0 11408 0 -1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_509
timestamp 1679235063
transform 1 0 16560 0 -1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_510
timestamp 1679235063
transform 1 0 21712 0 -1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_511
timestamp 1679235063
transform 1 0 3680 0 1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_512
timestamp 1679235063
transform 1 0 8832 0 1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_513
timestamp 1679235063
transform 1 0 13984 0 1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_514
timestamp 1679235063
transform 1 0 19136 0 1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_515
timestamp 1679235063
transform 1 0 24288 0 1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_516
timestamp 1679235063
transform 1 0 6256 0 -1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_517
timestamp 1679235063
transform 1 0 11408 0 -1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_518
timestamp 1679235063
transform 1 0 16560 0 -1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_519
timestamp 1679235063
transform 1 0 21712 0 -1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_520
timestamp 1679235063
transform 1 0 3680 0 1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_521
timestamp 1679235063
transform 1 0 8832 0 1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_522
timestamp 1679235063
transform 1 0 13984 0 1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_523
timestamp 1679235063
transform 1 0 19136 0 1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_524
timestamp 1679235063
transform 1 0 24288 0 1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_525
timestamp 1679235063
transform 1 0 6256 0 -1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_526
timestamp 1679235063
transform 1 0 11408 0 -1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_527
timestamp 1679235063
transform 1 0 16560 0 -1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_528
timestamp 1679235063
transform 1 0 21712 0 -1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_529
timestamp 1679235063
transform 1 0 3680 0 1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_530
timestamp 1679235063
transform 1 0 8832 0 1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_531
timestamp 1679235063
transform 1 0 13984 0 1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_532
timestamp 1679235063
transform 1 0 19136 0 1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_533
timestamp 1679235063
transform 1 0 24288 0 1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_534
timestamp 1679235063
transform 1 0 6256 0 -1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_535
timestamp 1679235063
transform 1 0 11408 0 -1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_536
timestamp 1679235063
transform 1 0 16560 0 -1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_537
timestamp 1679235063
transform 1 0 21712 0 -1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_538
timestamp 1679235063
transform 1 0 3680 0 1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_539
timestamp 1679235063
transform 1 0 8832 0 1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_540
timestamp 1679235063
transform 1 0 13984 0 1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_541
timestamp 1679235063
transform 1 0 19136 0 1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_542
timestamp 1679235063
transform 1 0 24288 0 1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_543
timestamp 1679235063
transform 1 0 6256 0 -1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_544
timestamp 1679235063
transform 1 0 11408 0 -1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_545
timestamp 1679235063
transform 1 0 16560 0 -1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_546
timestamp 1679235063
transform 1 0 21712 0 -1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_547
timestamp 1679235063
transform 1 0 3680 0 1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_548
timestamp 1679235063
transform 1 0 8832 0 1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_549
timestamp 1679235063
transform 1 0 13984 0 1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_550
timestamp 1679235063
transform 1 0 19136 0 1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_551
timestamp 1679235063
transform 1 0 24288 0 1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_552
timestamp 1679235063
transform 1 0 6256 0 -1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_553
timestamp 1679235063
transform 1 0 11408 0 -1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_554
timestamp 1679235063
transform 1 0 16560 0 -1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_555
timestamp 1679235063
transform 1 0 21712 0 -1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_556
timestamp 1679235063
transform 1 0 3680 0 1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_557
timestamp 1679235063
transform 1 0 8832 0 1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_558
timestamp 1679235063
transform 1 0 13984 0 1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_559
timestamp 1679235063
transform 1 0 19136 0 1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_560
timestamp 1679235063
transform 1 0 24288 0 1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_561
timestamp 1679235063
transform 1 0 6256 0 -1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_562
timestamp 1679235063
transform 1 0 11408 0 -1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_563
timestamp 1679235063
transform 1 0 16560 0 -1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_564
timestamp 1679235063
transform 1 0 21712 0 -1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_565
timestamp 1679235063
transform 1 0 3680 0 1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_566
timestamp 1679235063
transform 1 0 8832 0 1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_567
timestamp 1679235063
transform 1 0 13984 0 1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_568
timestamp 1679235063
transform 1 0 19136 0 1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_569
timestamp 1679235063
transform 1 0 24288 0 1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_570
timestamp 1679235063
transform 1 0 6256 0 -1 47872
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_571
timestamp 1679235063
transform 1 0 11408 0 -1 47872
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_572
timestamp 1679235063
transform 1 0 16560 0 -1 47872
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_573
timestamp 1679235063
transform 1 0 21712 0 -1 47872
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_574
timestamp 1679235063
transform 1 0 3680 0 1 47872
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_575
timestamp 1679235063
transform 1 0 8832 0 1 47872
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_576
timestamp 1679235063
transform 1 0 13984 0 1 47872
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_577
timestamp 1679235063
transform 1 0 19136 0 1 47872
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_578
timestamp 1679235063
transform 1 0 24288 0 1 47872
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_579
timestamp 1679235063
transform 1 0 6256 0 -1 48960
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_580
timestamp 1679235063
transform 1 0 11408 0 -1 48960
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_581
timestamp 1679235063
transform 1 0 16560 0 -1 48960
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_582
timestamp 1679235063
transform 1 0 21712 0 -1 48960
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_583
timestamp 1679235063
transform 1 0 3680 0 1 48960
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_584
timestamp 1679235063
transform 1 0 8832 0 1 48960
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_585
timestamp 1679235063
transform 1 0 13984 0 1 48960
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_586
timestamp 1679235063
transform 1 0 19136 0 1 48960
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_587
timestamp 1679235063
transform 1 0 24288 0 1 48960
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_588
timestamp 1679235063
transform 1 0 6256 0 -1 50048
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_589
timestamp 1679235063
transform 1 0 11408 0 -1 50048
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_590
timestamp 1679235063
transform 1 0 16560 0 -1 50048
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_591
timestamp 1679235063
transform 1 0 21712 0 -1 50048
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_592
timestamp 1679235063
transform 1 0 3680 0 1 50048
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_593
timestamp 1679235063
transform 1 0 8832 0 1 50048
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_594
timestamp 1679235063
transform 1 0 13984 0 1 50048
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_595
timestamp 1679235063
transform 1 0 19136 0 1 50048
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_596
timestamp 1679235063
transform 1 0 24288 0 1 50048
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_597
timestamp 1679235063
transform 1 0 6256 0 -1 51136
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_598
timestamp 1679235063
transform 1 0 11408 0 -1 51136
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_599
timestamp 1679235063
transform 1 0 16560 0 -1 51136
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_600
timestamp 1679235063
transform 1 0 21712 0 -1 51136
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_601
timestamp 1679235063
transform 1 0 3680 0 1 51136
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_602
timestamp 1679235063
transform 1 0 8832 0 1 51136
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_603
timestamp 1679235063
transform 1 0 13984 0 1 51136
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_604
timestamp 1679235063
transform 1 0 19136 0 1 51136
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_605
timestamp 1679235063
transform 1 0 24288 0 1 51136
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_606
timestamp 1679235063
transform 1 0 6256 0 -1 52224
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_607
timestamp 1679235063
transform 1 0 11408 0 -1 52224
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_608
timestamp 1679235063
transform 1 0 16560 0 -1 52224
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_609
timestamp 1679235063
transform 1 0 21712 0 -1 52224
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_610
timestamp 1679235063
transform 1 0 3680 0 1 52224
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_611
timestamp 1679235063
transform 1 0 8832 0 1 52224
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_612
timestamp 1679235063
transform 1 0 13984 0 1 52224
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_613
timestamp 1679235063
transform 1 0 19136 0 1 52224
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_614
timestamp 1679235063
transform 1 0 24288 0 1 52224
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_615
timestamp 1679235063
transform 1 0 6256 0 -1 53312
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_616
timestamp 1679235063
transform 1 0 11408 0 -1 53312
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_617
timestamp 1679235063
transform 1 0 16560 0 -1 53312
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_618
timestamp 1679235063
transform 1 0 21712 0 -1 53312
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_619
timestamp 1679235063
transform 1 0 3680 0 1 53312
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_620
timestamp 1679235063
transform 1 0 8832 0 1 53312
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_621
timestamp 1679235063
transform 1 0 13984 0 1 53312
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_622
timestamp 1679235063
transform 1 0 19136 0 1 53312
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_623
timestamp 1679235063
transform 1 0 24288 0 1 53312
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_624
timestamp 1679235063
transform 1 0 3680 0 -1 54400
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_625
timestamp 1679235063
transform 1 0 6256 0 -1 54400
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_626
timestamp 1679235063
transform 1 0 8832 0 -1 54400
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_627
timestamp 1679235063
transform 1 0 11408 0 -1 54400
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_628
timestamp 1679235063
transform 1 0 13984 0 -1 54400
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_629
timestamp 1679235063
transform 1 0 16560 0 -1 54400
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_630
timestamp 1679235063
transform 1 0 19136 0 -1 54400
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_631
timestamp 1679235063
transform 1 0 21712 0 -1 54400
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_632
timestamp 1679235063
transform 1 0 24288 0 -1 54400
box -38 -48 130 592
<< labels >>
flabel metal4 s 7944 2128 8264 54448 0 FreeSans 1920 90 0 0 VGND
port 0 nsew ground bidirectional
flabel metal4 s 17944 2128 18264 54448 0 FreeSans 1920 90 0 0 VGND
port 0 nsew ground bidirectional
flabel metal4 s 2944 2128 3264 54448 0 FreeSans 1920 90 0 0 VPWR
port 1 nsew power bidirectional
flabel metal4 s 12944 2128 13264 54448 0 FreeSans 1920 90 0 0 VPWR
port 1 nsew power bidirectional
flabel metal4 s 22944 2128 23264 54448 0 FreeSans 1920 90 0 0 VPWR
port 1 nsew power bidirectional
flabel metal3 s 0 55360 800 55480 0 FreeSans 480 0 0 0 ccff_head
port 2 nsew signal input
flabel metal3 s 0 1504 800 1624 0 FreeSans 480 0 0 0 ccff_head_0
port 3 nsew signal input
flabel metal3 s 26200 688 27000 808 0 FreeSans 480 0 0 0 ccff_tail
port 4 nsew signal tristate
flabel metal2 s 1490 56200 1546 57000 0 FreeSans 224 90 0 0 ccff_tail_0
port 5 nsew signal tristate
flabel metal3 s 26200 25984 27000 26104 0 FreeSans 480 0 0 0 chanx_right_in[0]
port 6 nsew signal input
flabel metal3 s 26200 34144 27000 34264 0 FreeSans 480 0 0 0 chanx_right_in[10]
port 7 nsew signal input
flabel metal3 s 26200 34960 27000 35080 0 FreeSans 480 0 0 0 chanx_right_in[11]
port 8 nsew signal input
flabel metal3 s 26200 35776 27000 35896 0 FreeSans 480 0 0 0 chanx_right_in[12]
port 9 nsew signal input
flabel metal3 s 26200 36592 27000 36712 0 FreeSans 480 0 0 0 chanx_right_in[13]
port 10 nsew signal input
flabel metal3 s 26200 37408 27000 37528 0 FreeSans 480 0 0 0 chanx_right_in[14]
port 11 nsew signal input
flabel metal3 s 26200 38224 27000 38344 0 FreeSans 480 0 0 0 chanx_right_in[15]
port 12 nsew signal input
flabel metal3 s 26200 39040 27000 39160 0 FreeSans 480 0 0 0 chanx_right_in[16]
port 13 nsew signal input
flabel metal3 s 26200 39856 27000 39976 0 FreeSans 480 0 0 0 chanx_right_in[17]
port 14 nsew signal input
flabel metal3 s 26200 40672 27000 40792 0 FreeSans 480 0 0 0 chanx_right_in[18]
port 15 nsew signal input
flabel metal3 s 26200 41488 27000 41608 0 FreeSans 480 0 0 0 chanx_right_in[19]
port 16 nsew signal input
flabel metal3 s 26200 26800 27000 26920 0 FreeSans 480 0 0 0 chanx_right_in[1]
port 17 nsew signal input
flabel metal3 s 26200 42304 27000 42424 0 FreeSans 480 0 0 0 chanx_right_in[20]
port 18 nsew signal input
flabel metal3 s 26200 43120 27000 43240 0 FreeSans 480 0 0 0 chanx_right_in[21]
port 19 nsew signal input
flabel metal3 s 26200 43936 27000 44056 0 FreeSans 480 0 0 0 chanx_right_in[22]
port 20 nsew signal input
flabel metal3 s 26200 44752 27000 44872 0 FreeSans 480 0 0 0 chanx_right_in[23]
port 21 nsew signal input
flabel metal3 s 26200 45568 27000 45688 0 FreeSans 480 0 0 0 chanx_right_in[24]
port 22 nsew signal input
flabel metal3 s 26200 46384 27000 46504 0 FreeSans 480 0 0 0 chanx_right_in[25]
port 23 nsew signal input
flabel metal3 s 26200 47200 27000 47320 0 FreeSans 480 0 0 0 chanx_right_in[26]
port 24 nsew signal input
flabel metal3 s 26200 48016 27000 48136 0 FreeSans 480 0 0 0 chanx_right_in[27]
port 25 nsew signal input
flabel metal3 s 26200 48832 27000 48952 0 FreeSans 480 0 0 0 chanx_right_in[28]
port 26 nsew signal input
flabel metal3 s 26200 49648 27000 49768 0 FreeSans 480 0 0 0 chanx_right_in[29]
port 27 nsew signal input
flabel metal3 s 26200 27616 27000 27736 0 FreeSans 480 0 0 0 chanx_right_in[2]
port 28 nsew signal input
flabel metal3 s 26200 28432 27000 28552 0 FreeSans 480 0 0 0 chanx_right_in[3]
port 29 nsew signal input
flabel metal3 s 26200 29248 27000 29368 0 FreeSans 480 0 0 0 chanx_right_in[4]
port 30 nsew signal input
flabel metal3 s 26200 30064 27000 30184 0 FreeSans 480 0 0 0 chanx_right_in[5]
port 31 nsew signal input
flabel metal3 s 26200 30880 27000 31000 0 FreeSans 480 0 0 0 chanx_right_in[6]
port 32 nsew signal input
flabel metal3 s 26200 31696 27000 31816 0 FreeSans 480 0 0 0 chanx_right_in[7]
port 33 nsew signal input
flabel metal3 s 26200 32512 27000 32632 0 FreeSans 480 0 0 0 chanx_right_in[8]
port 34 nsew signal input
flabel metal3 s 26200 33328 27000 33448 0 FreeSans 480 0 0 0 chanx_right_in[9]
port 35 nsew signal input
flabel metal3 s 26200 1504 27000 1624 0 FreeSans 480 0 0 0 chanx_right_out[0]
port 36 nsew signal tristate
flabel metal3 s 26200 9664 27000 9784 0 FreeSans 480 0 0 0 chanx_right_out[10]
port 37 nsew signal tristate
flabel metal3 s 26200 10480 27000 10600 0 FreeSans 480 0 0 0 chanx_right_out[11]
port 38 nsew signal tristate
flabel metal3 s 26200 11296 27000 11416 0 FreeSans 480 0 0 0 chanx_right_out[12]
port 39 nsew signal tristate
flabel metal3 s 26200 12112 27000 12232 0 FreeSans 480 0 0 0 chanx_right_out[13]
port 40 nsew signal tristate
flabel metal3 s 26200 12928 27000 13048 0 FreeSans 480 0 0 0 chanx_right_out[14]
port 41 nsew signal tristate
flabel metal3 s 26200 13744 27000 13864 0 FreeSans 480 0 0 0 chanx_right_out[15]
port 42 nsew signal tristate
flabel metal3 s 26200 14560 27000 14680 0 FreeSans 480 0 0 0 chanx_right_out[16]
port 43 nsew signal tristate
flabel metal3 s 26200 15376 27000 15496 0 FreeSans 480 0 0 0 chanx_right_out[17]
port 44 nsew signal tristate
flabel metal3 s 26200 16192 27000 16312 0 FreeSans 480 0 0 0 chanx_right_out[18]
port 45 nsew signal tristate
flabel metal3 s 26200 17008 27000 17128 0 FreeSans 480 0 0 0 chanx_right_out[19]
port 46 nsew signal tristate
flabel metal3 s 26200 2320 27000 2440 0 FreeSans 480 0 0 0 chanx_right_out[1]
port 47 nsew signal tristate
flabel metal3 s 26200 17824 27000 17944 0 FreeSans 480 0 0 0 chanx_right_out[20]
port 48 nsew signal tristate
flabel metal3 s 26200 18640 27000 18760 0 FreeSans 480 0 0 0 chanx_right_out[21]
port 49 nsew signal tristate
flabel metal3 s 26200 19456 27000 19576 0 FreeSans 480 0 0 0 chanx_right_out[22]
port 50 nsew signal tristate
flabel metal3 s 26200 20272 27000 20392 0 FreeSans 480 0 0 0 chanx_right_out[23]
port 51 nsew signal tristate
flabel metal3 s 26200 21088 27000 21208 0 FreeSans 480 0 0 0 chanx_right_out[24]
port 52 nsew signal tristate
flabel metal3 s 26200 21904 27000 22024 0 FreeSans 480 0 0 0 chanx_right_out[25]
port 53 nsew signal tristate
flabel metal3 s 26200 22720 27000 22840 0 FreeSans 480 0 0 0 chanx_right_out[26]
port 54 nsew signal tristate
flabel metal3 s 26200 23536 27000 23656 0 FreeSans 480 0 0 0 chanx_right_out[27]
port 55 nsew signal tristate
flabel metal3 s 26200 24352 27000 24472 0 FreeSans 480 0 0 0 chanx_right_out[28]
port 56 nsew signal tristate
flabel metal3 s 26200 25168 27000 25288 0 FreeSans 480 0 0 0 chanx_right_out[29]
port 57 nsew signal tristate
flabel metal3 s 26200 3136 27000 3256 0 FreeSans 480 0 0 0 chanx_right_out[2]
port 58 nsew signal tristate
flabel metal3 s 26200 3952 27000 4072 0 FreeSans 480 0 0 0 chanx_right_out[3]
port 59 nsew signal tristate
flabel metal3 s 26200 4768 27000 4888 0 FreeSans 480 0 0 0 chanx_right_out[4]
port 60 nsew signal tristate
flabel metal3 s 26200 5584 27000 5704 0 FreeSans 480 0 0 0 chanx_right_out[5]
port 61 nsew signal tristate
flabel metal3 s 26200 6400 27000 6520 0 FreeSans 480 0 0 0 chanx_right_out[6]
port 62 nsew signal tristate
flabel metal3 s 26200 7216 27000 7336 0 FreeSans 480 0 0 0 chanx_right_out[7]
port 63 nsew signal tristate
flabel metal3 s 26200 8032 27000 8152 0 FreeSans 480 0 0 0 chanx_right_out[8]
port 64 nsew signal tristate
flabel metal3 s 26200 8848 27000 8968 0 FreeSans 480 0 0 0 chanx_right_out[9]
port 65 nsew signal tristate
flabel metal2 s 1674 0 1730 800 0 FreeSans 224 90 0 0 chany_bottom_in[0]
port 66 nsew signal input
flabel metal2 s 5354 0 5410 800 0 FreeSans 224 90 0 0 chany_bottom_in[10]
port 67 nsew signal input
flabel metal2 s 5722 0 5778 800 0 FreeSans 224 90 0 0 chany_bottom_in[11]
port 68 nsew signal input
flabel metal2 s 6090 0 6146 800 0 FreeSans 224 90 0 0 chany_bottom_in[12]
port 69 nsew signal input
flabel metal2 s 6458 0 6514 800 0 FreeSans 224 90 0 0 chany_bottom_in[13]
port 70 nsew signal input
flabel metal2 s 6826 0 6882 800 0 FreeSans 224 90 0 0 chany_bottom_in[14]
port 71 nsew signal input
flabel metal2 s 7194 0 7250 800 0 FreeSans 224 90 0 0 chany_bottom_in[15]
port 72 nsew signal input
flabel metal2 s 7562 0 7618 800 0 FreeSans 224 90 0 0 chany_bottom_in[16]
port 73 nsew signal input
flabel metal2 s 7930 0 7986 800 0 FreeSans 224 90 0 0 chany_bottom_in[17]
port 74 nsew signal input
flabel metal2 s 8298 0 8354 800 0 FreeSans 224 90 0 0 chany_bottom_in[18]
port 75 nsew signal input
flabel metal2 s 8666 0 8722 800 0 FreeSans 224 90 0 0 chany_bottom_in[19]
port 76 nsew signal input
flabel metal2 s 2042 0 2098 800 0 FreeSans 224 90 0 0 chany_bottom_in[1]
port 77 nsew signal input
flabel metal2 s 9034 0 9090 800 0 FreeSans 224 90 0 0 chany_bottom_in[20]
port 78 nsew signal input
flabel metal2 s 9402 0 9458 800 0 FreeSans 224 90 0 0 chany_bottom_in[21]
port 79 nsew signal input
flabel metal2 s 9770 0 9826 800 0 FreeSans 224 90 0 0 chany_bottom_in[22]
port 80 nsew signal input
flabel metal2 s 10138 0 10194 800 0 FreeSans 224 90 0 0 chany_bottom_in[23]
port 81 nsew signal input
flabel metal2 s 10506 0 10562 800 0 FreeSans 224 90 0 0 chany_bottom_in[24]
port 82 nsew signal input
flabel metal2 s 10874 0 10930 800 0 FreeSans 224 90 0 0 chany_bottom_in[25]
port 83 nsew signal input
flabel metal2 s 11242 0 11298 800 0 FreeSans 224 90 0 0 chany_bottom_in[26]
port 84 nsew signal input
flabel metal2 s 11610 0 11666 800 0 FreeSans 224 90 0 0 chany_bottom_in[27]
port 85 nsew signal input
flabel metal2 s 11978 0 12034 800 0 FreeSans 224 90 0 0 chany_bottom_in[28]
port 86 nsew signal input
flabel metal2 s 12346 0 12402 800 0 FreeSans 224 90 0 0 chany_bottom_in[29]
port 87 nsew signal input
flabel metal2 s 2410 0 2466 800 0 FreeSans 224 90 0 0 chany_bottom_in[2]
port 88 nsew signal input
flabel metal2 s 2778 0 2834 800 0 FreeSans 224 90 0 0 chany_bottom_in[3]
port 89 nsew signal input
flabel metal2 s 3146 0 3202 800 0 FreeSans 224 90 0 0 chany_bottom_in[4]
port 90 nsew signal input
flabel metal2 s 3514 0 3570 800 0 FreeSans 224 90 0 0 chany_bottom_in[5]
port 91 nsew signal input
flabel metal2 s 3882 0 3938 800 0 FreeSans 224 90 0 0 chany_bottom_in[6]
port 92 nsew signal input
flabel metal2 s 4250 0 4306 800 0 FreeSans 224 90 0 0 chany_bottom_in[7]
port 93 nsew signal input
flabel metal2 s 4618 0 4674 800 0 FreeSans 224 90 0 0 chany_bottom_in[8]
port 94 nsew signal input
flabel metal2 s 4986 0 5042 800 0 FreeSans 224 90 0 0 chany_bottom_in[9]
port 95 nsew signal input
flabel metal2 s 12714 0 12770 800 0 FreeSans 224 90 0 0 chany_bottom_out[0]
port 96 nsew signal tristate
flabel metal2 s 16394 0 16450 800 0 FreeSans 224 90 0 0 chany_bottom_out[10]
port 97 nsew signal tristate
flabel metal2 s 16762 0 16818 800 0 FreeSans 224 90 0 0 chany_bottom_out[11]
port 98 nsew signal tristate
flabel metal2 s 17130 0 17186 800 0 FreeSans 224 90 0 0 chany_bottom_out[12]
port 99 nsew signal tristate
flabel metal2 s 17498 0 17554 800 0 FreeSans 224 90 0 0 chany_bottom_out[13]
port 100 nsew signal tristate
flabel metal2 s 17866 0 17922 800 0 FreeSans 224 90 0 0 chany_bottom_out[14]
port 101 nsew signal tristate
flabel metal2 s 18234 0 18290 800 0 FreeSans 224 90 0 0 chany_bottom_out[15]
port 102 nsew signal tristate
flabel metal2 s 18602 0 18658 800 0 FreeSans 224 90 0 0 chany_bottom_out[16]
port 103 nsew signal tristate
flabel metal2 s 18970 0 19026 800 0 FreeSans 224 90 0 0 chany_bottom_out[17]
port 104 nsew signal tristate
flabel metal2 s 19338 0 19394 800 0 FreeSans 224 90 0 0 chany_bottom_out[18]
port 105 nsew signal tristate
flabel metal2 s 19706 0 19762 800 0 FreeSans 224 90 0 0 chany_bottom_out[19]
port 106 nsew signal tristate
flabel metal2 s 13082 0 13138 800 0 FreeSans 224 90 0 0 chany_bottom_out[1]
port 107 nsew signal tristate
flabel metal2 s 20074 0 20130 800 0 FreeSans 224 90 0 0 chany_bottom_out[20]
port 108 nsew signal tristate
flabel metal2 s 20442 0 20498 800 0 FreeSans 224 90 0 0 chany_bottom_out[21]
port 109 nsew signal tristate
flabel metal2 s 20810 0 20866 800 0 FreeSans 224 90 0 0 chany_bottom_out[22]
port 110 nsew signal tristate
flabel metal2 s 21178 0 21234 800 0 FreeSans 224 90 0 0 chany_bottom_out[23]
port 111 nsew signal tristate
flabel metal2 s 21546 0 21602 800 0 FreeSans 224 90 0 0 chany_bottom_out[24]
port 112 nsew signal tristate
flabel metal2 s 21914 0 21970 800 0 FreeSans 224 90 0 0 chany_bottom_out[25]
port 113 nsew signal tristate
flabel metal2 s 22282 0 22338 800 0 FreeSans 224 90 0 0 chany_bottom_out[26]
port 114 nsew signal tristate
flabel metal2 s 22650 0 22706 800 0 FreeSans 224 90 0 0 chany_bottom_out[27]
port 115 nsew signal tristate
flabel metal2 s 23018 0 23074 800 0 FreeSans 224 90 0 0 chany_bottom_out[28]
port 116 nsew signal tristate
flabel metal2 s 23386 0 23442 800 0 FreeSans 224 90 0 0 chany_bottom_out[29]
port 117 nsew signal tristate
flabel metal2 s 13450 0 13506 800 0 FreeSans 224 90 0 0 chany_bottom_out[2]
port 118 nsew signal tristate
flabel metal2 s 13818 0 13874 800 0 FreeSans 224 90 0 0 chany_bottom_out[3]
port 119 nsew signal tristate
flabel metal2 s 14186 0 14242 800 0 FreeSans 224 90 0 0 chany_bottom_out[4]
port 120 nsew signal tristate
flabel metal2 s 14554 0 14610 800 0 FreeSans 224 90 0 0 chany_bottom_out[5]
port 121 nsew signal tristate
flabel metal2 s 14922 0 14978 800 0 FreeSans 224 90 0 0 chany_bottom_out[6]
port 122 nsew signal tristate
flabel metal2 s 15290 0 15346 800 0 FreeSans 224 90 0 0 chany_bottom_out[7]
port 123 nsew signal tristate
flabel metal2 s 15658 0 15714 800 0 FreeSans 224 90 0 0 chany_bottom_out[8]
port 124 nsew signal tristate
flabel metal2 s 16026 0 16082 800 0 FreeSans 224 90 0 0 chany_bottom_out[9]
port 125 nsew signal tristate
flabel metal2 s 12898 56200 12954 57000 0 FreeSans 224 90 0 0 chany_top_in_0[0]
port 126 nsew signal input
flabel metal2 s 16578 56200 16634 57000 0 FreeSans 224 90 0 0 chany_top_in_0[10]
port 127 nsew signal input
flabel metal2 s 16946 56200 17002 57000 0 FreeSans 224 90 0 0 chany_top_in_0[11]
port 128 nsew signal input
flabel metal2 s 17314 56200 17370 57000 0 FreeSans 224 90 0 0 chany_top_in_0[12]
port 129 nsew signal input
flabel metal2 s 17682 56200 17738 57000 0 FreeSans 224 90 0 0 chany_top_in_0[13]
port 130 nsew signal input
flabel metal2 s 18050 56200 18106 57000 0 FreeSans 224 90 0 0 chany_top_in_0[14]
port 131 nsew signal input
flabel metal2 s 18418 56200 18474 57000 0 FreeSans 224 90 0 0 chany_top_in_0[15]
port 132 nsew signal input
flabel metal2 s 18786 56200 18842 57000 0 FreeSans 224 90 0 0 chany_top_in_0[16]
port 133 nsew signal input
flabel metal2 s 19154 56200 19210 57000 0 FreeSans 224 90 0 0 chany_top_in_0[17]
port 134 nsew signal input
flabel metal2 s 19522 56200 19578 57000 0 FreeSans 224 90 0 0 chany_top_in_0[18]
port 135 nsew signal input
flabel metal2 s 19890 56200 19946 57000 0 FreeSans 224 90 0 0 chany_top_in_0[19]
port 136 nsew signal input
flabel metal2 s 13266 56200 13322 57000 0 FreeSans 224 90 0 0 chany_top_in_0[1]
port 137 nsew signal input
flabel metal2 s 20258 56200 20314 57000 0 FreeSans 224 90 0 0 chany_top_in_0[20]
port 138 nsew signal input
flabel metal2 s 20626 56200 20682 57000 0 FreeSans 224 90 0 0 chany_top_in_0[21]
port 139 nsew signal input
flabel metal2 s 20994 56200 21050 57000 0 FreeSans 224 90 0 0 chany_top_in_0[22]
port 140 nsew signal input
flabel metal2 s 21362 56200 21418 57000 0 FreeSans 224 90 0 0 chany_top_in_0[23]
port 141 nsew signal input
flabel metal2 s 21730 56200 21786 57000 0 FreeSans 224 90 0 0 chany_top_in_0[24]
port 142 nsew signal input
flabel metal2 s 22098 56200 22154 57000 0 FreeSans 224 90 0 0 chany_top_in_0[25]
port 143 nsew signal input
flabel metal2 s 22466 56200 22522 57000 0 FreeSans 224 90 0 0 chany_top_in_0[26]
port 144 nsew signal input
flabel metal2 s 22834 56200 22890 57000 0 FreeSans 224 90 0 0 chany_top_in_0[27]
port 145 nsew signal input
flabel metal2 s 23202 56200 23258 57000 0 FreeSans 224 90 0 0 chany_top_in_0[28]
port 146 nsew signal input
flabel metal2 s 23570 56200 23626 57000 0 FreeSans 224 90 0 0 chany_top_in_0[29]
port 147 nsew signal input
flabel metal2 s 13634 56200 13690 57000 0 FreeSans 224 90 0 0 chany_top_in_0[2]
port 148 nsew signal input
flabel metal2 s 14002 56200 14058 57000 0 FreeSans 224 90 0 0 chany_top_in_0[3]
port 149 nsew signal input
flabel metal2 s 14370 56200 14426 57000 0 FreeSans 224 90 0 0 chany_top_in_0[4]
port 150 nsew signal input
flabel metal2 s 14738 56200 14794 57000 0 FreeSans 224 90 0 0 chany_top_in_0[5]
port 151 nsew signal input
flabel metal2 s 15106 56200 15162 57000 0 FreeSans 224 90 0 0 chany_top_in_0[6]
port 152 nsew signal input
flabel metal2 s 15474 56200 15530 57000 0 FreeSans 224 90 0 0 chany_top_in_0[7]
port 153 nsew signal input
flabel metal2 s 15842 56200 15898 57000 0 FreeSans 224 90 0 0 chany_top_in_0[8]
port 154 nsew signal input
flabel metal2 s 16210 56200 16266 57000 0 FreeSans 224 90 0 0 chany_top_in_0[9]
port 155 nsew signal input
flabel metal2 s 1858 56200 1914 57000 0 FreeSans 224 90 0 0 chany_top_out_0[0]
port 156 nsew signal tristate
flabel metal2 s 5538 56200 5594 57000 0 FreeSans 224 90 0 0 chany_top_out_0[10]
port 157 nsew signal tristate
flabel metal2 s 5906 56200 5962 57000 0 FreeSans 224 90 0 0 chany_top_out_0[11]
port 158 nsew signal tristate
flabel metal2 s 6274 56200 6330 57000 0 FreeSans 224 90 0 0 chany_top_out_0[12]
port 159 nsew signal tristate
flabel metal2 s 6642 56200 6698 57000 0 FreeSans 224 90 0 0 chany_top_out_0[13]
port 160 nsew signal tristate
flabel metal2 s 7010 56200 7066 57000 0 FreeSans 224 90 0 0 chany_top_out_0[14]
port 161 nsew signal tristate
flabel metal2 s 7378 56200 7434 57000 0 FreeSans 224 90 0 0 chany_top_out_0[15]
port 162 nsew signal tristate
flabel metal2 s 7746 56200 7802 57000 0 FreeSans 224 90 0 0 chany_top_out_0[16]
port 163 nsew signal tristate
flabel metal2 s 8114 56200 8170 57000 0 FreeSans 224 90 0 0 chany_top_out_0[17]
port 164 nsew signal tristate
flabel metal2 s 8482 56200 8538 57000 0 FreeSans 224 90 0 0 chany_top_out_0[18]
port 165 nsew signal tristate
flabel metal2 s 8850 56200 8906 57000 0 FreeSans 224 90 0 0 chany_top_out_0[19]
port 166 nsew signal tristate
flabel metal2 s 2226 56200 2282 57000 0 FreeSans 224 90 0 0 chany_top_out_0[1]
port 167 nsew signal tristate
flabel metal2 s 9218 56200 9274 57000 0 FreeSans 224 90 0 0 chany_top_out_0[20]
port 168 nsew signal tristate
flabel metal2 s 9586 56200 9642 57000 0 FreeSans 224 90 0 0 chany_top_out_0[21]
port 169 nsew signal tristate
flabel metal2 s 9954 56200 10010 57000 0 FreeSans 224 90 0 0 chany_top_out_0[22]
port 170 nsew signal tristate
flabel metal2 s 10322 56200 10378 57000 0 FreeSans 224 90 0 0 chany_top_out_0[23]
port 171 nsew signal tristate
flabel metal2 s 10690 56200 10746 57000 0 FreeSans 224 90 0 0 chany_top_out_0[24]
port 172 nsew signal tristate
flabel metal2 s 11058 56200 11114 57000 0 FreeSans 224 90 0 0 chany_top_out_0[25]
port 173 nsew signal tristate
flabel metal2 s 11426 56200 11482 57000 0 FreeSans 224 90 0 0 chany_top_out_0[26]
port 174 nsew signal tristate
flabel metal2 s 11794 56200 11850 57000 0 FreeSans 224 90 0 0 chany_top_out_0[27]
port 175 nsew signal tristate
flabel metal2 s 12162 56200 12218 57000 0 FreeSans 224 90 0 0 chany_top_out_0[28]
port 176 nsew signal tristate
flabel metal2 s 12530 56200 12586 57000 0 FreeSans 224 90 0 0 chany_top_out_0[29]
port 177 nsew signal tristate
flabel metal2 s 2594 56200 2650 57000 0 FreeSans 224 90 0 0 chany_top_out_0[2]
port 178 nsew signal tristate
flabel metal2 s 2962 56200 3018 57000 0 FreeSans 224 90 0 0 chany_top_out_0[3]
port 179 nsew signal tristate
flabel metal2 s 3330 56200 3386 57000 0 FreeSans 224 90 0 0 chany_top_out_0[4]
port 180 nsew signal tristate
flabel metal2 s 3698 56200 3754 57000 0 FreeSans 224 90 0 0 chany_top_out_0[5]
port 181 nsew signal tristate
flabel metal2 s 4066 56200 4122 57000 0 FreeSans 224 90 0 0 chany_top_out_0[6]
port 182 nsew signal tristate
flabel metal2 s 4434 56200 4490 57000 0 FreeSans 224 90 0 0 chany_top_out_0[7]
port 183 nsew signal tristate
flabel metal2 s 4802 56200 4858 57000 0 FreeSans 224 90 0 0 chany_top_out_0[8]
port 184 nsew signal tristate
flabel metal2 s 5170 56200 5226 57000 0 FreeSans 224 90 0 0 chany_top_out_0[9]
port 185 nsew signal tristate
flabel metal3 s 0 13744 800 13864 0 FreeSans 480 0 0 0 gfpga_pad_io_soc_dir[0]
port 186 nsew signal tristate
flabel metal3 s 0 16192 800 16312 0 FreeSans 480 0 0 0 gfpga_pad_io_soc_dir[1]
port 187 nsew signal tristate
flabel metal3 s 0 18640 800 18760 0 FreeSans 480 0 0 0 gfpga_pad_io_soc_dir[2]
port 188 nsew signal tristate
flabel metal3 s 0 21088 800 21208 0 FreeSans 480 0 0 0 gfpga_pad_io_soc_dir[3]
port 189 nsew signal tristate
flabel metal3 s 0 33328 800 33448 0 FreeSans 480 0 0 0 gfpga_pad_io_soc_in[0]
port 190 nsew signal input
flabel metal3 s 0 35776 800 35896 0 FreeSans 480 0 0 0 gfpga_pad_io_soc_in[1]
port 191 nsew signal input
flabel metal3 s 0 38224 800 38344 0 FreeSans 480 0 0 0 gfpga_pad_io_soc_in[2]
port 192 nsew signal input
flabel metal3 s 0 40672 800 40792 0 FreeSans 480 0 0 0 gfpga_pad_io_soc_in[3]
port 193 nsew signal input
flabel metal3 s 0 23536 800 23656 0 FreeSans 480 0 0 0 gfpga_pad_io_soc_out[0]
port 194 nsew signal tristate
flabel metal3 s 0 25984 800 26104 0 FreeSans 480 0 0 0 gfpga_pad_io_soc_out[1]
port 195 nsew signal tristate
flabel metal3 s 0 28432 800 28552 0 FreeSans 480 0 0 0 gfpga_pad_io_soc_out[2]
port 196 nsew signal tristate
flabel metal3 s 0 30880 800 31000 0 FreeSans 480 0 0 0 gfpga_pad_io_soc_out[3]
port 197 nsew signal tristate
flabel metal3 s 0 43120 800 43240 0 FreeSans 480 0 0 0 isol_n
port 198 nsew signal input
flabel metal2 s 23754 0 23810 800 0 FreeSans 224 90 0 0 prog_clk
port 199 nsew signal input
flabel metal2 s 24122 0 24178 800 0 FreeSans 224 90 0 0 prog_reset
port 200 nsew signal input
flabel metal2 s 24490 0 24546 800 0 FreeSans 224 90 0 0 reset
port 201 nsew signal input
flabel metal3 s 26200 50464 27000 50584 0 FreeSans 480 0 0 0 right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_
port 202 nsew signal input
flabel metal3 s 26200 51280 27000 51400 0 FreeSans 480 0 0 0 right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_
port 203 nsew signal input
flabel metal3 s 26200 52096 27000 52216 0 FreeSans 480 0 0 0 right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_
port 204 nsew signal input
flabel metal3 s 26200 52912 27000 53032 0 FreeSans 480 0 0 0 right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_
port 205 nsew signal input
flabel metal3 s 26200 53728 27000 53848 0 FreeSans 480 0 0 0 right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_4_
port 206 nsew signal input
flabel metal3 s 26200 54544 27000 54664 0 FreeSans 480 0 0 0 right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_5_
port 207 nsew signal input
flabel metal3 s 26200 55360 27000 55480 0 FreeSans 480 0 0 0 right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_6_
port 208 nsew signal input
flabel metal3 s 26200 56176 27000 56296 0 FreeSans 480 0 0 0 right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_7_
port 209 nsew signal input
flabel metal3 s 0 3952 800 4072 0 FreeSans 480 0 0 0 right_width_0_height_0_subtile_0__pin_inpad_0_
port 210 nsew signal tristate
flabel metal3 s 0 6400 800 6520 0 FreeSans 480 0 0 0 right_width_0_height_0_subtile_1__pin_inpad_0_
port 211 nsew signal tristate
flabel metal3 s 0 8848 800 8968 0 FreeSans 480 0 0 0 right_width_0_height_0_subtile_2__pin_inpad_0_
port 212 nsew signal tristate
flabel metal3 s 0 11296 800 11416 0 FreeSans 480 0 0 0 right_width_0_height_0_subtile_3__pin_inpad_0_
port 213 nsew signal tristate
flabel metal2 s 24858 0 24914 800 0 FreeSans 224 90 0 0 test_enable
port 214 nsew signal input
flabel metal3 s 0 45568 800 45688 0 FreeSans 480 0 0 0 top_left_grid_right_width_0_height_0_subtile_0__pin_inpad_0_
port 215 nsew signal input
flabel metal3 s 0 48016 800 48136 0 FreeSans 480 0 0 0 top_left_grid_right_width_0_height_0_subtile_1__pin_inpad_0_
port 216 nsew signal input
flabel metal3 s 0 50464 800 50584 0 FreeSans 480 0 0 0 top_left_grid_right_width_0_height_0_subtile_2__pin_inpad_0_
port 217 nsew signal input
flabel metal3 s 0 52912 800 53032 0 FreeSans 480 0 0 0 top_left_grid_right_width_0_height_0_subtile_3__pin_inpad_0_
port 218 nsew signal input
rlabel metal1 13478 54400 13478 54400 0 VGND
rlabel metal1 13478 53856 13478 53856 0 VPWR
rlabel metal1 5888 21454 5888 21454 0 cby_0__1_.cby_0__1_.ccff_tail
rlabel metal1 2070 27948 2070 27948 0 cby_0__1_.cby_0__1_.left_grid_right_width_0_height_0_subtile_0__pin_outpad_0_
rlabel metal1 4048 20570 4048 20570 0 cby_0__1_.cby_0__1_.left_grid_right_width_0_height_0_subtile_1__pin_outpad_0_
rlabel metal1 3082 20570 3082 20570 0 cby_0__1_.cby_0__1_.left_grid_right_width_0_height_0_subtile_2__pin_outpad_0_
rlabel metal1 1886 21556 1886 21556 0 cby_0__1_.cby_0__1_.left_grid_right_width_0_height_0_subtile_3__pin_outpad_0_
rlabel metal1 7728 23834 7728 23834 0 cby_0__1_.cby_0__1_.mem_right_ipin_0.ccff_tail
rlabel metal2 6808 17612 6808 17612 0 cby_0__1_.cby_0__1_.mem_right_ipin_0.mem_out\[0\]
rlabel metal1 9568 22066 9568 22066 0 cby_0__1_.cby_0__1_.mem_right_ipin_0.mem_out\[1\]
rlabel metal1 8970 20978 8970 20978 0 cby_0__1_.cby_0__1_.mem_right_ipin_0.mem_out\[2\]
rlabel metal2 8234 15878 8234 15878 0 cby_0__1_.cby_0__1_.mem_right_ipin_1.ccff_tail
rlabel metal2 11730 21862 11730 21862 0 cby_0__1_.cby_0__1_.mem_right_ipin_1.mem_out\[0\]
rlabel metal1 12144 18802 12144 18802 0 cby_0__1_.cby_0__1_.mem_right_ipin_1.mem_out\[1\]
rlabel metal1 10350 16626 10350 16626 0 cby_0__1_.cby_0__1_.mem_right_ipin_1.mem_out\[2\]
rlabel metal1 6026 18190 6026 18190 0 cby_0__1_.cby_0__1_.mem_right_ipin_2.ccff_tail
rlabel metal1 16767 12274 16767 12274 0 cby_0__1_.cby_0__1_.mem_right_ipin_2.mem_out\[0\]
rlabel metal1 11960 19278 11960 19278 0 cby_0__1_.cby_0__1_.mem_right_ipin_2.mem_out\[1\]
rlabel metal1 6141 17170 6141 17170 0 cby_0__1_.cby_0__1_.mem_right_ipin_2.mem_out\[2\]
rlabel metal1 12374 19244 12374 19244 0 cby_0__1_.cby_0__1_.mem_right_ipin_3.mem_out\[0\]
rlabel metal2 9890 18666 9890 18666 0 cby_0__1_.cby_0__1_.mem_right_ipin_3.mem_out\[1\]
rlabel metal1 7498 19686 7498 19686 0 cby_0__1_.cby_0__1_.mem_right_ipin_3.mem_out\[2\]
rlabel metal1 11960 19686 11960 19686 0 cby_0__1_.cby_0__1_.mux_right_ipin_0.sky130_fd_sc_hd__mux2_1_0_X
rlabel metal1 7176 21862 7176 21862 0 cby_0__1_.cby_0__1_.mux_right_ipin_0.sky130_fd_sc_hd__mux2_1_10_X
rlabel metal2 6486 24786 6486 24786 0 cby_0__1_.cby_0__1_.mux_right_ipin_0.sky130_fd_sc_hd__mux2_1_11_X
rlabel metal1 12926 18938 12926 18938 0 cby_0__1_.cby_0__1_.mux_right_ipin_0.sky130_fd_sc_hd__mux2_1_1_X
rlabel metal2 14306 19856 14306 19856 0 cby_0__1_.cby_0__1_.mux_right_ipin_0.sky130_fd_sc_hd__mux2_1_2_X
rlabel metal1 11914 20910 11914 20910 0 cby_0__1_.cby_0__1_.mux_right_ipin_0.sky130_fd_sc_hd__mux2_1_3_X
rlabel metal1 10074 19482 10074 19482 0 cby_0__1_.cby_0__1_.mux_right_ipin_0.sky130_fd_sc_hd__mux2_1_4_X
rlabel metal2 11270 20468 11270 20468 0 cby_0__1_.cby_0__1_.mux_right_ipin_0.sky130_fd_sc_hd__mux2_1_5_X
rlabel metal1 10396 20842 10396 20842 0 cby_0__1_.cby_0__1_.mux_right_ipin_0.sky130_fd_sc_hd__mux2_1_6_X
rlabel metal1 8602 21930 8602 21930 0 cby_0__1_.cby_0__1_.mux_right_ipin_0.sky130_fd_sc_hd__mux2_1_7_X
rlabel metal1 7820 21998 7820 21998 0 cby_0__1_.cby_0__1_.mux_right_ipin_0.sky130_fd_sc_hd__mux2_1_8_X
rlabel metal1 8050 24038 8050 24038 0 cby_0__1_.cby_0__1_.mux_right_ipin_0.sky130_fd_sc_hd__mux2_1_9_X
rlabel metal1 14352 12410 14352 12410 0 cby_0__1_.cby_0__1_.mux_right_ipin_1.sky130_fd_sc_hd__mux2_1_0_X
rlabel metal2 9154 16320 9154 16320 0 cby_0__1_.cby_0__1_.mux_right_ipin_1.sky130_fd_sc_hd__mux2_1_10_X
rlabel metal2 6440 16796 6440 16796 0 cby_0__1_.cby_0__1_.mux_right_ipin_1.sky130_fd_sc_hd__mux2_1_11_X
rlabel metal1 14260 14382 14260 14382 0 cby_0__1_.cby_0__1_.mux_right_ipin_1.sky130_fd_sc_hd__mux2_1_1_X
rlabel metal2 12558 20332 12558 20332 0 cby_0__1_.cby_0__1_.mux_right_ipin_1.sky130_fd_sc_hd__mux2_1_2_X
rlabel metal2 14030 18530 14030 18530 0 cby_0__1_.cby_0__1_.mux_right_ipin_1.sky130_fd_sc_hd__mux2_1_3_X
rlabel metal1 10626 16218 10626 16218 0 cby_0__1_.cby_0__1_.mux_right_ipin_1.sky130_fd_sc_hd__mux2_1_4_X
rlabel metal2 11086 15504 11086 15504 0 cby_0__1_.cby_0__1_.mux_right_ipin_1.sky130_fd_sc_hd__mux2_1_5_X
rlabel metal1 11270 18870 11270 18870 0 cby_0__1_.cby_0__1_.mux_right_ipin_1.sky130_fd_sc_hd__mux2_1_6_X
rlabel metal2 9614 16320 9614 16320 0 cby_0__1_.cby_0__1_.mux_right_ipin_1.sky130_fd_sc_hd__mux2_1_7_X
rlabel metal2 9338 16966 9338 16966 0 cby_0__1_.cby_0__1_.mux_right_ipin_1.sky130_fd_sc_hd__mux2_1_8_X
rlabel metal2 10350 16286 10350 16286 0 cby_0__1_.cby_0__1_.mux_right_ipin_1.sky130_fd_sc_hd__mux2_1_9_X
rlabel metal1 16330 12410 16330 12410 0 cby_0__1_.cby_0__1_.mux_right_ipin_2.sky130_fd_sc_hd__mux2_1_0_X
rlabel metal2 7130 18122 7130 18122 0 cby_0__1_.cby_0__1_.mux_right_ipin_2.sky130_fd_sc_hd__mux2_1_10_X
rlabel metal1 4784 18394 4784 18394 0 cby_0__1_.cby_0__1_.mux_right_ipin_2.sky130_fd_sc_hd__mux2_1_11_X
rlabel metal1 13110 12954 13110 12954 0 cby_0__1_.cby_0__1_.mux_right_ipin_2.sky130_fd_sc_hd__mux2_1_1_X
rlabel metal2 12742 20536 12742 20536 0 cby_0__1_.cby_0__1_.mux_right_ipin_2.sky130_fd_sc_hd__mux2_1_2_X
rlabel metal2 12098 18326 12098 18326 0 cby_0__1_.cby_0__1_.mux_right_ipin_2.sky130_fd_sc_hd__mux2_1_3_X
rlabel metal1 10028 19822 10028 19822 0 cby_0__1_.cby_0__1_.mux_right_ipin_2.sky130_fd_sc_hd__mux2_1_4_X
rlabel metal1 7866 17068 7866 17068 0 cby_0__1_.cby_0__1_.mux_right_ipin_2.sky130_fd_sc_hd__mux2_1_5_X
rlabel metal1 8510 17306 8510 17306 0 cby_0__1_.cby_0__1_.mux_right_ipin_2.sky130_fd_sc_hd__mux2_1_6_X
rlabel metal2 7590 18836 7590 18836 0 cby_0__1_.cby_0__1_.mux_right_ipin_2.sky130_fd_sc_hd__mux2_1_7_X
rlabel metal1 8280 17646 8280 17646 0 cby_0__1_.cby_0__1_.mux_right_ipin_2.sky130_fd_sc_hd__mux2_1_8_X
rlabel metal1 5750 18122 5750 18122 0 cby_0__1_.cby_0__1_.mux_right_ipin_2.sky130_fd_sc_hd__mux2_1_9_X
rlabel metal1 11454 18258 11454 18258 0 cby_0__1_.cby_0__1_.mux_right_ipin_3.sky130_fd_sc_hd__mux2_1_0_X
rlabel metal1 6118 21658 6118 21658 0 cby_0__1_.cby_0__1_.mux_right_ipin_3.sky130_fd_sc_hd__mux2_1_10_X
rlabel metal1 4278 21658 4278 21658 0 cby_0__1_.cby_0__1_.mux_right_ipin_3.sky130_fd_sc_hd__mux2_1_11_X
rlabel metal1 11822 18394 11822 18394 0 cby_0__1_.cby_0__1_.mux_right_ipin_3.sky130_fd_sc_hd__mux2_1_1_X
rlabel metal2 12374 20468 12374 20468 0 cby_0__1_.cby_0__1_.mux_right_ipin_3.sky130_fd_sc_hd__mux2_1_2_X
rlabel metal1 11316 24582 11316 24582 0 cby_0__1_.cby_0__1_.mux_right_ipin_3.sky130_fd_sc_hd__mux2_1_3_X
rlabel metal1 9568 17306 9568 17306 0 cby_0__1_.cby_0__1_.mux_right_ipin_3.sky130_fd_sc_hd__mux2_1_4_X
rlabel metal1 10396 18394 10396 18394 0 cby_0__1_.cby_0__1_.mux_right_ipin_3.sky130_fd_sc_hd__mux2_1_5_X
rlabel metal1 8372 19822 8372 19822 0 cby_0__1_.cby_0__1_.mux_right_ipin_3.sky130_fd_sc_hd__mux2_1_6_X
rlabel metal1 7682 20570 7682 20570 0 cby_0__1_.cby_0__1_.mux_right_ipin_3.sky130_fd_sc_hd__mux2_1_7_X
rlabel metal1 7130 21658 7130 21658 0 cby_0__1_.cby_0__1_.mux_right_ipin_3.sky130_fd_sc_hd__mux2_1_8_X
rlabel metal1 7406 20026 7406 20026 0 cby_0__1_.cby_0__1_.mux_right_ipin_3.sky130_fd_sc_hd__mux2_1_9_X
rlabel metal2 4830 24820 4830 24820 0 cby_0__1_.grid_io_left_left_0__1_.logical_tile_io_mode_io__0.ccff_tail
rlabel metal2 2254 27200 2254 27200 0 cby_0__1_.grid_io_left_left_0__1_.logical_tile_io_mode_io__0.gfpga_pad_io_soc_dir
rlabel metal1 3611 29274 3611 29274 0 cby_0__1_.grid_io_left_left_0__1_.logical_tile_io_mode_io__0.logical_tile_io_mode_physical__iopad_0.io_0_.SOC_DIR_N
rlabel metal1 5060 24718 5060 24718 0 cby_0__1_.grid_io_left_left_0__1_.logical_tile_io_mode_io__1.ccff_tail
rlabel metal1 1932 24718 1932 24718 0 cby_0__1_.grid_io_left_left_0__1_.logical_tile_io_mode_io__1.gfpga_pad_io_soc_dir
rlabel metal1 4025 27370 4025 27370 0 cby_0__1_.grid_io_left_left_0__1_.logical_tile_io_mode_io__1.logical_tile_io_mode_physical__iopad_0.io_0_.SOC_DIR_N
rlabel metal2 5934 19788 5934 19788 0 cby_0__1_.grid_io_left_left_0__1_.logical_tile_io_mode_io__2.ccff_tail
rlabel metal1 1932 23018 1932 23018 0 cby_0__1_.grid_io_left_left_0__1_.logical_tile_io_mode_io__2.gfpga_pad_io_soc_dir
rlabel via1 3519 26010 3519 26010 0 cby_0__1_.grid_io_left_left_0__1_.logical_tile_io_mode_io__2.logical_tile_io_mode_physical__iopad_0.io_0_.SOC_DIR_N
rlabel metal1 2300 17238 2300 17238 0 cby_0__1_.grid_io_left_left_0__1_.logical_tile_io_mode_io__3.gfpga_pad_io_soc_dir
rlabel metal1 3749 23834 3749 23834 0 cby_0__1_.grid_io_left_left_0__1_.logical_tile_io_mode_io__3.logical_tile_io_mode_physical__iopad_0.io_0_.SOC_DIR_N
rlabel metal3 1740 55420 1740 55420 0 ccff_head
rlabel metal1 2484 3910 2484 3910 0 ccff_head_0
rlabel metal1 19274 6188 19274 6188 0 ccff_tail
rlabel metal1 1794 49266 1794 49266 0 ccff_tail_0
rlabel metal2 22586 25415 22586 25415 0 chanx_right_in[0]
rlabel via2 25346 34187 25346 34187 0 chanx_right_in[10]
rlabel metal2 24702 35513 24702 35513 0 chanx_right_in[11]
rlabel metal2 24886 35921 24886 35921 0 chanx_right_in[12]
rlabel metal1 24380 38250 24380 38250 0 chanx_right_in[13]
rlabel metal1 22402 36788 22402 36788 0 chanx_right_in[14]
rlabel metal2 25346 39695 25346 39695 0 chanx_right_in[15]
rlabel metal2 24058 39797 24058 39797 0 chanx_right_in[16]
rlabel via2 24173 40052 24173 40052 0 chanx_right_in[17]
rlabel metal3 25584 40732 25584 40732 0 chanx_right_in[18]
rlabel metal1 21482 42126 21482 42126 0 chanx_right_in[19]
rlabel metal1 21482 25908 21482 25908 0 chanx_right_in[1]
rlabel metal2 23230 42517 23230 42517 0 chanx_right_in[20]
rlabel metal1 24564 44302 24564 44302 0 chanx_right_in[21]
rlabel metal2 24518 44693 24518 44693 0 chanx_right_in[22]
rlabel metal1 24932 46954 24932 46954 0 chanx_right_in[23]
rlabel metal2 24426 46359 24426 46359 0 chanx_right_in[24]
rlabel metal1 25024 47974 25024 47974 0 chanx_right_in[25]
rlabel via1 25530 47617 25530 47617 0 chanx_right_in[26]
rlabel metal2 24518 48909 24518 48909 0 chanx_right_in[27]
rlabel metal2 25346 49045 25346 49045 0 chanx_right_in[28]
rlabel metal2 25346 49997 25346 49997 0 chanx_right_in[29]
rlabel metal2 24150 28407 24150 28407 0 chanx_right_in[2]
rlabel metal2 25254 28339 25254 28339 0 chanx_right_in[3]
rlabel via2 25530 29291 25530 29291 0 chanx_right_in[4]
rlabel metal2 25346 29869 25346 29869 0 chanx_right_in[5]
rlabel metal2 25346 31127 25346 31127 0 chanx_right_in[6]
rlabel via2 25346 31773 25346 31773 0 chanx_right_in[7]
rlabel metal2 25346 32725 25346 32725 0 chanx_right_in[8]
rlabel metal1 25392 32402 25392 32402 0 chanx_right_in[9]
rlabel metal3 25676 9724 25676 9724 0 chanx_right_out[10]
rlabel metal2 24702 10013 24702 10013 0 chanx_right_out[11]
rlabel metal2 24794 10965 24794 10965 0 chanx_right_out[12]
rlabel metal2 25162 11985 25162 11985 0 chanx_right_out[13]
rlabel metal3 25676 12988 25676 12988 0 chanx_right_out[14]
rlabel metal2 24794 13277 24794 13277 0 chanx_right_out[15]
rlabel metal2 25162 14297 25162 14297 0 chanx_right_out[16]
rlabel metal3 25676 15436 25676 15436 0 chanx_right_out[17]
rlabel metal2 24702 15589 24702 15589 0 chanx_right_out[18]
rlabel metal3 25584 17068 25584 17068 0 chanx_right_out[19]
rlabel metal3 24020 2380 24020 2380 0 chanx_right_out[1]
rlabel metal1 23368 18190 23368 18190 0 chanx_right_out[20]
rlabel metal2 24702 17901 24702 17901 0 chanx_right_out[21]
rlabel metal2 24794 18853 24794 18853 0 chanx_right_out[22]
rlabel metal1 24426 19890 24426 19890 0 chanx_right_out[23]
rlabel metal1 23368 20502 23368 20502 0 chanx_right_out[24]
rlabel metal1 24380 20978 24380 20978 0 chanx_right_out[25]
rlabel metal1 23874 20366 23874 20366 0 chanx_right_out[26]
rlabel metal2 23874 23341 23874 23341 0 chanx_right_out[27]
rlabel metal1 24380 24242 24380 24242 0 chanx_right_out[28]
rlabel metal2 25162 25517 25162 25517 0 chanx_right_out[29]
rlabel metal3 24572 3196 24572 3196 0 chanx_right_out[2]
rlabel metal1 19182 5270 19182 5270 0 chanx_right_out[3]
rlabel metal2 23368 4828 23368 4828 0 chanx_right_out[4]
rlabel metal2 24794 5389 24794 5389 0 chanx_right_out[5]
rlabel metal3 26090 6460 26090 6460 0 chanx_right_out[6]
rlabel metal3 25584 7276 25584 7276 0 chanx_right_out[7]
rlabel metal2 25162 7769 25162 7769 0 chanx_right_out[8]
rlabel metal2 25162 8721 25162 8721 0 chanx_right_out[9]
rlabel metal1 1840 3502 1840 3502 0 chany_bottom_in[0]
rlabel metal1 5198 3026 5198 3026 0 chany_bottom_in[10]
rlabel metal1 5934 2346 5934 2346 0 chany_bottom_in[11]
rlabel metal2 6118 2132 6118 2132 0 chany_bottom_in[12]
rlabel metal2 6486 1792 6486 1792 0 chany_bottom_in[13]
rlabel metal2 6854 1894 6854 1894 0 chany_bottom_in[14]
rlabel metal2 7222 1588 7222 1588 0 chany_bottom_in[15]
rlabel metal1 7636 2414 7636 2414 0 chany_bottom_in[16]
rlabel metal1 7820 3366 7820 3366 0 chany_bottom_in[17]
rlabel metal1 7912 3026 7912 3026 0 chany_bottom_in[18]
rlabel metal2 8694 2064 8694 2064 0 chany_bottom_in[19]
rlabel metal1 1978 3026 1978 3026 0 chany_bottom_in[1]
rlabel metal2 9062 1860 9062 1860 0 chany_bottom_in[20]
rlabel metal1 9292 3502 9292 3502 0 chany_bottom_in[21]
rlabel metal1 9844 3502 9844 3502 0 chany_bottom_in[22]
rlabel metal1 9890 2414 9890 2414 0 chany_bottom_in[23]
rlabel metal1 10442 2958 10442 2958 0 chany_bottom_in[24]
rlabel metal1 10948 3502 10948 3502 0 chany_bottom_in[25]
rlabel metal1 11500 3026 11500 3026 0 chany_bottom_in[26]
rlabel metal1 11684 4046 11684 4046 0 chany_bottom_in[27]
rlabel metal1 11914 2448 11914 2448 0 chany_bottom_in[28]
rlabel metal1 10350 2380 10350 2380 0 chany_bottom_in[29]
rlabel metal1 2024 2414 2024 2414 0 chany_bottom_in[2]
rlabel metal1 2668 3026 2668 3026 0 chany_bottom_in[3]
rlabel metal1 3312 2958 3312 2958 0 chany_bottom_in[4]
rlabel metal1 2990 2414 2990 2414 0 chany_bottom_in[5]
rlabel metal1 3588 2346 3588 2346 0 chany_bottom_in[6]
rlabel metal1 4140 2414 4140 2414 0 chany_bottom_in[7]
rlabel metal1 4692 2414 4692 2414 0 chany_bottom_in[8]
rlabel metal1 4876 3366 4876 3366 0 chany_bottom_in[9]
rlabel metal2 12742 2166 12742 2166 0 chany_bottom_out[0]
rlabel metal2 16422 2404 16422 2404 0 chany_bottom_out[10]
rlabel metal2 16790 1554 16790 1554 0 chany_bottom_out[11]
rlabel metal2 17158 1826 17158 1826 0 chany_bottom_out[12]
rlabel metal2 17526 2404 17526 2404 0 chany_bottom_out[13]
rlabel metal2 17894 1231 17894 1231 0 chany_bottom_out[14]
rlabel metal2 18262 959 18262 959 0 chany_bottom_out[15]
rlabel metal2 18630 1792 18630 1792 0 chany_bottom_out[16]
rlabel metal2 18998 2098 18998 2098 0 chany_bottom_out[17]
rlabel metal2 19366 2948 19366 2948 0 chany_bottom_out[18]
rlabel metal2 19734 1826 19734 1826 0 chany_bottom_out[19]
rlabel metal2 13110 823 13110 823 0 chany_bottom_out[1]
rlabel metal2 20102 2404 20102 2404 0 chany_bottom_out[20]
rlabel metal2 20470 3254 20470 3254 0 chany_bottom_out[21]
rlabel metal2 20838 1792 20838 1792 0 chany_bottom_out[22]
rlabel metal2 21206 2370 21206 2370 0 chany_bottom_out[23]
rlabel metal2 21574 3254 21574 3254 0 chany_bottom_out[24]
rlabel metal2 21942 3492 21942 3492 0 chany_bottom_out[25]
rlabel metal1 22448 7310 22448 7310 0 chany_bottom_out[26]
rlabel metal2 22678 1894 22678 1894 0 chany_bottom_out[27]
rlabel metal2 23046 1639 23046 1639 0 chany_bottom_out[28]
rlabel metal2 23414 1860 23414 1860 0 chany_bottom_out[29]
rlabel metal2 13478 2404 13478 2404 0 chany_bottom_out[2]
rlabel metal2 13846 1554 13846 1554 0 chany_bottom_out[3]
rlabel metal2 14214 1860 14214 1860 0 chany_bottom_out[4]
rlabel metal2 14582 1622 14582 1622 0 chany_bottom_out[5]
rlabel metal2 14950 2166 14950 2166 0 chany_bottom_out[6]
rlabel metal2 15318 1622 15318 1622 0 chany_bottom_out[7]
rlabel metal2 15686 1860 15686 1860 0 chany_bottom_out[8]
rlabel metal2 16054 2166 16054 2166 0 chany_bottom_out[9]
rlabel metal1 11914 54196 11914 54196 0 chany_top_in_0[0]
rlabel metal1 16652 53550 16652 53550 0 chany_top_in_0[10]
rlabel metal1 17296 54162 17296 54162 0 chany_top_in_0[11]
rlabel metal1 17480 53550 17480 53550 0 chany_top_in_0[12]
rlabel metal1 18078 54230 18078 54230 0 chany_top_in_0[13]
rlabel metal2 18262 56236 18262 56236 0 chany_top_in_0[14]
rlabel metal1 19458 54128 19458 54128 0 chany_top_in_0[15]
rlabel metal1 18952 53074 18952 53074 0 chany_top_in_0[16]
rlabel metal1 19320 53550 19320 53550 0 chany_top_in_0[17]
rlabel metal1 19872 54162 19872 54162 0 chany_top_in_0[18]
rlabel metal1 20102 53550 20102 53550 0 chany_top_in_0[19]
rlabel metal2 13294 55711 13294 55711 0 chany_top_in_0[1]
rlabel metal1 20424 53074 20424 53074 0 chany_top_in_0[20]
rlabel metal2 20654 55711 20654 55711 0 chany_top_in_0[21]
rlabel metal1 21068 53550 21068 53550 0 chany_top_in_0[22]
rlabel metal1 21712 54162 21712 54162 0 chany_top_in_0[23]
rlabel metal1 21896 53550 21896 53550 0 chany_top_in_0[24]
rlabel metal1 22218 53210 22218 53210 0 chany_top_in_0[25]
rlabel metal1 22632 54162 22632 54162 0 chany_top_in_0[26]
rlabel metal1 23092 53550 23092 53550 0 chany_top_in_0[27]
rlabel metal2 23230 55711 23230 55711 0 chany_top_in_0[28]
rlabel metal2 23598 55711 23598 55711 0 chany_top_in_0[29]
rlabel metal1 13754 53142 13754 53142 0 chany_top_in_0[2]
rlabel metal1 14168 53550 14168 53550 0 chany_top_in_0[3]
rlabel metal1 14536 53074 14536 53074 0 chany_top_in_0[4]
rlabel metal1 14674 54298 14674 54298 0 chany_top_in_0[5]
rlabel metal1 15410 54162 15410 54162 0 chany_top_in_0[6]
rlabel metal1 15594 53550 15594 53550 0 chany_top_in_0[7]
rlabel metal1 16008 53074 16008 53074 0 chany_top_in_0[8]
rlabel metal1 16721 54162 16721 54162 0 chany_top_in_0[9]
rlabel metal1 2714 52598 2714 52598 0 chany_top_out_0[0]
rlabel metal1 5566 53652 5566 53652 0 chany_top_out_0[10]
rlabel metal1 4600 54094 4600 54094 0 chany_top_out_0[11]
rlabel metal1 6072 53142 6072 53142 0 chany_top_out_0[12]
rlabel metal1 6624 52530 6624 52530 0 chany_top_out_0[13]
rlabel metal1 7314 51442 7314 51442 0 chany_top_out_0[14]
rlabel metal1 6992 53618 6992 53618 0 chany_top_out_0[15]
rlabel metal2 7774 54376 7774 54376 0 chany_top_out_0[16]
rlabel metal2 7958 56236 7958 56236 0 chany_top_out_0[17]
rlabel metal2 8510 54070 8510 54070 0 chany_top_out_0[18]
rlabel metal1 8648 53618 8648 53618 0 chany_top_out_0[19]
rlabel metal1 2852 52666 2852 52666 0 chany_top_out_0[1]
rlabel metal1 9200 53142 9200 53142 0 chany_top_out_0[20]
rlabel metal2 9660 53550 9660 53550 0 chany_top_out_0[21]
rlabel metal1 9982 54264 9982 54264 0 chany_top_out_0[22]
rlabel metal2 10350 55711 10350 55711 0 chany_top_out_0[23]
rlabel metal1 10994 52530 10994 52530 0 chany_top_out_0[24]
rlabel metal2 11086 54920 11086 54920 0 chany_top_out_0[25]
rlabel metal1 11224 54230 11224 54230 0 chany_top_out_0[26]
rlabel metal1 12098 53006 12098 53006 0 chany_top_out_0[27]
rlabel metal1 12466 53618 12466 53618 0 chany_top_out_0[28]
rlabel metal1 12696 54094 12696 54094 0 chany_top_out_0[29]
rlabel metal2 2714 52972 2714 52972 0 chany_top_out_0[2]
rlabel metal2 2990 55711 2990 55711 0 chany_top_out_0[3]
rlabel metal2 3358 54070 3358 54070 0 chany_top_out_0[4]
rlabel metal1 3496 52530 3496 52530 0 chany_top_out_0[5]
rlabel metal2 4186 52972 4186 52972 0 chany_top_out_0[6]
rlabel metal1 4232 53142 4232 53142 0 chany_top_out_0[7]
rlabel metal2 4830 55711 4830 55711 0 chany_top_out_0[8]
rlabel metal1 5474 53210 5474 53210 0 chany_top_out_0[9]
rlabel metal1 20378 43282 20378 43282 0 clknet_0_prog_clk
rlabel metal1 5428 16626 5428 16626 0 clknet_4_0_0_prog_clk
rlabel metal1 6302 38386 6302 38386 0 clknet_4_10_0_prog_clk
rlabel metal1 13110 44404 13110 44404 0 clknet_4_11_0_prog_clk
rlabel metal1 16882 38964 16882 38964 0 clknet_4_12_0_prog_clk
rlabel metal1 23460 33422 23460 33422 0 clknet_4_13_0_prog_clk
rlabel metal2 16882 44642 16882 44642 0 clknet_4_14_0_prog_clk
rlabel metal1 18262 45322 18262 45322 0 clknet_4_15_0_prog_clk
rlabel metal1 8924 18802 8924 18802 0 clknet_4_1_0_prog_clk
rlabel metal1 4094 22066 4094 22066 0 clknet_4_2_0_prog_clk
rlabel metal2 9246 26656 9246 26656 0 clknet_4_3_0_prog_clk
rlabel metal1 17986 11764 17986 11764 0 clknet_4_4_0_prog_clk
rlabel metal1 20286 12274 20286 12274 0 clknet_4_5_0_prog_clk
rlabel metal1 14076 20910 14076 20910 0 clknet_4_6_0_prog_clk
rlabel metal1 20976 21998 20976 21998 0 clknet_4_7_0_prog_clk
rlabel metal1 7682 32436 7682 32436 0 clknet_4_8_0_prog_clk
rlabel metal1 13892 33490 13892 33490 0 clknet_4_9_0_prog_clk
rlabel metal3 1004 13804 1004 13804 0 gfpga_pad_io_soc_dir[0]
rlabel metal3 1004 16252 1004 16252 0 gfpga_pad_io_soc_dir[1]
rlabel metal3 1004 18700 1004 18700 0 gfpga_pad_io_soc_dir[2]
rlabel metal3 1004 21148 1004 21148 0 gfpga_pad_io_soc_dir[3]
rlabel metal1 1564 33490 1564 33490 0 gfpga_pad_io_soc_in[0]
rlabel metal1 1932 36142 1932 36142 0 gfpga_pad_io_soc_in[1]
rlabel metal1 1564 38318 1564 38318 0 gfpga_pad_io_soc_in[2]
rlabel metal1 1564 41106 1564 41106 0 gfpga_pad_io_soc_in[3]
rlabel metal3 1786 23596 1786 23596 0 gfpga_pad_io_soc_out[0]
rlabel metal1 2990 23222 2990 23222 0 gfpga_pad_io_soc_out[1]
rlabel metal2 2898 26605 2898 26605 0 gfpga_pad_io_soc_out[2]
rlabel metal2 2806 29461 2806 29461 0 gfpga_pad_io_soc_out[3]
rlabel metal1 1518 43282 1518 43282 0 isol_n
rlabel metal1 2852 52870 2852 52870 0 net1
rlabel metal1 19918 38828 19918 38828 0 net10
rlabel metal1 18538 41480 18538 41480 0 net100
rlabel metal1 20056 43826 20056 43826 0 net101
rlabel metal1 17572 41582 17572 41582 0 net102
rlabel metal2 22034 44268 22034 44268 0 net103
rlabel metal3 23805 53244 23805 53244 0 net104
rlabel metal1 23782 53958 23782 53958 0 net105
rlabel metal3 22517 52972 22517 52972 0 net106
rlabel metal1 18124 6290 18124 6290 0 net107
rlabel metal1 1794 49130 1794 49130 0 net108
rlabel metal1 22586 9690 22586 9690 0 net109
rlabel metal1 20746 41650 20746 41650 0 net11
rlabel metal1 23920 9554 23920 9554 0 net110
rlabel metal2 23966 12750 23966 12750 0 net111
rlabel metal1 23368 11730 23368 11730 0 net112
rlabel metal1 22678 13362 22678 13362 0 net113
rlabel metal1 23690 12818 23690 12818 0 net114
rlabel metal1 23920 13906 23920 13906 0 net115
rlabel metal2 22770 17612 22770 17612 0 net116
rlabel metal1 24564 19686 24564 19686 0 net117
rlabel metal1 24472 21862 24472 21862 0 net118
rlabel metal1 22770 5882 22770 5882 0 net119
rlabel metal1 21022 41106 21022 41106 0 net12
rlabel metal1 23000 18258 23000 18258 0 net120
rlabel metal2 23966 21148 23966 21148 0 net121
rlabel metal1 24288 18258 24288 18258 0 net122
rlabel metal1 24104 19822 24104 19822 0 net123
rlabel metal2 22218 25228 22218 25228 0 net124
rlabel metal1 24058 20910 24058 20910 0 net125
rlabel metal1 24564 20434 24564 20434 0 net126
rlabel metal1 22862 23052 22862 23052 0 net127
rlabel metal1 22862 24140 22862 24140 0 net128
rlabel metal1 24380 22746 24380 22746 0 net129
rlabel metal1 18952 41990 18952 41990 0 net13
rlabel metal1 23598 4794 23598 4794 0 net130
rlabel metal2 17802 4964 17802 4964 0 net131
rlabel metal1 23230 7854 23230 7854 0 net132
rlabel metal2 23966 7004 23966 7004 0 net133
rlabel metal1 23138 6766 23138 6766 0 net134
rlabel metal1 23736 6290 23736 6290 0 net135
rlabel metal1 20286 7276 20286 7276 0 net136
rlabel metal1 23690 8466 23690 8466 0 net137
rlabel metal1 13110 3502 13110 3502 0 net138
rlabel metal1 16790 4114 16790 4114 0 net139
rlabel metal1 17204 25330 17204 25330 0 net14
rlabel metal1 19458 2482 19458 2482 0 net140
rlabel metal1 18308 3026 18308 3026 0 net141
rlabel metal1 19090 4114 19090 4114 0 net142
rlabel metal1 18538 3502 18538 3502 0 net143
rlabel metal1 19734 2618 19734 2618 0 net144
rlabel metal1 19090 4590 19090 4590 0 net145
rlabel metal1 20240 3638 20240 3638 0 net146
rlabel metal1 19274 5202 19274 5202 0 net147
rlabel metal1 21160 8330 21160 8330 0 net148
rlabel metal2 12650 4284 12650 4284 0 net149
rlabel metal1 19274 32538 19274 32538 0 net15
rlabel metal1 21022 4114 21022 4114 0 net150
rlabel metal1 20516 13226 20516 13226 0 net151
rlabel metal1 22172 12614 22172 12614 0 net152
rlabel metal1 23368 4114 23368 4114 0 net153
rlabel metal1 21528 5678 21528 5678 0 net154
rlabel metal1 21712 11254 21712 11254 0 net155
rlabel metal1 22126 7412 22126 7412 0 net156
rlabel metal1 20378 7718 20378 7718 0 net157
rlabel metal1 20470 6630 20470 6630 0 net158
rlabel metal1 18676 7242 18676 7242 0 net159
rlabel metal1 21206 31926 21206 31926 0 net16
rlabel metal2 13616 13158 13616 13158 0 net160
rlabel metal1 12374 10506 12374 10506 0 net161
rlabel metal1 14398 12070 14398 12070 0 net162
rlabel metal1 14628 13838 14628 13838 0 net163
rlabel metal2 15134 3842 15134 3842 0 net164
rlabel metal2 16974 6154 16974 6154 0 net165
rlabel metal1 16836 3026 16836 3026 0 net166
rlabel metal1 16606 3502 16606 3502 0 net167
rlabel metal1 2898 49810 2898 49810 0 net168
rlabel metal1 3358 53550 3358 53550 0 net169
rlabel metal1 16468 35530 16468 35530 0 net17
rlabel metal1 3312 54162 3312 54162 0 net170
rlabel metal1 5658 53074 5658 53074 0 net171
rlabel metal1 5566 52462 5566 52462 0 net172
rlabel metal2 7176 47668 7176 47668 0 net173
rlabel metal1 6210 53550 6210 53550 0 net174
rlabel metal2 7222 51761 7222 51761 0 net175
rlabel metal1 6670 43350 6670 43350 0 net176
rlabel metal1 7636 51986 7636 51986 0 net177
rlabel metal1 8234 53550 8234 53550 0 net178
rlabel metal1 3496 50286 3496 50286 0 net179
rlabel metal1 12834 37094 12834 37094 0 net18
rlabel metal1 8786 53074 8786 53074 0 net180
rlabel metal1 10580 45050 10580 45050 0 net181
rlabel metal1 8832 54094 8832 54094 0 net182
rlabel metal1 9614 49878 9614 49878 0 net183
rlabel metal1 10212 50966 10212 50966 0 net184
rlabel metal1 10396 53550 10396 53550 0 net185
rlabel metal1 10120 51578 10120 51578 0 net186
rlabel metal1 11822 52122 11822 52122 0 net187
rlabel metal2 12650 53108 12650 53108 0 net188
rlabel metal2 12374 53142 12374 53142 0 net189
rlabel metal2 23690 38233 23690 38233 0 net19
rlabel metal2 4186 46342 4186 46342 0 net190
rlabel metal1 2254 51340 2254 51340 0 net191
rlabel metal1 3772 51986 3772 51986 0 net192
rlabel metal1 3542 52462 3542 52462 0 net193
rlabel metal2 4370 46614 4370 46614 0 net194
rlabel metal1 2990 53040 2990 53040 0 net195
rlabel metal1 4922 51986 4922 51986 0 net196
rlabel metal1 6118 51374 6118 51374 0 net197
rlabel metal1 2070 16966 2070 16966 0 net198
rlabel metal1 2024 16558 2024 16558 0 net199
rlabel metal1 2208 3978 2208 3978 0 net2
rlabel metal1 21344 34646 21344 34646 0 net20
rlabel metal2 1794 20298 1794 20298 0 net200
rlabel metal1 1840 20910 1840 20910 0 net201
rlabel metal2 25346 1989 25346 1989 0 net202
rlabel metal2 17710 21216 17710 21216 0 net203
rlabel metal2 12374 27438 12374 27438 0 net204
rlabel metal2 22402 34272 22402 34272 0 net205
rlabel metal1 24978 23120 24978 23120 0 net206
rlabel metal2 15410 38080 15410 38080 0 net207
rlabel metal2 15778 24276 15778 24276 0 net208
rlabel metal1 21390 28526 21390 28526 0 net209
rlabel metal1 17434 41650 17434 41650 0 net21
rlabel metal1 17020 36074 17020 36074 0 net210
rlabel metal1 17986 36890 17986 36890 0 net211
rlabel metal1 16744 37978 16744 37978 0 net212
rlabel metal1 14582 38386 14582 38386 0 net213
rlabel metal1 13846 36890 13846 36890 0 net214
rlabel metal1 23368 39338 23368 39338 0 net215
rlabel metal2 12466 32062 12466 32062 0 net216
rlabel metal1 11270 30226 11270 30226 0 net217
rlabel metal1 11454 26010 11454 26010 0 net218
rlabel metal2 9522 27200 9522 27200 0 net219
rlabel metal1 17526 43418 17526 43418 0 net22
rlabel metal1 7360 25262 7360 25262 0 net220
rlabel metal1 8924 24242 8924 24242 0 net221
rlabel metal2 11730 23188 11730 23188 0 net222
rlabel metal1 12880 21658 12880 21658 0 net223
rlabel metal2 7498 9214 7498 9214 0 net224
rlabel metal2 17618 11968 17618 11968 0 net225
rlabel metal2 20930 34068 20930 34068 0 net226
rlabel metal1 16928 12886 16928 12886 0 net227
rlabel metal1 18722 14450 18722 14450 0 net228
rlabel metal2 21298 15810 21298 15810 0 net229
rlabel metal1 18446 42330 18446 42330 0 net23
rlabel metal1 22816 16082 22816 16082 0 net230
rlabel metal2 19550 16320 19550 16320 0 net231
rlabel metal1 21942 12886 21942 12886 0 net232
rlabel metal2 19550 10880 19550 10880 0 net233
rlabel metal1 20884 13906 20884 13906 0 net234
rlabel metal1 22540 35802 22540 35802 0 net235
rlabel metal1 21942 41242 21942 41242 0 net236
rlabel metal1 9752 37162 9752 37162 0 net237
rlabel metal1 8096 31314 8096 31314 0 net238
rlabel metal1 7360 32538 7360 32538 0 net239
rlabel metal1 21114 41038 21114 41038 0 net24
rlabel metal1 13708 42194 13708 42194 0 net240
rlabel metal2 9798 33150 9798 33150 0 net241
rlabel metal2 5566 32980 5566 32980 0 net242
rlabel metal1 8970 39066 8970 39066 0 net243
rlabel metal2 11730 38454 11730 38454 0 net244
rlabel metal1 10442 38318 10442 38318 0 net245
rlabel metal1 15088 36074 15088 36074 0 net246
rlabel metal1 10028 32334 10028 32334 0 net247
rlabel metal1 10304 24786 10304 24786 0 net248
rlabel metal1 11546 20434 11546 20434 0 net249
rlabel metal1 13386 30566 13386 30566 0 net25
rlabel metal1 8924 17714 8924 17714 0 net250
rlabel metal2 9614 23392 9614 23392 0 net251
rlabel metal1 16836 21522 16836 21522 0 net252
rlabel metal1 12052 25194 12052 25194 0 net253
rlabel metal2 19826 26622 19826 26622 0 net254
rlabel metal1 22908 25874 22908 25874 0 net255
rlabel metal1 17848 29546 17848 29546 0 net256
rlabel metal1 17940 46002 17940 46002 0 net257
rlabel metal2 6854 38318 6854 38318 0 net258
rlabel metal1 15863 27642 15863 27642 0 net259
rlabel metal1 17434 32402 17434 32402 0 net26
rlabel metal2 18630 16830 18630 16830 0 net260
rlabel metal2 20010 18088 20010 18088 0 net261
rlabel metal1 8786 40086 8786 40086 0 net262
rlabel metal2 15042 43112 15042 43112 0 net263
rlabel metal2 12834 44030 12834 44030 0 net264
rlabel metal1 20976 21658 20976 21658 0 net265
rlabel metal1 20976 17306 20976 17306 0 net266
rlabel metal1 15180 12750 15180 12750 0 net267
rlabel metal2 9982 30124 9982 30124 0 net268
rlabel metal1 17848 17850 17848 17850 0 net269
rlabel metal2 21114 28243 21114 28243 0 net27
rlabel metal1 18584 11662 18584 11662 0 net270
rlabel metal2 12098 12444 12098 12444 0 net271
rlabel metal2 14122 38624 14122 38624 0 net272
rlabel metal1 15962 31450 15962 31450 0 net273
rlabel metal1 5750 39066 5750 39066 0 net274
rlabel metal1 14352 39950 14352 39950 0 net275
rlabel metal1 19688 44506 19688 44506 0 net276
rlabel metal2 4278 24990 4278 24990 0 net277
rlabel metal2 13662 18700 13662 18700 0 net278
rlabel metal2 6854 24174 6854 24174 0 net279
rlabel metal1 19872 38998 19872 38998 0 net28
rlabel metal1 4692 22950 4692 22950 0 net280
rlabel metal1 16560 14042 16560 14042 0 net281
rlabel metal1 19918 12104 19918 12104 0 net282
rlabel metal2 21574 44438 21574 44438 0 net283
rlabel metal1 9660 25194 9660 25194 0 net284
rlabel metal2 12466 46376 12466 46376 0 net285
rlabel metal1 10396 11866 10396 11866 0 net286
rlabel metal1 20746 11866 20746 11866 0 net287
rlabel metal1 14122 11662 14122 11662 0 net288
rlabel metal2 6854 18462 6854 18462 0 net289
rlabel metal2 15962 36448 15962 36448 0 net29
rlabel metal1 19320 34986 19320 34986 0 net290
rlabel metal2 25254 35428 25254 35428 0 net291
rlabel metal2 8418 15470 8418 15470 0 net292
rlabel metal1 16146 15130 16146 15130 0 net293
rlabel metal2 7866 42398 7866 42398 0 net294
rlabel metal1 20516 46002 20516 46002 0 net295
rlabel metal2 16054 47464 16054 47464 0 net296
rlabel metal2 22034 16796 22034 16796 0 net297
rlabel metal2 12466 23987 12466 23987 0 net298
rlabel metal1 20700 25330 20700 25330 0 net299
rlabel metal1 20424 24242 20424 24242 0 net3
rlabel metal2 21482 34969 21482 34969 0 net30
rlabel metal2 22218 18700 22218 18700 0 net300
rlabel metal1 23230 22542 23230 22542 0 net301
rlabel metal1 14858 20366 14858 20366 0 net302
rlabel metal2 19182 14484 19182 14484 0 net303
rlabel metal1 15226 30158 15226 30158 0 net304
rlabel metal1 14582 25976 14582 25976 0 net305
rlabel metal1 23920 18802 23920 18802 0 net306
rlabel metal1 16100 45390 16100 45390 0 net307
rlabel metal1 23920 31994 23920 31994 0 net308
rlabel metal2 23782 42398 23782 42398 0 net309
rlabel metal1 15410 37774 15410 37774 0 net31
rlabel metal1 14858 35258 14858 35258 0 net310
rlabel metal1 21344 20570 21344 20570 0 net311
rlabel metal1 4922 23834 4922 23834 0 net312
rlabel metal1 10902 28186 10902 28186 0 net313
rlabel metal2 25254 39508 25254 39508 0 net314
rlabel metal1 7958 21590 7958 21590 0 net315
rlabel metal1 22770 25466 22770 25466 0 net316
rlabel metal1 7813 28934 7813 28934 0 net317
rlabel metal1 7912 32470 7912 32470 0 net318
rlabel metal2 9798 34884 9798 34884 0 net319
rlabel metal1 12880 38930 12880 38930 0 net32
rlabel metal2 22310 14892 22310 14892 0 net320
rlabel metal1 18170 35598 18170 35598 0 net321
rlabel metal2 6762 26860 6762 26860 0 net322
rlabel metal1 25208 26554 25208 26554 0 net323
rlabel metal1 23092 45390 23092 45390 0 net324
rlabel metal1 9154 18598 9154 18598 0 net325
rlabel metal1 7774 39610 7774 39610 0 net326
rlabel metal2 11178 46784 11178 46784 0 net327
rlabel metal1 21942 33864 21942 33864 0 net328
rlabel metal1 16882 34714 16882 34714 0 net329
rlabel metal1 3726 3638 3726 3638 0 net33
rlabel metal2 18630 40868 18630 40868 0 net330
rlabel metal2 5842 34476 5842 34476 0 net331
rlabel metal2 11086 34986 11086 34986 0 net332
rlabel metal2 6854 28254 6854 28254 0 net333
rlabel metal1 18032 46478 18032 46478 0 net334
rlabel metal1 19228 42262 19228 42262 0 net335
rlabel metal1 16054 33082 16054 33082 0 net336
rlabel metal2 16146 32980 16146 32980 0 net337
rlabel metal2 12466 35190 12466 35190 0 net338
rlabel metal1 14950 22406 14950 22406 0 net339
rlabel metal2 5198 4352 5198 4352 0 net34
rlabel metal2 16514 46308 16514 46308 0 net340
rlabel metal2 13386 41242 13386 41242 0 net341
rlabel metal2 9154 14110 9154 14110 0 net342
rlabel metal1 23782 38862 23782 38862 0 net343
rlabel metal2 6578 35292 6578 35292 0 net344
rlabel metal1 19044 43214 19044 43214 0 net345
rlabel metal2 7774 20060 7774 20060 0 net346
rlabel metal1 10810 42602 10810 42602 0 net347
rlabel metal1 22862 42330 22862 42330 0 net348
rlabel metal1 16008 40698 16008 40698 0 net349
rlabel metal2 5934 7480 5934 7480 0 net35
rlabel metal2 6026 38114 6026 38114 0 net350
rlabel metal1 5566 17306 5566 17306 0 net351
rlabel metal1 23920 44914 23920 44914 0 net352
rlabel metal2 10534 28832 10534 28832 0 net353
rlabel metal1 10396 13498 10396 13498 0 net354
rlabel metal2 13570 27166 13570 27166 0 net355
rlabel metal1 7123 16762 7123 16762 0 net356
rlabel metal1 17894 24106 17894 24106 0 net357
rlabel metal1 18630 33592 18630 33592 0 net358
rlabel metal1 25162 37230 25162 37230 0 net359
rlabel metal2 16146 3876 16146 3876 0 net36
rlabel metal2 8602 15062 8602 15062 0 net360
rlabel metal1 23966 37434 23966 37434 0 net361
rlabel metal1 17204 38998 17204 38998 0 net362
rlabel metal1 19734 22066 19734 22066 0 net363
rlabel metal1 9844 31858 9844 31858 0 net364
rlabel metal1 24564 41786 24564 41786 0 net365
rlabel metal1 15088 41038 15088 41038 0 net366
rlabel metal1 19366 21454 19366 21454 0 net367
rlabel metal2 11270 25500 11270 25500 0 net368
rlabel metal1 8096 21114 8096 21114 0 net369
rlabel metal1 6394 3706 6394 3706 0 net37
rlabel metal2 23966 43248 23966 43248 0 net370
rlabel metal1 6348 21114 6348 21114 0 net371
rlabel metal3 8349 19244 8349 19244 0 net38
rlabel metal1 7406 2618 7406 2618 0 net39
rlabel metal1 15180 33626 15180 33626 0 net4
rlabel metal1 11132 2414 11132 2414 0 net40
rlabel metal1 7820 3706 7820 3706 0 net41
rlabel metal1 7544 3162 7544 3162 0 net42
rlabel metal2 8510 3655 8510 3655 0 net43
rlabel metal1 3956 2890 3956 2890 0 net44
rlabel metal1 11408 5678 11408 5678 0 net45
rlabel metal1 9430 3706 9430 3706 0 net46
rlabel metal1 12098 9622 12098 9622 0 net47
rlabel metal1 10442 2618 10442 2618 0 net48
rlabel metal1 11270 5814 11270 5814 0 net49
rlabel metal1 22540 30702 22540 30702 0 net5
rlabel metal1 13018 3434 13018 3434 0 net50
rlabel via2 11914 3179 11914 3179 0 net51
rlabel metal2 16882 11798 16882 11798 0 net52
rlabel metal1 13754 2618 13754 2618 0 net53
rlabel metal1 11730 2550 11730 2550 0 net54
rlabel metal2 1886 7514 1886 7514 0 net55
rlabel metal2 2714 4386 2714 4386 0 net56
rlabel metal1 5658 2958 5658 2958 0 net57
rlabel metal2 2622 3434 2622 3434 0 net58
rlabel metal1 4094 2618 4094 2618 0 net59
rlabel metal1 20286 32470 20286 32470 0 net6
rlabel metal1 5888 2550 5888 2550 0 net60
rlabel metal2 5014 7650 5014 7650 0 net61
rlabel metal1 5428 3706 5428 3706 0 net62
rlabel metal1 12880 40494 12880 40494 0 net63
rlabel metal3 17319 52564 17319 52564 0 net64
rlabel metal1 11592 21862 11592 21862 0 net65
rlabel metal1 17940 47770 17940 47770 0 net66
rlabel metal1 19090 41446 19090 41446 0 net67
rlabel metal2 18538 50626 18538 50626 0 net68
rlabel metal1 19320 47702 19320 47702 0 net69
rlabel metal1 20286 37196 20286 37196 0 net7
rlabel metal2 18630 49980 18630 49980 0 net70
rlabel metal1 18538 11118 18538 11118 0 net71
rlabel via2 19366 44693 19366 44693 0 net72
rlabel metal1 21160 46682 21160 46682 0 net73
rlabel metal3 13777 52564 13777 52564 0 net74
rlabel metal1 20286 46682 20286 46682 0 net75
rlabel metal2 21942 43231 21942 43231 0 net76
rlabel metal1 21390 44166 21390 44166 0 net77
rlabel metal1 22172 12818 22172 12818 0 net78
rlabel metal1 21390 53414 21390 53414 0 net79
rlabel metal1 20746 36856 20746 36856 0 net8
rlabel metal2 22494 50048 22494 50048 0 net80
rlabel metal1 21068 11050 21068 11050 0 net81
rlabel metal1 22770 53686 22770 53686 0 net82
rlabel metal1 22954 52870 22954 52870 0 net83
rlabel metal1 23368 45934 23368 45934 0 net84
rlabel via3 14053 52564 14053 52564 0 net85
rlabel metal2 14536 44506 14536 44506 0 net86
rlabel metal1 14950 43418 14950 43418 0 net87
rlabel metal1 16514 44166 16514 44166 0 net88
rlabel metal3 15847 53924 15847 53924 0 net89
rlabel metal1 19918 36244 19918 36244 0 net9
rlabel metal3 15571 52564 15571 52564 0 net90
rlabel metal2 15962 50320 15962 50320 0 net91
rlabel metal1 10488 17170 10488 17170 0 net92
rlabel metal1 2530 33286 2530 33286 0 net93
rlabel metal2 1610 32300 1610 32300 0 net94
rlabel metal1 2760 38182 2760 38182 0 net95
rlabel metal1 2622 40902 2622 40902 0 net96
rlabel metal2 6854 18938 6854 18938 0 net97
rlabel metal2 6762 19571 6762 19571 0 net98
rlabel metal1 16192 17306 16192 17306 0 net99
rlabel metal2 23782 2115 23782 2115 0 prog_clk
rlabel metal2 23598 3230 23598 3230 0 prog_reset
rlabel metal2 25070 50711 25070 50711 0 right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_
rlabel metal2 25530 51561 25530 51561 0 right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_
rlabel metal2 24794 52309 24794 52309 0 right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_
rlabel metal2 25070 53023 25070 53023 0 right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_
rlabel metal2 25070 53975 25070 53975 0 right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_4_
rlabel metal1 24886 53550 24886 53550 0 right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_5_
rlabel metal3 25538 55420 25538 55420 0 right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_6_
rlabel metal3 25446 56236 25446 56236 0 right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_7_
rlabel metal3 1786 4012 1786 4012 0 right_width_0_height_0_subtile_0__pin_inpad_0_
rlabel metal3 1878 6460 1878 6460 0 right_width_0_height_0_subtile_1__pin_inpad_0_
rlabel metal3 1786 8908 1786 8908 0 right_width_0_height_0_subtile_2__pin_inpad_0_
rlabel metal3 1740 11356 1740 11356 0 right_width_0_height_0_subtile_3__pin_inpad_0_
rlabel metal1 20608 15130 20608 15130 0 sb_0__1_.mem_bottom_track_1.ccff_head
rlabel metal1 20056 21658 20056 21658 0 sb_0__1_.mem_bottom_track_1.ccff_tail
rlabel metal1 20700 21862 20700 21862 0 sb_0__1_.mem_bottom_track_1.mem_out\[0\]
rlabel metal1 17940 21454 17940 21454 0 sb_0__1_.mem_bottom_track_1.mem_out\[1\]
rlabel metal1 16790 24378 16790 24378 0 sb_0__1_.mem_bottom_track_11.ccff_head
rlabel metal1 15226 27098 15226 27098 0 sb_0__1_.mem_bottom_track_11.ccff_tail
rlabel metal1 18446 34442 18446 34442 0 sb_0__1_.mem_bottom_track_11.mem_out\[0\]
rlabel metal2 14766 28628 14766 28628 0 sb_0__1_.mem_bottom_track_11.mem_out\[1\]
rlabel metal2 22126 24922 22126 24922 0 sb_0__1_.mem_bottom_track_13.ccff_tail
rlabel metal1 21160 34374 21160 34374 0 sb_0__1_.mem_bottom_track_13.mem_out\[0\]
rlabel metal2 20930 28832 20930 28832 0 sb_0__1_.mem_bottom_track_13.mem_out\[1\]
rlabel metal1 24288 24582 24288 24582 0 sb_0__1_.mem_bottom_track_21.ccff_tail
rlabel metal1 20148 30770 20148 30770 0 sb_0__1_.mem_bottom_track_21.mem_out\[0\]
rlabel metal1 23690 27506 23690 27506 0 sb_0__1_.mem_bottom_track_21.mem_out\[1\]
rlabel metal2 16330 29308 16330 29308 0 sb_0__1_.mem_bottom_track_29.ccff_tail
rlabel metal1 20194 29240 20194 29240 0 sb_0__1_.mem_bottom_track_29.mem_out\[0\]
rlabel metal1 17894 32266 17894 32266 0 sb_0__1_.mem_bottom_track_29.mem_out\[1\]
rlabel metal1 21160 20434 21160 20434 0 sb_0__1_.mem_bottom_track_3.ccff_tail
rlabel metal1 20240 27506 20240 27506 0 sb_0__1_.mem_bottom_track_3.mem_out\[0\]
rlabel metal1 19090 20842 19090 20842 0 sb_0__1_.mem_bottom_track_3.mem_out\[1\]
rlabel metal1 14950 32878 14950 32878 0 sb_0__1_.mem_bottom_track_37.ccff_tail
rlabel metal1 16514 31994 16514 31994 0 sb_0__1_.mem_bottom_track_37.mem_out\[0\]
rlabel metal1 14720 33286 14720 33286 0 sb_0__1_.mem_bottom_track_37.mem_out\[1\]
rlabel metal2 20102 34000 20102 34000 0 sb_0__1_.mem_bottom_track_45.ccff_tail
rlabel metal1 18262 34986 18262 34986 0 sb_0__1_.mem_bottom_track_45.mem_out\[0\]
rlabel metal1 21252 34918 21252 34918 0 sb_0__1_.mem_bottom_track_45.mem_out\[1\]
rlabel metal2 23414 21828 23414 21828 0 sb_0__1_.mem_bottom_track_5.ccff_tail
rlabel metal1 22816 22066 22816 22066 0 sb_0__1_.mem_bottom_track_5.mem_out\[0\]
rlabel metal1 24012 21454 24012 21454 0 sb_0__1_.mem_bottom_track_5.mem_out\[1\]
rlabel metal1 15732 37774 15732 37774 0 sb_0__1_.mem_bottom_track_53.mem_out\[0\]
rlabel metal2 17434 29325 17434 29325 0 sb_0__1_.mem_bottom_track_7.mem_out\[0\]
rlabel metal1 18538 24718 18538 24718 0 sb_0__1_.mem_bottom_track_7.mem_out\[1\]
rlabel metal2 18630 39270 18630 39270 0 sb_0__1_.mem_right_track_0.ccff_head
rlabel metal1 23046 31790 23046 31790 0 sb_0__1_.mem_right_track_0.ccff_tail
rlabel metal1 20838 33966 20838 33966 0 sb_0__1_.mem_right_track_0.mem_out\[0\]
rlabel metal1 23138 31858 23138 31858 0 sb_0__1_.mem_right_track_0.mem_out\[1\]
rlabel metal1 23276 40562 23276 40562 0 sb_0__1_.mem_right_track_10.ccff_head
rlabel metal1 20884 42058 20884 42058 0 sb_0__1_.mem_right_track_10.ccff_tail
rlabel metal1 21206 45390 21206 45390 0 sb_0__1_.mem_right_track_10.mem_out\[0\]
rlabel metal1 21022 42534 21022 42534 0 sb_0__1_.mem_right_track_10.mem_out\[1\]
rlabel metal1 20056 43078 20056 43078 0 sb_0__1_.mem_right_track_12.ccff_tail
rlabel metal1 20930 45050 20930 45050 0 sb_0__1_.mem_right_track_12.mem_out\[0\]
rlabel metal1 18768 36686 18768 36686 0 sb_0__1_.mem_right_track_12.mem_out\[1\]
rlabel metal1 18768 44166 18768 44166 0 sb_0__1_.mem_right_track_14.ccff_tail
rlabel metal1 19734 47022 19734 47022 0 sb_0__1_.mem_right_track_14.mem_out\[0\]
rlabel metal1 18722 41616 18722 41616 0 sb_0__1_.mem_right_track_14.mem_out\[1\]
rlabel metal1 16882 44744 16882 44744 0 sb_0__1_.mem_right_track_16.ccff_tail
rlabel metal2 18722 47838 18722 47838 0 sb_0__1_.mem_right_track_16.mem_out\[0\]
rlabel metal1 17618 43860 17618 43860 0 sb_0__1_.mem_right_track_16.mem_out\[1\]
rlabel metal1 16698 40018 16698 40018 0 sb_0__1_.mem_right_track_18.ccff_tail
rlabel metal1 16928 45458 16928 45458 0 sb_0__1_.mem_right_track_18.mem_out\[0\]
rlabel metal1 15870 43758 15870 43758 0 sb_0__1_.mem_right_track_18.mem_out\[1\]
rlabel metal1 25024 42670 25024 42670 0 sb_0__1_.mem_right_track_2.ccff_tail
rlabel metal2 21896 42636 21896 42636 0 sb_0__1_.mem_right_track_2.mem_out\[0\]
rlabel metal1 23460 39474 23460 39474 0 sb_0__1_.mem_right_track_2.mem_out\[1\]
rlabel metal1 14030 34102 14030 34102 0 sb_0__1_.mem_right_track_20.ccff_tail
rlabel metal1 15088 43146 15088 43146 0 sb_0__1_.mem_right_track_20.mem_out\[0\]
rlabel metal1 11914 36720 11914 36720 0 sb_0__1_.mem_right_track_20.mem_out\[1\]
rlabel via1 13018 30685 13018 30685 0 sb_0__1_.mem_right_track_22.ccff_tail
rlabel metal1 13570 35530 13570 35530 0 sb_0__1_.mem_right_track_22.mem_out\[0\]
rlabel metal1 13662 34476 13662 34476 0 sb_0__1_.mem_right_track_22.mem_out\[1\]
rlabel metal1 13202 25840 13202 25840 0 sb_0__1_.mem_right_track_24.ccff_tail
rlabel metal1 13662 28152 13662 28152 0 sb_0__1_.mem_right_track_24.mem_out\[0\]
rlabel metal2 8786 28254 8786 28254 0 sb_0__1_.mem_right_track_26.ccff_tail
rlabel metal1 14858 30804 14858 30804 0 sb_0__1_.mem_right_track_26.mem_out\[0\]
rlabel metal1 9522 26826 9522 26826 0 sb_0__1_.mem_right_track_28.ccff_tail
rlabel metal1 8464 28186 8464 28186 0 sb_0__1_.mem_right_track_28.mem_out\[0\]
rlabel metal1 13294 24820 13294 24820 0 sb_0__1_.mem_right_track_30.ccff_tail
rlabel metal1 12811 28594 12811 28594 0 sb_0__1_.mem_right_track_30.mem_out\[0\]
rlabel metal1 14214 24174 14214 24174 0 sb_0__1_.mem_right_track_32.ccff_tail
rlabel metal1 11914 26962 11914 26962 0 sb_0__1_.mem_right_track_32.mem_out\[0\]
rlabel metal1 16284 21114 16284 21114 0 sb_0__1_.mem_right_track_34.ccff_tail
rlabel metal2 14674 24718 14674 24718 0 sb_0__1_.mem_right_track_34.mem_out\[0\]
rlabel metal1 10810 12954 10810 12954 0 sb_0__1_.mem_right_track_36.ccff_tail
rlabel metal1 14398 20570 14398 20570 0 sb_0__1_.mem_right_track_36.mem_out\[0\]
rlabel metal2 9338 17306 9338 17306 0 sb_0__1_.mem_right_track_36.mem_out\[1\]
rlabel via1 14306 12274 14306 12274 0 sb_0__1_.mem_right_track_38.ccff_tail
rlabel metal2 11730 13294 11730 13294 0 sb_0__1_.mem_right_track_38.mem_out\[0\]
rlabel metal2 24058 34476 24058 34476 0 sb_0__1_.mem_right_track_4.ccff_tail
rlabel metal1 24426 40494 24426 40494 0 sb_0__1_.mem_right_track_4.mem_out\[0\]
rlabel metal1 22402 34986 22402 34986 0 sb_0__1_.mem_right_track_4.mem_out\[1\]
rlabel metal2 17066 13056 17066 13056 0 sb_0__1_.mem_right_track_40.ccff_tail
rlabel metal1 14812 11118 14812 11118 0 sb_0__1_.mem_right_track_40.mem_out\[0\]
rlabel metal1 17894 15674 17894 15674 0 sb_0__1_.mem_right_track_44.ccff_tail
rlabel metal2 15686 14790 15686 14790 0 sb_0__1_.mem_right_track_44.mem_out\[0\]
rlabel metal1 20332 18122 20332 18122 0 sb_0__1_.mem_right_track_46.ccff_tail
rlabel metal2 16882 17306 16882 17306 0 sb_0__1_.mem_right_track_46.mem_out\[0\]
rlabel metal1 24150 17850 24150 17850 0 sb_0__1_.mem_right_track_48.ccff_tail
rlabel metal2 21482 18836 21482 18836 0 sb_0__1_.mem_right_track_48.mem_out\[0\]
rlabel metal1 21850 18802 21850 18802 0 sb_0__1_.mem_right_track_50.ccff_tail
rlabel metal1 22218 19278 22218 19278 0 sb_0__1_.mem_right_track_50.mem_out\[0\]
rlabel metal2 22126 13770 22126 13770 0 sb_0__1_.mem_right_track_52.ccff_tail
rlabel metal2 24610 15946 24610 15946 0 sb_0__1_.mem_right_track_52.mem_out\[0\]
rlabel metal2 19734 11050 19734 11050 0 sb_0__1_.mem_right_track_54.ccff_tail
rlabel via1 18722 12206 18722 12206 0 sb_0__1_.mem_right_track_54.mem_out\[0\]
rlabel metal1 18722 13906 18722 13906 0 sb_0__1_.mem_right_track_56.mem_out\[0\]
rlabel metal1 24656 37638 24656 37638 0 sb_0__1_.mem_right_track_6.ccff_tail
rlabel metal1 20194 32980 20194 32980 0 sb_0__1_.mem_right_track_6.mem_out\[0\]
rlabel metal1 24518 36890 24518 36890 0 sb_0__1_.mem_right_track_6.mem_out\[1\]
rlabel metal2 21482 39202 21482 39202 0 sb_0__1_.mem_right_track_8.mem_out\[0\]
rlabel metal1 22494 42772 22494 42772 0 sb_0__1_.mem_right_track_8.mem_out\[1\]
rlabel metal1 11638 46886 11638 46886 0 sb_0__1_.mem_top_track_0.ccff_tail
rlabel metal1 17296 42058 17296 42058 0 sb_0__1_.mem_top_track_0.mem_out\[0\]
rlabel metal1 12466 44268 12466 44268 0 sb_0__1_.mem_top_track_0.mem_out\[1\]
rlabel metal2 7774 39440 7774 39440 0 sb_0__1_.mem_top_track_10.ccff_head
rlabel metal1 6072 35802 6072 35802 0 sb_0__1_.mem_top_track_10.ccff_tail
rlabel metal1 17664 37638 17664 37638 0 sb_0__1_.mem_top_track_10.mem_out\[0\]
rlabel metal2 7038 37298 7038 37298 0 sb_0__1_.mem_top_track_10.mem_out\[1\]
rlabel metal1 7636 33490 7636 33490 0 sb_0__1_.mem_top_track_12.ccff_tail
rlabel metal2 8602 32402 8602 32402 0 sb_0__1_.mem_top_track_12.mem_out\[0\]
rlabel metal1 8280 32946 8280 32946 0 sb_0__1_.mem_top_track_12.mem_out\[1\]
rlabel metal1 13800 45390 13800 45390 0 sb_0__1_.mem_top_track_2.ccff_tail
rlabel metal1 17802 43214 17802 43214 0 sb_0__1_.mem_top_track_2.mem_out\[0\]
rlabel metal1 14720 42126 14720 42126 0 sb_0__1_.mem_top_track_2.mem_out\[1\]
rlabel metal1 9568 34714 9568 34714 0 sb_0__1_.mem_top_track_20.ccff_tail
rlabel metal1 14030 32334 14030 32334 0 sb_0__1_.mem_top_track_20.mem_out\[0\]
rlabel metal1 13386 35088 13386 35088 0 sb_0__1_.mem_top_track_20.mem_out\[1\]
rlabel metal1 5382 38964 5382 38964 0 sb_0__1_.mem_top_track_28.ccff_tail
rlabel metal2 13386 34612 13386 34612 0 sb_0__1_.mem_top_track_28.mem_out\[0\]
rlabel metal1 7360 35258 7360 35258 0 sb_0__1_.mem_top_track_28.mem_out\[1\]
rlabel metal1 9062 41718 9062 41718 0 sb_0__1_.mem_top_track_36.ccff_tail
rlabel metal1 8142 39406 8142 39406 0 sb_0__1_.mem_top_track_36.mem_out\[0\]
rlabel metal1 12834 38828 12834 38828 0 sb_0__1_.mem_top_track_36.mem_out\[1\]
rlabel metal1 9384 41242 9384 41242 0 sb_0__1_.mem_top_track_4.ccff_tail
rlabel metal1 14444 41446 14444 41446 0 sb_0__1_.mem_top_track_4.mem_out\[0\]
rlabel metal1 12650 41582 12650 41582 0 sb_0__1_.mem_top_track_4.mem_out\[1\]
rlabel metal1 13248 42738 13248 42738 0 sb_0__1_.mem_top_track_44.ccff_tail
rlabel metal1 12834 39032 12834 39032 0 sb_0__1_.mem_top_track_44.mem_out\[0\]
rlabel metal1 16560 42806 16560 42806 0 sb_0__1_.mem_top_track_52.mem_out\[0\]
rlabel metal1 16974 39406 16974 39406 0 sb_0__1_.mem_top_track_52.mem_out\[1\]
rlabel metal2 17526 38114 17526 38114 0 sb_0__1_.mem_top_track_6.mem_out\[0\]
rlabel metal1 8970 37434 8970 37434 0 sb_0__1_.mem_top_track_6.mem_out\[1\]
rlabel metal1 19458 7412 19458 7412 0 sb_0__1_.mux_bottom_track_1.out
rlabel metal2 18354 26928 18354 26928 0 sb_0__1_.mux_bottom_track_1.sky130_fd_sc_hd__mux2_1_0_X
rlabel metal1 18584 32198 18584 32198 0 sb_0__1_.mux_bottom_track_1.sky130_fd_sc_hd__mux2_1_1_X
rlabel metal1 15548 22474 15548 22474 0 sb_0__1_.mux_bottom_track_1.sky130_fd_sc_hd__mux2_1_2_X
rlabel metal1 17848 22066 17848 22066 0 sb_0__1_.mux_bottom_track_1.sky130_fd_sc_hd__mux2_1_3_X
rlabel metal1 17342 21658 17342 21658 0 sb_0__1_.mux_bottom_track_1.sky130_fd_sc_hd__mux2_1_4_X
rlabel metal1 17112 21862 17112 21862 0 sb_0__1_.mux_bottom_track_1.sky130_fd_sc_hd__mux2_1_5_X
rlabel metal1 16882 7446 16882 7446 0 sb_0__1_.mux_bottom_track_11.out
rlabel metal1 17250 31926 17250 31926 0 sb_0__1_.mux_bottom_track_11.sky130_fd_sc_hd__mux2_1_0_X
rlabel metal1 17158 29206 17158 29206 0 sb_0__1_.mux_bottom_track_11.sky130_fd_sc_hd__mux2_1_1_X
rlabel metal1 13478 26452 13478 26452 0 sb_0__1_.mux_bottom_track_11.sky130_fd_sc_hd__mux2_1_2_X
rlabel metal2 13386 25840 13386 25840 0 sb_0__1_.mux_bottom_track_11.sky130_fd_sc_hd__mux2_1_3_X
rlabel metal1 15272 25262 15272 25262 0 sb_0__1_.mux_bottom_track_11.sky130_fd_sc_hd__mux2_1_4_X
rlabel metal1 14904 25262 14904 25262 0 sb_0__1_.mux_bottom_track_11.sky130_fd_sc_hd__mux2_1_5_X
rlabel metal1 15272 17646 15272 17646 0 sb_0__1_.mux_bottom_track_11.sky130_fd_sc_hd__mux2_1_6_X
rlabel metal1 18998 9622 18998 9622 0 sb_0__1_.mux_bottom_track_13.out
rlabel metal1 19182 29682 19182 29682 0 sb_0__1_.mux_bottom_track_13.sky130_fd_sc_hd__mux2_1_0_X
rlabel metal1 20286 29614 20286 29614 0 sb_0__1_.mux_bottom_track_13.sky130_fd_sc_hd__mux2_1_1_X
rlabel metal1 18998 26418 18998 26418 0 sb_0__1_.mux_bottom_track_13.sky130_fd_sc_hd__mux2_1_2_X
rlabel metal1 20010 24786 20010 24786 0 sb_0__1_.mux_bottom_track_13.sky130_fd_sc_hd__mux2_1_3_X
rlabel metal1 19734 24922 19734 24922 0 sb_0__1_.mux_bottom_track_13.sky130_fd_sc_hd__mux2_1_4_X
rlabel metal1 18538 19346 18538 19346 0 sb_0__1_.mux_bottom_track_13.sky130_fd_sc_hd__mux2_1_5_X
rlabel metal1 21114 8534 21114 8534 0 sb_0__1_.mux_bottom_track_21.out
rlabel metal2 20746 30022 20746 30022 0 sb_0__1_.mux_bottom_track_21.sky130_fd_sc_hd__mux2_1_0_X
rlabel metal2 22034 31824 22034 31824 0 sb_0__1_.mux_bottom_track_21.sky130_fd_sc_hd__mux2_1_1_X
rlabel metal1 22402 26010 22402 26010 0 sb_0__1_.mux_bottom_track_21.sky130_fd_sc_hd__mux2_1_2_X
rlabel metal2 21942 26622 21942 26622 0 sb_0__1_.mux_bottom_track_21.sky130_fd_sc_hd__mux2_1_3_X
rlabel metal2 22402 24922 22402 24922 0 sb_0__1_.mux_bottom_track_21.sky130_fd_sc_hd__mux2_1_4_X
rlabel metal2 21712 19652 21712 19652 0 sb_0__1_.mux_bottom_track_21.sky130_fd_sc_hd__mux2_1_5_X
rlabel metal1 17250 9622 17250 9622 0 sb_0__1_.mux_bottom_track_29.out
rlabel metal1 17250 32334 17250 32334 0 sb_0__1_.mux_bottom_track_29.sky130_fd_sc_hd__mux2_1_0_X
rlabel metal1 20194 37128 20194 37128 0 sb_0__1_.mux_bottom_track_29.sky130_fd_sc_hd__mux2_1_1_X
rlabel metal1 17802 29274 17802 29274 0 sb_0__1_.mux_bottom_track_29.sky130_fd_sc_hd__mux2_1_2_X
rlabel metal1 17158 32198 17158 32198 0 sb_0__1_.mux_bottom_track_29.sky130_fd_sc_hd__mux2_1_3_X
rlabel metal1 16836 28526 16836 28526 0 sb_0__1_.mux_bottom_track_29.sky130_fd_sc_hd__mux2_1_4_X
rlabel metal1 16468 20910 16468 20910 0 sb_0__1_.mux_bottom_track_29.sky130_fd_sc_hd__mux2_1_5_X
rlabel metal1 17940 6766 17940 6766 0 sb_0__1_.mux_bottom_track_3.out
rlabel metal2 19734 26656 19734 26656 0 sb_0__1_.mux_bottom_track_3.sky130_fd_sc_hd__mux2_1_0_X
rlabel metal1 19734 31926 19734 31926 0 sb_0__1_.mux_bottom_track_3.sky130_fd_sc_hd__mux2_1_1_X
rlabel metal1 19320 20570 19320 20570 0 sb_0__1_.mux_bottom_track_3.sky130_fd_sc_hd__mux2_1_2_X
rlabel metal1 19228 20434 19228 20434 0 sb_0__1_.mux_bottom_track_3.sky130_fd_sc_hd__mux2_1_3_X
rlabel metal1 16468 13906 16468 13906 0 sb_0__1_.mux_bottom_track_3.sky130_fd_sc_hd__mux2_1_4_X
rlabel metal1 11500 19414 11500 19414 0 sb_0__1_.mux_bottom_track_37.out
rlabel metal2 16054 36108 16054 36108 0 sb_0__1_.mux_bottom_track_37.sky130_fd_sc_hd__mux2_1_0_X
rlabel metal1 17756 34646 17756 34646 0 sb_0__1_.mux_bottom_track_37.sky130_fd_sc_hd__mux2_1_1_X
rlabel metal1 15410 34714 15410 34714 0 sb_0__1_.mux_bottom_track_37.sky130_fd_sc_hd__mux2_1_2_X
rlabel metal2 13386 28934 13386 28934 0 sb_0__1_.mux_bottom_track_37.sky130_fd_sc_hd__mux2_1_3_X
rlabel metal1 12834 22610 12834 22610 0 sb_0__1_.mux_bottom_track_37.sky130_fd_sc_hd__mux2_1_4_X
rlabel metal1 17710 10030 17710 10030 0 sb_0__1_.mux_bottom_track_45.out
rlabel metal2 21390 37468 21390 37468 0 sb_0__1_.mux_bottom_track_45.sky130_fd_sc_hd__mux2_1_0_X
rlabel metal1 20470 36006 20470 36006 0 sb_0__1_.mux_bottom_track_45.sky130_fd_sc_hd__mux2_1_1_X
rlabel metal1 21850 33286 21850 33286 0 sb_0__1_.mux_bottom_track_45.sky130_fd_sc_hd__mux2_1_2_X
rlabel metal1 19090 19822 19090 19822 0 sb_0__1_.mux_bottom_track_45.sky130_fd_sc_hd__mux2_1_3_X
rlabel metal1 18170 12138 18170 12138 0 sb_0__1_.mux_bottom_track_5.out
rlabel metal1 21390 29036 21390 29036 0 sb_0__1_.mux_bottom_track_5.sky130_fd_sc_hd__mux2_1_0_X
rlabel metal1 22724 26282 22724 26282 0 sb_0__1_.mux_bottom_track_5.sky130_fd_sc_hd__mux2_1_1_X
rlabel metal1 25070 23188 25070 23188 0 sb_0__1_.mux_bottom_track_5.sky130_fd_sc_hd__mux2_1_2_X
rlabel metal2 22494 23936 22494 23936 0 sb_0__1_.mux_bottom_track_5.sky130_fd_sc_hd__mux2_1_3_X
rlabel metal1 22494 21522 22494 21522 0 sb_0__1_.mux_bottom_track_5.sky130_fd_sc_hd__mux2_1_4_X
rlabel metal1 21528 14994 21528 14994 0 sb_0__1_.mux_bottom_track_5.sky130_fd_sc_hd__mux2_1_5_X
rlabel metal1 9798 18394 9798 18394 0 sb_0__1_.mux_bottom_track_53.out
rlabel metal2 14214 37978 14214 37978 0 sb_0__1_.mux_bottom_track_53.sky130_fd_sc_hd__mux2_1_0_X
rlabel metal2 11730 37468 11730 37468 0 sb_0__1_.mux_bottom_track_53.sky130_fd_sc_hd__mux2_1_1_X
rlabel metal1 11270 37094 11270 37094 0 sb_0__1_.mux_bottom_track_53.sky130_fd_sc_hd__mux2_1_2_X
rlabel metal1 17986 8534 17986 8534 0 sb_0__1_.mux_bottom_track_7.out
rlabel metal1 18308 27438 18308 27438 0 sb_0__1_.mux_bottom_track_7.sky130_fd_sc_hd__mux2_1_0_X
rlabel metal1 19688 32198 19688 32198 0 sb_0__1_.mux_bottom_track_7.sky130_fd_sc_hd__mux2_1_1_X
rlabel metal1 16192 24786 16192 24786 0 sb_0__1_.mux_bottom_track_7.sky130_fd_sc_hd__mux2_1_2_X
rlabel metal2 15410 24310 15410 24310 0 sb_0__1_.mux_bottom_track_7.sky130_fd_sc_hd__mux2_1_3_X
rlabel metal1 17526 23834 17526 23834 0 sb_0__1_.mux_bottom_track_7.sky130_fd_sc_hd__mux2_1_4_X
rlabel metal2 17250 24208 17250 24208 0 sb_0__1_.mux_bottom_track_7.sky130_fd_sc_hd__mux2_1_5_X
rlabel metal1 16376 19822 16376 19822 0 sb_0__1_.mux_bottom_track_7.sky130_fd_sc_hd__mux2_1_6_X
rlabel metal2 24794 25500 24794 25500 0 sb_0__1_.mux_right_track_0.out
rlabel metal2 20930 32300 20930 32300 0 sb_0__1_.mux_right_track_0.sky130_fd_sc_hd__mux2_1_0_X
rlabel metal1 22172 32742 22172 32742 0 sb_0__1_.mux_right_track_0.sky130_fd_sc_hd__mux2_1_1_X
rlabel metal1 22678 31926 22678 31926 0 sb_0__1_.mux_right_track_0.sky130_fd_sc_hd__mux2_1_2_X
rlabel metal2 22586 29172 22586 29172 0 sb_0__1_.mux_right_track_0.sky130_fd_sc_hd__mux2_1_3_X
rlabel metal2 24794 29036 24794 29036 0 sb_0__1_.mux_right_track_0.sky130_fd_sc_hd__mux2_1_4_X
rlabel metal1 23092 32198 23092 32198 0 sb_0__1_.mux_right_track_10.out
rlabel metal1 20194 41582 20194 41582 0 sb_0__1_.mux_right_track_10.sky130_fd_sc_hd__mux2_1_0_X
rlabel metal1 20332 40154 20332 40154 0 sb_0__1_.mux_right_track_10.sky130_fd_sc_hd__mux2_1_1_X
rlabel metal1 20378 37978 20378 37978 0 sb_0__1_.mux_right_track_10.sky130_fd_sc_hd__mux2_1_2_X
rlabel metal2 16238 37094 16238 37094 0 sb_0__1_.mux_right_track_10.sky130_fd_sc_hd__mux2_1_3_X
rlabel metal2 20286 35088 20286 35088 0 sb_0__1_.mux_right_track_10.sky130_fd_sc_hd__mux2_1_4_X
rlabel metal1 22586 32198 22586 32198 0 sb_0__1_.mux_right_track_12.out
rlabel metal1 19780 46342 19780 46342 0 sb_0__1_.mux_right_track_12.sky130_fd_sc_hd__mux2_1_0_X
rlabel metal1 19642 40154 19642 40154 0 sb_0__1_.mux_right_track_12.sky130_fd_sc_hd__mux2_1_1_X
rlabel metal1 19550 39814 19550 39814 0 sb_0__1_.mux_right_track_12.sky130_fd_sc_hd__mux2_1_2_X
rlabel metal1 19458 39984 19458 39984 0 sb_0__1_.mux_right_track_12.sky130_fd_sc_hd__mux2_1_3_X
rlabel metal1 21942 32198 21942 32198 0 sb_0__1_.mux_right_track_14.out
rlabel metal1 18492 41650 18492 41650 0 sb_0__1_.mux_right_track_14.sky130_fd_sc_hd__mux2_1_0_X
rlabel metal1 18308 41446 18308 41446 0 sb_0__1_.mux_right_track_14.sky130_fd_sc_hd__mux2_1_1_X
rlabel metal1 16422 38522 16422 38522 0 sb_0__1_.mux_right_track_14.sky130_fd_sc_hd__mux2_1_2_X
rlabel metal2 18262 40103 18262 40103 0 sb_0__1_.mux_right_track_14.sky130_fd_sc_hd__mux2_1_3_X
rlabel metal1 21160 31722 21160 31722 0 sb_0__1_.mux_right_track_16.out
rlabel metal1 17802 47430 17802 47430 0 sb_0__1_.mux_right_track_16.sky130_fd_sc_hd__mux2_1_0_X
rlabel metal1 17158 43622 17158 43622 0 sb_0__1_.mux_right_track_16.sky130_fd_sc_hd__mux2_1_1_X
rlabel metal1 15686 39610 15686 39610 0 sb_0__1_.mux_right_track_16.sky130_fd_sc_hd__mux2_1_2_X
rlabel metal1 20148 32402 20148 32402 0 sb_0__1_.mux_right_track_16.sky130_fd_sc_hd__mux2_1_3_X
rlabel metal1 20861 30022 20861 30022 0 sb_0__1_.mux_right_track_18.out
rlabel metal1 16790 41582 16790 41582 0 sb_0__1_.mux_right_track_18.sky130_fd_sc_hd__mux2_1_0_X
rlabel metal1 16514 37298 16514 37298 0 sb_0__1_.mux_right_track_18.sky130_fd_sc_hd__mux2_1_1_X
rlabel metal1 13064 36890 13064 36890 0 sb_0__1_.mux_right_track_18.sky130_fd_sc_hd__mux2_1_2_X
rlabel metal2 16192 34442 16192 34442 0 sb_0__1_.mux_right_track_18.sky130_fd_sc_hd__mux2_1_3_X
rlabel metal1 24656 29206 24656 29206 0 sb_0__1_.mux_right_track_2.out
rlabel metal1 22954 41650 22954 41650 0 sb_0__1_.mux_right_track_2.sky130_fd_sc_hd__mux2_1_0_X
rlabel metal1 22080 39610 22080 39610 0 sb_0__1_.mux_right_track_2.sky130_fd_sc_hd__mux2_1_1_X
rlabel metal1 20332 36890 20332 36890 0 sb_0__1_.mux_right_track_2.sky130_fd_sc_hd__mux2_1_2_X
rlabel metal1 24426 41718 24426 41718 0 sb_0__1_.mux_right_track_2.sky130_fd_sc_hd__mux2_1_3_X
rlabel metal1 24426 39338 24426 39338 0 sb_0__1_.mux_right_track_2.sky130_fd_sc_hd__mux2_1_4_X
rlabel metal2 24794 36618 24794 36618 0 sb_0__1_.mux_right_track_2.sky130_fd_sc_hd__mux2_1_5_X
rlabel metal1 22678 21896 22678 21896 0 sb_0__1_.mux_right_track_20.out
rlabel metal1 14904 43078 14904 43078 0 sb_0__1_.mux_right_track_20.sky130_fd_sc_hd__mux2_1_0_X
rlabel metal1 14628 32946 14628 32946 0 sb_0__1_.mux_right_track_20.sky130_fd_sc_hd__mux2_1_1_X
rlabel metal2 14674 32368 14674 32368 0 sb_0__1_.mux_right_track_20.sky130_fd_sc_hd__mux2_1_2_X
rlabel metal1 16514 33014 16514 33014 0 sb_0__1_.mux_right_track_20.sky130_fd_sc_hd__mux2_1_3_X
rlabel metal1 23782 19754 23782 19754 0 sb_0__1_.mux_right_track_22.out
rlabel metal2 13570 37570 13570 37570 0 sb_0__1_.mux_right_track_22.sky130_fd_sc_hd__mux2_1_0_X
rlabel metal1 12926 34714 12926 34714 0 sb_0__1_.mux_right_track_22.sky130_fd_sc_hd__mux2_1_1_X
rlabel metal1 12673 30226 12673 30226 0 sb_0__1_.mux_right_track_22.sky130_fd_sc_hd__mux2_1_2_X
rlabel metal1 18308 23698 18308 23698 0 sb_0__1_.mux_right_track_22.sky130_fd_sc_hd__mux2_1_3_X
rlabel metal2 20470 20298 20470 20298 0 sb_0__1_.mux_right_track_24.out
rlabel metal1 13524 26010 13524 26010 0 sb_0__1_.mux_right_track_24.sky130_fd_sc_hd__mux2_1_0_X
rlabel metal2 11822 26248 11822 26248 0 sb_0__1_.mux_right_track_24.sky130_fd_sc_hd__mux2_1_1_X
rlabel metal1 18584 20910 18584 20910 0 sb_0__1_.mux_right_track_24.sky130_fd_sc_hd__mux2_1_2_X
rlabel metal3 21183 16524 21183 16524 0 sb_0__1_.mux_right_track_26.out
rlabel metal1 13662 27472 13662 27472 0 sb_0__1_.mux_right_track_26.sky130_fd_sc_hd__mux2_1_0_X
rlabel metal2 9154 27234 9154 27234 0 sb_0__1_.mux_right_track_26.sky130_fd_sc_hd__mux2_1_1_X
rlabel metal1 16330 22644 16330 22644 0 sb_0__1_.mux_right_track_26.sky130_fd_sc_hd__mux2_1_2_X
rlabel metal1 23046 17238 23046 17238 0 sb_0__1_.mux_right_track_28.out
rlabel metal1 10718 26010 10718 26010 0 sb_0__1_.mux_right_track_28.sky130_fd_sc_hd__mux2_1_0_X
rlabel metal1 9016 25466 9016 25466 0 sb_0__1_.mux_right_track_28.sky130_fd_sc_hd__mux2_1_1_X
rlabel metal1 12259 20230 12259 20230 0 sb_0__1_.mux_right_track_28.sky130_fd_sc_hd__mux2_1_2_X
rlabel metal1 20332 16558 20332 16558 0 sb_0__1_.mux_right_track_30.out
rlabel metal2 13478 26690 13478 26690 0 sb_0__1_.mux_right_track_30.sky130_fd_sc_hd__mux2_1_0_X
rlabel metal1 13386 24718 13386 24718 0 sb_0__1_.mux_right_track_30.sky130_fd_sc_hd__mux2_1_1_X
rlabel metal1 16146 19890 16146 19890 0 sb_0__1_.mux_right_track_30.sky130_fd_sc_hd__mux2_1_2_X
rlabel metal2 21942 14790 21942 14790 0 sb_0__1_.mux_right_track_32.out
rlabel metal1 14674 23154 14674 23154 0 sb_0__1_.mux_right_track_32.sky130_fd_sc_hd__mux2_1_0_X
rlabel metal1 13570 22984 13570 22984 0 sb_0__1_.mux_right_track_32.sky130_fd_sc_hd__mux2_1_1_X
rlabel metal1 17434 19346 17434 19346 0 sb_0__1_.mux_right_track_32.sky130_fd_sc_hd__mux2_1_2_X
rlabel metal2 21114 15198 21114 15198 0 sb_0__1_.mux_right_track_34.out
rlabel metal1 16514 21862 16514 21862 0 sb_0__1_.mux_right_track_34.sky130_fd_sc_hd__mux2_1_0_X
rlabel metal1 12466 21896 12466 21896 0 sb_0__1_.mux_right_track_34.sky130_fd_sc_hd__mux2_1_1_X
rlabel metal2 15962 21165 15962 21165 0 sb_0__1_.mux_right_track_34.sky130_fd_sc_hd__mux2_1_2_X
rlabel metal2 21758 11220 21758 11220 0 sb_0__1_.mux_right_track_36.out
rlabel metal2 9154 18887 9154 18887 0 sb_0__1_.mux_right_track_36.sky130_fd_sc_hd__mux2_1_0_X
rlabel metal1 9614 17034 9614 17034 0 sb_0__1_.mux_right_track_36.sky130_fd_sc_hd__mux2_1_1_X
rlabel metal2 7130 11186 7130 11186 0 sb_0__1_.mux_right_track_36.sky130_fd_sc_hd__mux2_1_2_X
rlabel metal1 16721 11118 16721 11118 0 sb_0__1_.mux_right_track_36.sky130_fd_sc_hd__mux2_1_3_X
rlabel metal1 21666 9554 21666 9554 0 sb_0__1_.mux_right_track_38.out
rlabel metal1 14076 13974 14076 13974 0 sb_0__1_.mux_right_track_38.sky130_fd_sc_hd__mux2_1_0_X
rlabel metal1 17526 11560 17526 11560 0 sb_0__1_.mux_right_track_38.sky130_fd_sc_hd__mux2_1_1_X
rlabel metal1 24702 25262 24702 25262 0 sb_0__1_.mux_right_track_4.out
rlabel metal1 22770 38386 22770 38386 0 sb_0__1_.mux_right_track_4.sky130_fd_sc_hd__mux2_1_0_X
rlabel metal2 22034 38114 22034 38114 0 sb_0__1_.mux_right_track_4.sky130_fd_sc_hd__mux2_1_1_X
rlabel metal1 22908 34034 22908 34034 0 sb_0__1_.mux_right_track_4.sky130_fd_sc_hd__mux2_1_2_X
rlabel metal2 20562 33762 20562 33762 0 sb_0__1_.mux_right_track_4.sky130_fd_sc_hd__mux2_1_3_X
rlabel metal1 23184 33830 23184 33830 0 sb_0__1_.mux_right_track_4.sky130_fd_sc_hd__mux2_1_4_X
rlabel metal1 23414 11152 23414 11152 0 sb_0__1_.mux_right_track_40.out
rlabel metal1 16606 13362 16606 13362 0 sb_0__1_.mux_right_track_40.sky130_fd_sc_hd__mux2_1_0_X
rlabel metal1 18400 11254 18400 11254 0 sb_0__1_.mux_right_track_40.sky130_fd_sc_hd__mux2_1_1_X
rlabel metal1 23414 9588 23414 9588 0 sb_0__1_.mux_right_track_44.out
rlabel metal1 17296 15130 17296 15130 0 sb_0__1_.mux_right_track_44.sky130_fd_sc_hd__mux2_1_0_X
rlabel metal1 21942 12206 21942 12206 0 sb_0__1_.mux_right_track_44.sky130_fd_sc_hd__mux2_1_1_X
rlabel metal2 24886 10642 24886 10642 0 sb_0__1_.mux_right_track_46.out
rlabel metal1 20608 16218 20608 16218 0 sb_0__1_.mux_right_track_46.sky130_fd_sc_hd__mux2_1_0_X
rlabel metal1 22862 12240 22862 12240 0 sb_0__1_.mux_right_track_46.sky130_fd_sc_hd__mux2_1_1_X
rlabel metal1 23598 8942 23598 8942 0 sb_0__1_.mux_right_track_48.out
rlabel metal1 22494 15980 22494 15980 0 sb_0__1_.mux_right_track_48.sky130_fd_sc_hd__mux2_1_0_X
rlabel metal2 23506 14042 23506 14042 0 sb_0__1_.mux_right_track_48.sky130_fd_sc_hd__mux2_1_1_X
rlabel metal1 23874 10030 23874 10030 0 sb_0__1_.mux_right_track_50.out
rlabel metal1 21436 26486 21436 26486 0 sb_0__1_.mux_right_track_50.sky130_fd_sc_hd__mux2_1_0_X
rlabel metal2 19182 17442 19182 17442 0 sb_0__1_.mux_right_track_50.sky130_fd_sc_hd__mux2_1_1_X
rlabel metal2 22448 17612 22448 17612 0 sb_0__1_.mux_right_track_50.sky130_fd_sc_hd__mux2_1_2_X
rlabel metal1 22908 4658 22908 4658 0 sb_0__1_.mux_right_track_52.out
rlabel metal2 21206 14280 21206 14280 0 sb_0__1_.mux_right_track_52.sky130_fd_sc_hd__mux2_1_0_X
rlabel metal1 21850 10642 21850 10642 0 sb_0__1_.mux_right_track_52.sky130_fd_sc_hd__mux2_1_1_X
rlabel metal1 23092 7718 23092 7718 0 sb_0__1_.mux_right_track_54.out
rlabel metal1 18676 13498 18676 13498 0 sb_0__1_.mux_right_track_54.sky130_fd_sc_hd__mux2_1_0_X
rlabel metal1 21436 7854 21436 7854 0 sb_0__1_.mux_right_track_54.sky130_fd_sc_hd__mux2_1_1_X
rlabel metal1 23276 5610 23276 5610 0 sb_0__1_.mux_right_track_56.out
rlabel metal2 20562 14688 20562 14688 0 sb_0__1_.mux_right_track_56.sky130_fd_sc_hd__mux2_1_0_X
rlabel metal1 22080 10030 22080 10030 0 sb_0__1_.mux_right_track_56.sky130_fd_sc_hd__mux2_1_1_X
rlabel metal1 24518 27030 24518 27030 0 sb_0__1_.mux_right_track_6.out
rlabel metal1 25254 38318 25254 38318 0 sb_0__1_.mux_right_track_6.sky130_fd_sc_hd__mux2_1_0_X
rlabel metal1 21574 37128 21574 37128 0 sb_0__1_.mux_right_track_6.sky130_fd_sc_hd__mux2_1_1_X
rlabel metal2 22494 34340 22494 34340 0 sb_0__1_.mux_right_track_6.sky130_fd_sc_hd__mux2_1_2_X
rlabel metal1 23828 36142 23828 36142 0 sb_0__1_.mux_right_track_6.sky130_fd_sc_hd__mux2_1_3_X
rlabel metal2 23690 35734 23690 35734 0 sb_0__1_.mux_right_track_6.sky130_fd_sc_hd__mux2_1_4_X
rlabel metal1 23920 36278 23920 36278 0 sb_0__1_.mux_right_track_6.sky130_fd_sc_hd__mux2_1_5_X
rlabel metal1 24242 34510 24242 34510 0 sb_0__1_.mux_right_track_8.out
rlabel metal1 22540 42602 22540 42602 0 sb_0__1_.mux_right_track_8.sky130_fd_sc_hd__mux2_1_0_X
rlabel metal1 21574 40698 21574 40698 0 sb_0__1_.mux_right_track_8.sky130_fd_sc_hd__mux2_1_1_X
rlabel metal1 21298 41514 21298 41514 0 sb_0__1_.mux_right_track_8.sky130_fd_sc_hd__mux2_1_2_X
rlabel metal1 22264 40562 22264 40562 0 sb_0__1_.mux_right_track_8.sky130_fd_sc_hd__mux2_1_3_X
rlabel metal2 22862 40947 22862 40947 0 sb_0__1_.mux_right_track_8.sky130_fd_sc_hd__mux2_1_4_X
rlabel metal1 23782 34578 23782 34578 0 sb_0__1_.mux_right_track_8.sky130_fd_sc_hd__mux2_1_5_X
rlabel metal1 12282 51986 12282 51986 0 sb_0__1_.mux_top_track_0.out
rlabel metal1 9798 43418 9798 43418 0 sb_0__1_.mux_top_track_0.sky130_fd_sc_hd__mux2_1_0_X
rlabel metal1 17158 42296 17158 42296 0 sb_0__1_.mux_top_track_0.sky130_fd_sc_hd__mux2_1_1_X
rlabel metal1 14720 37094 14720 37094 0 sb_0__1_.mux_top_track_0.sky130_fd_sc_hd__mux2_1_2_X
rlabel metal1 9982 37298 9982 37298 0 sb_0__1_.mux_top_track_0.sky130_fd_sc_hd__mux2_1_3_X
rlabel metal1 11546 44506 11546 44506 0 sb_0__1_.mux_top_track_0.sky130_fd_sc_hd__mux2_1_4_X
rlabel metal2 11546 43860 11546 43860 0 sb_0__1_.mux_top_track_0.sky130_fd_sc_hd__mux2_1_5_X
rlabel metal2 10718 47668 10718 47668 0 sb_0__1_.mux_top_track_0.sky130_fd_sc_hd__mux2_1_6_X
rlabel metal1 8924 45050 8924 45050 0 sb_0__1_.mux_top_track_10.out
rlabel metal2 9706 39270 9706 39270 0 sb_0__1_.mux_top_track_10.sky130_fd_sc_hd__mux2_1_0_X
rlabel metal2 17342 36856 17342 36856 0 sb_0__1_.mux_top_track_10.sky130_fd_sc_hd__mux2_1_1_X
rlabel metal1 9430 33830 9430 33830 0 sb_0__1_.mux_top_track_10.sky130_fd_sc_hd__mux2_1_2_X
rlabel metal1 7866 33830 7866 33830 0 sb_0__1_.mux_top_track_10.sky130_fd_sc_hd__mux2_1_3_X
rlabel metal1 8694 38182 8694 38182 0 sb_0__1_.mux_top_track_10.sky130_fd_sc_hd__mux2_1_4_X
rlabel metal2 7866 36176 7866 36176 0 sb_0__1_.mux_top_track_10.sky130_fd_sc_hd__mux2_1_5_X
rlabel metal1 7636 38522 7636 38522 0 sb_0__1_.mux_top_track_10.sky130_fd_sc_hd__mux2_1_6_X
rlabel metal1 7820 43418 7820 43418 0 sb_0__1_.mux_top_track_12.out
rlabel metal1 12489 37094 12489 37094 0 sb_0__1_.mux_top_track_12.sky130_fd_sc_hd__mux2_1_0_X
rlabel metal2 16330 33983 16330 33983 0 sb_0__1_.mux_top_track_12.sky130_fd_sc_hd__mux2_1_1_X
rlabel metal1 7912 32810 7912 32810 0 sb_0__1_.mux_top_track_12.sky130_fd_sc_hd__mux2_1_2_X
rlabel metal2 10258 35088 10258 35088 0 sb_0__1_.mux_top_track_12.sky130_fd_sc_hd__mux2_1_3_X
rlabel metal2 7590 34544 7590 34544 0 sb_0__1_.mux_top_track_12.sky130_fd_sc_hd__mux2_1_4_X
rlabel metal1 7728 36346 7728 36346 0 sb_0__1_.mux_top_track_12.sky130_fd_sc_hd__mux2_1_5_X
rlabel metal1 12788 49402 12788 49402 0 sb_0__1_.mux_top_track_2.out
rlabel metal2 16974 42704 16974 42704 0 sb_0__1_.mux_top_track_2.sky130_fd_sc_hd__mux2_1_0_X
rlabel metal1 19090 42126 19090 42126 0 sb_0__1_.mux_top_track_2.sky130_fd_sc_hd__mux2_1_1_X
rlabel metal1 13432 42262 13432 42262 0 sb_0__1_.mux_top_track_2.sky130_fd_sc_hd__mux2_1_2_X
rlabel metal2 15318 43792 15318 43792 0 sb_0__1_.mux_top_track_2.sky130_fd_sc_hd__mux2_1_3_X
rlabel metal1 13248 42330 13248 42330 0 sb_0__1_.mux_top_track_2.sky130_fd_sc_hd__mux2_1_4_X
rlabel metal1 13340 45322 13340 45322 0 sb_0__1_.mux_top_track_2.sky130_fd_sc_hd__mux2_1_5_X
rlabel metal2 8418 47124 8418 47124 0 sb_0__1_.mux_top_track_20.out
rlabel metal1 13294 35156 13294 35156 0 sb_0__1_.mux_top_track_20.sky130_fd_sc_hd__mux2_1_0_X
rlabel metal1 14076 34918 14076 34918 0 sb_0__1_.mux_top_track_20.sky130_fd_sc_hd__mux2_1_1_X
rlabel metal1 9844 32742 9844 32742 0 sb_0__1_.mux_top_track_20.sky130_fd_sc_hd__mux2_1_2_X
rlabel metal2 11362 36550 11362 36550 0 sb_0__1_.mux_top_track_20.sky130_fd_sc_hd__mux2_1_3_X
rlabel metal2 9430 35462 9430 35462 0 sb_0__1_.mux_top_track_20.sky130_fd_sc_hd__mux2_1_4_X
rlabel metal1 9246 37978 9246 37978 0 sb_0__1_.mux_top_track_20.sky130_fd_sc_hd__mux2_1_5_X
rlabel metal2 5842 47396 5842 47396 0 sb_0__1_.mux_top_track_28.out
rlabel metal2 12558 36924 12558 36924 0 sb_0__1_.mux_top_track_28.sky130_fd_sc_hd__mux2_1_0_X
rlabel metal1 12742 33626 12742 33626 0 sb_0__1_.mux_top_track_28.sky130_fd_sc_hd__mux2_1_1_X
rlabel metal1 9062 36346 9062 36346 0 sb_0__1_.mux_top_track_28.sky130_fd_sc_hd__mux2_1_2_X
rlabel metal1 5336 32538 5336 32538 0 sb_0__1_.mux_top_track_28.sky130_fd_sc_hd__mux2_1_3_X
rlabel metal1 6302 44370 6302 44370 0 sb_0__1_.mux_top_track_28.sky130_fd_sc_hd__mux2_1_4_X
rlabel metal1 7406 46682 7406 46682 0 sb_0__1_.mux_top_track_36.out
rlabel metal1 12696 39066 12696 39066 0 sb_0__1_.mux_top_track_36.sky130_fd_sc_hd__mux2_1_0_X
rlabel metal1 12236 39066 12236 39066 0 sb_0__1_.mux_top_track_36.sky130_fd_sc_hd__mux2_1_1_X
rlabel metal1 9660 38794 9660 38794 0 sb_0__1_.mux_top_track_36.sky130_fd_sc_hd__mux2_1_2_X
rlabel metal1 9660 42330 9660 42330 0 sb_0__1_.mux_top_track_36.sky130_fd_sc_hd__mux2_1_3_X
rlabel metal1 11822 46682 11822 46682 0 sb_0__1_.mux_top_track_4.out
rlabel metal1 15272 41446 15272 41446 0 sb_0__1_.mux_top_track_4.sky130_fd_sc_hd__mux2_1_0_X
rlabel metal1 17250 36278 17250 36278 0 sb_0__1_.mux_top_track_4.sky130_fd_sc_hd__mux2_1_1_X
rlabel metal2 10902 35972 10902 35972 0 sb_0__1_.mux_top_track_4.sky130_fd_sc_hd__mux2_1_2_X
rlabel metal1 13064 40698 13064 40698 0 sb_0__1_.mux_top_track_4.sky130_fd_sc_hd__mux2_1_3_X
rlabel metal1 10580 39066 10580 39066 0 sb_0__1_.mux_top_track_4.sky130_fd_sc_hd__mux2_1_4_X
rlabel metal1 10488 41446 10488 41446 0 sb_0__1_.mux_top_track_4.sky130_fd_sc_hd__mux2_1_5_X
rlabel metal1 8096 52054 8096 52054 0 sb_0__1_.mux_top_track_44.out
rlabel metal1 15364 40154 15364 40154 0 sb_0__1_.mux_top_track_44.sky130_fd_sc_hd__mux2_1_0_X
rlabel metal1 10488 38522 10488 38522 0 sb_0__1_.mux_top_track_44.sky130_fd_sc_hd__mux2_1_1_X
rlabel metal2 11730 44982 11730 44982 0 sb_0__1_.mux_top_track_44.sky130_fd_sc_hd__mux2_1_2_X
rlabel metal1 8878 46070 8878 46070 0 sb_0__1_.mux_top_track_52.out
rlabel metal1 20194 39406 20194 39406 0 sb_0__1_.mux_top_track_52.sky130_fd_sc_hd__mux2_1_0_X
rlabel metal1 17802 39338 17802 39338 0 sb_0__1_.mux_top_track_52.sky130_fd_sc_hd__mux2_1_1_X
rlabel metal1 14766 36346 14766 36346 0 sb_0__1_.mux_top_track_52.sky130_fd_sc_hd__mux2_1_2_X
rlabel metal1 13432 45526 13432 45526 0 sb_0__1_.mux_top_track_52.sky130_fd_sc_hd__mux2_1_3_X
rlabel metal1 9890 51374 9890 51374 0 sb_0__1_.mux_top_track_6.out
rlabel metal1 9706 39474 9706 39474 0 sb_0__1_.mux_top_track_6.sky130_fd_sc_hd__mux2_1_0_X
rlabel metal1 17066 38522 17066 38522 0 sb_0__1_.mux_top_track_6.sky130_fd_sc_hd__mux2_1_1_X
rlabel metal2 11270 33728 11270 33728 0 sb_0__1_.mux_top_track_6.sky130_fd_sc_hd__mux2_1_2_X
rlabel metal1 7590 34918 7590 34918 0 sb_0__1_.mux_top_track_6.sky130_fd_sc_hd__mux2_1_3_X
rlabel metal1 9200 39610 9200 39610 0 sb_0__1_.mux_top_track_6.sky130_fd_sc_hd__mux2_1_4_X
rlabel metal1 9016 35258 9016 35258 0 sb_0__1_.mux_top_track_6.sky130_fd_sc_hd__mux2_1_5_X
rlabel metal1 7268 40154 7268 40154 0 sb_0__1_.mux_top_track_6.sky130_fd_sc_hd__mux2_1_6_X
rlabel metal1 12926 37162 12926 37162 0 top_left_grid_right_width_0_height_0_subtile_0__pin_inpad_0_
rlabel metal1 16997 43214 16997 43214 0 top_left_grid_right_width_0_height_0_subtile_1__pin_inpad_0_
rlabel metal3 1211 50524 1211 50524 0 top_left_grid_right_width_0_height_0_subtile_2__pin_inpad_0_
rlabel metal3 2062 52972 2062 52972 0 top_left_grid_right_width_0_height_0_subtile_3__pin_inpad_0_
<< properties >>
string FIXED_BBOX 0 0 27000 57000
<< end >>
