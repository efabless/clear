* NGSPICE file created from sb_1__2_.ext - technology: sky130A

* Black-box entry subcircuit for sky130_fd_sc_hd__tapvpwrvgnd_1 abstract view
.subckt sky130_fd_sc_hd__tapvpwrvgnd_1 VGND VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__diode_2 abstract view
.subckt sky130_fd_sc_hd__diode_2 DIODE VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__fill_2 abstract view
.subckt sky130_fd_sc_hd__fill_2 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dfxtp_1 abstract view
.subckt sky130_fd_sc_hd__dfxtp_1 CLK D VGND VNB VPB VPWR Q
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__mux2_1 abstract view
.subckt sky130_fd_sc_hd__mux2_1 A0 A1 S VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dfxtp_2 abstract view
.subckt sky130_fd_sc_hd__dfxtp_2 CLK D VGND VNB VPB VPWR Q
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__fill_1 abstract view
.subckt sky130_fd_sc_hd__fill_1 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_4 abstract view
.subckt sky130_fd_sc_hd__decap_4 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_3 abstract view
.subckt sky130_fd_sc_hd__decap_3 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_1 abstract view
.subckt sky130_fd_sc_hd__clkbuf_1 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__conb_1 abstract view
.subckt sky130_fd_sc_hd__conb_1 VGND VNB VPB VPWR HI LO
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__buf_2 abstract view
.subckt sky130_fd_sc_hd__buf_2 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__buf_6 abstract view
.subckt sky130_fd_sc_hd__buf_6 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__buf_8 abstract view
.subckt sky130_fd_sc_hd__buf_8 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_2 abstract view
.subckt sky130_fd_sc_hd__clkbuf_2 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dlymetal6s2s_1 abstract view
.subckt sky130_fd_sc_hd__dlymetal6s2s_1 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_8 abstract view
.subckt sky130_fd_sc_hd__decap_8 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_6 abstract view
.subckt sky130_fd_sc_hd__decap_6 VGND VNB VPB VPWR
.ends

.subckt sb_1__2_ SC_IN_BOT SC_OUT_BOT VGND VPWR bottom_left_grid_pin_42_ bottom_left_grid_pin_43_
+ bottom_left_grid_pin_44_ bottom_left_grid_pin_45_ bottom_left_grid_pin_46_ bottom_left_grid_pin_47_
+ bottom_left_grid_pin_48_ bottom_left_grid_pin_49_ ccff_head ccff_tail chanx_left_in[0]
+ chanx_left_in[10] chanx_left_in[11] chanx_left_in[12] chanx_left_in[13] chanx_left_in[14]
+ chanx_left_in[15] chanx_left_in[16] chanx_left_in[17] chanx_left_in[18] chanx_left_in[19]
+ chanx_left_in[1] chanx_left_in[2] chanx_left_in[3] chanx_left_in[4] chanx_left_in[5]
+ chanx_left_in[6] chanx_left_in[7] chanx_left_in[8] chanx_left_in[9] chanx_left_out[0]
+ chanx_left_out[10] chanx_left_out[11] chanx_left_out[12] chanx_left_out[13] chanx_left_out[14]
+ chanx_left_out[15] chanx_left_out[16] chanx_left_out[17] chanx_left_out[18] chanx_left_out[19]
+ chanx_left_out[1] chanx_left_out[2] chanx_left_out[3] chanx_left_out[4] chanx_left_out[5]
+ chanx_left_out[6] chanx_left_out[7] chanx_left_out[8] chanx_left_out[9] chanx_right_in[0]
+ chanx_right_in[10] chanx_right_in[11] chanx_right_in[12] chanx_right_in[13] chanx_right_in[14]
+ chanx_right_in[15] chanx_right_in[16] chanx_right_in[17] chanx_right_in[18] chanx_right_in[19]
+ chanx_right_in[1] chanx_right_in[2] chanx_right_in[3] chanx_right_in[4] chanx_right_in[5]
+ chanx_right_in[6] chanx_right_in[7] chanx_right_in[8] chanx_right_in[9] chanx_right_out[0]
+ chanx_right_out[10] chanx_right_out[11] chanx_right_out[12] chanx_right_out[13]
+ chanx_right_out[14] chanx_right_out[15] chanx_right_out[16] chanx_right_out[17]
+ chanx_right_out[18] chanx_right_out[19] chanx_right_out[1] chanx_right_out[2] chanx_right_out[3]
+ chanx_right_out[4] chanx_right_out[5] chanx_right_out[6] chanx_right_out[7] chanx_right_out[8]
+ chanx_right_out[9] chany_bottom_in[0] chany_bottom_in[10] chany_bottom_in[11] chany_bottom_in[12]
+ chany_bottom_in[13] chany_bottom_in[14] chany_bottom_in[15] chany_bottom_in[16]
+ chany_bottom_in[17] chany_bottom_in[18] chany_bottom_in[19] chany_bottom_in[1] chany_bottom_in[2]
+ chany_bottom_in[3] chany_bottom_in[4] chany_bottom_in[5] chany_bottom_in[6] chany_bottom_in[7]
+ chany_bottom_in[8] chany_bottom_in[9] chany_bottom_out[0] chany_bottom_out[10] chany_bottom_out[11]
+ chany_bottom_out[12] chany_bottom_out[13] chany_bottom_out[14] chany_bottom_out[15]
+ chany_bottom_out[16] chany_bottom_out[17] chany_bottom_out[18] chany_bottom_out[19]
+ chany_bottom_out[1] chany_bottom_out[2] chany_bottom_out[3] chany_bottom_out[4]
+ chany_bottom_out[5] chany_bottom_out[6] chany_bottom_out[7] chany_bottom_out[8]
+ chany_bottom_out[9] left_bottom_grid_pin_34_ left_bottom_grid_pin_35_ left_bottom_grid_pin_36_
+ left_bottom_grid_pin_37_ left_bottom_grid_pin_38_ left_bottom_grid_pin_39_ left_bottom_grid_pin_40_
+ left_bottom_grid_pin_41_ left_top_grid_pin_1_ prog_clk_0_S_in right_bottom_grid_pin_34_
+ right_bottom_grid_pin_35_ right_bottom_grid_pin_36_ right_bottom_grid_pin_37_ right_bottom_grid_pin_38_
+ right_bottom_grid_pin_39_ right_bottom_grid_pin_40_ right_bottom_grid_pin_41_ right_top_grid_pin_1_
XTAP_188 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_177 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_mem_right_track_0.sky130_fd_sc_hd__dfxtp_1_0__CLK prog_clk_0_FTB00/X VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_7_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmem_right_track_2.sky130_fd_sc_hd__dfxtp_1_0_ prog_clk_0_FTB00/X mux_right_track_0.mux_l4_in_0_/S
+ VGND VGND VPWR VPWR mux_right_track_2.mux_l1_in_1_/S sky130_fd_sc_hd__dfxtp_1
XFILLER_9_115 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_9_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_13_155 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_13_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmux_bottom_track_3.mux_l1_in_1_ input7/X input5/X mux_bottom_track_3.mux_l1_in_3_/S
+ VGND VGND VPWR VPWR mux_bottom_track_3.mux_l1_in_1_/X sky130_fd_sc_hd__mux2_1
XFILLER_3_67 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmem_left_track_17.sky130_fd_sc_hd__dfxtp_1_0_ prog_clk_0_FTB00/X mux_left_track_9.mux_l4_in_0_/S
+ VGND VGND VPWR VPWR mux_left_track_17.mux_l1_in_3_/S sky130_fd_sc_hd__dfxtp_2
XANTENNA_mux_bottom_track_11.mux_l1_in_0__A0 input3/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_10_114 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_12_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_12_76 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_12_87 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_5_151 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_5_140 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_mem_left_track_9.sky130_fd_sc_hd__dfxtp_1_0__CLK prog_clk_0_FTB00/X VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_062_ _062_/A VGND VGND VPWR VPWR _062_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_23_31 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_input55_A chany_bottom_in[13] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_2_187 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xmem_right_track_8.sky130_fd_sc_hd__dfxtp_1_1_ prog_clk_0_FTB00/X mux_right_track_8.mux_l1_in_0_/S
+ VGND VGND VPWR VPWR mux_right_track_8.mux_l2_in_3_/S sky130_fd_sc_hd__dfxtp_2
XFILLER_9_66 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_mem_bottom_track_27.sky130_fd_sc_hd__dfxtp_1_0__CLK prog_clk_0_FTB00/X VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_18_42 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_114_ _114_/A VGND VGND VPWR VPWR _114_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_22_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmem_bottom_track_25.sky130_fd_sc_hd__dfxtp_1_2_ prog_clk_0_FTB00/X mux_bottom_track_25.mux_l2_in_1_/S
+ VGND VGND VPWR VPWR mux_bottom_track_25.mux_l3_in_0_/S sky130_fd_sc_hd__dfxtp_1
XFILLER_29_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_29_128 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_29_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xmux_bottom_track_17.mux_l1_in_0_ input6/X _071_/A mux_bottom_track_17.mux_l1_in_1_/S
+ VGND VGND VPWR VPWR mux_bottom_track_17.mux_l1_in_0_/X sky130_fd_sc_hd__mux2_1
XANTENNA_mux_left_track_17.mux_l2_in_0__S mux_left_track_17.mux_l2_in_1_/S VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_4_205 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_20_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_29_52 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_29_30 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_28_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_input18_A chanx_left_in[16] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xmux_right_track_32.mux_l2_in_1__169 VGND VGND VPWR VPWR mux_right_track_32.mux_l2_in_1_/A0
+ mux_right_track_32.mux_l2_in_1__169/LO sky130_fd_sc_hd__conb_1
XFILLER_25_131 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_mem_bottom_track_19.sky130_fd_sc_hd__dfxtp_1_1__CLK prog_clk_0_FTB00/X VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_25_186 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_15_43 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_15_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_31_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_31_86 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xoutput97 _072_/X VGND VGND VPWR VPWR chanx_left_out[15] sky130_fd_sc_hd__buf_2
Xmux_bottom_track_3.sky130_fd_sc_hd__buf_4_0_ mux_bottom_track_3.mux_l3_in_0_/X VGND
+ VGND VPWR VPWR _098_/A sky130_fd_sc_hd__clkbuf_1
XANTENNA_mux_bottom_track_3.mux_l1_in_1__A0 input7/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_31_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_16_131 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_16_164 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_31_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_189 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_178 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_167 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_101 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_112 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_123 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_134 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_145 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_156 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_mem_right_track_24.sky130_fd_sc_hd__dfxtp_1_0__CLK prog_clk_0_FTB00/X VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mux_left_track_9.mux_l2_in_2__A0 input74/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mux_right_track_0.mux_l2_in_3__A1 _090_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_26_75 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_26_64 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_26_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_9_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_input85_A right_bottom_grid_pin_39_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xmux_bottom_track_3.mux_l1_in_0_ input3/X _062_/A mux_bottom_track_3.mux_l1_in_3_/S
+ VGND VGND VPWR VPWR mux_bottom_track_3.mux_l1_in_0_/X sky130_fd_sc_hd__mux2_1
XFILLER_3_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_3_24 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_3_13 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_mux_bottom_track_11.mux_l1_in_0__A1 _067_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_27_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_18_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_5_196 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_5_185 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_mem_right_track_16.sky130_fd_sc_hd__dfxtp_1_1__CLK prog_clk_0_FTB00/X VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mem_bottom_track_3.sky130_fd_sc_hd__dfxtp_1_1__CLK prog_clk_0_FTB00/X VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_23_43 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_23_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_061_ _061_/A VGND VGND VPWR VPWR _061_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_2_144 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_input48_A chanx_right_in[7] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xmem_right_track_8.sky130_fd_sc_hd__dfxtp_1_0_ prog_clk_0_FTB00/X mux_right_track_4.mux_l4_in_0_/S
+ VGND VGND VPWR VPWR mux_right_track_8.mux_l1_in_0_/S sky130_fd_sc_hd__dfxtp_1
Xmux_bottom_track_17.mux_l1_in_1__176 VGND VGND VPWR VPWR mux_bottom_track_17.mux_l1_in_1_/A0
+ mux_bottom_track_17.mux_l1_in_1__176/LO sky130_fd_sc_hd__conb_1
Xmux_left_track_9.sky130_fd_sc_hd__buf_4_0_ mux_left_track_9.mux_l4_in_0_/X VGND VGND
+ VPWR VPWR _061_/A sky130_fd_sc_hd__clkbuf_1
XANTENNA_mux_left_track_1.mux_l2_in_2__S mux_left_track_1.mux_l2_in_3_/S VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
X_113_ _113_/A VGND VGND VPWR VPWR _113_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_11_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmux_right_track_24.mux_l1_in_3__168 VGND VGND VPWR VPWR mux_right_track_24.mux_l1_in_3_/A0
+ mux_right_track_24.mux_l1_in_3__168/LO sky130_fd_sc_hd__conb_1
XANTENNA_mux_left_track_5.mux_l3_in_0__S mux_left_track_5.mux_l3_in_1_/S VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
Xmem_bottom_track_25.sky130_fd_sc_hd__dfxtp_1_1_ prog_clk_0_FTB00/X mux_bottom_track_25.mux_l1_in_0_/S
+ VGND VGND VPWR VPWR mux_bottom_track_25.mux_l2_in_1_/S sky130_fd_sc_hd__dfxtp_1
XFILLER_4_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_6_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_19_140 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_25_176 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_15_33 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_31_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_15_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xoutput98 _073_/X VGND VGND VPWR VPWR chanx_left_out[16] sky130_fd_sc_hd__buf_2
Xmux_right_track_8.mux_l2_in_3_ mux_right_track_8.mux_l2_in_3_/A0 _094_/A mux_right_track_8.mux_l2_in_3_/S
+ VGND VGND VPWR VPWR mux_right_track_8.mux_l2_in_3_/X sky130_fd_sc_hd__mux2_1
XANTENNA_input30_A chanx_left_in[9] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_179 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_168 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xmux_left_track_25.sky130_fd_sc_hd__buf_4_0_ mux_left_track_25.mux_l3_in_0_/X VGND
+ VGND VPWR VPWR _069_/A sky130_fd_sc_hd__clkbuf_1
XTAP_102 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_113 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_124 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_135 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_146 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_157 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_22_102 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmem_bottom_track_3.sky130_fd_sc_hd__dfxtp_1_2_ prog_clk_0_FTB00/X mux_bottom_track_3.mux_l2_in_1_/S
+ VGND VGND VPWR VPWR mem_bottom_track_5.delay_buf_2/X sky130_fd_sc_hd__dfxtp_1
XFILLER_22_157 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_26_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_26_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_13_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_input78_A left_bottom_grid_pin_41_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mux_left_track_33.mux_l1_in_1__S mux_left_track_33.mux_l1_in_2_/S VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_21_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_mux_right_track_32.mux_l2_in_1__S mux_right_track_32.mux_l2_in_1_/S VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mux_bottom_track_1.mux_l1_in_3__A1 _080_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_8_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmux_left_track_17.mux_l1_in_3__159 VGND VGND VPWR VPWR mux_left_track_17.mux_l1_in_3_/A0
+ mux_left_track_17.mux_l1_in_3__159/LO sky130_fd_sc_hd__conb_1
XFILLER_10_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_10_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmux_bottom_track_21.mux_l1_in_1__178 VGND VGND VPWR VPWR mux_bottom_track_21.mux_l1_in_1_/A0
+ mux_bottom_track_21.mux_l1_in_1__178/LO sky130_fd_sc_hd__conb_1
Xmux_right_track_8.mux_l4_in_0_ mux_right_track_8.mux_l3_in_1_/X mux_right_track_8.mux_l3_in_0_/X
+ mux_right_track_8.mux_l4_in_0_/S VGND VGND VPWR VPWR mux_right_track_8.mux_l4_in_0_/X
+ sky130_fd_sc_hd__mux2_1
XFILLER_23_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_3_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_060_ _060_/A VGND VGND VPWR VPWR _060_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_0_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_mem_left_track_3.sky130_fd_sc_hd__dfxtp_1_1__CLK prog_clk_0_FTB00/X VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_9_79 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_20_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_18_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_112_ _112_/A VGND VGND VPWR VPWR _112_/X sky130_fd_sc_hd__clkbuf_1
XANTENNA_input60_A chany_bottom_in[18] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xmux_right_track_8.mux_l3_in_1_ mux_right_track_8.mux_l2_in_3_/X mux_right_track_8.mux_l2_in_2_/X
+ mux_right_track_8.mux_l3_in_1_/S VGND VGND VPWR VPWR mux_right_track_8.mux_l3_in_1_/X
+ sky130_fd_sc_hd__mux2_1
Xmem_bottom_track_25.sky130_fd_sc_hd__dfxtp_1_0_ prog_clk_0_FTB00/X mux_bottom_track_23.mux_l2_in_0_/S
+ VGND VGND VPWR VPWR mux_bottom_track_25.mux_l1_in_0_/S sky130_fd_sc_hd__dfxtp_1
XANTENNA_mem_right_track_0.sky130_fd_sc_hd__dfxtp_1_3__CLK prog_clk_0_FTB00/X VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_28_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_mem_bottom_track_21.sky130_fd_sc_hd__dfxtp_1_1__CLK prog_clk_0_FTB00/X VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_28_185 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xmem_left_track_25.delay_buf_2 mem_left_track_25.delay_buf_2/X VGND VGND VPWR VPWR
+ mem_left_track_25.delay_buf_2/X sky130_fd_sc_hd__buf_6
XFILLER_6_58 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_13_5 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_25_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_25_144 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_25_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_31_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_31_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_31_22 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xoutput99 _074_/X VGND VGND VPWR VPWR chanx_left_out[17] sky130_fd_sc_hd__buf_2
XFILLER_0_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmux_right_track_8.mux_l2_in_2_ _084_/A input58/X mux_right_track_8.mux_l2_in_3_/S
+ VGND VGND VPWR VPWR mux_right_track_8.mux_l2_in_2_/X sky130_fd_sc_hd__mux2_1
XANTENNA_input23_A chanx_left_in[2] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_16_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_31_158 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_31_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_16_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_103 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_114 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_mem_left_track_9.sky130_fd_sc_hd__dfxtp_1_3__CLK prog_clk_0_FTB00/X VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_169 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_125 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_136 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_147 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_158 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xmem_bottom_track_3.sky130_fd_sc_hd__dfxtp_1_1_ prog_clk_0_FTB00/X mux_bottom_track_3.mux_l1_in_3_/S
+ VGND VGND VPWR VPWR mux_bottom_track_3.mux_l2_in_1_/S sky130_fd_sc_hd__dfxtp_1
XFILLER_9_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_13_136 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_mem_right_track_4.sky130_fd_sc_hd__dfxtp_1_0__CLK prog_clk_0_FTB00/X VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_10_106 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_10_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__064__A _064_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_5_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_12_13 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_33_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_24_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_mem_right_track_32.sky130_fd_sc_hd__dfxtp_1_2__CLK prog_clk_0_FTB00/X VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_4_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_mux_bottom_track_7.mux_l1_in_0__A0 input3/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_23_12 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_23_23 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_23_89 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_2_102 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xprog_clk_0_FTB00 prog_clk_0_S_in VGND VGND VPWR VPWR prog_clk_0_FTB00/X sky130_fd_sc_hd__buf_8
Xmem_bottom_track_9.sky130_fd_sc_hd__dfxtp_1_2_ prog_clk_0_FTB00/X mux_bottom_track_9.mux_l2_in_1_/S
+ VGND VGND VPWR VPWR mux_bottom_track_9.mux_l3_in_0_/S sky130_fd_sc_hd__dfxtp_1
XFILLER_9_14 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_9_25 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_9_36 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_9_47 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_111_ _111_/A VGND VGND VPWR VPWR _111_/X sky130_fd_sc_hd__clkbuf_1
XANTENNA_mux_bottom_track_5.mux_l1_in_2__A0 _083_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_input53_A chany_bottom_in[11] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xmux_right_track_8.mux_l3_in_0_ mux_right_track_8.mux_l2_in_1_/X mux_right_track_8.mux_l2_in_0_/X
+ mux_right_track_8.mux_l3_in_1_/S VGND VGND VPWR VPWR mux_right_track_8.mux_l3_in_0_/X
+ sky130_fd_sc_hd__mux2_1
XANTENNA_mem_left_track_25.sky130_fd_sc_hd__dfxtp_1_0__CLK prog_clk_0_FTB00/X VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__072__A _072_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_20_13 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_29_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_29_22 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_20_79 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_29_88 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_28_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_6_48 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_6_37 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_6_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_6_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_20_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_19_131 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_19_175 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_19_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_mux_bottom_track_13.mux_l1_in_1__A1 _088_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mux_right_track_0.mux_l2_in_2__S mux_right_track_0.mux_l2_in_3_/S VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_25_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_mux_left_track_1.mux_l3_in_0__S mux_left_track_1.mux_l3_in_1_/S VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__067__A _067_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_15_13 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_15_24 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xoutput89 _056_/X VGND VGND VPWR VPWR SC_OUT_BOT sky130_fd_sc_hd__buf_2
XFILLER_0_211 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xmux_right_track_8.mux_l2_in_1_ input70/X input63/X mux_right_track_8.mux_l2_in_3_/S
+ VGND VGND VPWR VPWR mux_right_track_8.mux_l2_in_1_/X sky130_fd_sc_hd__mux2_1
XANTENNA_input16_A chanx_left_in[14] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_16_156 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_16_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_104 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_115 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_126 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_137 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_148 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_159 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_mem_left_track_17.sky130_fd_sc_hd__dfxtp_1_1__CLK prog_clk_0_FTB00/X VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xmem_bottom_track_3.sky130_fd_sc_hd__dfxtp_1_0_ prog_clk_0_FTB00/X mem_bottom_track_3.delay_buf_2/X
+ VGND VGND VPWR VPWR mux_bottom_track_3.mux_l1_in_3_/S sky130_fd_sc_hd__dfxtp_2
XANTENNA_input8_A bottom_left_grid_pin_48_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_26_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_26_34 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_13_104 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_9_119 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_13_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_3_49 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_8_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_8_152 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_8_174 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_8_185 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmem_bottom_track_11.sky130_fd_sc_hd__dfxtp_1_2_ prog_clk_0_FTB00/X mux_bottom_track_11.mux_l2_in_1_/S
+ VGND VGND VPWR VPWR mux_bottom_track_11.mux_l3_in_0_/S sky130_fd_sc_hd__dfxtp_1
XFILLER_12_25 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_12_58 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__080__A _080_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_5_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_input83_A right_bottom_grid_pin_37_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_5_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_32_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_32_210 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_4_70 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_mux_bottom_track_7.mux_l1_in_0__A1 _064_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_23_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__075__A _075_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_23_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_2_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_2_136 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_2_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmem_bottom_track_9.sky130_fd_sc_hd__dfxtp_1_1_ prog_clk_0_FTB00/X mux_bottom_track_9.mux_l1_in_0_/S
+ VGND VGND VPWR VPWR mux_bottom_track_9.mux_l2_in_1_/S sky130_fd_sc_hd__dfxtp_1
XFILLER_0_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_14_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_1_191 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_mem_bottom_track_7.sky130_fd_sc_hd__dfxtp_1_1__CLK prog_clk_0_FTB00/X VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_18_13 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_18_24 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_18_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_110_ _110_/A VGND VGND VPWR VPWR _110_/X sky130_fd_sc_hd__clkbuf_1
XANTENNA_mux_bottom_track_5.mux_l1_in_2__A1 input8/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_input46_A chanx_right_in[5] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mux_bottom_track_21.mux_l1_in_1__A1 _094_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_1_60 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_20_25 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_20_36 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_29_67 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_29_34 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_29_12 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_28_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_28_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmem_bottom_track_7.delay_buf_2 mem_bottom_track_7.delay_buf_2/X VGND VGND VPWR VPWR
+ mem_bottom_track_7.delay_buf_2/X sky130_fd_sc_hd__buf_6
Xmux_bottom_track_11.sky130_fd_sc_hd__buf_4_0_ mux_bottom_track_11.mux_l3_in_0_/X
+ VGND VGND VPWR VPWR _102_/A sky130_fd_sc_hd__clkbuf_1
XFILLER_25_157 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_25_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_31_13 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__083__A _083_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_15_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_31_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_201 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_31_127 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_16_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_16_146 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_16_168 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xmux_right_track_8.mux_l2_in_0_ input87/X mux_right_track_8.mux_l1_in_0_/X mux_right_track_8.mux_l2_in_3_/S
+ VGND VGND VPWR VPWR mux_right_track_8.mux_l2_in_0_/X sky130_fd_sc_hd__mux2_1
XANTENNA_mux_right_track_8.mux_l2_in_1__A0 input70/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_105 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_116 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_127 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_138 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_149 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_22_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xrepeater151 repeater152/X VGND VGND VPWR VPWR repeater151/X sky130_fd_sc_hd__clkbuf_2
XFILLER_26_79 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_mux_right_track_4.mux_l1_in_6__A0 _092_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_9_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_21_182 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_3_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_3_28 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_12_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xmem_bottom_track_11.sky130_fd_sc_hd__dfxtp_1_1_ prog_clk_0_FTB00/X mux_bottom_track_11.mux_l1_in_0_/S
+ VGND VGND VPWR VPWR mux_bottom_track_11.mux_l2_in_1_/S sky130_fd_sc_hd__dfxtp_1
XFILLER_5_156 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_input76_A left_bottom_grid_pin_39_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mux_bottom_track_17.mux_l1_in_0__A0 input6/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__091__A _091_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xmem_bottom_track_9.sky130_fd_sc_hd__dfxtp_1_0_ prog_clk_0_FTB00/X mux_bottom_track_7.mux_l3_in_0_/S
+ VGND VGND VPWR VPWR mux_bottom_track_9.mux_l1_in_0_/S sky130_fd_sc_hd__dfxtp_1
Xmem_right_track_0.delay_buf input10/X VGND VGND VPWR VPWR input10/X sky130_fd_sc_hd__buf_6
XFILLER_18_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__086__A _086_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_input39_A chanx_right_in[17] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mem_bottom_track_11.sky130_fd_sc_hd__dfxtp_1_0__CLK prog_clk_0_FTB00/X VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_29_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_19_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_19_144 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_19_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_mem_right_track_4.sky130_fd_sc_hd__dfxtp_1_3__CLK prog_clk_0_FTB00/X VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_25_103 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_15_48 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_33_180 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_31_36 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_15_59 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_mem_bottom_track_25.sky130_fd_sc_hd__dfxtp_1_1__CLK prog_clk_0_FTB00/X VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_16_103 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_mux_right_track_8.mux_l2_in_1__A1 input63/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_31_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_106 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_117 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_128 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_139 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_0 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_30_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_7_60 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_7_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_26_14 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xrepeater152 repeater152/A VGND VGND VPWR VPWR repeater152/X sky130_fd_sc_hd__clkbuf_2
XANTENNA__094__A _094_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mem_left_track_33.sky130_fd_sc_hd__dfxtp_1_2__CLK prog_clk_0_FTB00/X VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mux_right_track_4.mux_l1_in_6__A1 _083_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_21_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmux_bottom_track_13.mux_l2_in_0_ mux_bottom_track_13.mux_l1_in_1_/X mux_bottom_track_13.mux_l1_in_0_/X
+ mux_bottom_track_13.mux_l2_in_0_/S VGND VGND VPWR VPWR mux_bottom_track_13.mux_l2_in_0_/X
+ sky130_fd_sc_hd__mux2_1
XANTENNA_input21_A chanx_left_in[19] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_8_132 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xmux_left_track_5.mux_l2_in_3__163 VGND VGND VPWR VPWR mux_left_track_5.mux_l2_in_3_/A0
+ mux_left_track_5.mux_l2_in_3__163/LO sky130_fd_sc_hd__conb_1
Xmem_bottom_track_11.sky130_fd_sc_hd__dfxtp_1_0_ prog_clk_0_FTB00/X mux_bottom_track_9.mux_l3_in_0_/S
+ VGND VGND VPWR VPWR mux_bottom_track_11.mux_l1_in_0_/S sky130_fd_sc_hd__dfxtp_1
Xmux_bottom_track_25.mux_l3_in_0_ mux_bottom_track_25.mux_l2_in_1_/X mux_bottom_track_25.mux_l2_in_0_/X
+ mux_bottom_track_25.mux_l3_in_0_/S VGND VGND VPWR VPWR mux_bottom_track_25.mux_l3_in_0_/X
+ sky130_fd_sc_hd__mux2_1
XFILLER_27_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_12_38 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xmux_right_track_8.mux_l1_in_0_ input83/X input88/X mux_right_track_8.mux_l1_in_0_/S
+ VGND VGND VPWR VPWR mux_right_track_8.mux_l1_in_0_/X sky130_fd_sc_hd__mux2_1
XANTENNA_input69_A chany_bottom_in[8] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_5_146 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_5_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_mux_bottom_track_17.mux_l1_in_0__A1 _071_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mem_right_track_8.sky130_fd_sc_hd__dfxtp_1_0__CLK prog_clk_0_FTB00/X VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mux_bottom_track_9.mux_l2_in_0__A0 _086_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_4_94 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmux_bottom_track_27.sky130_fd_sc_hd__buf_4_0_ mux_bottom_track_27.mux_l2_in_0_/X
+ VGND VGND VPWR VPWR _110_/A sky130_fd_sc_hd__clkbuf_1
XANTENNA_mem_left_track_1.sky130_fd_sc_hd__dfxtp_1_1__D mux_left_track_1.mux_l1_in_1_/S
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xmux_bottom_track_13.mux_l1_in_1_ mux_bottom_track_13.mux_l1_in_1_/A0 _088_/A mux_bottom_track_13.mux_l1_in_1_/S
+ VGND VGND VPWR VPWR mux_bottom_track_13.mux_l1_in_1_/X sky130_fd_sc_hd__mux2_1
Xmem_bottom_track_5.delay_buf_2 mem_bottom_track_5.delay_buf_2/X VGND VGND VPWR VPWR
+ mem_bottom_track_5.delay_buf_2/X sky130_fd_sc_hd__buf_6
Xmux_right_track_8.sky130_fd_sc_hd__buf_4_0_ mux_right_track_8.mux_l4_in_0_/X VGND
+ VGND VPWR VPWR _081_/A sky130_fd_sc_hd__clkbuf_1
Xmux_bottom_track_25.mux_l2_in_1_ mux_bottom_track_25.mux_l2_in_1_/A0 _096_/A mux_bottom_track_25.mux_l2_in_1_/S
+ VGND VGND VPWR VPWR mux_bottom_track_25.mux_l2_in_1_/X sky130_fd_sc_hd__mux2_1
Xmux_bottom_track_9.mux_l3_in_0_ mux_bottom_track_9.mux_l2_in_1_/X mux_bottom_track_9.mux_l2_in_0_/X
+ mux_bottom_track_9.mux_l3_in_0_/S VGND VGND VPWR VPWR mux_bottom_track_9.mux_l3_in_0_/X
+ sky130_fd_sc_hd__mux2_1
XANTENNA_mux_left_track_5.mux_l1_in_0__A0 _072_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xmux_bottom_track_25.mux_l2_in_1__180 VGND VGND VPWR VPWR mux_bottom_track_25.mux_l2_in_1_/A0
+ mux_bottom_track_25.mux_l2_in_1__180/LO sky130_fd_sc_hd__conb_1
Xmem_bottom_track_17.sky130_fd_sc_hd__dfxtp_1_1_ prog_clk_0_FTB00/X mux_bottom_track_17.mux_l1_in_1_/S
+ VGND VGND VPWR VPWR mux_bottom_track_17.mux_l2_in_0_/S sky130_fd_sc_hd__dfxtp_1
XFILLER_11_204 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_11_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_24_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_099_ _099_/A VGND VGND VPWR VPWR _099_/X sky130_fd_sc_hd__clkbuf_1
XANTENNA_mem_bottom_track_1.sky130_fd_sc_hd__dfxtp_1_2__CLK prog_clk_0_FTB00/X VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_20_49 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_28_145 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_28_134 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_28_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmux_bottom_track_9.mux_l2_in_1_ mux_bottom_track_9.mux_l2_in_1_/A0 input17/X mux_bottom_track_9.mux_l2_in_1_/S
+ VGND VGND VPWR VPWR mux_bottom_track_9.mux_l2_in_1_/X sky130_fd_sc_hd__mux2_1
XANTENNA_input51_A chany_bottom_in[0] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_10_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_19_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xmux_right_track_32.sky130_fd_sc_hd__buf_4_0_ mux_right_track_32.mux_l3_in_0_/X VGND
+ VGND VPWR VPWR _093_/A sky130_fd_sc_hd__clkbuf_1
XFILLER_25_148 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_25_115 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmux_right_track_4.mux_l1_in_6_ _092_/A _083_/A repeater152/X VGND VGND VPWR VPWR
+ mux_right_track_4.mux_l1_in_6_/X sky130_fd_sc_hd__mux2_1
XANTENNA_mem_right_track_24.sky130_fd_sc_hd__dfxtp_1_1__D mux_right_track_24.mux_l1_in_3_/S
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_21_70 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_21_92 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_107 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_118 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_129 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_30_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_26_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xrepeater153 repeater154/X VGND VGND VPWR VPWR repeater153/X sky130_fd_sc_hd__clkbuf_2
XFILLER_21_140 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_21_162 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_mux_bottom_track_25.mux_l1_in_0__A1 _076_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_input14_A chanx_left_in[12] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_12_162 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_input6_A bottom_left_grid_pin_46_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_26_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_26_210 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_5_103 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_5_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_5_136 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmux_left_track_3.mux_l2_in_3_ mux_left_track_3.mux_l2_in_3_/A0 input77/X mux_left_track_3.mux_l2_in_3_/S
+ VGND VGND VPWR VPWR mux_left_track_3.mux_l2_in_3_/X sky130_fd_sc_hd__mux2_1
Xmem_left_track_1.sky130_fd_sc_hd__dfxtp_1_3_ prog_clk_0_FTB00/X mux_left_track_1.mux_l3_in_1_/S
+ VGND VGND VPWR VPWR mux_left_track_1.mux_l4_in_0_/S sky130_fd_sc_hd__dfxtp_1
XANTENNA_mux_bottom_track_1.mux_l1_in_2__S mux_bottom_track_1.mux_l1_in_3_/S VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xmux_bottom_track_13.mux_l1_in_0_ input4/X _068_/A mux_bottom_track_13.mux_l1_in_1_/S
+ VGND VGND VPWR VPWR mux_bottom_track_13.mux_l1_in_0_/X sky130_fd_sc_hd__mux2_1
XFILLER_23_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_mux_left_track_33.mux_l3_in_0__S output90/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xmux_bottom_track_25.mux_l2_in_0_ input2/X mux_bottom_track_25.mux_l1_in_0_/X mux_bottom_track_25.mux_l2_in_1_/S
+ VGND VGND VPWR VPWR mux_bottom_track_25.mux_l2_in_0_/X sky130_fd_sc_hd__mux2_1
XANTENNA_input81_A right_bottom_grid_pin_35_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_13_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_29_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_mux_left_track_5.mux_l1_in_0__A1 _063_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xmux_bottom_track_15.mux_l1_in_1__175 VGND VGND VPWR VPWR mux_bottom_track_15.mux_l1_in_1_/A0
+ mux_bottom_track_15.mux_l1_in_1__175/LO sky130_fd_sc_hd__conb_1
XFILLER_18_38 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xmem_bottom_track_17.sky130_fd_sc_hd__dfxtp_1_0_ prog_clk_0_FTB00/X mux_bottom_track_15.mux_l2_in_0_/S
+ VGND VGND VPWR VPWR mux_bottom_track_17.mux_l1_in_1_/S sky130_fd_sc_hd__dfxtp_1
XFILLER_7_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_098_ _098_/A VGND VGND VPWR VPWR _098_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_6_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_mux_right_track_16.mux_l1_in_2__S mux_right_track_16.mux_l1_in_3_/S VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_1_30 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_29_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmux_left_track_3.mux_l4_in_0_ mux_left_track_3.mux_l3_in_1_/X mux_left_track_3.mux_l3_in_0_/X
+ mux_left_track_3.mux_l4_in_0_/S VGND VGND VPWR VPWR mux_left_track_3.mux_l4_in_0_/X
+ sky130_fd_sc_hd__mux2_1
XFILLER_29_48 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_28_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_28_102 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmux_bottom_track_9.mux_l2_in_0_ _086_/A mux_bottom_track_9.mux_l1_in_0_/X mux_bottom_track_9.mux_l2_in_1_/S
+ VGND VGND VPWR VPWR mux_bottom_track_9.mux_l2_in_0_/X sky130_fd_sc_hd__mux2_1
XFILLER_10_50 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_input44_A chanx_right_in[3] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mem_left_track_1.sky130_fd_sc_hd__dfxtp_1_2__CLK prog_clk_0_FTB00/X VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_19_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_19_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_25_127 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmux_right_track_4.mux_l1_in_5_ input59/X input52/X repeater152/A VGND VGND VPWR VPWR
+ mux_right_track_4.mux_l1_in_5_/X sky130_fd_sc_hd__mux2_1
XFILLER_31_108 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_24_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_108 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_119 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_mux_left_track_3.mux_l2_in_1__A1 input56/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_2 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xmux_left_track_3.mux_l3_in_1_ mux_left_track_3.mux_l2_in_3_/X mux_left_track_3.mux_l2_in_2_/X
+ mux_left_track_3.mux_l3_in_1_/S VGND VGND VPWR VPWR mux_left_track_3.mux_l3_in_1_/X
+ sky130_fd_sc_hd__mux2_1
XFILLER_15_171 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_15_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_30_174 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_30_163 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_30_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_7_40 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmem_bottom_track_3.delay_buf_2 mem_bottom_track_3.delay_buf_2/X VGND VGND VPWR VPWR
+ mem_bottom_track_3.delay_buf_2/X sky130_fd_sc_hd__buf_6
Xmux_left_track_5.sky130_fd_sc_hd__buf_4_0_ mux_left_track_5.mux_l4_in_0_/X VGND VGND
+ VPWR VPWR _059_/A sky130_fd_sc_hd__clkbuf_1
XFILLER_26_49 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_26_38 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xrepeater154 repeater154/A VGND VGND VPWR VPWR repeater154/X sky130_fd_sc_hd__clkbuf_2
XFILLER_13_108 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_21_174 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_16_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_mem_right_track_16.sky130_fd_sc_hd__dfxtp_1_2__D mux_right_track_16.mux_l2_in_1_/S
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_8_156 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_8_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_12_185 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmem_left_track_1.sky130_fd_sc_hd__dfxtp_1_2_ prog_clk_0_FTB00/X mux_left_track_1.mux_l2_in_3_/S
+ VGND VGND VPWR VPWR mux_left_track_1.mux_l3_in_1_/S sky130_fd_sc_hd__dfxtp_1
Xmux_left_track_3.mux_l2_in_2_ input75/X input73/X mux_left_track_3.mux_l2_in_3_/S
+ VGND VGND VPWR VPWR mux_left_track_3.mux_l2_in_2_/X sky130_fd_sc_hd__mux2_1
XFILLER_14_203 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_input74_A left_bottom_grid_pin_37_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mem_right_track_2.sky130_fd_sc_hd__dfxtp_1_1__CLK prog_clk_0_FTB00/X VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_1_173 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_1_140 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_mux_right_track_2.mux_l2_in_1__S mux_right_track_2.mux_l2_in_3_/S VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
Xmux_right_track_4.mux_l2_in_3_ mux_right_track_4.mux_l2_in_3_/A0 mux_right_track_4.mux_l1_in_6_/X
+ mux_right_track_4.mux_l2_in_3_/S VGND VGND VPWR VPWR mux_right_track_4.mux_l2_in_3_/X
+ sky130_fd_sc_hd__mux2_1
XANTENNA_mux_left_track_9.mux_l2_in_0__S mux_left_track_9.mux_l2_in_3_/S VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
X_097_ _097_/A VGND VGND VPWR VPWR _097_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_1_20 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_20_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_28_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xmux_bottom_track_25.mux_l1_in_0_ input41/X _076_/A mux_bottom_track_25.mux_l1_in_0_/S
+ VGND VGND VPWR VPWR mux_bottom_track_25.mux_l1_in_0_/X sky130_fd_sc_hd__mux2_1
XFILLER_10_40 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_input37_A chanx_right_in[15] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_19_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_19_103 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_mem_bottom_track_15.sky130_fd_sc_hd__dfxtp_1_0__CLK prog_clk_0_FTB00/X VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_33_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_33_172 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_15_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xmux_right_track_4.mux_l1_in_4_ input64/X input87/X repeater151/X VGND VGND VPWR VPWR
+ mux_right_track_4.mux_l1_in_4_/X sky130_fd_sc_hd__mux2_1
XFILLER_16_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_24_172 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_mux_bottom_track_19.mux_l1_in_1__A1 _092_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_109 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_mem_right_track_8.sky130_fd_sc_hd__dfxtp_1_3__CLK prog_clk_0_FTB00/X VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xmux_left_track_3.mux_l3_in_0_ mux_left_track_3.mux_l2_in_1_/X mux_left_track_3.mux_l2_in_0_/X
+ mux_left_track_3.mux_l3_in_1_/S VGND VGND VPWR VPWR mux_left_track_3.mux_l3_in_0_/X
+ sky130_fd_sc_hd__mux2_1
XFILLER_30_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_7_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmux_right_track_4.mux_l4_in_0_ mux_right_track_4.mux_l3_in_1_/X mux_right_track_4.mux_l3_in_0_/X
+ mux_right_track_4.mux_l4_in_0_/S VGND VGND VPWR VPWR mux_right_track_4.mux_l4_in_0_/X
+ sky130_fd_sc_hd__mux2_1
Xmux_bottom_track_9.mux_l1_in_0_ input2/X _066_/A mux_bottom_track_9.mux_l1_in_0_/S
+ VGND VGND VPWR VPWR mux_bottom_track_9.mux_l1_in_0_/X sky130_fd_sc_hd__mux2_1
XFILLER_21_186 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_32_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_32_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_32_71 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_8_124 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_12_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_mux_left_track_17.mux_l2_in_0__A0 mux_left_track_17.mux_l1_in_1_/X VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
Xmux_bottom_track_9.sky130_fd_sc_hd__buf_4_0_ mux_bottom_track_9.mux_l3_in_0_/X VGND
+ VGND VPWR VPWR _101_/A sky130_fd_sc_hd__clkbuf_1
XANTENNA_mux_right_track_24.mux_l1_in_0__S mux_right_track_24.mux_l1_in_3_/S VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_12_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xmem_left_track_1.sky130_fd_sc_hd__dfxtp_1_1_ prog_clk_0_FTB00/X mux_left_track_1.mux_l1_in_1_/S
+ VGND VGND VPWR VPWR mux_left_track_1.mux_l2_in_3_/S sky130_fd_sc_hd__dfxtp_2
Xmux_left_track_3.mux_l2_in_1_ input71/X input56/X mux_left_track_3.mux_l2_in_3_/S
+ VGND VGND VPWR VPWR mux_left_track_3.mux_l2_in_1_/X sky130_fd_sc_hd__mux2_1
XFILLER_32_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_mux_left_track_9.mux_l2_in_3__S mux_left_track_9.mux_l2_in_3_/S VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_4_42 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_4_31 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmux_right_track_4.mux_l3_in_1_ mux_right_track_4.mux_l2_in_3_/X mux_right_track_4.mux_l2_in_2_/X
+ mux_right_track_4.mux_l3_in_1_/S VGND VGND VPWR VPWR mux_right_track_4.mux_l3_in_1_/X
+ sky130_fd_sc_hd__mux2_1
XFILLER_4_75 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_4_64 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_4_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_13_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_input67_A chany_bottom_in[6] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mem_right_track_2.sky130_fd_sc_hd__dfxtp_1_2__D mux_right_track_2.mux_l2_in_3_/S
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_20_207 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_20_218 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xmem_right_track_4.sky130_fd_sc_hd__dfxtp_1_3_ prog_clk_0_FTB00/X mux_right_track_4.mux_l3_in_1_/S
+ VGND VGND VPWR VPWR mux_right_track_4.mux_l4_in_0_/S sky130_fd_sc_hd__dfxtp_1
Xmux_right_track_4.mux_l2_in_2_ mux_right_track_4.mux_l1_in_5_/X mux_right_track_4.mux_l1_in_4_/X
+ mux_right_track_4.mux_l2_in_3_/S VGND VGND VPWR VPWR mux_right_track_4.mux_l2_in_2_/X
+ sky130_fd_sc_hd__mux2_1
X_096_ _096_/A VGND VGND VPWR VPWR _096_/X sky130_fd_sc_hd__clkbuf_1
Xmem_bottom_track_1.delay_buf_2 mem_bottom_track_1.delay_buf_2/X VGND VGND VPWR VPWR
+ mem_bottom_track_1.delay_buf_2/X sky130_fd_sc_hd__buf_6
XFILLER_1_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_1_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_1_76 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_29_17 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_3_203 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_19_148 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_mux_right_track_24.mux_l1_in_3__S mux_right_track_24.mux_l1_in_3_/S VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_079_ _079_/A VGND VGND VPWR VPWR _079_/X sky130_fd_sc_hd__clkbuf_1
XANTENNA_mem_bottom_track_5.sky130_fd_sc_hd__dfxtp_1_2__CLK prog_clk_0_FTB00/X VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_25_107 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_33_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_33_151 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xmux_right_track_16.mux_l1_in_3_ mux_right_track_16.mux_l1_in_3_/A0 _095_/A mux_right_track_16.mux_l1_in_3_/S
+ VGND VGND VPWR VPWR mux_right_track_16.mux_l1_in_3_/X sky130_fd_sc_hd__mux2_1
XFILLER_31_18 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_mux_left_track_17.mux_l1_in_1__A1 input64/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xmux_right_track_4.mux_l1_in_3_ input86/X input85/X repeater151/X VGND VGND VPWR VPWR
+ mux_right_track_4.mux_l1_in_3_/X sky130_fd_sc_hd__mux2_1
XANTENNA_mux_left_track_17.mux_l1_in_0__S mux_left_track_17.mux_l1_in_3_/S VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_16_107 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_24_151 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_21_40 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_30_132 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_30_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_30_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_4 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_mux_right_track_16.mux_l2_in_0__S mux_right_track_16.mux_l2_in_1_/S VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_15_151 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_15_162 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_7_64 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_7_86 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_mem_left_track_33.sky130_fd_sc_hd__dfxtp_1_2__D mux_left_track_33.mux_l2_in_1_/S
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_26_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_21_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_21_198 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_29_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_29_210 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_8_103 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_32_50 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_8_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmem_left_track_1.sky130_fd_sc_hd__dfxtp_1_0_ prog_clk_0_FTB00/X mux_bottom_track_27.mux_l2_in_0_/S
+ VGND VGND VPWR VPWR mux_left_track_1.mux_l1_in_1_/S sky130_fd_sc_hd__dfxtp_1
Xmux_left_track_3.mux_l2_in_0_ mux_left_track_3.mux_l1_in_1_/X mux_left_track_3.mux_l1_in_0_/X
+ mux_left_track_3.mux_l2_in_3_/S VGND VGND VPWR VPWR mux_left_track_3.mux_l2_in_0_/X
+ sky130_fd_sc_hd__mux2_1
XFILLER_27_94 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_27_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_input12_A chanx_left_in[10] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xmux_right_track_16.mux_l3_in_0_ mux_right_track_16.mux_l2_in_1_/X mux_right_track_16.mux_l2_in_0_/X
+ mem_right_track_24.delay_buf_2/X VGND VGND VPWR VPWR mux_right_track_16.mux_l3_in_0_/X
+ sky130_fd_sc_hd__mux2_1
XFILLER_4_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmux_right_track_4.mux_l3_in_0_ mux_right_track_4.mux_l2_in_1_/X mux_right_track_4.mux_l2_in_0_/X
+ mux_right_track_4.mux_l3_in_1_/S VGND VGND VPWR VPWR mux_right_track_4.mux_l3_in_0_/X
+ sky130_fd_sc_hd__mux2_1
XANTENNA_input4_A bottom_left_grid_pin_44_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mux_left_track_33.mux_l1_in_1__A0 input61/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_1_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xmem_right_track_4.sky130_fd_sc_hd__dfxtp_1_2_ prog_clk_0_FTB00/X mux_right_track_4.mux_l2_in_3_/S
+ VGND VGND VPWR VPWR mux_right_track_4.mux_l3_in_1_/S sky130_fd_sc_hd__dfxtp_1
Xmux_left_track_3.mux_l1_in_1_ input68/X input51/X mux_left_track_3.mux_l1_in_1_/S
+ VGND VGND VPWR VPWR mux_left_track_3.mux_l1_in_1_/X sky130_fd_sc_hd__mux2_1
Xmux_right_track_16.mux_l2_in_1_ mux_right_track_16.mux_l1_in_3_/X mux_right_track_16.mux_l1_in_2_/X
+ mux_right_track_16.mux_l2_in_1_/S VGND VGND VPWR VPWR mux_right_track_16.mux_l2_in_1_/X
+ sky130_fd_sc_hd__mux2_1
XANTENNA_mux_left_track_17.mux_l1_in_3__S mux_left_track_17.mux_l1_in_3_/S VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_24_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_095_ _095_/A VGND VGND VPWR VPWR _095_/X sky130_fd_sc_hd__clkbuf_1
Xmux_right_track_4.mux_l2_in_1_ mux_right_track_4.mux_l1_in_3_/X mux_right_track_4.mux_l1_in_2_/X
+ mux_right_track_4.mux_l2_in_3_/S VGND VGND VPWR VPWR mux_right_track_4.mux_l2_in_1_/X
+ sky130_fd_sc_hd__mux2_1
XFILLER_27_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_28_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_28_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_10_20 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmux_bottom_track_11.mux_l2_in_1__173 VGND VGND VPWR VPWR mux_bottom_track_11.mux_l2_in_1_/A0
+ mux_bottom_track_11.mux_l2_in_1__173/LO sky130_fd_sc_hd__conb_1
XFILLER_27_171 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_19_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_078_ _078_/A VGND VGND VPWR VPWR _078_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_33_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_25_119 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_mux_left_track_5.mux_l2_in_0__S mux_left_track_5.mux_l2_in_3_/S VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
Xmux_right_track_16.mux_l1_in_2_ _086_/A input57/X mux_right_track_16.mux_l1_in_3_/S
+ VGND VGND VPWR VPWR mux_right_track_16.mux_l1_in_2_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_207 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xmux_right_track_4.mux_l1_in_2_ input84/X input83/X repeater151/X VGND VGND VPWR VPWR
+ mux_right_track_4.mux_l1_in_2_/X sky130_fd_sc_hd__mux2_1
XANTENNA_mem_left_track_5.sky130_fd_sc_hd__dfxtp_1_2__CLK prog_clk_0_FTB00/X VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mux_right_track_8.mux_l2_in_0__S mux_right_track_8.mux_l2_in_3_/S VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_21_52 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_21_63 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_21_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_input42_A chanx_right_in[1] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_5 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_7_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_21_122 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_21_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_29_200 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_mux_right_track_0.mux_l2_in_2__A0 _080_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_12_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_16_63 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_16_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_16_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmux_left_track_3.mux_l2_in_3__161 VGND VGND VPWR VPWR mux_left_track_3.mux_l2_in_3_/A0
+ mux_left_track_3.mux_l2_in_3__161/LO sky130_fd_sc_hd__conb_1
XFILLER_7_192 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_5_118 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_5_107 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_32_206 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_4_99 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_23_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_13_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_13_86 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_mux_left_track_33.mux_l1_in_1__A1 input54/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_9_210 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_9_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmem_right_track_4.sky130_fd_sc_hd__dfxtp_1_1_ prog_clk_0_FTB00/X repeater152/X VGND
+ VGND VPWR VPWR mux_right_track_4.mux_l2_in_3_/S sky130_fd_sc_hd__dfxtp_2
XANTENNA_mux_left_track_5.mux_l2_in_3__S mux_left_track_5.mux_l2_in_3_/S VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
Xmux_left_track_3.mux_l1_in_0_ _071_/A _062_/A mux_left_track_3.mux_l1_in_1_/S VGND
+ VGND VPWR VPWR mux_left_track_3.mux_l1_in_0_/X sky130_fd_sc_hd__mux2_1
Xmux_right_track_16.mux_l2_in_0_ mux_right_track_16.mux_l1_in_1_/X mux_right_track_16.mux_l1_in_0_/X
+ mux_right_track_16.mux_l2_in_1_/S VGND VGND VPWR VPWR mux_right_track_16.mux_l2_in_0_/X
+ sky130_fd_sc_hd__mux2_1
XANTENNA_mux_right_track_8.mux_l2_in_3__S mux_right_track_8.mux_l2_in_3_/S VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
Xmux_right_track_4.mux_l2_in_0_ mux_right_track_4.mux_l1_in_1_/X mux_right_track_4.mux_l1_in_0_/X
+ mux_right_track_4.mux_l2_in_3_/S VGND VGND VPWR VPWR mux_right_track_4.mux_l2_in_0_/X
+ sky130_fd_sc_hd__mux2_1
XFILLER_24_63 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_24_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_094_ _094_/A VGND VGND VPWR VPWR _094_/X sky130_fd_sc_hd__clkbuf_1
XANTENNA_input72_A left_bottom_grid_pin_35_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xmux_bottom_track_27.mux_l2_in_0__181 VGND VGND VPWR VPWR mux_bottom_track_27.mux_l2_in_0_/A0
+ mux_bottom_track_27.mux_l2_in_0__181/LO sky130_fd_sc_hd__conb_1
XFILLER_1_89 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_mem_left_track_17.sky130_fd_sc_hd__dfxtp_1_1__D mux_left_track_17.mux_l1_in_3_/S
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_10_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_10_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_10_87 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_19_30 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_19_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_077_ _077_/A VGND VGND VPWR VPWR _077_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_33_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_18_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmux_right_track_16.mux_l1_in_1_ input69/X input62/X mux_right_track_16.mux_l1_in_3_/S
+ VGND VGND VPWR VPWR mux_right_track_16.mux_l1_in_1_/X sky130_fd_sc_hd__mux2_1
Xmux_right_track_4.mux_l1_in_1_ input82/X input81/X repeater151/X VGND VGND VPWR VPWR
+ mux_right_track_4.mux_l1_in_1_/X sky130_fd_sc_hd__mux2_1
XFILLER_24_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_input35_A chanx_right_in[13] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mux_bottom_track_3.mux_l1_in_0__A0 input3/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_6 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_15_120 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_15_175 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_mem_bottom_track_19.sky130_fd_sc_hd__dfxtp_1_0__CLK prog_clk_0_FTB00/X VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_30_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_30_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_7_22 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_7_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_21_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xinput80 right_bottom_grid_pin_34_ VGND VGND VPWR VPWR input80/X sky130_fd_sc_hd__clkbuf_1
XANTENNA_mux_left_track_9.mux_l2_in_1__A0 input58/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mux_right_track_0.mux_l2_in_2__A1 input61/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_32_63 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_8_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_12_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_mux_right_track_24.mux_l2_in_1__S mux_right_track_24.mux_l2_in_1_/S VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xmux_right_track_2.mux_l2_in_3__167 VGND VGND VPWR VPWR mux_right_track_2.mux_l2_in_3_/A0
+ mux_right_track_2.mux_l2_in_3__167/LO sky130_fd_sc_hd__conb_1
XANTENNA_mem_left_track_5.sky130_fd_sc_hd__dfxtp_1_3__D mux_left_track_5.mux_l3_in_1_/S
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_4_130 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_mux_right_track_0.mux_l3_in_1__A1 mux_right_track_0.mux_l2_in_2_/X VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mem_right_track_16.sky130_fd_sc_hd__dfxtp_1_0__CLK prog_clk_0_FTB00/X VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_1_100 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_1_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_8_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_mem_bottom_track_3.sky130_fd_sc_hd__dfxtp_1_0__CLK prog_clk_0_FTB00/X VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xmem_right_track_4.sky130_fd_sc_hd__dfxtp_1_0_ prog_clk_0_FTB00/X mux_right_track_2.mux_l4_in_0_/S
+ VGND VGND VPWR VPWR repeater152/A sky130_fd_sc_hd__dfxtp_1
XFILLER_10_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_24_20 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_093_ _093_/A VGND VGND VPWR VPWR _093_/X sky130_fd_sc_hd__clkbuf_1
XANTENNA_input65_A chany_bottom_in[4] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_1_13 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_1_35 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_28_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_28_118 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xinput1 SC_IN_BOT VGND VGND VPWR VPWR _056_/A sky130_fd_sc_hd__clkbuf_1
Xmem_bottom_track_21.sky130_fd_sc_hd__dfxtp_1_1_ prog_clk_0_FTB00/X mux_bottom_track_21.mux_l1_in_1_/S
+ VGND VGND VPWR VPWR mux_bottom_track_21.mux_l2_in_0_/S sky130_fd_sc_hd__dfxtp_1
XTAP_90 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xmux_bottom_track_5.mux_l1_in_3_ mux_bottom_track_5.mux_l1_in_3_/A0 input28/X mux_bottom_track_5.mux_l1_in_3_/S
+ VGND VGND VPWR VPWR mux_bottom_track_5.mux_l1_in_3_/X sky130_fd_sc_hd__mux2_1
XFILLER_19_107 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_076_ _076_/A VGND VGND VPWR VPWR _076_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_32_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmux_bottom_track_23.sky130_fd_sc_hd__buf_4_0_ mux_bottom_track_23.mux_l2_in_0_/X
+ VGND VGND VPWR VPWR _108_/A sky130_fd_sc_hd__clkbuf_1
XFILLER_33_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmux_right_track_16.mux_l1_in_0_ input84/X input80/X mux_right_track_16.mux_l1_in_3_/S
+ VGND VGND VPWR VPWR mux_right_track_16.mux_l1_in_0_/X sky130_fd_sc_hd__mux2_1
Xmux_right_track_4.mux_l1_in_0_ input80/X input88/X repeater152/X VGND VGND VPWR VPWR
+ mux_right_track_4.mux_l1_in_0_/X sky130_fd_sc_hd__mux2_1
XFILLER_24_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_24_143 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmux_right_track_4.sky130_fd_sc_hd__buf_4_0_ mux_right_track_4.mux_l4_in_0_/X VGND
+ VGND VPWR VPWR _079_/A sky130_fd_sc_hd__clkbuf_1
XFILLER_24_176 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_mux_left_track_17.mux_l2_in_1__S mux_left_track_17.mux_l2_in_1_/S VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mux_bottom_track_3.mux_l1_in_0__A1 _062_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_input28_A chanx_left_in[7] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mem_bottom_track_9.sky130_fd_sc_hd__dfxtp_1_2__CLK prog_clk_0_FTB00/X VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xmux_left_track_25.mux_l1_in_3__160 VGND VGND VPWR VPWR mux_left_track_25.mux_l1_in_3_/A0
+ mux_left_track_25.mux_l1_in_3__160/LO sky130_fd_sc_hd__conb_1
XFILLER_30_146 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_30_124 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_30_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_30_179 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_30_157 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_7_45 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_7_78 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_059_ _059_/A VGND VGND VPWR VPWR _059_/X sky130_fd_sc_hd__clkbuf_1
XANTENNA_mem_right_track_0.delay_buf_A input10/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mux_left_track_9.mux_l2_in_1__A1 input70/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xinput70 chany_bottom_in[9] VGND VGND VPWR VPWR input70/X sky130_fd_sc_hd__clkbuf_1
Xinput81 right_bottom_grid_pin_35_ VGND VGND VPWR VPWR input81/X sky130_fd_sc_hd__clkbuf_1
XANTENNA_mux_left_track_1.mux_l2_in_0__S mux_left_track_1.mux_l2_in_3_/S VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
Xmux_bottom_track_17.sky130_fd_sc_hd__buf_4_0_ mux_bottom_track_17.mux_l2_in_0_/X
+ VGND VGND VPWR VPWR _105_/A sky130_fd_sc_hd__clkbuf_1
XFILLER_8_128 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_12_179 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmux_left_track_33.mux_l2_in_1__162 VGND VGND VPWR VPWR mux_left_track_33.mux_l2_in_1_/A0
+ mux_left_track_33.mux_l2_in_1__162/LO sky130_fd_sc_hd__conb_1
XANTENNA_mux_bottom_track_1.mux_l1_in_2__A1 input8/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xmux_bottom_track_5.mux_l3_in_0_ mux_bottom_track_5.mux_l2_in_1_/X mux_bottom_track_5.mux_l2_in_0_/X
+ mem_bottom_track_7.delay_buf_2/X VGND VGND VPWR VPWR mux_bottom_track_5.mux_l3_in_0_/X
+ sky130_fd_sc_hd__mux2_1
XFILLER_4_175 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_4_164 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_4_24 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_4_13 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_13_33 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_13_66 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_13_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_1_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_input10_A ccff_head VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xmux_bottom_track_5.mux_l2_in_1_ mux_bottom_track_5.mux_l1_in_3_/X mux_bottom_track_5.mux_l1_in_2_/X
+ mux_bottom_track_5.mux_l2_in_1_/S VGND VGND VPWR VPWR mux_bottom_track_5.mux_l2_in_1_/X
+ sky130_fd_sc_hd__mux2_1
Xmux_bottom_track_13.mux_l1_in_1__174 VGND VGND VPWR VPWR mux_bottom_track_13.mux_l1_in_1_/A0
+ mux_bottom_track_13.mux_l1_in_1__174/LO sky130_fd_sc_hd__conb_1
XANTENNA_mem_left_track_3.sky130_fd_sc_hd__dfxtp_1_0__CLK prog_clk_0_FTB00/X VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_input2_A bottom_left_grid_pin_42_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_24_87 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_092_ _092_/A VGND VGND VPWR VPWR _092_/X sky130_fd_sc_hd__clkbuf_1
XANTENNA_input58_A chany_bottom_in[16] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_1_25 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_1_47 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xinput2 bottom_left_grid_pin_42_ VGND VGND VPWR VPWR input2/X sky130_fd_sc_hd__clkbuf_2
Xmem_bottom_track_21.sky130_fd_sc_hd__dfxtp_1_0_ prog_clk_0_FTB00/X mux_bottom_track_19.mux_l2_in_0_/S
+ VGND VGND VPWR VPWR mux_bottom_track_21.mux_l1_in_1_/S sky130_fd_sc_hd__dfxtp_1
XANTENNA_mux_left_track_1.mux_l2_in_3__S mux_left_track_1.mux_l2_in_3_/S VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_91 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_80 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xmux_bottom_track_5.mux_l1_in_2_ _083_/A input8/X mux_bottom_track_5.mux_l1_in_3_/S
+ VGND VGND VPWR VPWR mux_bottom_track_5.mux_l1_in_2_/X sky130_fd_sc_hd__mux2_1
XFILLER_10_67 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_10_78 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_mem_right_track_0.sky130_fd_sc_hd__dfxtp_1_2__CLK prog_clk_0_FTB00/X VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_19_43 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_19_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_27_185 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_075_ _075_/A VGND VGND VPWR VPWR _075_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_25_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_18_130 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_mem_bottom_track_21.sky130_fd_sc_hd__dfxtp_1_0__CLK prog_clk_0_FTB00/X VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_33_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_33_155 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_33_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_33_122 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_mux_left_track_5.mux_l3_in_1__S mux_left_track_5.mux_l3_in_1_/S VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
Xmux_right_track_16.sky130_fd_sc_hd__buf_4_0_ mux_right_track_16.mux_l3_in_0_/X VGND
+ VGND VPWR VPWR _085_/A sky130_fd_sc_hd__clkbuf_1
XFILLER_24_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_24_155 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_21_22 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_21_66 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_8 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_15_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_15_155 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_15_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_058_ _058_/A VGND VGND VPWR VPWR _058_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_16_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmux_bottom_track_19.mux_l2_in_0_ mux_bottom_track_19.mux_l1_in_1_/X mux_bottom_track_19.mux_l1_in_0_/X
+ mux_bottom_track_19.mux_l2_in_0_/S VGND VGND VPWR VPWR mux_bottom_track_19.mux_l2_in_0_/X
+ sky130_fd_sc_hd__mux2_1
XFILLER_21_158 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_21_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xinput82 right_bottom_grid_pin_36_ VGND VGND VPWR VPWR input82/X sky130_fd_sc_hd__clkbuf_1
Xinput60 chany_bottom_in[18] VGND VGND VPWR VPWR input60/X sky130_fd_sc_hd__clkbuf_1
Xinput71 left_bottom_grid_pin_34_ VGND VGND VPWR VPWR input71/X sky130_fd_sc_hd__clkbuf_1
XANTENNA_mem_left_track_9.sky130_fd_sc_hd__dfxtp_1_2__CLK prog_clk_0_FTB00/X VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_8_107 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_12_158 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_16_33 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_32_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_32_43 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xmem_bottom_track_27.sky130_fd_sc_hd__dfxtp_1_1_ prog_clk_0_FTB00/X mux_bottom_track_27.mux_l1_in_0_/S
+ VGND VGND VPWR VPWR mux_bottom_track_27.mux_l2_in_0_/S sky130_fd_sc_hd__dfxtp_1
Xmux_bottom_track_21.mux_l2_in_0_ mux_bottom_track_21.mux_l1_in_1_/X mux_bottom_track_21.mux_l1_in_0_/X
+ mux_bottom_track_21.mux_l2_in_0_/S VGND VGND VPWR VPWR mux_bottom_track_21.mux_l2_in_0_/X
+ sky130_fd_sc_hd__mux2_1
XANTENNA_mem_bottom_track_13.sky130_fd_sc_hd__dfxtp_1_1__CLK prog_clk_0_FTB00/X VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_input40_A chanx_right_in[18] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_27_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_27_43 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_input88_A right_top_grid_pin_1_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mux_left_track_33.mux_l1_in_2__S mux_left_track_33.mux_l1_in_2_/S VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
Xmux_bottom_track_19.mux_l1_in_1_ mux_bottom_track_19.mux_l1_in_1_/A0 _092_/A mux_bottom_track_19.mux_l1_in_1_/S
+ VGND VGND VPWR VPWR mux_bottom_track_19.mux_l1_in_1_/X sky130_fd_sc_hd__mux2_1
XANTENNA_mem_bottom_track_1.sky130_fd_sc_hd__dfxtp_1_1__D mux_bottom_track_1.mux_l1_in_3_/S
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_14_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmux_bottom_track_21.mux_l1_in_1_ mux_bottom_track_21.mux_l1_in_1_/A0 _094_/A mux_bottom_track_21.mux_l1_in_1_/S
+ VGND VGND VPWR VPWR mux_bottom_track_21.mux_l1_in_1_/X sky130_fd_sc_hd__mux2_1
XFILLER_1_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_1_179 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_1_146 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_mem_right_track_32.sky130_fd_sc_hd__dfxtp_1_1__CLK prog_clk_0_FTB00/X VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xmux_bottom_track_5.mux_l2_in_0_ mux_bottom_track_5.mux_l1_in_1_/X mux_bottom_track_5.mux_l1_in_0_/X
+ mux_bottom_track_5.mux_l2_in_1_/S VGND VGND VPWR VPWR mux_bottom_track_5.mux_l2_in_0_/X
+ sky130_fd_sc_hd__mux2_1
Xmem_bottom_track_5.sky130_fd_sc_hd__dfxtp_1_2_ prog_clk_0_FTB00/X mux_bottom_track_5.mux_l2_in_1_/S
+ VGND VGND VPWR VPWR mem_bottom_track_7.delay_buf_2/X sky130_fd_sc_hd__dfxtp_1
Xmux_left_track_1.sky130_fd_sc_hd__buf_4_0_ mux_left_track_1.mux_l4_in_0_/X VGND VGND
+ VPWR VPWR _057_/A sky130_fd_sc_hd__clkbuf_1
XFILLER_24_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_091_ _091_/A VGND VGND VPWR VPWR _091_/X sky130_fd_sc_hd__clkbuf_1
XANTENNA_mux_bottom_track_5.mux_l1_in_1__A0 input6/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mux_bottom_track_21.mux_l1_in_0__A0 input8/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_92 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_81 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xinput3 bottom_left_grid_pin_43_ VGND VGND VPWR VPWR input3/X sky130_fd_sc_hd__clkbuf_2
XTAP_70 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_mux_right_track_2.mux_l2_in_3__A1 _091_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_3_219 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_3_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__062__A _062_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xmux_bottom_track_5.mux_l1_in_1_ input6/X input4/X mux_bottom_track_5.mux_l1_in_3_/S
+ VGND VGND VPWR VPWR mux_bottom_track_5.mux_l1_in_1_/X sky130_fd_sc_hd__mux2_1
XANTENNA_mem_right_track_24.sky130_fd_sc_hd__dfxtp_1_2__CLK prog_clk_0_FTB00/X VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_27_175 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_074_ _074_/A VGND VGND VPWR VPWR _074_/X sky130_fd_sc_hd__clkbuf_1
XANTENNA_input70_A chany_bottom_in[9] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_33_101 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_18_175 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_33_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmux_right_track_16.mux_l1_in_3__166 VGND VGND VPWR VPWR mux_right_track_16.mux_l1_in_3_/A0
+ mux_right_track_16.mux_l1_in_3__166/LO sky130_fd_sc_hd__conb_1
XANTENNA_mux_bottom_track_13.mux_l1_in_0__A1 _068_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_24_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_21_12 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_9 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_057_ _057_/A VGND VGND VPWR VPWR _057_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_21_115 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xinput61 chany_bottom_in[19] VGND VGND VPWR VPWR input61/X sky130_fd_sc_hd__clkbuf_1
Xinput72 left_bottom_grid_pin_35_ VGND VGND VPWR VPWR input72/X sky130_fd_sc_hd__clkbuf_1
Xinput50 chanx_right_in[9] VGND VGND VPWR VPWR _067_/A sky130_fd_sc_hd__clkbuf_2
Xinput83 right_bottom_grid_pin_37_ VGND VGND VPWR VPWR input83/X sky130_fd_sc_hd__clkbuf_1
XFILLER_29_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_prog_clk_0_FTB00_A prog_clk_0_S_in VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mux_left_track_1.mux_l1_in_0__A0 _070_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mem_left_track_17.sky130_fd_sc_hd__dfxtp_1_0__CLK prog_clk_0_FTB00/X VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_12_115 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_12_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_16_78 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_32_88 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xmem_bottom_track_27.sky130_fd_sc_hd__dfxtp_1_0_ prog_clk_0_FTB00/X mux_bottom_track_25.mux_l3_in_0_/S
+ VGND VGND VPWR VPWR mux_bottom_track_27.mux_l1_in_0_/S sky130_fd_sc_hd__dfxtp_1
XANTENNA_input33_A chanx_right_in[11] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_109_ _109_/A VGND VGND VPWR VPWR _109_/X sky130_fd_sc_hd__clkbuf_1
Xmux_left_track_9.mux_l2_in_3_ mux_left_track_9.mux_l2_in_3_/A0 input78/X mux_left_track_9.mux_l2_in_3_/S
+ VGND VGND VPWR VPWR mux_left_track_9.mux_l2_in_3_/X sky130_fd_sc_hd__mux2_1
XANTENNA__070__A _070_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_27_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_27_66 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_27_33 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_27_22 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmux_right_track_0.mux_l2_in_3_ mux_right_track_0.mux_l2_in_3_/A0 _090_/A mux_right_track_0.mux_l2_in_3_/S
+ VGND VGND VPWR VPWR mux_right_track_0.mux_l2_in_3_/X sky130_fd_sc_hd__mux2_1
XFILLER_4_199 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmux_bottom_track_19.mux_l1_in_0_ input7/X _072_/A mux_bottom_track_19.mux_l1_in_1_/S
+ VGND VGND VPWR VPWR mux_bottom_track_19.mux_l1_in_0_/X sky130_fd_sc_hd__mux2_1
XFILLER_31_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_31_210 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_mux_right_track_0.mux_l2_in_0__S mux_right_track_0.mux_l2_in_3_/S VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
Xmux_bottom_track_21.mux_l1_in_0_ input8/X _074_/A mux_bottom_track_21.mux_l1_in_1_/S
+ VGND VGND VPWR VPWR mux_bottom_track_21.mux_l1_in_0_/X sky130_fd_sc_hd__mux2_1
XFILLER_13_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_22_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmem_bottom_track_5.sky130_fd_sc_hd__dfxtp_1_1_ prog_clk_0_FTB00/X mux_bottom_track_5.mux_l1_in_3_/S
+ VGND VGND VPWR VPWR mux_bottom_track_5.mux_l2_in_1_/S sky130_fd_sc_hd__dfxtp_1
XFILLER_13_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_191 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_090_ _090_/A VGND VGND VPWR VPWR _090_/X sky130_fd_sc_hd__clkbuf_1
XANTENNA_mem_bottom_track_7.sky130_fd_sc_hd__dfxtp_1_0__CLK prog_clk_0_FTB00/X VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_6_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xmux_left_track_9.mux_l4_in_0_ mux_left_track_9.mux_l3_in_1_/X mux_left_track_9.mux_l3_in_0_/X
+ mux_left_track_9.mux_l4_in_0_/S VGND VGND VPWR VPWR mux_left_track_9.mux_l4_in_0_/X
+ sky130_fd_sc_hd__mux2_1
XANTENNA_mux_bottom_track_21.mux_l1_in_0__A1 _074_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xmux_bottom_track_5.sky130_fd_sc_hd__buf_4_0_ mux_bottom_track_5.mux_l3_in_0_/X VGND
+ VGND VPWR VPWR _099_/A sky130_fd_sc_hd__clkbuf_1
Xinput4 bottom_left_grid_pin_44_ VGND VGND VPWR VPWR input4/X sky130_fd_sc_hd__clkbuf_1
XTAP_82 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_71 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_93 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xmux_right_track_0.mux_l4_in_0_ mux_right_track_0.mux_l3_in_1_/X mux_right_track_0.mux_l3_in_0_/X
+ mux_right_track_0.mux_l4_in_0_/S VGND VGND VPWR VPWR mux_right_track_0.mux_l4_in_0_/X
+ sky130_fd_sc_hd__mux2_1
XFILLER_10_14 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_10_25 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_10_36 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xmux_bottom_track_5.mux_l1_in_0_ input2/X _063_/A mux_bottom_track_5.mux_l1_in_3_/S
+ VGND VGND VPWR VPWR mux_bottom_track_5.mux_l1_in_0_/X sky130_fd_sc_hd__mux2_1
XFILLER_27_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_27_143 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_27_132 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_27_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_19_78 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_27_198 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_073_ _073_/A VGND VGND VPWR VPWR _073_/X sky130_fd_sc_hd__clkbuf_1
XANTENNA_input63_A chany_bottom_in[2] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mux_bottom_track_3.mux_l1_in_3__A1 _082_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_33_146 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_33_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_18_143 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_18_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_24_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmux_left_track_9.mux_l3_in_1_ mux_left_track_9.mux_l2_in_3_/X mux_left_track_9.mux_l2_in_2_/X
+ mux_left_track_9.mux_l3_in_1_/S VGND VGND VPWR VPWR mux_left_track_9.mux_l3_in_1_/X
+ sky130_fd_sc_hd__mux2_1
XFILLER_15_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_15_124 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_30_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_30_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_056_ _056_/A VGND VGND VPWR VPWR _056_/X sky130_fd_sc_hd__clkbuf_1
Xmux_right_track_0.mux_l3_in_1_ mux_right_track_0.mux_l2_in_3_/X mux_right_track_0.mux_l2_in_2_/X
+ mux_right_track_0.mux_l3_in_1_/S VGND VGND VPWR VPWR mux_right_track_0.mux_l3_in_1_/X
+ sky130_fd_sc_hd__mux2_1
XANTENNA_mux_right_track_0.mux_l2_in_3__S mux_right_track_0.mux_l2_in_3_/S VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
Xinput84 right_bottom_grid_pin_38_ VGND VGND VPWR VPWR input84/X sky130_fd_sc_hd__clkbuf_1
Xinput62 chany_bottom_in[1] VGND VGND VPWR VPWR input62/X sky130_fd_sc_hd__clkbuf_1
Xinput51 chany_bottom_in[0] VGND VGND VPWR VPWR input51/X sky130_fd_sc_hd__clkbuf_1
Xinput73 left_bottom_grid_pin_36_ VGND VGND VPWR VPWR input73/X sky130_fd_sc_hd__clkbuf_1
Xinput40 chanx_right_in[18] VGND VGND VPWR VPWR _076_/A sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_29_205 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_mux_left_track_1.mux_l1_in_0__A1 _060_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_16_46 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__068__A _068_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mux_left_track_1.mux_l3_in_1__S mux_left_track_1.mux_l3_in_1_/S VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_32_67 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_32_23 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_12_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_input26_A chanx_left_in[5] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_108_ _108_/A VGND VGND VPWR VPWR _108_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_7_186 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_11_160 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_11_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmux_left_track_17.mux_l1_in_3_ mux_left_track_17.mux_l1_in_3_/A0 input75/X mux_left_track_17.mux_l1_in_3_/S
+ VGND VGND VPWR VPWR mux_left_track_17.mux_l1_in_3_/X sky130_fd_sc_hd__mux2_1
Xmux_left_track_9.mux_l2_in_2_ input74/X input79/X mux_left_track_9.mux_l2_in_3_/S
+ VGND VGND VPWR VPWR mux_left_track_9.mux_l2_in_2_/X sky130_fd_sc_hd__mux2_1
XANTENNA_mem_left_track_3.sky130_fd_sc_hd__dfxtp_1_3__CLK prog_clk_0_FTB00/X VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_17_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_17_219 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_4_134 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xmux_right_track_0.mux_l2_in_2_ _080_/A input61/X mux_right_track_0.mux_l2_in_3_/S
+ VGND VGND VPWR VPWR mux_right_track_0.mux_l2_in_2_/X sky130_fd_sc_hd__mux2_1
XFILLER_1_104 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xmux_left_track_33.sky130_fd_sc_hd__buf_4_0_ mux_left_track_33.mux_l3_in_0_/X VGND
+ VGND VPWR VPWR _073_/A sky130_fd_sc_hd__clkbuf_1
Xmem_bottom_track_5.sky130_fd_sc_hd__dfxtp_1_0_ prog_clk_0_FTB00/X mem_bottom_track_5.delay_buf_2/X
+ VGND VGND VPWR VPWR mux_bottom_track_5.mux_l1_in_3_/S sky130_fd_sc_hd__dfxtp_2
XANTENNA__076__A _076_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_10_214 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_24_24 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xmux_left_track_17.mux_l3_in_0_ mux_left_track_17.mux_l2_in_1_/X mux_left_track_17.mux_l2_in_0_/X
+ mem_left_track_25.delay_buf_2/X VGND VGND VPWR VPWR mux_left_track_17.mux_l3_in_0_/X
+ sky130_fd_sc_hd__mux2_1
XANTENNA_mux_left_track_33.mux_l2_in_0__S mux_left_track_33.mux_l2_in_1_/S VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
Xinput5 bottom_left_grid_pin_45_ VGND VGND VPWR VPWR input5/X sky130_fd_sc_hd__clkbuf_1
XTAP_83 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_72 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_94 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_19_35 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_27_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_19_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_072_ _072_/A VGND VGND VPWR VPWR _072_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_2_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_input56_A chany_bottom_in[14] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_18_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_33_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_2_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmux_left_track_17.mux_l2_in_1_ mux_left_track_17.mux_l1_in_3_/X mux_left_track_17.mux_l1_in_2_/X
+ mux_left_track_17.mux_l2_in_1_/S VGND VGND VPWR VPWR mux_left_track_17.mux_l2_in_1_/X
+ sky130_fd_sc_hd__mux2_1
XFILLER_24_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_mem_right_track_4.sky130_fd_sc_hd__dfxtp_1_2__CLK prog_clk_0_FTB00/X VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_24_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmux_left_track_9.mux_l3_in_0_ mux_left_track_9.mux_l2_in_1_/X mux_left_track_9.mux_l2_in_0_/X
+ mux_left_track_9.mux_l3_in_1_/S VGND VGND VPWR VPWR mux_left_track_9.mux_l3_in_0_/X
+ sky130_fd_sc_hd__mux2_1
Xoutput150 _106_/X VGND VGND VPWR VPWR chany_bottom_out[9] sky130_fd_sc_hd__buf_2
XFILLER_30_128 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_30_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_30_106 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_15_103 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_15_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_15_158 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_7_49 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_7_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_mem_bottom_track_25.sky130_fd_sc_hd__dfxtp_1_0__CLK prog_clk_0_FTB00/X VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_23_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmux_right_track_0.mux_l3_in_0_ mux_right_track_0.mux_l2_in_1_/X mux_right_track_0.mux_l2_in_0_/X
+ mux_right_track_0.mux_l3_in_1_/S VGND VGND VPWR VPWR mux_right_track_0.mux_l3_in_0_/X
+ sky130_fd_sc_hd__mux2_1
XFILLER_14_191 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xinput63 chany_bottom_in[2] VGND VGND VPWR VPWR input63/X sky130_fd_sc_hd__clkbuf_1
Xinput74 left_bottom_grid_pin_37_ VGND VGND VPWR VPWR input74/X sky130_fd_sc_hd__dlymetal6s2s_1
Xinput52 chany_bottom_in[10] VGND VGND VPWR VPWR input52/X sky130_fd_sc_hd__clkbuf_1
Xinput85 right_bottom_grid_pin_39_ VGND VGND VPWR VPWR input85/X sky130_fd_sc_hd__clkbuf_1
Xinput30 chanx_left_in[9] VGND VGND VPWR VPWR _087_/A sky130_fd_sc_hd__dlymetal6s2s_1
Xinput41 chanx_right_in[19] VGND VGND VPWR VPWR input41/X sky130_fd_sc_hd__clkbuf_1
XANTENNA_mux_bottom_track_9.mux_l1_in_0__A0 input2/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_16_14 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_16_25 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_16_58 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_32_13 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__084__A _084_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_20_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_input19_A chanx_left_in[17] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mem_left_track_33.sky130_fd_sc_hd__dfxtp_1_1__CLK prog_clk_0_FTB00/X VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_107_ _107_/A VGND VGND VPWR VPWR _107_/X sky130_fd_sc_hd__clkbuf_1
Xmux_left_track_17.mux_l1_in_2_ input71/X input59/X mux_left_track_17.mux_l1_in_3_/S
+ VGND VGND VPWR VPWR mux_left_track_17.mux_l1_in_2_/X sky130_fd_sc_hd__mux2_1
XFILLER_7_198 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_14_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xmux_right_track_0.mux_l2_in_3__165 VGND VGND VPWR VPWR mux_right_track_0.mux_l2_in_3_/A0
+ mux_right_track_0.mux_l2_in_3__165/LO sky130_fd_sc_hd__conb_1
Xmux_left_track_9.mux_l2_in_1_ input58/X input70/X mux_left_track_9.mux_l2_in_3_/S
+ VGND VGND VPWR VPWR mux_left_track_9.mux_l2_in_1_/X sky130_fd_sc_hd__mux2_1
XFILLER_27_79 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_mux_bottom_track_7.mux_l1_in_2__A0 _084_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mem_bottom_track_17.sky130_fd_sc_hd__dfxtp_1_1__CLK prog_clk_0_FTB00/X VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_4_157 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xmux_right_track_0.mux_l2_in_1_ input54/X mux_right_track_0.mux_l1_in_2_/X mux_right_track_0.mux_l2_in_3_/S
+ VGND VGND VPWR VPWR mux_right_track_0.mux_l2_in_1_/X sky130_fd_sc_hd__mux2_1
XANTENNA_mem_left_track_9.sky130_fd_sc_hd__dfxtp_1_2__D mux_left_track_9.mux_l2_in_3_/S
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mem_left_track_25.sky130_fd_sc_hd__dfxtp_1_2__CLK prog_clk_0_FTB00/X VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_input86_A right_bottom_grid_pin_40_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mux_bottom_track_15.mux_l1_in_1__A1 _090_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mem_right_track_8.sky130_fd_sc_hd__dfxtp_1_2__D mux_right_track_8.mux_l2_in_3_/S
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xmux_right_track_0.mux_l1_in_2_ input66/X input87/X mux_right_track_0.mux_l1_in_2_/S
+ VGND VGND VPWR VPWR mux_right_track_0.mux_l1_in_2_/X sky130_fd_sc_hd__mux2_1
XANTENNA__092__A _092_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xmem_bottom_track_13.sky130_fd_sc_hd__dfxtp_1_1_ prog_clk_0_FTB00/X mux_bottom_track_13.mux_l1_in_1_/S
+ VGND VGND VPWR VPWR mux_bottom_track_13.mux_l2_in_0_/S sky130_fd_sc_hd__dfxtp_1
Xinput6 bottom_left_grid_pin_46_ VGND VGND VPWR VPWR input6/X sky130_fd_sc_hd__clkbuf_1
XTAP_84 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_73 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_95 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_19_14 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_19_25 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__087__A _087_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mem_bottom_track_1.sky130_fd_sc_hd__dfxtp_1_1__CLK prog_clk_0_FTB00/X VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_071_ _071_/A VGND VGND VPWR VPWR _071_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_2_211 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_input49_A chanx_right_in[8] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_18_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_18_134 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_33_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_33_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_2_50 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xmux_left_track_17.mux_l2_in_0_ mux_left_track_17.mux_l1_in_1_/X mux_left_track_17.mux_l1_in_0_/X
+ mux_left_track_17.mux_l2_in_1_/S VGND VGND VPWR VPWR mux_left_track_17.mux_l2_in_0_/X
+ sky130_fd_sc_hd__mux2_1
XFILLER_32_192 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xmux_right_track_24.mux_l1_in_3_ mux_right_track_24.mux_l1_in_3_/A0 _096_/A mux_right_track_24.mux_l1_in_3_/S
+ VGND VGND VPWR VPWR mux_right_track_24.mux_l1_in_3_/X sky130_fd_sc_hd__mux2_1
Xoutput140 _115_/X VGND VGND VPWR VPWR chany_bottom_out[18] sky130_fd_sc_hd__buf_2
XFILLER_21_59 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xinput31 chanx_right_in[0] VGND VGND VPWR VPWR _115_/A sky130_fd_sc_hd__clkbuf_1
Xinput20 chanx_left_in[18] VGND VGND VPWR VPWR _096_/A sky130_fd_sc_hd__clkbuf_2
Xinput86 right_bottom_grid_pin_40_ VGND VGND VPWR VPWR input86/X sky130_fd_sc_hd__clkbuf_1
Xinput53 chany_bottom_in[11] VGND VGND VPWR VPWR input53/X sky130_fd_sc_hd__clkbuf_1
Xinput64 chany_bottom_in[3] VGND VGND VPWR VPWR input64/X sky130_fd_sc_hd__clkbuf_1
Xinput75 left_bottom_grid_pin_38_ VGND VGND VPWR VPWR input75/X sky130_fd_sc_hd__clkbuf_1
Xinput42 chanx_right_in[1] VGND VGND VPWR VPWR _114_/A sky130_fd_sc_hd__clkbuf_1
XANTENNA_mux_bottom_track_9.mux_l1_in_0__A1 _066_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_32_58 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_20_151 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_7_122 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_106_ _106_/A VGND VGND VPWR VPWR _106_/X sky130_fd_sc_hd__clkbuf_1
Xmux_left_track_17.mux_l1_in_1_ input52/X input64/X mux_left_track_17.mux_l1_in_3_/S
+ VGND VGND VPWR VPWR mux_left_track_17.mux_l1_in_1_/X sky130_fd_sc_hd__mux2_1
XFILLER_7_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmux_left_track_9.mux_l2_in_0_ input63/X mux_left_track_9.mux_l1_in_0_/X mux_left_track_9.mux_l2_in_3_/S
+ VGND VGND VPWR VPWR mux_left_track_9.mux_l2_in_0_/X sky130_fd_sc_hd__mux2_1
XFILLER_8_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_25_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__095__A _095_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mux_bottom_track_7.mux_l1_in_2__A1 input9/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_4_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_4_103 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmux_right_track_0.mux_l2_in_0_ mux_right_track_0.mux_l1_in_1_/X mux_right_track_0.mux_l1_in_0_/X
+ mux_right_track_0.mux_l2_in_3_/S VGND VGND VPWR VPWR mux_right_track_0.mux_l2_in_0_/X
+ sky130_fd_sc_hd__mux2_1
XANTENNA_mux_bottom_track_23.mux_l1_in_1__A1 _095_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_input31_A chanx_right_in[0] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xmux_right_track_24.mux_l3_in_0_ mux_right_track_24.mux_l2_in_1_/X mux_right_track_24.mux_l2_in_0_/X
+ mux_right_track_24.mux_l3_in_0_/S VGND VGND VPWR VPWR mux_right_track_24.mux_l3_in_0_/X
+ sky130_fd_sc_hd__mux2_1
XFILLER_16_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_17_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_33_90 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_13_16 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_13_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_13_38 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_13_49 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_input79_A left_top_grid_pin_1_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_5_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_24_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_6_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmux_right_track_0.mux_l1_in_1_ input85/X input83/X mux_right_track_0.mux_l1_in_2_/S
+ VGND VGND VPWR VPWR mux_right_track_0.mux_l1_in_1_/X sky130_fd_sc_hd__mux2_1
XANTENNA_mem_left_track_1.sky130_fd_sc_hd__dfxtp_1_2__D mux_left_track_1.mux_l2_in_3_/S
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xmem_bottom_track_13.sky130_fd_sc_hd__dfxtp_1_0_ prog_clk_0_FTB00/X mux_bottom_track_11.mux_l3_in_0_/S
+ VGND VGND VPWR VPWR mux_bottom_track_13.mux_l1_in_1_/S sky130_fd_sc_hd__dfxtp_1
Xmux_right_track_24.mux_l2_in_1_ mux_right_track_24.mux_l1_in_3_/X mux_right_track_24.mux_l1_in_2_/X
+ mux_right_track_24.mux_l2_in_1_/S VGND VGND VPWR VPWR mux_right_track_24.mux_l2_in_1_/X
+ sky130_fd_sc_hd__mux2_1
XFILLER_30_91 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_85 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_74 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xinput7 bottom_left_grid_pin_47_ VGND VGND VPWR VPWR input7/X sky130_fd_sc_hd__dlymetal6s2s_1
XTAP_96 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_070_ _070_/A VGND VGND VPWR VPWR _070_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_2_201 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_mem_right_track_0.sky130_fd_sc_hd__dfxtp_1_2__D mux_right_track_0.mux_l2_in_3_/S
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mux_bottom_track_1.mux_l1_in_0__S mux_bottom_track_1.mux_l1_in_3_/S VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_25_91 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_mem_left_track_1.sky130_fd_sc_hd__dfxtp_1_1__CLK prog_clk_0_FTB00/X VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_24_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_24_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_32_182 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_32_171 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_32_160 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmux_right_track_24.mux_l1_in_2_ _087_/A input56/X mux_right_track_24.mux_l1_in_3_/S
+ VGND VGND VPWR VPWR mux_right_track_24.mux_l1_in_2_/X sky130_fd_sc_hd__mux2_1
XFILLER_21_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xoutput130 _086_/X VGND VGND VPWR VPWR chanx_right_out[9] sky130_fd_sc_hd__buf_2
Xoutput141 _116_/X VGND VGND VPWR VPWR chany_bottom_out[19] sky130_fd_sc_hd__buf_2
XFILLER_15_116 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_mux_bottom_track_19.mux_l1_in_0__A0 input7/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_23_171 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_input61_A chany_bottom_in[19] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xmem_bottom_track_19.sky130_fd_sc_hd__dfxtp_1_1_ prog_clk_0_FTB00/X mux_bottom_track_19.mux_l1_in_1_/S
+ VGND VGND VPWR VPWR mux_bottom_track_19.mux_l2_in_0_/S sky130_fd_sc_hd__dfxtp_1
Xmem_right_track_32.sky130_fd_sc_hd__dfxtp_1_2_ prog_clk_0_FTB00/X mux_right_track_32.mux_l2_in_1_/S
+ VGND VGND VPWR VPWR mem_bottom_track_1.delay_buf_2/X sky130_fd_sc_hd__dfxtp_1
Xinput10 ccff_head VGND VGND VPWR VPWR input10/X sky130_fd_sc_hd__dlymetal6s2s_1
Xinput54 chany_bottom_in[12] VGND VGND VPWR VPWR input54/X sky130_fd_sc_hd__dlymetal6s2s_1
Xinput43 chanx_right_in[2] VGND VGND VPWR VPWR _060_/A sky130_fd_sc_hd__clkbuf_2
Xinput32 chanx_right_in[10] VGND VGND VPWR VPWR _068_/A sky130_fd_sc_hd__dlymetal6s2s_1
Xinput21 chanx_left_in[19] VGND VGND VPWR VPWR input21/X sky130_fd_sc_hd__clkbuf_1
XFILLER_21_119 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xinput87 right_bottom_grid_pin_41_ VGND VGND VPWR VPWR input87/X sky130_fd_sc_hd__clkbuf_1
Xinput65 chany_bottom_in[4] VGND VGND VPWR VPWR input65/X sky130_fd_sc_hd__clkbuf_1
Xinput76 left_bottom_grid_pin_39_ VGND VGND VPWR VPWR input76/X sky130_fd_sc_hd__clkbuf_1
X_105_ _105_/A VGND VGND VPWR VPWR _105_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_7_145 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_11_152 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_11_185 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_mem_right_track_24.sky130_fd_sc_hd__dfxtp_1_2__D mux_right_track_24.mux_l2_in_1_/S
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xmux_left_track_17.mux_l1_in_0_ _075_/A _066_/A mux_left_track_17.mux_l1_in_3_/S VGND
+ VGND VPWR VPWR mux_left_track_17.mux_l1_in_0_/X sky130_fd_sc_hd__mux2_1
XANTENNA_mux_right_track_16.mux_l1_in_0__S mux_right_track_16.mux_l1_in_3_/S VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mux_left_track_1.mux_l2_in_2__A1 input74/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xmux_bottom_track_7.mux_l1_in_3__156 VGND VGND VPWR VPWR mux_bottom_track_7.mux_l1_in_3_/A0
+ mux_bottom_track_7.mux_l1_in_3__156/LO sky130_fd_sc_hd__conb_1
XFILLER_27_37 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_25_200 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_4_126 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_input24_A chanx_left_in[3] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xmux_right_track_0.sky130_fd_sc_hd__buf_4_0_ mux_right_track_0.mux_l4_in_0_/X VGND
+ VGND VPWR VPWR _077_/A sky130_fd_sc_hd__clkbuf_1
XFILLER_1_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmux_bottom_track_1.mux_l1_in_3_ mux_bottom_track_1.mux_l1_in_3_/A0 _080_/A mux_bottom_track_1.mux_l1_in_3_/S
+ VGND VGND VPWR VPWR mux_bottom_track_1.mux_l1_in_3_/X sky130_fd_sc_hd__mux2_1
XFILLER_13_203 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_mem_bottom_track_11.sky130_fd_sc_hd__dfxtp_1_2__CLK prog_clk_0_FTB00/X VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xmux_left_track_9.mux_l1_in_0_ _074_/A _064_/A mux_left_track_9.mux_l1_in_0_/S VGND
+ VGND VPWR VPWR mux_left_track_9.mux_l1_in_0_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_151 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_28_91 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_173 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_mux_bottom_track_1.mux_l1_in_3__S mux_bottom_track_1.mux_l1_in_3_/S VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_5_40 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_mem_right_track_2.sky130_fd_sc_hd__dfxtp_1_0__CLK prog_clk_0_FTB00/X VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xmux_bottom_track_13.sky130_fd_sc_hd__buf_4_0_ mux_bottom_track_13.mux_l2_in_0_/X
+ VGND VGND VPWR VPWR _103_/A sky130_fd_sc_hd__clkbuf_1
Xmux_right_track_0.mux_l1_in_0_ input81/X input88/X mux_right_track_0.mux_l1_in_2_/S
+ VGND VGND VPWR VPWR mux_right_track_0.mux_l1_in_0_/X sky130_fd_sc_hd__mux2_1
XFILLER_24_38 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xmux_right_track_24.mux_l2_in_0_ mux_right_track_24.mux_l1_in_1_/X mux_right_track_24.mux_l1_in_0_/X
+ mux_right_track_24.mux_l2_in_1_/S VGND VGND VPWR VPWR mux_right_track_24.mux_l2_in_0_/X
+ sky130_fd_sc_hd__mux2_1
XFILLER_14_71 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_30_70 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_5_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_14_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xinput8 bottom_left_grid_pin_48_ VGND VGND VPWR VPWR input8/X sky130_fd_sc_hd__dlymetal6s2s_1
XTAP_86 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_75 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_97 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xmem_left_track_3.sky130_fd_sc_hd__dfxtp_1_3_ prog_clk_0_FTB00/X mux_left_track_3.mux_l3_in_1_/S
+ VGND VGND VPWR VPWR mux_left_track_3.mux_l4_in_0_/S sky130_fd_sc_hd__dfxtp_1
XANTENNA_mux_bottom_track_27.mux_l1_in_0__A0 input3/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_33_106 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_18_103 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_18_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_18_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_mux_right_track_8.mux_l2_in_3__A1 _094_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mux_right_track_16.mux_l1_in_3__S mux_right_track_16.mux_l1_in_3_/S VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xmux_bottom_track_1.mux_l3_in_0_ mux_bottom_track_1.mux_l2_in_1_/X mux_bottom_track_1.mux_l2_in_0_/X
+ mem_bottom_track_3.delay_buf_2/X VGND VGND VPWR VPWR mux_bottom_track_1.mux_l3_in_0_/X
+ sky130_fd_sc_hd__mux2_1
Xmux_right_track_24.mux_l1_in_1_ input68/X input51/X mux_right_track_24.mux_l1_in_3_/S
+ VGND VGND VPWR VPWR mux_right_track_24.mux_l1_in_1_/X sky130_fd_sc_hd__mux2_1
XFILLER_24_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_mux_left_track_17.mux_l1_in_0__A0 _075_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_21_17 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xoutput120 _095_/X VGND VGND VPWR VPWR chanx_right_out[18] sky130_fd_sc_hd__buf_2
Xoutput142 _098_/X VGND VGND VPWR VPWR chany_bottom_out[1] sky130_fd_sc_hd__buf_2
Xoutput131 _097_/X VGND VGND VPWR VPWR chany_bottom_out[0] sky130_fd_sc_hd__buf_2
XFILLER_15_128 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_mux_bottom_track_19.mux_l1_in_0__A1 _072_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_input54_A chany_bottom_in[12] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xmem_bottom_track_19.sky130_fd_sc_hd__dfxtp_1_0_ prog_clk_0_FTB00/X mux_bottom_track_17.mux_l2_in_0_/S
+ VGND VGND VPWR VPWR mux_bottom_track_19.mux_l1_in_1_/S sky130_fd_sc_hd__dfxtp_1
Xmem_right_track_32.sky130_fd_sc_hd__dfxtp_1_1_ prog_clk_0_FTB00/X mux_right_track_32.mux_l1_in_1_/S
+ VGND VGND VPWR VPWR mux_right_track_32.mux_l2_in_1_/S sky130_fd_sc_hd__dfxtp_1
Xinput88 right_top_grid_pin_1_ VGND VGND VPWR VPWR input88/X sky130_fd_sc_hd__clkbuf_1
Xinput77 left_bottom_grid_pin_40_ VGND VGND VPWR VPWR input77/X sky130_fd_sc_hd__clkbuf_1
Xinput22 chanx_left_in[1] VGND VGND VPWR VPWR input22/X sky130_fd_sc_hd__clkbuf_1
Xinput11 chanx_left_in[0] VGND VGND VPWR VPWR _116_/A sky130_fd_sc_hd__clkbuf_1
Xinput55 chany_bottom_in[13] VGND VGND VPWR VPWR input55/X sky130_fd_sc_hd__clkbuf_1
Xinput66 chany_bottom_in[5] VGND VGND VPWR VPWR input66/X sky130_fd_sc_hd__dlymetal6s2s_1
Xinput44 chanx_right_in[3] VGND VGND VPWR VPWR _113_/A sky130_fd_sc_hd__clkbuf_1
Xinput33 chanx_right_in[11] VGND VGND VPWR VPWR _111_/A sky130_fd_sc_hd__clkbuf_1
XFILLER_14_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_mem_right_track_8.sky130_fd_sc_hd__dfxtp_1_2__CLK prog_clk_0_FTB00/X VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_32_38 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_32_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_12_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_104_ _104_/A VGND VGND VPWR VPWR _104_/X sky130_fd_sc_hd__clkbuf_1
Xmux_bottom_track_1.mux_l2_in_1_ mux_bottom_track_1.mux_l1_in_3_/X mux_bottom_track_1.mux_l1_in_2_/X
+ mux_bottom_track_1.mux_l2_in_1_/S VGND VGND VPWR VPWR mux_bottom_track_1.mux_l2_in_1_/X
+ sky130_fd_sc_hd__mux2_1
XFILLER_11_142 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_11_164 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_22_60 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_22_71 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmux_right_track_8.mux_l2_in_3__171 VGND VGND VPWR VPWR mux_right_track_8.mux_l2_in_3_/A0
+ mux_right_track_8.mux_l2_in_3__171/LO sky130_fd_sc_hd__conb_1
XFILLER_21_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmux_left_track_5.mux_l1_in_6_ input78/X input77/X repeater153/X VGND VGND VPWR VPWR
+ mux_left_track_5.mux_l1_in_6_/X sky130_fd_sc_hd__mux2_1
XFILLER_4_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_input17_A chanx_left_in[15] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_31_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_22_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_input9_A bottom_left_grid_pin_49_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xmux_bottom_track_1.mux_l1_in_2_ input22/X input8/X mux_bottom_track_1.mux_l1_in_3_/S
+ VGND VGND VPWR VPWR mux_bottom_track_1.mux_l1_in_2_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_185 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_163 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_5_30 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmem_right_track_0.sky130_fd_sc_hd__dfxtp_1_3_ prog_clk_0_FTB00/X mux_right_track_0.mux_l3_in_1_/S
+ VGND VGND VPWR VPWR mux_right_track_0.mux_l4_in_0_/S sky130_fd_sc_hd__dfxtp_1
XANTENNA_input84_A right_bottom_grid_pin_38_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_30_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xinput9 bottom_left_grid_pin_49_ VGND VGND VPWR VPWR input9/X sky130_fd_sc_hd__dlymetal6s2s_1
XTAP_87 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xmem_left_track_3.sky130_fd_sc_hd__dfxtp_1_2_ prog_clk_0_FTB00/X mux_left_track_3.mux_l2_in_3_/S
+ VGND VGND VPWR VPWR mux_left_track_3.mux_l3_in_1_/S sky130_fd_sc_hd__dfxtp_1
XTAP_76 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_98 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_mux_right_track_2.mux_l2_in_2__S mux_right_track_2.mux_l2_in_3_/S VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mux_left_track_25.mux_l1_in_0__A0 _076_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xmux_bottom_track_15.mux_l2_in_0_ mux_bottom_track_15.mux_l1_in_1_/X mux_bottom_track_15.mux_l1_in_0_/X
+ mux_bottom_track_15.mux_l2_in_0_/S VGND VGND VPWR VPWR mux_bottom_track_15.mux_l2_in_0_/X
+ sky130_fd_sc_hd__mux2_1
XFILLER_27_115 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_19_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_18_115 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_33_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_33_118 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_60 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_26_192 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_18_126 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_mux_left_track_9.mux_l2_in_1__S mux_left_track_9.mux_l2_in_3_/S VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mem_left_track_3.sky130_fd_sc_hd__dfxtp_1_0__D mux_left_track_1.mux_l4_in_0_/S
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_2_75 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_2_64 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_mux_left_track_17.mux_l1_in_0__A1 _066_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xmux_right_track_24.mux_l1_in_0_ input85/X input81/X mux_right_track_24.mux_l1_in_3_/S
+ VGND VGND VPWR VPWR mux_right_track_24.mux_l1_in_0_/X sky130_fd_sc_hd__mux2_1
XFILLER_24_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xoutput121 _096_/X VGND VGND VPWR VPWR chanx_right_out[19] sky130_fd_sc_hd__buf_2
Xoutput110 _066_/X VGND VGND VPWR VPWR chanx_left_out[9] sky130_fd_sc_hd__buf_2
Xoutput132 _107_/X VGND VGND VPWR VPWR chany_bottom_out[10] sky130_fd_sc_hd__buf_2
Xoutput143 _099_/X VGND VGND VPWR VPWR chany_bottom_out[2] sky130_fd_sc_hd__buf_2
XANTENNA_mem_bottom_track_5.sky130_fd_sc_hd__dfxtp_1_1__CLK prog_clk_0_FTB00/X VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mux_right_track_16.mux_l1_in_3__A1 _095_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_15_107 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_11_84 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_input47_A chanx_right_in[6] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xmem_right_track_32.sky130_fd_sc_hd__dfxtp_1_0_ prog_clk_0_FTB00/X mux_right_track_24.mux_l3_in_0_/S
+ VGND VGND VPWR VPWR mux_right_track_32.mux_l1_in_1_/S sky130_fd_sc_hd__dfxtp_1
XFILLER_14_151 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmux_bottom_track_15.mux_l1_in_1_ mux_bottom_track_15.mux_l1_in_1_/A0 _090_/A mux_bottom_track_15.mux_l1_in_1_/S
+ VGND VGND VPWR VPWR mux_bottom_track_15.mux_l1_in_1_/X sky130_fd_sc_hd__mux2_1
Xinput23 chanx_left_in[2] VGND VGND VPWR VPWR _080_/A sky130_fd_sc_hd__clkbuf_2
Xinput67 chany_bottom_in[6] VGND VGND VPWR VPWR input67/X sky130_fd_sc_hd__clkbuf_1
Xinput78 left_bottom_grid_pin_41_ VGND VGND VPWR VPWR input78/X sky130_fd_sc_hd__dlymetal6s2s_1
Xinput56 chany_bottom_in[14] VGND VGND VPWR VPWR input56/X sky130_fd_sc_hd__dlymetal6s2s_1
Xinput45 chanx_right_in[4] VGND VGND VPWR VPWR _062_/A sky130_fd_sc_hd__dlymetal6s2s_1
Xinput12 chanx_left_in[10] VGND VGND VPWR VPWR _088_/A sky130_fd_sc_hd__clkbuf_2
Xinput34 chanx_right_in[12] VGND VGND VPWR VPWR _070_/A sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_20_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_20_143 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_20_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_20_176 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmem_left_track_9.sky130_fd_sc_hd__dfxtp_1_3_ prog_clk_0_FTB00/X mux_left_track_9.mux_l3_in_1_/S
+ VGND VGND VPWR VPWR mux_left_track_9.mux_l4_in_0_/S sky130_fd_sc_hd__dfxtp_1
XFILLER_28_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_11_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_103_ _103_/A VGND VGND VPWR VPWR _103_/X sky130_fd_sc_hd__clkbuf_1
Xmux_bottom_track_1.mux_l2_in_0_ mux_bottom_track_1.mux_l1_in_1_/X mux_bottom_track_1.mux_l1_in_0_/X
+ mux_bottom_track_1.mux_l2_in_1_/S VGND VGND VPWR VPWR mux_bottom_track_1.mux_l2_in_0_/X
+ sky130_fd_sc_hd__mux2_1
XFILLER_22_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xmux_left_track_5.mux_l1_in_5_ input76/X input75/X repeater154/X VGND VGND VPWR VPWR
+ mux_left_track_5.mux_l1_in_5_/X sky130_fd_sc_hd__mux2_1
XFILLER_19_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_8_52 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_8_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_mux_bottom_track_25.mux_l2_in_1__A1 _096_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_17_72 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_mux_right_track_24.mux_l1_in_1__S mux_right_track_24.mux_l1_in_3_/S VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mux_left_track_5.mux_l1_in_2__A1 input57/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_1_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xmux_bottom_track_1.mux_l1_in_1_ input6/X input4/X mux_bottom_track_1.mux_l1_in_3_/S
+ VGND VGND VPWR VPWR mux_bottom_track_1.mux_l1_in_1_/X sky130_fd_sc_hd__mux2_1
XANTENNA_mux_left_track_33.mux_l1_in_0__A0 input66/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_28_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_28_71 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_5_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_5_20 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmem_right_track_0.sky130_fd_sc_hd__dfxtp_1_2_ prog_clk_0_FTB00/X mux_right_track_0.mux_l2_in_3_/S
+ VGND VGND VPWR VPWR mux_right_track_0.mux_l3_in_1_/S sky130_fd_sc_hd__dfxtp_1
XFILLER_30_50 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_input77_A left_bottom_grid_pin_40_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_88 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_77 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xmem_left_track_3.sky130_fd_sc_hd__dfxtp_1_1_ prog_clk_0_FTB00/X mux_left_track_3.mux_l1_in_1_/S
+ VGND VGND VPWR VPWR mux_left_track_3.mux_l2_in_3_/S sky130_fd_sc_hd__dfxtp_1
XTAP_99 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_mux_left_track_25.mux_l1_in_0__A1 _067_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mux_right_track_24.mux_l1_in_3__A1 _096_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_27_127 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_18_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_61 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_25_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_25_72 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_25_61 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_50 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_mux_right_track_0.mux_l1_in_2__A0 input66/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_2_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_17_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xoutput100 _075_/X VGND VGND VPWR VPWR chanx_left_out[18] sky130_fd_sc_hd__buf_2
Xoutput144 _100_/X VGND VGND VPWR VPWR chany_bottom_out[3] sky130_fd_sc_hd__buf_2
Xoutput133 _108_/X VGND VGND VPWR VPWR chany_bottom_out[11] sky130_fd_sc_hd__buf_2
Xmux_left_track_5.mux_l2_in_3_ mux_left_track_5.mux_l2_in_3_/A0 mux_left_track_5.mux_l1_in_6_/X
+ mux_left_track_5.mux_l2_in_3_/S VGND VGND VPWR VPWR mux_left_track_5.mux_l2_in_3_/X
+ sky130_fd_sc_hd__mux2_1
Xoutput111 _077_/X VGND VGND VPWR VPWR chanx_right_out[0] sky130_fd_sc_hd__buf_2
Xoutput122 _078_/X VGND VGND VPWR VPWR chanx_right_out[1] sky130_fd_sc_hd__buf_2
XFILLER_23_163 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_2_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_11_63 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_11_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_mem_left_track_5.sky130_fd_sc_hd__dfxtp_1_1__CLK prog_clk_0_FTB00/X VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xinput13 chanx_left_in[11] VGND VGND VPWR VPWR input13/X sky130_fd_sc_hd__clkbuf_1
Xmux_bottom_track_15.mux_l1_in_0_ input5/X _070_/A mux_bottom_track_15.mux_l1_in_1_/S
+ VGND VGND VPWR VPWR mux_bottom_track_15.mux_l1_in_0_/X sky130_fd_sc_hd__mux2_1
Xinput79 left_top_grid_pin_1_ VGND VGND VPWR VPWR input79/X sky130_fd_sc_hd__clkbuf_1
Xinput24 chanx_left_in[3] VGND VGND VPWR VPWR input24/X sky130_fd_sc_hd__clkbuf_1
Xinput46 chanx_right_in[5] VGND VGND VPWR VPWR _063_/A sky130_fd_sc_hd__clkbuf_2
Xinput68 chany_bottom_in[7] VGND VGND VPWR VPWR input68/X sky130_fd_sc_hd__clkbuf_1
Xinput57 chany_bottom_in[15] VGND VGND VPWR VPWR input57/X sky130_fd_sc_hd__clkbuf_2
Xinput35 chanx_right_in[13] VGND VGND VPWR VPWR _071_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_32_18 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmux_bottom_track_27.mux_l2_in_0_ mux_bottom_track_27.mux_l2_in_0_/A0 mux_bottom_track_27.mux_l1_in_0_/X
+ mux_bottom_track_27.mux_l2_in_0_/S VGND VGND VPWR VPWR mux_bottom_track_27.mux_l2_in_0_/X
+ sky130_fd_sc_hd__mux2_1
XFILLER_20_199 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xmem_left_track_9.sky130_fd_sc_hd__dfxtp_1_2_ prog_clk_0_FTB00/X mux_left_track_9.mux_l2_in_3_/S
+ VGND VGND VPWR VPWR mux_left_track_9.mux_l3_in_1_/S sky130_fd_sc_hd__dfxtp_1
XANTENNA_mux_right_track_0.mux_l2_in_1__A0 input54/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xmux_bottom_track_1.sky130_fd_sc_hd__buf_4_0_ mux_bottom_track_1.mux_l3_in_0_/X VGND
+ VGND VPWR VPWR _097_/A sky130_fd_sc_hd__clkbuf_1
XFILLER_7_104 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_mux_left_track_17.mux_l1_in_1__S mux_left_track_17.mux_l1_in_3_/S VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
X_102_ _102_/A VGND VGND VPWR VPWR _102_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_7_115 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_7_126 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_mux_right_track_16.mux_l2_in_1__S mux_right_track_16.mux_l2_in_1_/S VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xmux_left_track_5.mux_l1_in_4_ input74/X input73/X repeater153/X VGND VGND VPWR VPWR
+ mux_left_track_5.mux_l1_in_4_/X sky130_fd_sc_hd__mux2_1
XFILLER_8_42 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_mem_right_track_2.sky130_fd_sc_hd__dfxtp_1_3__CLK prog_clk_0_FTB00/X VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mux_left_track_1.mux_l1_in_0__S mux_left_track_1.mux_l1_in_1_/S VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mem_bottom_track_23.sky130_fd_sc_hd__dfxtp_1_1__CLK prog_clk_0_FTB00/X VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_31_206 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_16_214 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_17_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_17_84 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_33_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xmux_left_track_5.mux_l4_in_0_ mux_left_track_5.mux_l3_in_1_/X mux_left_track_5.mux_l3_in_0_/X
+ mux_left_track_5.mux_l4_in_0_/S VGND VGND VPWR VPWR mux_left_track_5.mux_l4_in_0_/X
+ sky130_fd_sc_hd__mux2_1
Xmux_bottom_track_1.mux_l1_in_0_ input2/X _060_/A mux_bottom_track_1.mux_l1_in_3_/S
+ VGND VGND VPWR VPWR mux_bottom_track_1.mux_l1_in_0_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_input22_A chanx_left_in[1] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mux_left_track_33.mux_l1_in_0__A1 _068_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_output90_A output90/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_8_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmem_right_track_0.sky130_fd_sc_hd__dfxtp_1_1_ prog_clk_0_FTB00/X mux_right_track_0.mux_l1_in_2_/S
+ VGND VGND VPWR VPWR mux_right_track_0.mux_l2_in_3_/S sky130_fd_sc_hd__dfxtp_2
Xmux_left_track_5.mux_l3_in_1_ mux_left_track_5.mux_l2_in_3_/X mux_left_track_5.mux_l2_in_2_/X
+ mux_left_track_5.mux_l3_in_1_/S VGND VGND VPWR VPWR mux_left_track_5.mux_l3_in_1_/X
+ sky130_fd_sc_hd__mux2_1
XFILLER_30_95 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_30_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_29_191 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_89 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_78 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xmem_left_track_3.sky130_fd_sc_hd__dfxtp_1_0_ prog_clk_0_FTB00/X mux_left_track_1.mux_l4_in_0_/S
+ VGND VGND VPWR VPWR mux_left_track_3.mux_l1_in_1_/S sky130_fd_sc_hd__dfxtp_1
XFILLER_27_106 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_26_172 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_25_95 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_40 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_25_40 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_24_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xoutput101 _076_/X VGND VGND VPWR VPWR chanx_left_out[19] sky130_fd_sc_hd__buf_2
Xoutput112 _087_/X VGND VGND VPWR VPWR chanx_right_out[10] sky130_fd_sc_hd__buf_2
Xoutput134 _109_/X VGND VGND VPWR VPWR chany_bottom_out[12] sky130_fd_sc_hd__buf_2
Xoutput145 _101_/X VGND VGND VPWR VPWR chany_bottom_out[4] sky130_fd_sc_hd__buf_2
Xmux_left_track_5.mux_l2_in_2_ mux_left_track_5.mux_l1_in_5_/X mux_left_track_5.mux_l1_in_4_/X
+ mux_left_track_5.mux_l2_in_3_/S VGND VGND VPWR VPWR mux_left_track_5.mux_l2_in_2_/X
+ sky130_fd_sc_hd__mux2_1
Xoutput123 _079_/X VGND VGND VPWR VPWR chanx_right_out[2] sky130_fd_sc_hd__buf_2
XFILLER_23_175 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_23_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_11_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xinput25 chanx_left_in[4] VGND VGND VPWR VPWR _082_/A sky130_fd_sc_hd__clkbuf_2
Xinput14 chanx_left_in[12] VGND VGND VPWR VPWR _090_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_14_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xinput36 chanx_right_in[14] VGND VGND VPWR VPWR _072_/A sky130_fd_sc_hd__clkbuf_2
Xinput58 chany_bottom_in[16] VGND VGND VPWR VPWR input58/X sky130_fd_sc_hd__clkbuf_1
Xinput69 chany_bottom_in[8] VGND VGND VPWR VPWR input69/X sky130_fd_sc_hd__clkbuf_1
Xinput47 chanx_right_in[6] VGND VGND VPWR VPWR _064_/A sky130_fd_sc_hd__clkbuf_2
XANTENNA_mux_left_track_5.mux_l2_in_1__S mux_left_track_5.mux_l2_in_3_/S VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_20_101 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_9_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xmem_left_track_9.sky130_fd_sc_hd__dfxtp_1_1_ prog_clk_0_FTB00/X mux_left_track_9.mux_l1_in_0_/S
+ VGND VGND VPWR VPWR mux_left_track_9.mux_l2_in_3_/S sky130_fd_sc_hd__dfxtp_2
XFILLER_20_134 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_mux_left_track_9.mux_l2_in_0__A0 input63/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mux_right_track_8.mux_l2_in_1__S mux_right_track_8.mux_l2_in_3_/S VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
X_101_ _101_/A VGND VGND VPWR VPWR _101_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_11_134 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_11_156 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_11_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_22_52 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_input52_A chany_bottom_in[10] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_22_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_19_201 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xmux_left_track_5.mux_l1_in_3_ input72/X input71/X repeater154/X VGND VGND VPWR VPWR
+ mux_left_track_5.mux_l1_in_3_/X sky130_fd_sc_hd__mux2_1
XANTENNA_mux_bottom_track_1.mux_l1_in_1__A0 input6/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_6_171 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_4_108 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_33_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_3_185 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_mux_bottom_track_23.sky130_fd_sc_hd__buf_4_0__A mux_bottom_track_23.mux_l2_in_0_/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xmux_bottom_track_27.mux_l1_in_0_ input3/X input37/X mux_bottom_track_27.mux_l1_in_0_/S
+ VGND VGND VPWR VPWR mux_bottom_track_27.mux_l1_in_0_/X sky130_fd_sc_hd__mux2_1
Xmux_left_track_17.sky130_fd_sc_hd__buf_4_0_ mux_left_track_17.mux_l3_in_0_/X VGND
+ VGND VPWR VPWR _065_/A sky130_fd_sc_hd__clkbuf_1
XFILLER_0_122 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_28_40 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_input15_A chanx_left_in[13] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_10_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmem_right_track_0.sky130_fd_sc_hd__dfxtp_1_0_ prog_clk_0_FTB00/X input10/X VGND VGND
+ VPWR VPWR mux_right_track_0.mux_l1_in_2_/S sky130_fd_sc_hd__dfxtp_1
XANTENNA_input7_A bottom_left_grid_pin_47_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xmux_left_track_5.mux_l3_in_0_ mux_left_track_5.mux_l2_in_1_/X mux_left_track_5.mux_l2_in_0_/X
+ mux_left_track_5.mux_l3_in_1_/S VGND VGND VPWR VPWR mux_left_track_5.mux_l3_in_0_/X
+ sky130_fd_sc_hd__mux2_1
XFILLER_14_31 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_14_42 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_5_214 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_79 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_68 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_30 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_18_107 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_63 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_52 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_input82_A right_bottom_grid_pin_36_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_mem_left_track_17.sky130_fd_sc_hd__dfxtp_1_2__D mux_left_track_17.mux_l2_in_1_/S
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_32_187 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmux_left_track_5.mux_l2_in_1_ mux_left_track_5.mux_l1_in_3_/X mux_left_track_5.mux_l1_in_2_/X
+ mux_left_track_5.mux_l2_in_3_/S VGND VGND VPWR VPWR mux_left_track_5.mux_l2_in_1_/X
+ sky130_fd_sc_hd__mux2_1
Xoutput113 _088_/X VGND VGND VPWR VPWR chanx_right_out[11] sky130_fd_sc_hd__buf_2
Xoutput135 _110_/X VGND VGND VPWR VPWR chany_bottom_out[13] sky130_fd_sc_hd__buf_2
Xoutput146 _102_/X VGND VGND VPWR VPWR chany_bottom_out[5] sky130_fd_sc_hd__buf_2
Xmem_right_track_24.sky130_fd_sc_hd__dfxtp_1_2_ prog_clk_0_FTB00/X mux_right_track_24.mux_l2_in_1_/S
+ VGND VGND VPWR VPWR mux_right_track_24.mux_l3_in_0_/S sky130_fd_sc_hd__dfxtp_1
Xoutput102 _058_/X VGND VGND VPWR VPWR chanx_left_out[1] sky130_fd_sc_hd__buf_2
Xoutput124 _080_/X VGND VGND VPWR VPWR chanx_right_out[3] sky130_fd_sc_hd__buf_2
XFILLER_14_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_14_143 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xinput59 chany_bottom_in[17] VGND VGND VPWR VPWR input59/X sky130_fd_sc_hd__clkbuf_1
Xinput26 chanx_left_in[5] VGND VGND VPWR VPWR _083_/A sky130_fd_sc_hd__clkbuf_2
Xinput48 chanx_right_in[7] VGND VGND VPWR VPWR _112_/A sky130_fd_sc_hd__clkbuf_1
XFILLER_14_187 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xinput15 chanx_left_in[13] VGND VGND VPWR VPWR _091_/A sky130_fd_sc_hd__dlymetal6s2s_1
Xinput37 chanx_right_in[15] VGND VGND VPWR VPWR input37/X sky130_fd_sc_hd__clkbuf_1
XANTENNA_mem_bottom_track_9.sky130_fd_sc_hd__dfxtp_1_1__CLK prog_clk_0_FTB00/X VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_20_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmem_left_track_9.sky130_fd_sc_hd__dfxtp_1_0_ prog_clk_0_FTB00/X mux_left_track_5.mux_l4_in_0_/S
+ VGND VGND VPWR VPWR mux_left_track_9.mux_l1_in_0_/S sky130_fd_sc_hd__dfxtp_1
X_100_ _100_/A VGND VGND VPWR VPWR _100_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_11_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_22_42 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_22_75 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_input45_A chanx_right_in[4] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xmux_left_track_5.mux_l1_in_2_ input79/X input57/X repeater153/X VGND VGND VPWR VPWR
+ mux_left_track_5.mux_l1_in_2_/X sky130_fd_sc_hd__mux2_1
XFILLER_6_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_6_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_8_66 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_8_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xmux_left_track_25.mux_l1_in_3_ mux_left_track_25.mux_l1_in_3_/A0 input76/X mux_left_track_25.mux_l1_in_3_/S
+ VGND VGND VPWR VPWR mux_left_track_25.mux_l1_in_3_/X sky130_fd_sc_hd__mux2_1
Xmem_left_track_33.sky130_fd_sc_hd__dfxtp_1_2_ prog_clk_0_FTB00/X mux_left_track_33.mux_l2_in_1_/S
+ VGND VGND VPWR VPWR output90/A sky130_fd_sc_hd__dfxtp_1
XFILLER_33_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_3_164 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_3_131 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_145 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_28_63 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_28_52 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_5_78 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_5_67 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_14_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_14_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_14_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_30_31 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmux_left_track_25.mux_l3_in_0_ mux_left_track_25.mux_l2_in_1_/X mux_left_track_25.mux_l2_in_0_/X
+ mux_left_track_25.mux_l3_in_0_/S VGND VGND VPWR VPWR mux_left_track_25.mux_l3_in_0_/X
+ sky130_fd_sc_hd__mux2_1
XTAP_69 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_207 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_mux_right_track_2.mux_l2_in_2__A0 _082_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_64 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_26_163 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_26_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_25_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_20 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_31 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_18_119 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_42 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_input75_A left_bottom_grid_pin_38_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mem_right_track_0.sky130_fd_sc_hd__dfxtp_1_1__CLK prog_clk_0_FTB00/X VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_32_144 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_17_185 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xoutput114 _089_/X VGND VGND VPWR VPWR chanx_right_out[12] sky130_fd_sc_hd__buf_2
Xmem_right_track_24.sky130_fd_sc_hd__dfxtp_1_1_ prog_clk_0_FTB00/X mux_right_track_24.mux_l1_in_3_/S
+ VGND VGND VPWR VPWR mux_right_track_24.mux_l2_in_1_/S sky130_fd_sc_hd__dfxtp_1
Xmux_left_track_5.mux_l2_in_0_ mux_left_track_5.mux_l1_in_1_/X mux_left_track_5.mux_l1_in_0_/X
+ mux_left_track_5.mux_l2_in_3_/S VGND VGND VPWR VPWR mux_left_track_5.mux_l2_in_0_/X
+ sky130_fd_sc_hd__mux2_1
Xoutput103 _059_/X VGND VGND VPWR VPWR chanx_left_out[2] sky130_fd_sc_hd__buf_2
Xoutput125 _081_/X VGND VGND VPWR VPWR chanx_right_out[4] sky130_fd_sc_hd__buf_2
Xoutput136 _111_/X VGND VGND VPWR VPWR chany_bottom_out[14] sky130_fd_sc_hd__buf_2
Xoutput147 _103_/X VGND VGND VPWR VPWR chany_bottom_out[6] sky130_fd_sc_hd__buf_2
Xmux_left_track_25.mux_l2_in_1_ mux_left_track_25.mux_l1_in_3_/X mux_left_track_25.mux_l1_in_2_/X
+ mux_left_track_25.mux_l2_in_1_/S VGND VGND VPWR VPWR mux_left_track_25.mux_l2_in_1_/X
+ sky130_fd_sc_hd__mux2_1
XFILLER_23_144 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_11_33 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_11_88 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xinput27 chanx_left_in[6] VGND VGND VPWR VPWR _084_/A sky130_fd_sc_hd__clkbuf_2
Xinput49 chanx_right_in[8] VGND VGND VPWR VPWR _066_/A sky130_fd_sc_hd__clkbuf_2
Xinput16 chanx_left_in[14] VGND VGND VPWR VPWR _092_/A sky130_fd_sc_hd__clkbuf_2
Xinput38 chanx_right_in[16] VGND VGND VPWR VPWR _074_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_20_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_20_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_20_158 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_input38_A chanx_right_in[16] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mem_left_track_9.sky130_fd_sc_hd__dfxtp_1_1__CLK prog_clk_0_FTB00/X VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xmux_left_track_5.mux_l1_in_1_ input69/X input62/X repeater154/A VGND VGND VPWR VPWR
+ mux_left_track_5.mux_l1_in_1_/X sky130_fd_sc_hd__mux2_1
Xmem_bottom_track_23.sky130_fd_sc_hd__dfxtp_1_1_ prog_clk_0_FTB00/X mux_bottom_track_23.mux_l1_in_1_/S
+ VGND VGND VPWR VPWR mux_bottom_track_23.mux_l2_in_0_/S sky130_fd_sc_hd__dfxtp_1
XFILLER_8_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xmux_left_track_25.mux_l1_in_2_ input72/X input60/X mux_left_track_25.mux_l1_in_3_/S
+ VGND VGND VPWR VPWR mux_left_track_25.mux_l1_in_2_/X sky130_fd_sc_hd__mux2_1
XANTENNA_mem_bottom_track_13.sky130_fd_sc_hd__dfxtp_1_0__CLK prog_clk_0_FTB00/X VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_25_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_25_206 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmux_bottom_track_5.mux_l1_in_3__155 VGND VGND VPWR VPWR mux_bottom_track_5.mux_l1_in_3_/A0
+ mux_bottom_track_5.mux_l1_in_3__155/LO sky130_fd_sc_hd__conb_1
XANTENNA_mux_left_track_1.mux_l2_in_1__S mux_left_track_1.mux_l2_in_3_/S VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_17_43 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_33_31 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_17_76 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmem_left_track_33.sky130_fd_sc_hd__dfxtp_1_1_ prog_clk_0_FTB00/X mux_left_track_33.mux_l1_in_2_/S
+ VGND VGND VPWR VPWR mux_left_track_33.mux_l2_in_1_/S sky130_fd_sc_hd__dfxtp_1
XFILLER_3_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_3_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_mux_bottom_track_11.mux_l2_in_0__A0 _087_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mem_bottom_track_27.sky130_fd_sc_hd__dfxtp_1_1__CLK prog_clk_0_FTB00/X VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_13_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_179 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_157 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_8_213 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_5_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_5_35 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmem_bottom_track_1.sky130_fd_sc_hd__dfxtp_1_2_ prog_clk_0_FTB00/X mux_bottom_track_1.mux_l2_in_1_/S
+ VGND VGND VPWR VPWR mem_bottom_track_3.delay_buf_2/X sky130_fd_sc_hd__dfxtp_1
XANTENNA_mem_right_track_32.sky130_fd_sc_hd__dfxtp_1_0__CLK prog_clk_0_FTB00/X VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_30_87 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_30_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_mux_bottom_track_5.mux_l1_in_0__A0 input2/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_29_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_29_150 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_input20_A chanx_left_in[18] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_26_131 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_25_87 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_10 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_43 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_mux_left_track_33.mux_l1_in_0__S mux_left_track_33.mux_l1_in_2_/S VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_input68_A chany_bottom_in[7] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mem_right_track_24.sky130_fd_sc_hd__dfxtp_1_1__CLK prog_clk_0_FTB00/X VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_17_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xoutput115 _090_/X VGND VGND VPWR VPWR chanx_right_out[13] sky130_fd_sc_hd__buf_2
Xoutput137 _112_/X VGND VGND VPWR VPWR chany_bottom_out[15] sky130_fd_sc_hd__buf_2
Xoutput148 _104_/X VGND VGND VPWR VPWR chany_bottom_out[7] sky130_fd_sc_hd__buf_2
XANTENNA_mux_right_track_32.mux_l2_in_0__S mux_right_track_32.mux_l2_in_1_/S VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xmem_right_track_24.sky130_fd_sc_hd__dfxtp_1_0_ prog_clk_0_FTB00/X mem_right_track_24.delay_buf_2/X
+ VGND VGND VPWR VPWR mux_right_track_24.mux_l1_in_3_/S sky130_fd_sc_hd__dfxtp_2
Xoutput104 _060_/X VGND VGND VPWR VPWR chanx_left_out[3] sky130_fd_sc_hd__buf_2
Xoutput126 _082_/X VGND VGND VPWR VPWR chanx_right_out[5] sky130_fd_sc_hd__buf_2
Xmux_left_track_25.mux_l2_in_0_ mux_left_track_25.mux_l1_in_1_/X mux_left_track_25.mux_l1_in_0_/X
+ mux_left_track_25.mux_l2_in_1_/S VGND VGND VPWR VPWR mux_left_track_25.mux_l2_in_0_/X
+ sky130_fd_sc_hd__mux2_1
XFILLER_23_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_23_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_23_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_11_78 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_14_101 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xinput28 chanx_left_in[7] VGND VGND VPWR VPWR input28/X sky130_fd_sc_hd__clkbuf_1
Xinput17 chanx_left_in[15] VGND VGND VPWR VPWR input17/X sky130_fd_sc_hd__clkbuf_1
Xinput39 chanx_right_in[17] VGND VGND VPWR VPWR _075_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_9_171 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_28_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmux_left_track_1.mux_l2_in_3__158 VGND VGND VPWR VPWR mux_left_track_1.mux_l2_in_3_/A0
+ mux_left_track_1.mux_l2_in_3__158/LO sky130_fd_sc_hd__conb_1
Xmux_bottom_track_11.mux_l3_in_0_ mux_bottom_track_11.mux_l2_in_1_/X mux_bottom_track_11.mux_l2_in_0_/X
+ mux_bottom_track_11.mux_l3_in_0_/S VGND VGND VPWR VPWR mux_bottom_track_11.mux_l3_in_0_/X
+ sky130_fd_sc_hd__mux2_1
XFILLER_7_108 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_7_119 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_11_148 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_22_22 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmem_bottom_track_23.sky130_fd_sc_hd__dfxtp_1_0_ prog_clk_0_FTB00/X mux_bottom_track_21.mux_l2_in_0_/S
+ VGND VGND VPWR VPWR mux_bottom_track_23.mux_l1_in_1_/S sky130_fd_sc_hd__dfxtp_1
XANTENNA_mem_right_track_16.sky130_fd_sc_hd__dfxtp_1_2__CLK prog_clk_0_FTB00/X VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xmux_left_track_5.mux_l1_in_0_ _072_/A _063_/A repeater153/X VGND VGND VPWR VPWR mux_left_track_5.mux_l1_in_0_/X
+ sky130_fd_sc_hd__mux2_1
Xmem_right_track_16.delay_buf_2 mux_right_track_8.mux_l4_in_0_/S VGND VGND VPWR VPWR
+ mux_right_track_8.mux_l4_in_0_/S sky130_fd_sc_hd__buf_6
X_089_ _089_/A VGND VGND VPWR VPWR _089_/X sky130_fd_sc_hd__clkbuf_1
Xmux_left_track_25.mux_l1_in_1_ input53/X input65/X mux_left_track_25.mux_l1_in_3_/S
+ VGND VGND VPWR VPWR mux_left_track_25.mux_l1_in_1_/X sky130_fd_sc_hd__mux2_1
XANTENNA_mem_bottom_track_3.sky130_fd_sc_hd__dfxtp_1_2__CLK prog_clk_0_FTB00/X VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xmux_bottom_track_3.mux_l1_in_3__182 VGND VGND VPWR VPWR mux_bottom_track_3.mux_l1_in_3_/A0
+ mux_bottom_track_3.mux_l1_in_3__182/LO sky130_fd_sc_hd__conb_1
XANTENNA__060__A _060_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_17_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_17_88 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_33_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_33_43 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmem_left_track_33.sky130_fd_sc_hd__dfxtp_1_0_ prog_clk_0_FTB00/X mux_left_track_25.mux_l3_in_0_/S
+ VGND VGND VPWR VPWR mux_left_track_33.mux_l1_in_2_/S sky130_fd_sc_hd__dfxtp_1
XANTENNA_input50_A chanx_right_in[9] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xmux_right_track_32.mux_l3_in_0_ mux_right_track_32.mux_l2_in_1_/X mux_right_track_32.mux_l2_in_0_/X
+ mem_bottom_track_1.delay_buf_2/X VGND VGND VPWR VPWR mux_right_track_32.mux_l3_in_0_/X
+ sky130_fd_sc_hd__mux2_1
XFILLER_30_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmux_bottom_track_11.mux_l2_in_1_ mux_bottom_track_11.mux_l2_in_1_/A0 input21/X mux_bottom_track_11.mux_l2_in_1_/S
+ VGND VGND VPWR VPWR mux_bottom_track_11.mux_l2_in_1_/X sky130_fd_sc_hd__mux2_1
XFILLER_21_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_28_87 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_12_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_5_25 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmem_bottom_track_1.sky130_fd_sc_hd__dfxtp_1_1_ prog_clk_0_FTB00/X mux_bottom_track_1.mux_l1_in_3_/S
+ VGND VGND VPWR VPWR mux_bottom_track_1.mux_l2_in_1_/S sky130_fd_sc_hd__dfxtp_1
XFILLER_30_22 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmux_right_track_32.mux_l2_in_1_ mux_right_track_32.mux_l2_in_1_/A0 _088_/A mux_right_track_32.mux_l2_in_1_/S
+ VGND VGND VPWR VPWR mux_right_track_32.mux_l2_in_1_/X sky130_fd_sc_hd__mux2_1
XFILLER_30_66 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_mux_bottom_track_5.mux_l1_in_0__A1 _063_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_29_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_input13_A chanx_left_in[11] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xmux_bottom_track_9.mux_l2_in_1__157 VGND VGND VPWR VPWR mux_bottom_track_9.mux_l2_in_1_/A0
+ mux_bottom_track_9.mux_l2_in_1__157/LO sky130_fd_sc_hd__conb_1
XFILLER_26_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_input5_A bottom_left_grid_pin_45_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_66 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_26_187 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_26_176 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_25_99 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_22 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_33 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_25_22 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_25_33 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_25_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_2_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_2_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_mux_bottom_track_3.mux_l1_in_2__A1 input9/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_17_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xoutput116 _091_/X VGND VGND VPWR VPWR chanx_right_out[14] sky130_fd_sc_hd__buf_2
Xoutput127 _083_/X VGND VGND VPWR VPWR chanx_right_out[6] sky130_fd_sc_hd__buf_2
Xoutput138 _113_/X VGND VGND VPWR VPWR chany_bottom_out[16] sky130_fd_sc_hd__buf_2
Xoutput149 _105_/X VGND VGND VPWR VPWR chany_bottom_out[8] sky130_fd_sc_hd__buf_2
Xoutput105 _061_/X VGND VGND VPWR VPWR chanx_left_out[4] sky130_fd_sc_hd__buf_2
Xmem_bottom_track_7.sky130_fd_sc_hd__dfxtp_1_2_ prog_clk_0_FTB00/X mux_bottom_track_7.mux_l2_in_1_/S
+ VGND VGND VPWR VPWR mux_bottom_track_7.mux_l3_in_0_/S sky130_fd_sc_hd__dfxtp_1
XFILLER_11_13 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_11_24 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__063__A _063_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_190 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_input80_A right_bottom_grid_pin_34_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xinput18 chanx_left_in[16] VGND VGND VPWR VPWR _094_/A sky130_fd_sc_hd__dlymetal6s2s_1
Xinput29 chanx_left_in[8] VGND VGND VPWR VPWR _086_/A sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_28_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_20_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_20_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_11_116 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_11_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_mux_right_track_4.mux_l1_in_4__A0 input64/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_22_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_19_205 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_10_160 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmux_left_track_25.mux_l1_in_0_ _076_/A _067_/A mux_left_track_25.mux_l1_in_3_/S VGND
+ VGND VPWR VPWR mux_left_track_25.mux_l1_in_0_/X sky130_fd_sc_hd__mux2_1
X_088_ _088_/A VGND VGND VPWR VPWR _088_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_6_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_19_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_mem_left_track_3.sky130_fd_sc_hd__dfxtp_1_2__CLK prog_clk_0_FTB00/X VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_3_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_input43_A chanx_right_in[2] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xmux_bottom_track_7.mux_l1_in_3_ mux_bottom_track_7.mux_l1_in_3_/A0 input13/X mux_bottom_track_7.mux_l1_in_3_/S
+ VGND VGND VPWR VPWR mux_bottom_track_7.mux_l1_in_3_/X sky130_fd_sc_hd__mux2_1
Xmux_bottom_track_11.mux_l2_in_0_ _087_/A mux_bottom_track_11.mux_l1_in_0_/X mux_bottom_track_11.mux_l2_in_1_/S
+ VGND VGND VPWR VPWR mux_bottom_track_11.mux_l2_in_0_/X sky130_fd_sc_hd__mux2_1
XANTENNA__071__A _071_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xmem_bottom_track_1.sky130_fd_sc_hd__dfxtp_1_0_ prog_clk_0_FTB00/X mem_bottom_track_1.delay_buf_2/X
+ VGND VGND VPWR VPWR mux_bottom_track_1.mux_l1_in_3_/S sky130_fd_sc_hd__dfxtp_2
Xmux_bottom_track_25.sky130_fd_sc_hd__buf_4_0_ mux_bottom_track_25.mux_l3_in_0_/X
+ VGND VGND VPWR VPWR _109_/A sky130_fd_sc_hd__clkbuf_1
XANTENNA_mux_right_track_0.mux_l2_in_1__S mux_right_track_0.mux_l2_in_3_/S VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__066__A _066_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_30_12 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmux_right_track_32.mux_l2_in_0_ mux_right_track_32.mux_l1_in_1_/X mux_right_track_32.mux_l1_in_0_/X
+ mux_right_track_32.mux_l2_in_1_/S VGND VGND VPWR VPWR mux_right_track_32.mux_l2_in_0_/X
+ sky130_fd_sc_hd__mux2_1
XPHY_12 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_67 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_26_199 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmux_bottom_track_7.mux_l3_in_0_ mux_bottom_track_7.mux_l2_in_1_/X mux_bottom_track_7.mux_l2_in_0_/X
+ mux_bottom_track_7.mux_l3_in_0_/S VGND VGND VPWR VPWR mux_bottom_track_7.mux_l3_in_0_/X
+ sky130_fd_sc_hd__mux2_1
XPHY_23 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_34 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_45 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xmux_bottom_track_19.sky130_fd_sc_hd__buf_4_0_ mux_bottom_track_19.mux_l2_in_0_/X
+ VGND VGND VPWR VPWR _106_/A sky130_fd_sc_hd__clkbuf_1
XFILLER_2_38 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_1_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_17_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_17_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xoutput117 _092_/X VGND VGND VPWR VPWR chanx_right_out[15] sky130_fd_sc_hd__buf_2
Xoutput128 _084_/X VGND VGND VPWR VPWR chanx_right_out[7] sky130_fd_sc_hd__buf_2
Xoutput139 _114_/X VGND VGND VPWR VPWR chany_bottom_out[17] sky130_fd_sc_hd__buf_2
Xoutput106 _062_/X VGND VGND VPWR VPWR chanx_left_out[5] sky130_fd_sc_hd__buf_2
Xmem_bottom_track_7.sky130_fd_sc_hd__dfxtp_1_1_ prog_clk_0_FTB00/X mux_bottom_track_7.mux_l1_in_3_/S
+ VGND VGND VPWR VPWR mux_bottom_track_7.mux_l2_in_1_/S sky130_fd_sc_hd__dfxtp_1
Xmux_right_track_32.mux_l1_in_1_ input55/X input67/X mux_right_track_32.mux_l1_in_1_/S
+ VGND VGND VPWR VPWR mux_right_track_32.mux_l1_in_1_/X sky130_fd_sc_hd__mux2_1
XFILLER_31_191 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_191 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_180 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_114 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_14_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_14_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_mem_right_track_4.sky130_fd_sc_hd__dfxtp_1_1__CLK prog_clk_0_FTB00/X VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xinput19 chanx_left_in[17] VGND VGND VPWR VPWR _095_/A sky130_fd_sc_hd__dlymetal6s2s_1
XANTENNA_input73_A left_bottom_grid_pin_36_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_20_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmux_bottom_track_7.mux_l2_in_1_ mux_bottom_track_7.mux_l1_in_3_/X mux_bottom_track_7.mux_l1_in_2_/X
+ mux_bottom_track_7.mux_l2_in_1_/S VGND VGND VPWR VPWR mux_bottom_track_7.mux_l2_in_1_/X
+ sky130_fd_sc_hd__mux2_1
XANTENNA__074__A _074_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_11_106 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_22_13 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_22_79 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_8_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_087_ _087_/A VGND VGND VPWR VPWR _087_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_6_143 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_8_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_10_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_mem_left_track_33.sky130_fd_sc_hd__dfxtp_1_0__CLK prog_clk_0_FTB00/X VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_17_13 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_33_23 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_17_24 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_mux_bottom_track_7.mux_l1_in_1__A0 input7/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_33_67 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_mux_bottom_track_23.mux_l1_in_0__A0 input9/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_3_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_input36_A chanx_right_in[14] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xmux_right_track_24.sky130_fd_sc_hd__buf_4_0_ mux_right_track_24.mux_l3_in_0_/X VGND
+ VGND VPWR VPWR _089_/A sky130_fd_sc_hd__clkbuf_1
XANTENNA_mem_bottom_track_17.sky130_fd_sc_hd__dfxtp_1_0__CLK prog_clk_0_FTB00/X VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xmux_bottom_track_7.mux_l1_in_2_ _084_/A input9/X mux_bottom_track_7.mux_l1_in_3_/S
+ VGND VGND VPWR VPWR mux_bottom_track_7.mux_l1_in_2_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_28_67 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_28_23 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_12_201 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_12_212 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_mem_left_track_25.sky130_fd_sc_hd__dfxtp_1_1__CLK prog_clk_0_FTB00/X VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mux_bottom_track_15.mux_l1_in_0__A1 _070_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xmux_left_track_1.mux_l2_in_3_ mux_left_track_1.mux_l2_in_3_/A0 input78/X mux_left_track_1.mux_l2_in_3_/S
+ VGND VGND VPWR VPWR mux_left_track_1.mux_l2_in_3_/X sky130_fd_sc_hd__mux2_1
XFILLER_30_46 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_30_35 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__082__A _082_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_29_120 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmux_bottom_track_11.mux_l1_in_0_ input3/X _067_/A mux_bottom_track_11.mux_l1_in_0_/S
+ VGND VGND VPWR VPWR mux_bottom_track_11.mux_l1_in_0_/X sky130_fd_sc_hd__mux2_1
XANTENNA_mux_left_track_3.mux_l1_in_0__A0 _071_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xmux_bottom_track_23.mux_l2_in_0_ mux_bottom_track_23.mux_l1_in_1_/X mux_bottom_track_23.mux_l1_in_0_/X
+ mux_bottom_track_23.mux_l2_in_0_/S VGND VGND VPWR VPWR mux_bottom_track_23.mux_l2_in_0_/X
+ sky130_fd_sc_hd__mux2_1
XFILLER_26_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_13 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_24 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_35 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xmem_right_track_16.sky130_fd_sc_hd__dfxtp_1_2_ prog_clk_0_FTB00/X mux_right_track_16.mux_l2_in_1_/S
+ VGND VGND VPWR VPWR mem_right_track_24.delay_buf_2/X sky130_fd_sc_hd__dfxtp_1
XPHY_46 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_25_13 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_25_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_9_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_mux_left_track_33.mux_l2_in_1__S mux_left_track_33.mux_l2_in_1_/S VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mem_left_track_17.sky130_fd_sc_hd__dfxtp_1_2__CLK prog_clk_0_FTB00/X VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_32_115 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_32_104 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_mem_bottom_track_1.sky130_fd_sc_hd__dfxtp_1_0__CLK prog_clk_0_FTB00/X VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_17_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xoutput107 _063_/X VGND VGND VPWR VPWR chanx_left_out[6] sky130_fd_sc_hd__buf_2
Xoutput118 _093_/X VGND VGND VPWR VPWR chanx_right_out[16] sky130_fd_sc_hd__buf_2
Xoutput129 _085_/X VGND VGND VPWR VPWR chanx_right_out[8] sky130_fd_sc_hd__buf_2
Xmem_bottom_track_7.sky130_fd_sc_hd__dfxtp_1_0_ prog_clk_0_FTB00/X mem_bottom_track_7.delay_buf_2/X
+ VGND VGND VPWR VPWR mux_bottom_track_7.mux_l1_in_3_/S sky130_fd_sc_hd__dfxtp_2
Xmux_right_track_32.mux_l1_in_0_ input86/X input82/X mux_right_track_32.mux_l1_in_1_/S
+ VGND VGND VPWR VPWR mux_right_track_32.mux_l1_in_0_/X sky130_fd_sc_hd__mux2_1
XFILLER_23_115 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_23_126 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_11_59 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_192 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_181 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_170 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xmux_left_track_1.mux_l4_in_0_ mux_left_track_1.mux_l3_in_1_/X mux_left_track_1.mux_l3_in_0_/X
+ mux_left_track_1.mux_l4_in_0_/S VGND VGND VPWR VPWR mux_left_track_1.mux_l4_in_0_/X
+ sky130_fd_sc_hd__mux2_1
XANTENNA_input66_A chany_bottom_in[5] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xmux_bottom_track_23.mux_l1_in_1_ mux_bottom_track_23.mux_l1_in_1_/A0 _095_/A mux_bottom_track_23.mux_l1_in_1_/S
+ VGND VGND VPWR VPWR mux_bottom_track_23.mux_l1_in_1_/X sky130_fd_sc_hd__mux2_1
XFILLER_9_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_20_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_9_163 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_28_207 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_3_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmux_bottom_track_7.mux_l2_in_0_ mux_bottom_track_7.mux_l1_in_1_/X mux_bottom_track_7.mux_l1_in_0_/X
+ mux_bottom_track_7.mux_l2_in_1_/S VGND VGND VPWR VPWR mux_bottom_track_7.mux_l2_in_0_/X
+ sky130_fd_sc_hd__mux2_1
Xmux_left_track_9.mux_l2_in_3__164 VGND VGND VPWR VPWR mux_left_track_9.mux_l2_in_3_/A0
+ mux_left_track_9.mux_l2_in_3__164/LO sky130_fd_sc_hd__conb_1
XANTENNA__090__A _090_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_8_38 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_086_ _086_/A VGND VGND VPWR VPWR _086_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_6_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_6_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_33_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmem_left_track_25.sky130_fd_sc_hd__dfxtp_1_2_ prog_clk_0_FTB00/X mux_left_track_25.mux_l2_in_1_/S
+ VGND VGND VPWR VPWR mux_left_track_25.mux_l3_in_0_/S sky130_fd_sc_hd__dfxtp_1
XFILLER_33_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmux_left_track_3.sky130_fd_sc_hd__buf_4_0_ mux_left_track_3.mux_l4_in_0_/X VGND VGND
+ VPWR VPWR _058_/A sky130_fd_sc_hd__clkbuf_1
XFILLER_17_47 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_33_35 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_33_13 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmux_left_track_1.mux_l3_in_1_ mux_left_track_1.mux_l2_in_3_/X mux_left_track_1.mux_l2_in_2_/X
+ mux_left_track_1.mux_l3_in_1_/S VGND VGND VPWR VPWR mux_left_track_1.mux_l3_in_1_/X
+ sky130_fd_sc_hd__mux2_1
XFILLER_24_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_33_79 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_mux_bottom_track_23.mux_l1_in_0__A1 _075_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_15_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_input29_A chanx_left_in[8] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_30_213 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_mem_bottom_track_7.sky130_fd_sc_hd__dfxtp_1_2__CLK prog_clk_0_FTB00/X VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xmux_bottom_track_7.mux_l1_in_1_ input7/X input5/X mux_bottom_track_7.mux_l1_in_3_/S
+ VGND VGND VPWR VPWR mux_bottom_track_7.mux_l1_in_1_/X sky130_fd_sc_hd__mux2_1
X_069_ _069_/A VGND VGND VPWR VPWR _069_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_28_13 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_28_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xmux_left_track_1.mux_l2_in_2_ input76/X input74/X mux_left_track_1.mux_l2_in_3_/S
+ VGND VGND VPWR VPWR mux_left_track_1.mux_l2_in_2_/X sky130_fd_sc_hd__mux2_1
XFILLER_14_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_14_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_30_58 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_6_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_mux_left_track_3.mux_l1_in_0__A1 _062_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_58 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xmem_left_track_17.delay_buf_2 mux_left_track_9.mux_l4_in_0_/S VGND VGND VPWR VPWR
+ mux_left_track_9.mux_l4_in_0_/S sky130_fd_sc_hd__buf_6
XFILLER_26_168 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_26_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_26_102 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_14 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_25 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xmem_right_track_16.sky130_fd_sc_hd__dfxtp_1_1_ prog_clk_0_FTB00/X mux_right_track_16.mux_l1_in_3_/S
+ VGND VGND VPWR VPWR mux_right_track_16.mux_l2_in_1_/S sky130_fd_sc_hd__dfxtp_1
XPHY_36 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_47 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_input11_A chanx_left_in[0] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_32_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_32_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_32_127 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_mux_right_track_8.mux_l2_in_2__A0 _084_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_25_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xoutput119 _094_/X VGND VGND VPWR VPWR chanx_right_out[17] sky130_fd_sc_hd__buf_2
XFILLER_31_90 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xoutput108 _064_/X VGND VGND VPWR VPWR chanx_left_out[7] sky130_fd_sc_hd__buf_2
Xoutput90 output90/A VGND VGND VPWR VPWR ccff_tail sky130_fd_sc_hd__buf_2
Xmux_right_track_2.mux_l2_in_3_ mux_right_track_2.mux_l2_in_3_/A0 _091_/A mux_right_track_2.mux_l2_in_3_/S
+ VGND VGND VPWR VPWR mux_right_track_2.mux_l2_in_3_/X sky130_fd_sc_hd__mux2_1
XFILLER_11_38 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_11_49 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_193 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__088__A _088_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_182 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_input3_A bottom_left_grid_pin_43_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_171 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_160 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_mem_left_track_1.sky130_fd_sc_hd__dfxtp_1_0__CLK prog_clk_0_FTB00/X VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_14_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_input59_A chany_bottom_in[17] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xmux_bottom_track_23.mux_l1_in_0_ input9/X _075_/A mux_bottom_track_23.mux_l1_in_1_/S
+ VGND VGND VPWR VPWR mux_bottom_track_23.mux_l1_in_0_/X sky130_fd_sc_hd__mux2_1
XFILLER_9_175 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xmem_bottom_track_15.sky130_fd_sc_hd__dfxtp_1_1_ prog_clk_0_FTB00/X mux_bottom_track_15.mux_l1_in_1_/S
+ VGND VGND VPWR VPWR mux_bottom_track_15.mux_l2_in_0_/S sky130_fd_sc_hd__dfxtp_1
XFILLER_13_171 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_13_182 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_3_72 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_22_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_22_48 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_10_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_085_ _085_/A VGND VGND VPWR VPWR _085_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_6_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmem_left_track_25.sky130_fd_sc_hd__dfxtp_1_1_ prog_clk_0_FTB00/X mux_left_track_25.mux_l1_in_3_/S
+ VGND VGND VPWR VPWR mux_left_track_25.mux_l2_in_1_/S sky130_fd_sc_hd__dfxtp_1
XFILLER_26_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_mem_right_track_32.sky130_fd_sc_hd__dfxtp_1_2__D mux_right_track_32.mux_l2_in_1_/S
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_17_59 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_33_47 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xmux_left_track_1.mux_l3_in_0_ mux_left_track_1.mux_l2_in_1_/X mux_left_track_1.mux_l2_in_0_/X
+ mux_left_track_1.mux_l3_in_1_/S VGND VGND VPWR VPWR mux_left_track_1.mux_l3_in_0_/X
+ sky130_fd_sc_hd__mux2_1
XFILLER_3_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_mem_right_track_0.sky130_fd_sc_hd__dfxtp_1_0__D input10/X VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XFILLER_30_203 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmux_right_track_2.mux_l4_in_0_ mux_right_track_2.mux_l3_in_1_/X mux_right_track_2.mux_l3_in_0_/X
+ mux_right_track_2.mux_l4_in_0_/S VGND VGND VPWR VPWR mux_right_track_2.mux_l4_in_0_/X
+ sky130_fd_sc_hd__mux2_1
Xmux_bottom_track_7.mux_l1_in_0_ input3/X _064_/A mux_bottom_track_7.mux_l1_in_3_/S
+ VGND VGND VPWR VPWR mux_bottom_track_7.mux_l1_in_0_/X sky130_fd_sc_hd__mux2_1
Xmux_bottom_track_7.sky130_fd_sc_hd__buf_4_0_ mux_bottom_track_7.mux_l3_in_0_/X VGND
+ VGND VPWR VPWR _100_/A sky130_fd_sc_hd__clkbuf_1
X_068_ _068_/A VGND VGND VPWR VPWR _068_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_0_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_9_71 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__096__A _096_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_input41_A chanx_right_in[19] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mem_bottom_track_11.sky130_fd_sc_hd__dfxtp_1_1__CLK prog_clk_0_FTB00/X VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xmux_left_track_1.mux_l2_in_1_ input72/X input79/X mux_left_track_1.mux_l2_in_3_/S
+ VGND VGND VPWR VPWR mux_left_track_1.mux_l2_in_1_/X sky130_fd_sc_hd__mux2_1
XANTENNA_mux_left_track_1.mux_l4_in_0__S mux_left_track_1.mux_l4_in_0_/S VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_30_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_29_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_29_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xmux_right_track_2.mux_l3_in_1_ mux_right_track_2.mux_l2_in_3_/X mux_right_track_2.mux_l2_in_2_/X
+ mux_right_track_2.mux_l3_in_1_/S VGND VGND VPWR VPWR mux_right_track_2.mux_l3_in_1_/X
+ sky130_fd_sc_hd__mux2_1
XFILLER_4_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_mem_bottom_track_25.sky130_fd_sc_hd__dfxtp_1_2__CLK prog_clk_0_FTB00/X VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_6_72 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_59 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_26_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_37 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xmem_right_track_16.sky130_fd_sc_hd__dfxtp_1_0_ prog_clk_0_FTB00/X mux_right_track_8.mux_l4_in_0_/S
+ VGND VGND VPWR VPWR mux_right_track_16.mux_l1_in_3_/S sky130_fd_sc_hd__dfxtp_2
XPHY_48 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_25_37 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_25_48 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_mem_left_track_1.sky130_fd_sc_hd__dfxtp_1_3__D mux_left_track_1.mux_l3_in_1_/S
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_1_202 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_17_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_mux_right_track_8.mux_l2_in_2__A1 input58/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_25_180 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_15_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xoutput109 _065_/X VGND VGND VPWR VPWR chanx_left_out[8] sky130_fd_sc_hd__buf_2
Xoutput91 _057_/X VGND VGND VPWR VPWR chanx_left_out[0] sky130_fd_sc_hd__buf_2
Xmux_right_track_2.mux_l2_in_2_ _082_/A input60/X mux_right_track_2.mux_l2_in_3_/S
+ VGND VGND VPWR VPWR mux_right_track_2.mux_l2_in_2_/X sky130_fd_sc_hd__mux2_1
XTAP_150 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_183 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_172 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_161 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_mux_right_track_16.mux_l1_in_2__A0 _086_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_22_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_mux_bottom_track_1.mux_l1_in_1__S mux_bottom_track_1.mux_l1_in_3_/S VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xmem_bottom_track_15.sky130_fd_sc_hd__dfxtp_1_0_ prog_clk_0_FTB00/X mux_bottom_track_13.mux_l2_in_0_/S
+ VGND VGND VPWR VPWR mux_bottom_track_15.mux_l1_in_1_/S sky130_fd_sc_hd__dfxtp_1
XFILLER_20_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_3_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_22_38 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_9 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_mem_right_track_8.sky130_fd_sc_hd__dfxtp_1_1__CLK prog_clk_0_FTB00/X VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_19_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_6_102 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_6_124 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_10_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_10_164 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_084_ _084_/A VGND VGND VPWR VPWR _084_/X sky130_fd_sc_hd__clkbuf_1
XANTENNA_mux_bottom_track_17.mux_l1_in_1__A1 _091_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_input71_A left_bottom_grid_pin_34_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_12_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmem_left_track_25.sky130_fd_sc_hd__dfxtp_1_0_ prog_clk_0_FTB00/X mem_left_track_25.delay_buf_2/X
+ VGND VGND VPWR VPWR mux_left_track_25.mux_l1_in_3_/S sky130_fd_sc_hd__dfxtp_2
XANTENNA_mux_bottom_track_25.mux_l2_in_0__A0 input2/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_17_38 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_3_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_15_212 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_23_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_067_ _067_/A VGND VGND VPWR VPWR _067_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_2_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_mux_right_track_16.mux_l1_in_1__S mux_right_track_16.mux_l1_in_3_/S VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_63 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_9_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmux_bottom_track_19.mux_l1_in_1__177 VGND VGND VPWR VPWR mux_bottom_track_19.mux_l1_in_1_/A0
+ mux_bottom_track_19.mux_l1_in_1__177/LO sky130_fd_sc_hd__conb_1
XANTENNA_input34_A chanx_right_in[12] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_18_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xmux_left_track_1.mux_l2_in_0_ mux_left_track_1.mux_l1_in_1_/X mux_left_track_1.mux_l1_in_0_/X
+ mux_left_track_1.mux_l2_in_3_/S VGND VGND VPWR VPWR mux_left_track_1.mux_l2_in_0_/X
+ sky130_fd_sc_hd__mux2_1
XFILLER_29_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_29_101 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmux_right_track_2.mux_l3_in_0_ mux_right_track_2.mux_l2_in_1_/X mux_right_track_2.mux_l2_in_0_/X
+ mux_right_track_2.mux_l3_in_1_/S VGND VGND VPWR VPWR mux_right_track_2.mux_l3_in_0_/X
+ sky130_fd_sc_hd__mux2_1
XFILLER_20_60 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_29_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_mux_right_track_24.mux_l1_in_2__A0 _087_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_26_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_16 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_38 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_49 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_17_115 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_17_148 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmux_left_track_1.mux_l1_in_1_ input55/X input67/X mux_left_track_1.mux_l1_in_1_/S
+ VGND VGND VPWR VPWR mux_left_track_1.mux_l1_in_1_/X sky130_fd_sc_hd__mux2_1
XANTENNA_mem_right_track_16.sky130_fd_sc_hd__dfxtp_1_1__D mux_right_track_16.mux_l1_in_3_/S
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xoutput92 _067_/X VGND VGND VPWR VPWR chanx_left_out[10] sky130_fd_sc_hd__buf_2
XFILLER_16_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_31_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmux_right_track_2.mux_l2_in_1_ input53/X input65/X mux_right_track_2.mux_l2_in_3_/S
+ VGND VGND VPWR VPWR mux_right_track_2.mux_l2_in_1_/X sky130_fd_sc_hd__mux2_1
XFILLER_11_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_184 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_173 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_162 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_140 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_151 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_mux_right_track_16.mux_l1_in_2__A1 input57/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mem_bottom_track_5.sky130_fd_sc_hd__dfxtp_1_0__CLK prog_clk_0_FTB00/X VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_9_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_27_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmem_left_track_5.sky130_fd_sc_hd__dfxtp_1_3_ prog_clk_0_FTB00/X mux_left_track_5.mux_l3_in_1_/S
+ VGND VGND VPWR VPWR mux_left_track_5.mux_l4_in_0_/S sky130_fd_sc_hd__dfxtp_1
X_083_ _083_/A VGND VGND VPWR VPWR _083_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_10_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_10_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_10_132 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_10_187 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_12_50 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_12_72 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_input64_A chany_bottom_in[3] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_18_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmux_bottom_track_23.mux_l1_in_1__179 VGND VGND VPWR VPWR mux_bottom_track_23.mux_l1_in_1_/A0
+ mux_bottom_track_23.mux_l1_in_1__179/LO sky130_fd_sc_hd__conb_1
XANTENNA_mux_right_track_2.mux_l2_in_0__S mux_right_track_2.mux_l2_in_3_/S VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_5_191 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_5_180 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_17_28 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_33_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_3_106 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_066_ _066_/A VGND VGND VPWR VPWR _066_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_31_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_75 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_9_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_21_216 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_28_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_12_216 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_input27_A chanx_left_in[6] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_30_17 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_mem_left_track_1.sky130_fd_sc_hd__dfxtp_1_3__CLK prog_clk_0_FTB00/X VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_29_124 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_29_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xmux_left_track_33.mux_l3_in_0_ mux_left_track_33.mux_l2_in_1_/X mux_left_track_33.mux_l2_in_0_/X
+ output90/A VGND VGND VPWR VPWR mux_left_track_33.mux_l3_in_0_/X sky130_fd_sc_hd__mux2_1
XFILLER_20_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_6_63 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_6_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_mux_right_track_24.mux_l1_in_2__A1 input56/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_26_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_26_127 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_17 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_28 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_25_171 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xmux_left_track_1.mux_l1_in_0_ _070_/A _060_/A mux_left_track_1.mux_l1_in_1_/S VGND
+ VGND VPWR VPWR mux_left_track_1.mux_l1_in_0_/X sky130_fd_sc_hd__mux2_1
XFILLER_31_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xoutput93 _068_/X VGND VGND VPWR VPWR chanx_left_out[11] sky130_fd_sc_hd__buf_2
XANTENNA_mux_right_track_2.mux_l2_in_3__S mux_right_track_2.mux_l2_in_3_/S VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_31_163 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_16_160 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_23_119 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xmux_right_track_2.mux_l2_in_0_ mux_right_track_2.mux_l1_in_1_/X mux_right_track_2.mux_l1_in_0_/X
+ mux_right_track_2.mux_l2_in_3_/S VGND VGND VPWR VPWR mux_right_track_2.mux_l2_in_0_/X
+ sky130_fd_sc_hd__mux2_1
XTAP_185 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_174 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_163 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_130 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_141 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_152 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xmux_left_track_33.mux_l2_in_1_ mux_left_track_33.mux_l2_in_1_/A0 mux_left_track_33.mux_l1_in_2_/X
+ mux_left_track_33.mux_l2_in_1_/S VGND VGND VPWR VPWR mux_left_track_33.mux_l2_in_1_/X
+ sky130_fd_sc_hd__mux2_1
XFILLER_14_119 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmem_right_track_2.sky130_fd_sc_hd__dfxtp_1_3_ prog_clk_0_FTB00/X mux_right_track_2.mux_l3_in_1_/S
+ VGND VGND VPWR VPWR mux_right_track_2.mux_l4_in_0_/S sky130_fd_sc_hd__dfxtp_1
XANTENNA_mux_left_track_9.mux_l2_in_2__S mux_left_track_9.mux_l2_in_3_/S VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_26_60 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_9_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_9_145 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_9_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_mem_left_track_5.sky130_fd_sc_hd__dfxtp_1_0__CLK prog_clk_0_FTB00/X VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_22_18 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_input1_A SC_IN_BOT VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xmem_left_track_5.sky130_fd_sc_hd__dfxtp_1_2_ prog_clk_0_FTB00/X mux_left_track_5.mux_l2_in_3_/S
+ VGND VGND VPWR VPWR mux_left_track_5.mux_l3_in_1_/S sky130_fd_sc_hd__dfxtp_1
Xmux_right_track_4.mux_l2_in_3__170 VGND VGND VPWR VPWR mux_right_track_4.mux_l2_in_3_/A0
+ mux_right_track_4.mux_l2_in_3__170/LO sky130_fd_sc_hd__conb_1
XFILLER_12_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_082_ _082_/A VGND VGND VPWR VPWR _082_/X sky130_fd_sc_hd__clkbuf_1
XANTENNA_input57_A chany_bottom_in[15] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_33_203 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmux_right_track_2.mux_l1_in_1_ input86/X input84/X mux_right_track_2.mux_l1_in_1_/S
+ VGND VGND VPWR VPWR mux_right_track_2.mux_l1_in_1_/X sky130_fd_sc_hd__mux2_1
XFILLER_18_200 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_18_211 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmux_left_track_33.mux_l1_in_2_ input77/X input73/X mux_left_track_33.mux_l1_in_2_/S
+ VGND VGND VPWR VPWR mux_left_track_33.mux_l1_in_2_/X sky130_fd_sc_hd__mux2_1
XFILLER_33_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_24_203 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_mem_right_track_2.sky130_fd_sc_hd__dfxtp_1_2__CLK prog_clk_0_FTB00/X VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_065_ _065_/A VGND VGND VPWR VPWR _065_/X sky130_fd_sc_hd__clkbuf_1
XANTENNA_mem_bottom_track_23.sky130_fd_sc_hd__dfxtp_1_0__CLK prog_clk_0_FTB00/X VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_24_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_7_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_mux_right_track_24.mux_l1_in_2__S mux_right_track_24.mux_l1_in_3_/S VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mem_bottom_track_15.sky130_fd_sc_hd__dfxtp_1_1__CLK prog_clk_0_FTB00/X VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_6_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_mem_left_track_33.sky130_fd_sc_hd__dfxtp_1_1__D mux_left_track_33.mux_l1_in_2_/S
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_26_106 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_18 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_25_18 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_1_216 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_mux_right_track_32.mux_l2_in_1__A1 _088_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_15_73 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_15_84 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_31_94 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_mux_left_track_9.mux_l1_in_0__A0 _074_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_input87_A right_bottom_grid_pin_41_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xoutput94 _069_/X VGND VGND VPWR VPWR chanx_left_out[12] sky130_fd_sc_hd__buf_2
XFILLER_16_150 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_23_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_16_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_186 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_175 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_164 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_120 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_131 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_142 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_153 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xmux_left_track_33.mux_l2_in_0_ mux_left_track_33.mux_l1_in_1_/X mux_left_track_33.mux_l1_in_0_/X
+ mux_left_track_33.mux_l2_in_1_/S VGND VGND VPWR VPWR mux_left_track_33.mux_l2_in_0_/X
+ sky130_fd_sc_hd__mux2_1
XFILLER_22_120 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_22_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmem_right_track_2.sky130_fd_sc_hd__dfxtp_1_2_ prog_clk_0_FTB00/X mux_right_track_2.mux_l2_in_3_/S
+ VGND VGND VPWR VPWR mux_right_track_2.mux_l3_in_1_/S sky130_fd_sc_hd__dfxtp_1
XFILLER_26_94 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_26_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_13_186 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xmux_bottom_track_21.sky130_fd_sc_hd__buf_4_0_ mux_bottom_track_21.mux_l2_in_0_/X
+ VGND VGND VPWR VPWR _107_/A sky130_fd_sc_hd__clkbuf_1
XFILLER_9_179 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_3_87 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_3_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmux_bottom_track_3.mux_l1_in_3_ mux_bottom_track_3.mux_l1_in_3_/A0 _082_/A mux_bottom_track_3.mux_l1_in_3_/S
+ VGND VGND VPWR VPWR mux_bottom_track_3.mux_l1_in_3_/X sky130_fd_sc_hd__mux2_1
Xmem_left_track_17.sky130_fd_sc_hd__dfxtp_1_2_ prog_clk_0_FTB00/X mux_left_track_17.mux_l2_in_1_/S
+ VGND VGND VPWR VPWR mem_left_track_25.delay_buf_2/X sky130_fd_sc_hd__dfxtp_1
XANTENNA_mux_right_track_32.mux_l3_in_0__A1 mux_right_track_32.mux_l2_in_0_/X VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xmux_right_track_2.sky130_fd_sc_hd__buf_4_0_ mux_right_track_2.mux_l4_in_0_/X VGND
+ VGND VPWR VPWR _078_/A sky130_fd_sc_hd__clkbuf_1
Xmem_left_track_5.sky130_fd_sc_hd__dfxtp_1_1_ prog_clk_0_FTB00/X repeater154/A VGND
+ VGND VPWR VPWR mux_left_track_5.mux_l2_in_3_/S sky130_fd_sc_hd__dfxtp_2
X_081_ _081_/A VGND VGND VPWR VPWR _081_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_6_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_10_145 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_33_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmux_right_track_2.mux_l1_in_0_ input82/X input80/X mux_right_track_2.mux_l1_in_1_/S
+ VGND VGND VPWR VPWR mux_right_track_2.mux_l1_in_0_/X sky130_fd_sc_hd__mux2_1
Xmux_left_track_33.mux_l1_in_1_ input61/X input54/X mux_left_track_33.mux_l1_in_2_/S
+ VGND VGND VPWR VPWR mux_left_track_33.mux_l1_in_1_/X sky130_fd_sc_hd__mux2_1
XANTENNA_mux_bottom_track_1.mux_l1_in_0__A0 input2/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xmux_bottom_track_1.mux_l1_in_3__172 VGND VGND VPWR VPWR mux_bottom_track_1.mux_l1_in_3_/A0
+ mux_bottom_track_1.mux_l1_in_3__172/LO sky130_fd_sc_hd__conb_1
XANTENNA_mux_left_track_5.mux_l1_in_4__A0 input74/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_33_18 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_24_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmux_bottom_track_15.sky130_fd_sc_hd__buf_4_0_ mux_bottom_track_15.mux_l2_in_0_/X
+ VGND VGND VPWR VPWR _104_/A sky130_fd_sc_hd__clkbuf_1
XANTENNA_mux_left_track_17.mux_l1_in_2__S mux_left_track_17.mux_l1_in_3_/S VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_23_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_23_73 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_064_ _064_/A VGND VGND VPWR VPWR _064_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_2_174 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_2_130 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_9_20 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmem_right_track_8.sky130_fd_sc_hd__dfxtp_1_3_ prog_clk_0_FTB00/X mux_right_track_8.mux_l3_in_1_/S
+ VGND VGND VPWR VPWR mux_right_track_8.mux_l4_in_0_/S sky130_fd_sc_hd__dfxtp_1
XFILLER_9_75 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_28_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_28_18 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_mux_left_track_1.mux_l1_in_1__S mux_left_track_1.mux_l1_in_1_/S VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
Xmux_bottom_track_3.mux_l3_in_0_ mux_bottom_track_3.mux_l2_in_1_/X mux_bottom_track_3.mux_l2_in_0_/X
+ mem_bottom_track_5.delay_buf_2/X VGND VGND VPWR VPWR mux_bottom_track_3.mux_l3_in_0_/X
+ sky130_fd_sc_hd__mux2_1
XFILLER_18_73 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_116_ _116_/A VGND VGND VPWR VPWR _116_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_28_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_input32_A chanx_right_in[10] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_6_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmux_bottom_track_3.mux_l2_in_1_ mux_bottom_track_3.mux_l1_in_3_/X mux_bottom_track_3.mux_l1_in_2_/X
+ mux_bottom_track_3.mux_l2_in_1_/S VGND VGND VPWR VPWR mux_bottom_track_3.mux_l2_in_1_/X
+ sky130_fd_sc_hd__mux2_1
XPHY_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_17_107 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_17_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_25_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_25_162 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_25_140 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_15_52 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_31_73 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_31_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_31_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_31_40 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_mux_left_track_9.mux_l1_in_0__A1 _064_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xoutput95 _070_/X VGND VGND VPWR VPWR chanx_left_out[13] sky130_fd_sc_hd__buf_2
XFILLER_16_173 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_31_143 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_110 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_121 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_132 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_187 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_176 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_165 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_143 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_154 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_22_176 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmem_right_track_2.sky130_fd_sc_hd__dfxtp_1_1_ prog_clk_0_FTB00/X mux_right_track_2.mux_l1_in_1_/S
+ VGND VGND VPWR VPWR mux_right_track_2.mux_l2_in_3_/S sky130_fd_sc_hd__dfxtp_2
XFILLER_13_132 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmux_bottom_track_3.mux_l1_in_2_ input24/X input9/X mux_bottom_track_3.mux_l1_in_3_/S
+ VGND VGND VPWR VPWR mux_bottom_track_3.mux_l1_in_2_/X sky130_fd_sc_hd__mux2_1
XFILLER_3_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_3_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_3_33 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xmem_left_track_17.sky130_fd_sc_hd__dfxtp_1_1_ prog_clk_0_FTB00/X mux_left_track_17.mux_l1_in_3_/S
+ VGND VGND VPWR VPWR mux_left_track_17.mux_l2_in_1_/S sky130_fd_sc_hd__dfxtp_1
Xmem_right_track_24.delay_buf_2 mem_right_track_24.delay_buf_2/X VGND VGND VPWR VPWR
+ mem_right_track_24.delay_buf_2/X sky130_fd_sc_hd__buf_6
Xmem_left_track_5.sky130_fd_sc_hd__dfxtp_1_0_ prog_clk_0_FTB00/X mux_left_track_3.mux_l4_in_0_/S
+ VGND VGND VPWR VPWR repeater154/A sky130_fd_sc_hd__dfxtp_1
XANTENNA_mem_bottom_track_9.sky130_fd_sc_hd__dfxtp_1_0__CLK prog_clk_0_FTB00/X VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_6_106 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_10_157 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_10_168 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_080_ _080_/A VGND VGND VPWR VPWR _080_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_6_128 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xmux_left_track_33.mux_l1_in_0_ input66/X _068_/A mux_left_track_33.mux_l1_in_2_/S
+ VGND VGND VPWR VPWR mux_left_track_33.mux_l1_in_0_/X sky130_fd_sc_hd__mux2_1
XANTENNA_mux_bottom_track_1.mux_l1_in_0__A1 _060_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_5_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_mux_left_track_5.mux_l2_in_2__S mux_left_track_5.mux_l2_in_3_/S VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mux_right_track_8.mux_l2_in_2__S mux_right_track_8.mux_l2_in_3_/S VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_30_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_15_216 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xmux_bottom_track_17.mux_l2_in_0_ mux_bottom_track_17.mux_l1_in_1_/X mux_bottom_track_17.mux_l1_in_0_/X
+ mux_bottom_track_17.mux_l2_in_0_/S VGND VGND VPWR VPWR mux_bottom_track_17.mux_l2_in_0_/X
+ sky130_fd_sc_hd__mux2_1
XFILLER_23_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_063_ _063_/A VGND VGND VPWR VPWR _063_/X sky130_fd_sc_hd__clkbuf_1
XANTENNA_input62_A chany_bottom_in[1] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_2_164 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_2_120 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_9_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_9_87 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmem_right_track_8.sky130_fd_sc_hd__dfxtp_1_2_ prog_clk_0_FTB00/X mux_right_track_8.mux_l2_in_3_/S
+ VGND VGND VPWR VPWR mux_right_track_8.mux_l3_in_1_/S sky130_fd_sc_hd__dfxtp_1
XFILLER_18_52 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_18_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_115_ _115_/A VGND VGND VPWR VPWR _115_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_29_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xmux_bottom_track_17.mux_l1_in_1_ mux_bottom_track_17.mux_l1_in_1_/A0 _091_/A mux_bottom_track_17.mux_l1_in_1_/S
+ VGND VGND VPWR VPWR mux_bottom_track_17.mux_l1_in_1_/X sky130_fd_sc_hd__mux2_1
XFILLER_20_20 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_20_64 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_20_75 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_29_84 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_input25_A chanx_left_in[4] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xmux_bottom_track_3.mux_l2_in_0_ mux_bottom_track_3.mux_l1_in_1_/X mux_bottom_track_3.mux_l1_in_0_/X
+ mux_bottom_track_3.mux_l2_in_1_/S VGND VGND VPWR VPWR mux_bottom_track_3.mux_l2_in_0_/X
+ sky130_fd_sc_hd__mux2_1
XANTENNA_mem_left_track_5.sky130_fd_sc_hd__dfxtp_1_3__CLK prog_clk_0_FTB00/X VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_19_171 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_25_152 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xoutput96 _071_/X VGND VGND VPWR VPWR chanx_left_out[14] sky130_fd_sc_hd__buf_2
XFILLER_31_122 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_16_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_16_185 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_mux_right_track_24.mux_l2_in_0__S mux_right_track_24.mux_l2_in_1_/S VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_166 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_100 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_111 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_mem_left_track_5.sky130_fd_sc_hd__dfxtp_1_2__D mux_left_track_5.mux_l2_in_3_/S
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_122 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_133 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_144 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_155 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
.ends

