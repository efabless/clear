VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO cbx_1__2_
  CLASS BLOCK ;
  FOREIGN cbx_1__2_ ;
  ORIGIN 0.000 0.000 ;
  SIZE 100.000 BY 86.000 ;
  PIN IO_ISOL_N
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 5.610 82.000 5.890 86.000 ;
    END
  END IO_ISOL_N
  PIN SC_IN_BOT
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 84.730 0.000 85.010 4.000 ;
    END
  END SC_IN_BOT
  PIN SC_IN_TOP
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 16.650 82.000 16.930 86.000 ;
    END
  END SC_IN_TOP
  PIN SC_OUT_BOT
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 88.870 0.000 89.150 4.000 ;
    END
  END SC_OUT_BOT
  PIN SC_OUT_TOP
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 27.690 82.000 27.970 86.000 ;
    END
  END SC_OUT_TOP
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 26.960 10.640 28.560 73.680 ;
    END
    PORT
      LAYER met4 ;
        RECT 49.200 10.640 50.800 73.680 ;
    END
    PORT
      LAYER met4 ;
        RECT 71.440 10.640 73.040 73.680 ;
    END
  END VGND
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 15.840 10.640 17.440 73.680 ;
    END
    PORT
      LAYER met4 ;
        RECT 38.080 10.640 39.680 73.680 ;
    END
    PORT
      LAYER met4 ;
        RECT 60.320 10.640 61.920 73.680 ;
    END
    PORT
      LAYER met4 ;
        RECT 82.560 10.640 84.160 73.680 ;
    END
  END VPWR
  PIN bottom_grid_pin_0_
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 10.210 0.000 10.490 4.000 ;
    END
  END bottom_grid_pin_0_
  PIN bottom_grid_pin_10_
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 51.610 0.000 51.890 4.000 ;
    END
  END bottom_grid_pin_10_
  PIN bottom_grid_pin_11_
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 55.750 0.000 56.030 4.000 ;
    END
  END bottom_grid_pin_11_
  PIN bottom_grid_pin_12_
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 59.890 0.000 60.170 4.000 ;
    END
  END bottom_grid_pin_12_
  PIN bottom_grid_pin_13_
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 64.030 0.000 64.310 4.000 ;
    END
  END bottom_grid_pin_13_
  PIN bottom_grid_pin_14_
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 68.170 0.000 68.450 4.000 ;
    END
  END bottom_grid_pin_14_
  PIN bottom_grid_pin_15_
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 72.310 0.000 72.590 4.000 ;
    END
  END bottom_grid_pin_15_
  PIN bottom_grid_pin_1_
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 14.350 0.000 14.630 4.000 ;
    END
  END bottom_grid_pin_1_
  PIN bottom_grid_pin_2_
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 18.490 0.000 18.770 4.000 ;
    END
  END bottom_grid_pin_2_
  PIN bottom_grid_pin_3_
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 22.630 0.000 22.910 4.000 ;
    END
  END bottom_grid_pin_3_
  PIN bottom_grid_pin_4_
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 26.770 0.000 27.050 4.000 ;
    END
  END bottom_grid_pin_4_
  PIN bottom_grid_pin_5_
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 30.910 0.000 31.190 4.000 ;
    END
  END bottom_grid_pin_5_
  PIN bottom_grid_pin_6_
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 35.050 0.000 35.330 4.000 ;
    END
  END bottom_grid_pin_6_
  PIN bottom_grid_pin_7_
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 39.190 0.000 39.470 4.000 ;
    END
  END bottom_grid_pin_7_
  PIN bottom_grid_pin_8_
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 43.330 0.000 43.610 4.000 ;
    END
  END bottom_grid_pin_8_
  PIN bottom_grid_pin_9_
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 47.470 0.000 47.750 4.000 ;
    END
  END bottom_grid_pin_9_
  PIN bottom_width_0_height_0__pin_0_
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 76.450 0.000 76.730 4.000 ;
    END
  END bottom_width_0_height_0__pin_0_
  PIN bottom_width_0_height_0__pin_1_lower
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 80.590 0.000 80.870 4.000 ;
    END
  END bottom_width_0_height_0__pin_1_lower
  PIN bottom_width_0_height_0__pin_1_upper
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 6.070 0.000 6.350 4.000 ;
    END
  END bottom_width_0_height_0__pin_1_upper
  PIN ccff_head
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 38.730 82.000 39.010 86.000 ;
    END
  END ccff_head
  PIN ccff_tail
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 49.770 82.000 50.050 86.000 ;
    END
  END ccff_tail
  PIN chanx_left_in[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 44.240 4.000 44.840 ;
    END
  END chanx_left_in[0]
  PIN chanx_left_in[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 64.640 4.000 65.240 ;
    END
  END chanx_left_in[10]
  PIN chanx_left_in[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 66.680 4.000 67.280 ;
    END
  END chanx_left_in[11]
  PIN chanx_left_in[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 68.720 4.000 69.320 ;
    END
  END chanx_left_in[12]
  PIN chanx_left_in[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 70.760 4.000 71.360 ;
    END
  END chanx_left_in[13]
  PIN chanx_left_in[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 72.800 4.000 73.400 ;
    END
  END chanx_left_in[14]
  PIN chanx_left_in[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 74.840 4.000 75.440 ;
    END
  END chanx_left_in[15]
  PIN chanx_left_in[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 76.880 4.000 77.480 ;
    END
  END chanx_left_in[16]
  PIN chanx_left_in[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 78.920 4.000 79.520 ;
    END
  END chanx_left_in[17]
  PIN chanx_left_in[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 80.960 4.000 81.560 ;
    END
  END chanx_left_in[18]
  PIN chanx_left_in[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 83.000 4.000 83.600 ;
    END
  END chanx_left_in[19]
  PIN chanx_left_in[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 46.280 4.000 46.880 ;
    END
  END chanx_left_in[1]
  PIN chanx_left_in[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 48.320 4.000 48.920 ;
    END
  END chanx_left_in[2]
  PIN chanx_left_in[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 50.360 4.000 50.960 ;
    END
  END chanx_left_in[3]
  PIN chanx_left_in[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 52.400 4.000 53.000 ;
    END
  END chanx_left_in[4]
  PIN chanx_left_in[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 54.440 4.000 55.040 ;
    END
  END chanx_left_in[5]
  PIN chanx_left_in[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 56.480 4.000 57.080 ;
    END
  END chanx_left_in[6]
  PIN chanx_left_in[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 58.520 4.000 59.120 ;
    END
  END chanx_left_in[7]
  PIN chanx_left_in[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 60.560 4.000 61.160 ;
    END
  END chanx_left_in[8]
  PIN chanx_left_in[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 62.600 4.000 63.200 ;
    END
  END chanx_left_in[9]
  PIN chanx_left_out[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 3.440 4.000 4.040 ;
    END
  END chanx_left_out[0]
  PIN chanx_left_out[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 23.840 4.000 24.440 ;
    END
  END chanx_left_out[10]
  PIN chanx_left_out[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 25.880 4.000 26.480 ;
    END
  END chanx_left_out[11]
  PIN chanx_left_out[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 27.920 4.000 28.520 ;
    END
  END chanx_left_out[12]
  PIN chanx_left_out[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 29.960 4.000 30.560 ;
    END
  END chanx_left_out[13]
  PIN chanx_left_out[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 32.000 4.000 32.600 ;
    END
  END chanx_left_out[14]
  PIN chanx_left_out[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 34.040 4.000 34.640 ;
    END
  END chanx_left_out[15]
  PIN chanx_left_out[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 36.080 4.000 36.680 ;
    END
  END chanx_left_out[16]
  PIN chanx_left_out[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 38.120 4.000 38.720 ;
    END
  END chanx_left_out[17]
  PIN chanx_left_out[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 40.160 4.000 40.760 ;
    END
  END chanx_left_out[18]
  PIN chanx_left_out[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 42.200 4.000 42.800 ;
    END
  END chanx_left_out[19]
  PIN chanx_left_out[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 5.480 4.000 6.080 ;
    END
  END chanx_left_out[1]
  PIN chanx_left_out[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 7.520 4.000 8.120 ;
    END
  END chanx_left_out[2]
  PIN chanx_left_out[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 9.560 4.000 10.160 ;
    END
  END chanx_left_out[3]
  PIN chanx_left_out[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 11.600 4.000 12.200 ;
    END
  END chanx_left_out[4]
  PIN chanx_left_out[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 13.640 4.000 14.240 ;
    END
  END chanx_left_out[5]
  PIN chanx_left_out[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 15.680 4.000 16.280 ;
    END
  END chanx_left_out[6]
  PIN chanx_left_out[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 17.720 4.000 18.320 ;
    END
  END chanx_left_out[7]
  PIN chanx_left_out[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 19.760 4.000 20.360 ;
    END
  END chanx_left_out[8]
  PIN chanx_left_out[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 21.800 4.000 22.400 ;
    END
  END chanx_left_out[9]
  PIN chanx_right_in[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 96.000 43.560 100.000 44.160 ;
    END
  END chanx_right_in[0]
  PIN chanx_right_in[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 96.000 63.960 100.000 64.560 ;
    END
  END chanx_right_in[10]
  PIN chanx_right_in[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 96.000 66.000 100.000 66.600 ;
    END
  END chanx_right_in[11]
  PIN chanx_right_in[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 96.000 68.040 100.000 68.640 ;
    END
  END chanx_right_in[12]
  PIN chanx_right_in[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 96.000 70.080 100.000 70.680 ;
    END
  END chanx_right_in[13]
  PIN chanx_right_in[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 96.000 72.120 100.000 72.720 ;
    END
  END chanx_right_in[14]
  PIN chanx_right_in[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 96.000 74.160 100.000 74.760 ;
    END
  END chanx_right_in[15]
  PIN chanx_right_in[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 96.000 76.200 100.000 76.800 ;
    END
  END chanx_right_in[16]
  PIN chanx_right_in[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 96.000 78.240 100.000 78.840 ;
    END
  END chanx_right_in[17]
  PIN chanx_right_in[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 96.000 80.280 100.000 80.880 ;
    END
  END chanx_right_in[18]
  PIN chanx_right_in[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 96.000 82.320 100.000 82.920 ;
    END
  END chanx_right_in[19]
  PIN chanx_right_in[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 96.000 45.600 100.000 46.200 ;
    END
  END chanx_right_in[1]
  PIN chanx_right_in[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 96.000 47.640 100.000 48.240 ;
    END
  END chanx_right_in[2]
  PIN chanx_right_in[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 96.000 49.680 100.000 50.280 ;
    END
  END chanx_right_in[3]
  PIN chanx_right_in[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 96.000 51.720 100.000 52.320 ;
    END
  END chanx_right_in[4]
  PIN chanx_right_in[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 96.000 53.760 100.000 54.360 ;
    END
  END chanx_right_in[5]
  PIN chanx_right_in[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 96.000 55.800 100.000 56.400 ;
    END
  END chanx_right_in[6]
  PIN chanx_right_in[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 96.000 57.840 100.000 58.440 ;
    END
  END chanx_right_in[7]
  PIN chanx_right_in[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 96.000 59.880 100.000 60.480 ;
    END
  END chanx_right_in[8]
  PIN chanx_right_in[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 96.000 61.920 100.000 62.520 ;
    END
  END chanx_right_in[9]
  PIN chanx_right_out[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 96.000 2.760 100.000 3.360 ;
    END
  END chanx_right_out[0]
  PIN chanx_right_out[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 96.000 23.160 100.000 23.760 ;
    END
  END chanx_right_out[10]
  PIN chanx_right_out[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 96.000 25.200 100.000 25.800 ;
    END
  END chanx_right_out[11]
  PIN chanx_right_out[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 96.000 27.240 100.000 27.840 ;
    END
  END chanx_right_out[12]
  PIN chanx_right_out[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 96.000 29.280 100.000 29.880 ;
    END
  END chanx_right_out[13]
  PIN chanx_right_out[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 96.000 31.320 100.000 31.920 ;
    END
  END chanx_right_out[14]
  PIN chanx_right_out[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 96.000 33.360 100.000 33.960 ;
    END
  END chanx_right_out[15]
  PIN chanx_right_out[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 96.000 35.400 100.000 36.000 ;
    END
  END chanx_right_out[16]
  PIN chanx_right_out[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 96.000 37.440 100.000 38.040 ;
    END
  END chanx_right_out[17]
  PIN chanx_right_out[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 96.000 39.480 100.000 40.080 ;
    END
  END chanx_right_out[18]
  PIN chanx_right_out[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 96.000 41.520 100.000 42.120 ;
    END
  END chanx_right_out[19]
  PIN chanx_right_out[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 96.000 4.800 100.000 5.400 ;
    END
  END chanx_right_out[1]
  PIN chanx_right_out[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 96.000 6.840 100.000 7.440 ;
    END
  END chanx_right_out[2]
  PIN chanx_right_out[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 96.000 8.880 100.000 9.480 ;
    END
  END chanx_right_out[3]
  PIN chanx_right_out[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 96.000 10.920 100.000 11.520 ;
    END
  END chanx_right_out[4]
  PIN chanx_right_out[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 96.000 12.960 100.000 13.560 ;
    END
  END chanx_right_out[5]
  PIN chanx_right_out[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 96.000 15.000 100.000 15.600 ;
    END
  END chanx_right_out[6]
  PIN chanx_right_out[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 96.000 17.040 100.000 17.640 ;
    END
  END chanx_right_out[7]
  PIN chanx_right_out[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 96.000 19.080 100.000 19.680 ;
    END
  END chanx_right_out[8]
  PIN chanx_right_out[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 96.000 21.120 100.000 21.720 ;
    END
  END chanx_right_out[9]
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_DIR
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 71.850 82.000 72.130 86.000 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_DIR
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_IN
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 82.890 82.000 83.170 86.000 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_IN
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_OUT
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 93.930 82.000 94.210 86.000 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_OUT
  PIN prog_clk_0_S_in
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 93.010 0.000 93.290 4.000 ;
    END
  END prog_clk_0_S_in
  PIN prog_clk_0_W_out
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1.400 4.000 2.000 ;
    END
  END prog_clk_0_W_out
  PIN top_grid_pin_0_
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 60.810 82.000 61.090 86.000 ;
    END
  END top_grid_pin_0_
  OBS
      LAYER li1 ;
        RECT 5.520 10.795 94.300 73.525 ;
      LAYER met1 ;
        RECT 4.670 7.520 96.990 76.800 ;
      LAYER met2 ;
        RECT 4.690 81.720 5.330 83.485 ;
        RECT 6.170 81.720 16.370 83.485 ;
        RECT 17.210 81.720 27.410 83.485 ;
        RECT 28.250 81.720 38.450 83.485 ;
        RECT 39.290 81.720 49.490 83.485 ;
        RECT 50.330 81.720 60.530 83.485 ;
        RECT 61.370 81.720 71.570 83.485 ;
        RECT 72.410 81.720 82.610 83.485 ;
        RECT 83.450 81.720 93.650 83.485 ;
        RECT 94.490 81.720 96.960 83.485 ;
        RECT 4.690 4.280 96.960 81.720 ;
        RECT 4.690 1.515 5.790 4.280 ;
        RECT 6.630 1.515 9.930 4.280 ;
        RECT 10.770 1.515 14.070 4.280 ;
        RECT 14.910 1.515 18.210 4.280 ;
        RECT 19.050 1.515 22.350 4.280 ;
        RECT 23.190 1.515 26.490 4.280 ;
        RECT 27.330 1.515 30.630 4.280 ;
        RECT 31.470 1.515 34.770 4.280 ;
        RECT 35.610 1.515 38.910 4.280 ;
        RECT 39.750 1.515 43.050 4.280 ;
        RECT 43.890 1.515 47.190 4.280 ;
        RECT 48.030 1.515 51.330 4.280 ;
        RECT 52.170 1.515 55.470 4.280 ;
        RECT 56.310 1.515 59.610 4.280 ;
        RECT 60.450 1.515 63.750 4.280 ;
        RECT 64.590 1.515 67.890 4.280 ;
        RECT 68.730 1.515 72.030 4.280 ;
        RECT 72.870 1.515 76.170 4.280 ;
        RECT 77.010 1.515 80.310 4.280 ;
        RECT 81.150 1.515 84.450 4.280 ;
        RECT 85.290 1.515 88.590 4.280 ;
        RECT 89.430 1.515 92.730 4.280 ;
        RECT 93.570 1.515 96.960 4.280 ;
      LAYER met3 ;
        RECT 4.400 83.320 96.000 83.465 ;
        RECT 4.400 82.600 95.600 83.320 ;
        RECT 4.000 81.960 95.600 82.600 ;
        RECT 4.400 81.920 95.600 81.960 ;
        RECT 4.400 81.280 96.000 81.920 ;
        RECT 4.400 80.560 95.600 81.280 ;
        RECT 4.000 79.920 95.600 80.560 ;
        RECT 4.400 79.880 95.600 79.920 ;
        RECT 4.400 79.240 96.000 79.880 ;
        RECT 4.400 78.520 95.600 79.240 ;
        RECT 4.000 77.880 95.600 78.520 ;
        RECT 4.400 77.840 95.600 77.880 ;
        RECT 4.400 77.200 96.000 77.840 ;
        RECT 4.400 76.480 95.600 77.200 ;
        RECT 4.000 75.840 95.600 76.480 ;
        RECT 4.400 75.800 95.600 75.840 ;
        RECT 4.400 75.160 96.000 75.800 ;
        RECT 4.400 74.440 95.600 75.160 ;
        RECT 4.000 73.800 95.600 74.440 ;
        RECT 4.400 73.760 95.600 73.800 ;
        RECT 4.400 73.120 96.000 73.760 ;
        RECT 4.400 72.400 95.600 73.120 ;
        RECT 4.000 71.760 95.600 72.400 ;
        RECT 4.400 71.720 95.600 71.760 ;
        RECT 4.400 71.080 96.000 71.720 ;
        RECT 4.400 70.360 95.600 71.080 ;
        RECT 4.000 69.720 95.600 70.360 ;
        RECT 4.400 69.680 95.600 69.720 ;
        RECT 4.400 69.040 96.000 69.680 ;
        RECT 4.400 68.320 95.600 69.040 ;
        RECT 4.000 67.680 95.600 68.320 ;
        RECT 4.400 67.640 95.600 67.680 ;
        RECT 4.400 67.000 96.000 67.640 ;
        RECT 4.400 66.280 95.600 67.000 ;
        RECT 4.000 65.640 95.600 66.280 ;
        RECT 4.400 65.600 95.600 65.640 ;
        RECT 4.400 64.960 96.000 65.600 ;
        RECT 4.400 64.240 95.600 64.960 ;
        RECT 4.000 63.600 95.600 64.240 ;
        RECT 4.400 63.560 95.600 63.600 ;
        RECT 4.400 62.920 96.000 63.560 ;
        RECT 4.400 62.200 95.600 62.920 ;
        RECT 4.000 61.560 95.600 62.200 ;
        RECT 4.400 61.520 95.600 61.560 ;
        RECT 4.400 60.880 96.000 61.520 ;
        RECT 4.400 60.160 95.600 60.880 ;
        RECT 4.000 59.520 95.600 60.160 ;
        RECT 4.400 59.480 95.600 59.520 ;
        RECT 4.400 58.840 96.000 59.480 ;
        RECT 4.400 58.120 95.600 58.840 ;
        RECT 4.000 57.480 95.600 58.120 ;
        RECT 4.400 57.440 95.600 57.480 ;
        RECT 4.400 56.800 96.000 57.440 ;
        RECT 4.400 56.080 95.600 56.800 ;
        RECT 4.000 55.440 95.600 56.080 ;
        RECT 4.400 55.400 95.600 55.440 ;
        RECT 4.400 54.760 96.000 55.400 ;
        RECT 4.400 54.040 95.600 54.760 ;
        RECT 4.000 53.400 95.600 54.040 ;
        RECT 4.400 53.360 95.600 53.400 ;
        RECT 4.400 52.720 96.000 53.360 ;
        RECT 4.400 52.000 95.600 52.720 ;
        RECT 4.000 51.360 95.600 52.000 ;
        RECT 4.400 51.320 95.600 51.360 ;
        RECT 4.400 50.680 96.000 51.320 ;
        RECT 4.400 49.960 95.600 50.680 ;
        RECT 4.000 49.320 95.600 49.960 ;
        RECT 4.400 49.280 95.600 49.320 ;
        RECT 4.400 48.640 96.000 49.280 ;
        RECT 4.400 47.920 95.600 48.640 ;
        RECT 4.000 47.280 95.600 47.920 ;
        RECT 4.400 47.240 95.600 47.280 ;
        RECT 4.400 46.600 96.000 47.240 ;
        RECT 4.400 45.880 95.600 46.600 ;
        RECT 4.000 45.240 95.600 45.880 ;
        RECT 4.400 45.200 95.600 45.240 ;
        RECT 4.400 44.560 96.000 45.200 ;
        RECT 4.400 43.840 95.600 44.560 ;
        RECT 4.000 43.200 95.600 43.840 ;
        RECT 4.400 43.160 95.600 43.200 ;
        RECT 4.400 42.520 96.000 43.160 ;
        RECT 4.400 41.800 95.600 42.520 ;
        RECT 4.000 41.160 95.600 41.800 ;
        RECT 4.400 41.120 95.600 41.160 ;
        RECT 4.400 40.480 96.000 41.120 ;
        RECT 4.400 39.760 95.600 40.480 ;
        RECT 4.000 39.120 95.600 39.760 ;
        RECT 4.400 39.080 95.600 39.120 ;
        RECT 4.400 38.440 96.000 39.080 ;
        RECT 4.400 37.720 95.600 38.440 ;
        RECT 4.000 37.080 95.600 37.720 ;
        RECT 4.400 37.040 95.600 37.080 ;
        RECT 4.400 36.400 96.000 37.040 ;
        RECT 4.400 35.680 95.600 36.400 ;
        RECT 4.000 35.040 95.600 35.680 ;
        RECT 4.400 35.000 95.600 35.040 ;
        RECT 4.400 34.360 96.000 35.000 ;
        RECT 4.400 33.640 95.600 34.360 ;
        RECT 4.000 33.000 95.600 33.640 ;
        RECT 4.400 32.960 95.600 33.000 ;
        RECT 4.400 32.320 96.000 32.960 ;
        RECT 4.400 31.600 95.600 32.320 ;
        RECT 4.000 30.960 95.600 31.600 ;
        RECT 4.400 30.920 95.600 30.960 ;
        RECT 4.400 30.280 96.000 30.920 ;
        RECT 4.400 29.560 95.600 30.280 ;
        RECT 4.000 28.920 95.600 29.560 ;
        RECT 4.400 28.880 95.600 28.920 ;
        RECT 4.400 28.240 96.000 28.880 ;
        RECT 4.400 27.520 95.600 28.240 ;
        RECT 4.000 26.880 95.600 27.520 ;
        RECT 4.400 26.840 95.600 26.880 ;
        RECT 4.400 26.200 96.000 26.840 ;
        RECT 4.400 25.480 95.600 26.200 ;
        RECT 4.000 24.840 95.600 25.480 ;
        RECT 4.400 24.800 95.600 24.840 ;
        RECT 4.400 24.160 96.000 24.800 ;
        RECT 4.400 23.440 95.600 24.160 ;
        RECT 4.000 22.800 95.600 23.440 ;
        RECT 4.400 22.760 95.600 22.800 ;
        RECT 4.400 22.120 96.000 22.760 ;
        RECT 4.400 21.400 95.600 22.120 ;
        RECT 4.000 20.760 95.600 21.400 ;
        RECT 4.400 20.720 95.600 20.760 ;
        RECT 4.400 20.080 96.000 20.720 ;
        RECT 4.400 19.360 95.600 20.080 ;
        RECT 4.000 18.720 95.600 19.360 ;
        RECT 4.400 18.680 95.600 18.720 ;
        RECT 4.400 18.040 96.000 18.680 ;
        RECT 4.400 17.320 95.600 18.040 ;
        RECT 4.000 16.680 95.600 17.320 ;
        RECT 4.400 16.640 95.600 16.680 ;
        RECT 4.400 16.000 96.000 16.640 ;
        RECT 4.400 15.280 95.600 16.000 ;
        RECT 4.000 14.640 95.600 15.280 ;
        RECT 4.400 14.600 95.600 14.640 ;
        RECT 4.400 13.960 96.000 14.600 ;
        RECT 4.400 13.240 95.600 13.960 ;
        RECT 4.000 12.600 95.600 13.240 ;
        RECT 4.400 12.560 95.600 12.600 ;
        RECT 4.400 11.920 96.000 12.560 ;
        RECT 4.400 11.200 95.600 11.920 ;
        RECT 4.000 10.560 95.600 11.200 ;
        RECT 4.400 10.520 95.600 10.560 ;
        RECT 4.400 9.880 96.000 10.520 ;
        RECT 4.400 9.160 95.600 9.880 ;
        RECT 4.000 8.520 95.600 9.160 ;
        RECT 4.400 8.480 95.600 8.520 ;
        RECT 4.400 7.840 96.000 8.480 ;
        RECT 4.400 7.120 95.600 7.840 ;
        RECT 4.000 6.480 95.600 7.120 ;
        RECT 4.400 6.440 95.600 6.480 ;
        RECT 4.400 5.800 96.000 6.440 ;
        RECT 4.400 5.080 95.600 5.800 ;
        RECT 4.000 4.440 95.600 5.080 ;
        RECT 4.400 4.400 95.600 4.440 ;
        RECT 4.400 3.760 96.000 4.400 ;
        RECT 4.400 3.040 95.600 3.760 ;
        RECT 4.000 2.400 95.600 3.040 ;
        RECT 4.400 2.360 95.600 2.400 ;
        RECT 4.400 1.535 96.000 2.360 ;
      LAYER met4 ;
        RECT 12.255 74.080 88.945 80.745 ;
        RECT 12.255 11.735 15.440 74.080 ;
        RECT 17.840 11.735 26.560 74.080 ;
        RECT 28.960 11.735 37.680 74.080 ;
        RECT 40.080 11.735 48.800 74.080 ;
        RECT 51.200 11.735 59.920 74.080 ;
        RECT 62.320 11.735 71.040 74.080 ;
        RECT 73.440 11.735 82.160 74.080 ;
        RECT 84.560 11.735 88.945 74.080 ;
  END
END cbx_1__2_
END LIBRARY

