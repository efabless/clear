magic
tech sky130A
magscale 1 2
timestamp 1656942746
<< viali >>
rect 9413 20417 9447 20451
rect 9965 20417 9999 20451
rect 20361 20417 20395 20451
rect 20637 20417 20671 20451
rect 21281 20349 21315 20383
rect 9229 20281 9263 20315
rect 9597 20281 9631 20315
rect 8309 20213 8343 20247
rect 9781 20213 9815 20247
rect 2789 20009 2823 20043
rect 7757 20009 7791 20043
rect 8677 20009 8711 20043
rect 10793 20009 10827 20043
rect 14473 20009 14507 20043
rect 9229 19941 9263 19975
rect 9597 19941 9631 19975
rect 13737 19941 13771 19975
rect 8125 19873 8159 19907
rect 21557 19873 21591 19907
rect 2973 19805 3007 19839
rect 7205 19805 7239 19839
rect 7573 19805 7607 19839
rect 8401 19805 8435 19839
rect 8493 19805 8527 19839
rect 9413 19805 9447 19839
rect 9781 19805 9815 19839
rect 9873 19805 9907 19839
rect 10241 19805 10275 19839
rect 10609 19805 10643 19839
rect 13001 19805 13035 19839
rect 13553 19805 13587 19839
rect 14105 19805 14139 19839
rect 14289 19805 14323 19839
rect 14657 19805 14691 19839
rect 16313 19805 16347 19839
rect 7113 19737 7147 19771
rect 9045 19737 9079 19771
rect 12734 19737 12768 19771
rect 16129 19737 16163 19771
rect 21290 19737 21324 19771
rect 6929 19669 6963 19703
rect 7389 19669 7423 19703
rect 10057 19669 10091 19703
rect 10425 19669 10459 19703
rect 11621 19669 11655 19703
rect 13093 19669 13127 19703
rect 13277 19669 13311 19703
rect 16497 19669 16531 19703
rect 20177 19669 20211 19703
rect 8309 19465 8343 19499
rect 9413 19465 9447 19499
rect 9873 19465 9907 19499
rect 11529 19465 11563 19499
rect 13001 19465 13035 19499
rect 19349 19465 19383 19499
rect 20913 19465 20947 19499
rect 21557 19465 21591 19499
rect 12642 19397 12676 19431
rect 14473 19397 14507 19431
rect 8125 19329 8159 19363
rect 8769 19329 8803 19363
rect 9229 19329 9263 19363
rect 9689 19329 9723 19363
rect 10057 19329 10091 19363
rect 12909 19329 12943 19363
rect 14114 19329 14148 19363
rect 20473 19329 20507 19363
rect 20729 19329 20763 19363
rect 8953 19261 8987 19295
rect 14381 19261 14415 19295
rect 8585 19125 8619 19159
rect 9137 19125 9171 19159
rect 10333 19125 10367 19159
rect 21005 18921 21039 18955
rect 8953 18785 8987 18819
rect 9413 18785 9447 18819
rect 13553 18785 13587 18819
rect 20913 18785 20947 18819
rect 8125 18717 8159 18751
rect 8769 18717 8803 18751
rect 9229 18717 9263 18751
rect 10057 18717 10091 18751
rect 11538 18717 11572 18751
rect 11805 18717 11839 18751
rect 11897 18717 11931 18751
rect 13461 18717 13495 18751
rect 13829 18717 13863 18751
rect 14749 18717 14783 18751
rect 16313 18717 16347 18751
rect 16681 18717 16715 18751
rect 18153 18717 18187 18751
rect 12142 18649 12176 18683
rect 14994 18649 15028 18683
rect 17886 18649 17920 18683
rect 20646 18649 20680 18683
rect 8309 18581 8343 18615
rect 8585 18581 8619 18615
rect 10241 18581 10275 18615
rect 10425 18581 10459 18615
rect 13277 18581 13311 18615
rect 16129 18581 16163 18615
rect 16773 18581 16807 18615
rect 18245 18581 18279 18615
rect 19533 18581 19567 18615
rect 2145 18377 2179 18411
rect 8033 18377 8067 18411
rect 8677 18377 8711 18411
rect 14657 18377 14691 18411
rect 15117 18377 15151 18411
rect 16681 18377 16715 18411
rect 18153 18377 18187 18411
rect 21097 18377 21131 18411
rect 4813 18309 4847 18343
rect 5549 18309 5583 18343
rect 2329 18241 2363 18275
rect 8585 18241 8619 18275
rect 9658 18241 9692 18275
rect 9781 18241 9815 18275
rect 12642 18241 12676 18275
rect 12909 18241 12943 18275
rect 14206 18241 14240 18275
rect 14473 18241 14507 18275
rect 16230 18241 16264 18275
rect 16497 18241 16531 18275
rect 17794 18241 17828 18275
rect 18061 18241 18095 18275
rect 19266 18241 19300 18275
rect 19533 18241 19567 18275
rect 19625 18241 19659 18275
rect 19881 18241 19915 18275
rect 4997 18173 5031 18207
rect 5641 18173 5675 18207
rect 5825 18173 5859 18207
rect 8861 18173 8895 18207
rect 9413 18173 9447 18207
rect 10057 18173 10091 18207
rect 11529 18105 11563 18139
rect 21005 18105 21039 18139
rect 5181 18037 5215 18071
rect 6101 18037 6135 18071
rect 7941 18037 7975 18071
rect 8217 18037 8251 18071
rect 11345 18037 11379 18071
rect 13093 18037 13127 18071
rect 2789 17833 2823 17867
rect 3801 17833 3835 17867
rect 8585 17833 8619 17867
rect 13461 17833 13495 17867
rect 18061 17833 18095 17867
rect 18245 17833 18279 17867
rect 19717 17833 19751 17867
rect 21281 17833 21315 17867
rect 13185 17765 13219 17799
rect 5181 17697 5215 17731
rect 5365 17697 5399 17731
rect 6469 17697 6503 17731
rect 6745 17697 6779 17731
rect 8033 17697 8067 17731
rect 11713 17697 11747 17731
rect 13645 17697 13679 17731
rect 16497 17697 16531 17731
rect 19809 17697 19843 17731
rect 2973 17629 3007 17663
rect 8217 17629 8251 17663
rect 9505 17629 9539 17663
rect 9781 17629 9815 17663
rect 16753 17629 16787 17663
rect 20065 17629 20099 17663
rect 4905 17561 4939 17595
rect 6285 17561 6319 17595
rect 8125 17561 8159 17595
rect 11980 17561 12014 17595
rect 5457 17493 5491 17527
rect 5825 17493 5859 17527
rect 5917 17493 5951 17527
rect 6377 17493 6411 17527
rect 7757 17493 7791 17527
rect 9873 17493 9907 17527
rect 13093 17493 13127 17527
rect 17877 17493 17911 17527
rect 21189 17493 21223 17527
rect 2237 17289 2271 17323
rect 3985 17289 4019 17323
rect 4445 17289 4479 17323
rect 4537 17289 4571 17323
rect 4905 17289 4939 17323
rect 5457 17289 5491 17323
rect 5917 17289 5951 17323
rect 6929 17289 6963 17323
rect 7389 17289 7423 17323
rect 7941 17289 7975 17323
rect 8309 17289 8343 17323
rect 9137 17289 9171 17323
rect 9229 17289 9263 17323
rect 9597 17289 9631 17323
rect 20545 17289 20579 17323
rect 3433 17221 3467 17255
rect 3893 17221 3927 17255
rect 7021 17221 7055 17255
rect 7849 17221 7883 17255
rect 8677 17221 8711 17255
rect 10057 17221 10091 17255
rect 10701 17221 10735 17255
rect 12664 17221 12698 17255
rect 14473 17221 14507 17255
rect 2421 17153 2455 17187
rect 2789 17153 2823 17187
rect 3157 17153 3191 17187
rect 3709 17153 3743 17187
rect 5549 17153 5583 17187
rect 9965 17153 9999 17187
rect 10425 17153 10459 17187
rect 13268 17153 13302 17187
rect 16230 17153 16264 17187
rect 16497 17153 16531 17187
rect 17794 17153 17828 17187
rect 19237 17153 19271 17187
rect 4353 17085 4387 17119
rect 4997 17085 5031 17119
rect 5273 17085 5307 17119
rect 6837 17085 6871 17119
rect 7757 17085 7791 17119
rect 9413 17085 9447 17119
rect 10241 17085 10275 17119
rect 12909 17085 12943 17119
rect 13001 17085 13035 17119
rect 18061 17085 18095 17119
rect 18153 17085 18187 17119
rect 18981 17085 19015 17119
rect 2973 17017 3007 17051
rect 8769 17017 8803 17051
rect 15117 17017 15151 17051
rect 2605 16949 2639 16983
rect 6009 16949 6043 16983
rect 8401 16949 8435 16983
rect 10977 16949 11011 16983
rect 11529 16949 11563 16983
rect 14381 16949 14415 16983
rect 16681 16949 16715 16983
rect 20361 16949 20395 16983
rect 3893 16745 3927 16779
rect 6561 16745 6595 16779
rect 14381 16745 14415 16779
rect 15853 16745 15887 16779
rect 16589 16745 16623 16779
rect 18337 16745 18371 16779
rect 20821 16745 20855 16779
rect 21281 16745 21315 16779
rect 3341 16609 3375 16643
rect 4169 16609 4203 16643
rect 6193 16609 6227 16643
rect 7573 16609 7607 16643
rect 7757 16609 7791 16643
rect 8125 16609 8159 16643
rect 9689 16609 9723 16643
rect 9873 16609 9907 16643
rect 10977 16609 11011 16643
rect 11621 16609 11655 16643
rect 13553 16609 13587 16643
rect 15761 16609 15795 16643
rect 18245 16609 18279 16643
rect 20637 16609 20671 16643
rect 2789 16541 2823 16575
rect 3065 16541 3099 16575
rect 3617 16541 3651 16575
rect 6377 16541 6411 16575
rect 9229 16541 9263 16575
rect 9505 16541 9539 16575
rect 9965 16541 9999 16575
rect 13277 16541 13311 16575
rect 20370 16541 20404 16575
rect 4353 16473 4387 16507
rect 7021 16473 7055 16507
rect 7481 16473 7515 16507
rect 8309 16473 8343 16507
rect 10793 16473 10827 16507
rect 11253 16473 11287 16507
rect 13010 16473 13044 16507
rect 13461 16473 13495 16507
rect 15494 16473 15528 16507
rect 16037 16473 16071 16507
rect 17978 16473 18012 16507
rect 4261 16405 4295 16439
rect 4721 16405 4755 16439
rect 4905 16405 4939 16439
rect 5549 16405 5583 16439
rect 5917 16405 5951 16439
rect 6009 16405 6043 16439
rect 7113 16405 7147 16439
rect 8217 16405 8251 16439
rect 8677 16405 8711 16439
rect 10333 16405 10367 16439
rect 10425 16405 10459 16439
rect 10885 16405 10919 16439
rect 11897 16405 11931 16439
rect 16865 16405 16899 16439
rect 19257 16405 19291 16439
rect 21465 16405 21499 16439
rect 4077 16201 4111 16235
rect 4353 16201 4387 16235
rect 5273 16201 5307 16235
rect 6101 16201 6135 16235
rect 7757 16201 7791 16235
rect 10609 16201 10643 16235
rect 11069 16201 11103 16235
rect 3065 16133 3099 16167
rect 3617 16133 3651 16167
rect 6929 16133 6963 16167
rect 9781 16133 9815 16167
rect 11529 16133 11563 16167
rect 19441 16133 19475 16167
rect 3341 16065 3375 16099
rect 3893 16065 3927 16099
rect 5733 16065 5767 16099
rect 6837 16065 6871 16099
rect 7849 16065 7883 16099
rect 10057 16065 10091 16099
rect 10701 16065 10735 16099
rect 13286 16065 13320 16099
rect 14953 16065 14987 16099
rect 15485 16065 15519 16099
rect 18990 16065 19024 16099
rect 19257 16065 19291 16099
rect 21198 16065 21232 16099
rect 21465 16065 21499 16099
rect 4905 15997 4939 16031
rect 5549 15997 5583 16031
rect 5641 15997 5675 16031
rect 6745 15997 6779 16031
rect 7665 15997 7699 16031
rect 10517 15997 10551 16031
rect 11161 15997 11195 16031
rect 13553 15997 13587 16031
rect 15209 15997 15243 16031
rect 15301 15997 15335 16031
rect 7297 15929 7331 15963
rect 8861 15929 8895 15963
rect 12173 15929 12207 15963
rect 6377 15861 6411 15895
rect 8217 15861 8251 15895
rect 8309 15861 8343 15895
rect 9229 15861 9263 15895
rect 9413 15861 9447 15895
rect 10149 15861 10183 15895
rect 13737 15861 13771 15895
rect 13829 15861 13863 15895
rect 17877 15861 17911 15895
rect 20085 15861 20119 15895
rect 1961 15657 1995 15691
rect 2329 15657 2363 15691
rect 2697 15657 2731 15691
rect 3617 15657 3651 15691
rect 5181 15657 5215 15691
rect 6009 15657 6043 15691
rect 6101 15657 6135 15691
rect 8953 15657 8987 15691
rect 9965 15657 9999 15691
rect 10241 15657 10275 15691
rect 8401 15589 8435 15623
rect 15853 15589 15887 15623
rect 4353 15521 4387 15555
rect 4629 15521 4663 15555
rect 5457 15521 5491 15555
rect 6561 15521 6595 15555
rect 6745 15521 6779 15555
rect 7757 15521 7791 15555
rect 7941 15521 7975 15555
rect 9413 15521 9447 15555
rect 9505 15521 9539 15555
rect 10885 15521 10919 15555
rect 2145 15453 2179 15487
rect 2513 15453 2547 15487
rect 2881 15453 2915 15487
rect 4813 15453 4847 15487
rect 6469 15453 6503 15487
rect 10609 15453 10643 15487
rect 13369 15453 13403 15487
rect 15229 15453 15263 15487
rect 15485 15453 15519 15487
rect 15669 15453 15703 15487
rect 16129 15453 16163 15487
rect 17601 15453 17635 15487
rect 19901 15453 19935 15487
rect 20085 15453 20119 15487
rect 21557 15453 21591 15487
rect 3893 15385 3927 15419
rect 5641 15385 5675 15419
rect 7573 15385 7607 15419
rect 9781 15385 9815 15419
rect 13124 15385 13158 15419
rect 16374 15385 16408 15419
rect 21290 15385 21324 15419
rect 3433 15317 3467 15351
rect 4169 15317 4203 15351
rect 4721 15317 4755 15351
rect 5549 15317 5583 15351
rect 8033 15317 8067 15351
rect 9321 15317 9355 15351
rect 10701 15317 10735 15351
rect 11069 15317 11103 15351
rect 11989 15317 12023 15351
rect 13553 15317 13587 15351
rect 14105 15317 14139 15351
rect 17509 15317 17543 15351
rect 20177 15317 20211 15351
rect 1961 15113 1995 15147
rect 2697 15113 2731 15147
rect 3341 15113 3375 15147
rect 4077 15113 4111 15147
rect 4169 15113 4203 15147
rect 5917 15113 5951 15147
rect 7481 15113 7515 15147
rect 7849 15113 7883 15147
rect 8217 15113 8251 15147
rect 8953 15113 8987 15147
rect 9045 15113 9079 15147
rect 9505 15113 9539 15147
rect 10609 15113 10643 15147
rect 11069 15113 11103 15147
rect 11621 15113 11655 15147
rect 13921 15113 13955 15147
rect 16681 15113 16715 15147
rect 2513 15045 2547 15079
rect 4905 15045 4939 15079
rect 7665 15045 7699 15079
rect 8309 15045 8343 15079
rect 21290 15045 21324 15079
rect 2145 14977 2179 15011
rect 2881 14977 2915 15011
rect 3249 14977 3283 15011
rect 4997 14977 5031 15011
rect 7113 14977 7147 15011
rect 9873 14977 9907 15011
rect 10977 14977 11011 15011
rect 13205 14977 13239 15011
rect 13461 14977 13495 15011
rect 15034 14977 15068 15011
rect 15301 14977 15335 15011
rect 15393 14977 15427 15011
rect 17794 14977 17828 15011
rect 19818 14977 19852 15011
rect 20085 14977 20119 15011
rect 21557 14977 21591 15011
rect 3157 14909 3191 14943
rect 3893 14909 3927 14943
rect 4721 14909 4755 14943
rect 5457 14909 5491 14943
rect 6101 14909 6135 14943
rect 6929 14909 6963 14943
rect 7021 14909 7055 14943
rect 8401 14909 8435 14943
rect 8769 14909 8803 14943
rect 9965 14909 9999 14943
rect 10149 14909 10183 14943
rect 11253 14909 11287 14943
rect 13645 14909 13679 14943
rect 18061 14909 18095 14943
rect 18153 14909 18187 14943
rect 4537 14841 4571 14875
rect 5733 14841 5767 14875
rect 16221 14841 16255 14875
rect 3709 14773 3743 14807
rect 5365 14773 5399 14807
rect 9413 14773 9447 14807
rect 10425 14773 10459 14807
rect 12081 14773 12115 14807
rect 18705 14773 18739 14807
rect 20177 14773 20211 14807
rect 3433 14569 3467 14603
rect 4629 14569 4663 14603
rect 6653 14569 6687 14603
rect 9873 14569 9907 14603
rect 15945 14569 15979 14603
rect 17693 14569 17727 14603
rect 21189 14569 21223 14603
rect 21465 14569 21499 14603
rect 3249 14501 3283 14535
rect 8401 14501 8435 14535
rect 3617 14433 3651 14467
rect 4077 14433 4111 14467
rect 5089 14433 5123 14467
rect 6101 14433 6135 14467
rect 6193 14433 6227 14467
rect 7481 14433 7515 14467
rect 8033 14433 8067 14467
rect 8217 14433 8251 14467
rect 9229 14433 9263 14467
rect 10609 14433 10643 14467
rect 13553 14433 13587 14467
rect 15853 14433 15887 14467
rect 17601 14433 17635 14467
rect 21097 14433 21131 14467
rect 4261 14365 4295 14399
rect 4721 14365 4755 14399
rect 5181 14365 5215 14399
rect 9505 14365 9539 14399
rect 10333 14365 10367 14399
rect 13286 14365 13320 14399
rect 15597 14365 15631 14399
rect 5273 14297 5307 14331
rect 9413 14297 9447 14331
rect 10425 14297 10459 14331
rect 17334 14297 17368 14331
rect 20830 14297 20864 14331
rect 4169 14229 4203 14263
rect 5641 14229 5675 14263
rect 6285 14229 6319 14263
rect 7573 14229 7607 14263
rect 7941 14229 7975 14263
rect 8585 14229 8619 14263
rect 9965 14229 9999 14263
rect 12173 14229 12207 14263
rect 13645 14229 13679 14263
rect 14473 14229 14507 14263
rect 16221 14229 16255 14263
rect 19717 14229 19751 14263
rect 4537 14025 4571 14059
rect 5365 14025 5399 14059
rect 5733 14025 5767 14059
rect 6377 14025 6411 14059
rect 7297 14025 7331 14059
rect 7757 14025 7791 14059
rect 10517 14025 10551 14059
rect 11069 14025 11103 14059
rect 11253 14025 11287 14059
rect 15117 14025 15151 14059
rect 18153 14025 18187 14059
rect 19717 14025 19751 14059
rect 21557 14025 21591 14059
rect 5917 13957 5951 13991
rect 6837 13957 6871 13991
rect 9229 13957 9263 13991
rect 16230 13957 16264 13991
rect 16926 13957 16960 13991
rect 19266 13957 19300 13991
rect 6745 13889 6779 13923
rect 7665 13889 7699 13923
rect 9689 13889 9723 13923
rect 12265 13889 12299 13923
rect 12521 13889 12555 13923
rect 16497 13889 16531 13923
rect 16681 13889 16715 13923
rect 19533 13889 19567 13923
rect 20177 13889 20211 13923
rect 20433 13889 20467 13923
rect 5089 13821 5123 13855
rect 5273 13821 5307 13855
rect 6101 13821 6135 13855
rect 6929 13821 6963 13855
rect 7849 13821 7883 13855
rect 9505 13821 9539 13855
rect 9597 13821 9631 13855
rect 10241 13821 10275 13855
rect 10425 13821 10459 13855
rect 10057 13753 10091 13787
rect 13645 13753 13679 13787
rect 18061 13753 18095 13787
rect 10885 13685 10919 13719
rect 13829 13685 13863 13719
rect 6101 13481 6135 13515
rect 7113 13481 7147 13515
rect 7941 13481 7975 13515
rect 13921 13481 13955 13515
rect 16129 13481 16163 13515
rect 21465 13481 21499 13515
rect 6193 13413 6227 13447
rect 8033 13413 8067 13447
rect 9413 13413 9447 13447
rect 11069 13413 11103 13447
rect 4721 13345 4755 13379
rect 6561 13345 6595 13379
rect 7297 13345 7331 13379
rect 7481 13345 7515 13379
rect 8677 13345 8711 13379
rect 9873 13345 9907 13379
rect 10057 13345 10091 13379
rect 10885 13345 10919 13379
rect 11713 13345 11747 13379
rect 2145 13277 2179 13311
rect 4997 13277 5031 13311
rect 10701 13277 10735 13311
rect 11529 13277 11563 13311
rect 12541 13277 12575 13311
rect 17509 13277 17543 13311
rect 19901 13277 19935 13311
rect 6653 13209 6687 13243
rect 12808 13209 12842 13243
rect 17242 13209 17276 13243
rect 20168 13209 20202 13243
rect 1961 13141 1995 13175
rect 6745 13141 6779 13175
rect 7573 13141 7607 13175
rect 8401 13141 8435 13175
rect 8493 13141 8527 13175
rect 9781 13141 9815 13175
rect 10241 13141 10275 13175
rect 10609 13141 10643 13175
rect 11437 13141 11471 13175
rect 14197 13141 14231 13175
rect 15945 13141 15979 13175
rect 17601 13141 17635 13175
rect 18153 13141 18187 13175
rect 21281 13141 21315 13175
rect 5089 12937 5123 12971
rect 5457 12937 5491 12971
rect 5917 12937 5951 12971
rect 6377 12937 6411 12971
rect 6745 12937 6779 12971
rect 7297 12937 7331 12971
rect 8585 12937 8619 12971
rect 9965 12937 9999 12971
rect 10425 12937 10459 12971
rect 18061 12937 18095 12971
rect 19533 12937 19567 12971
rect 21097 12937 21131 12971
rect 21373 12937 21407 12971
rect 3341 12869 3375 12903
rect 4261 12869 4295 12903
rect 10333 12869 10367 12903
rect 16926 12869 16960 12903
rect 3617 12801 3651 12835
rect 4537 12801 4571 12835
rect 4997 12801 5031 12835
rect 5825 12801 5859 12835
rect 6837 12801 6871 12835
rect 7573 12801 7607 12835
rect 8033 12801 8067 12835
rect 8953 12801 8987 12835
rect 13838 12801 13872 12835
rect 15310 12801 15344 12835
rect 15577 12801 15611 12835
rect 15669 12801 15703 12835
rect 16681 12801 16715 12835
rect 18409 12801 18443 12835
rect 20749 12801 20783 12835
rect 21005 12801 21039 12835
rect 5273 12733 5307 12767
rect 6101 12733 6135 12767
rect 7021 12733 7055 12767
rect 7757 12733 7791 12767
rect 7941 12733 7975 12767
rect 9045 12733 9079 12767
rect 9229 12733 9263 12767
rect 10609 12733 10643 12767
rect 14105 12733 14139 12767
rect 18153 12733 18187 12767
rect 4629 12665 4663 12699
rect 8401 12665 8435 12699
rect 12541 12597 12575 12631
rect 12725 12597 12759 12631
rect 14197 12597 14231 12631
rect 19625 12597 19659 12631
rect 1961 12393 1995 12427
rect 5641 12393 5675 12427
rect 7481 12393 7515 12427
rect 8401 12393 8435 12427
rect 10241 12393 10275 12427
rect 18153 12393 18187 12427
rect 18245 12393 18279 12427
rect 18429 12393 18463 12427
rect 19717 12393 19751 12427
rect 21281 12393 21315 12427
rect 8953 12325 8987 12359
rect 15301 12325 15335 12359
rect 5089 12257 5123 12291
rect 6285 12257 6319 12291
rect 8033 12257 8067 12291
rect 8585 12257 8619 12291
rect 9505 12257 9539 12291
rect 9781 12257 9815 12291
rect 10885 12257 10919 12291
rect 12449 12257 12483 12291
rect 12541 12257 12575 12291
rect 16681 12257 16715 12291
rect 16773 12257 16807 12291
rect 21189 12257 21223 12291
rect 2145 12189 2179 12223
rect 5365 12189 5399 12223
rect 10609 12189 10643 12223
rect 12182 12189 12216 12223
rect 16414 12189 16448 12223
rect 20922 12189 20956 12223
rect 10701 12121 10735 12155
rect 12786 12121 12820 12155
rect 17018 12121 17052 12155
rect 6009 12053 6043 12087
rect 6101 12053 6135 12087
rect 7297 12053 7331 12087
rect 7849 12053 7883 12087
rect 7941 12053 7975 12087
rect 9321 12053 9355 12087
rect 9413 12053 9447 12087
rect 11069 12053 11103 12087
rect 13921 12053 13955 12087
rect 14197 12053 14231 12087
rect 14381 12053 14415 12087
rect 19809 12053 19843 12087
rect 5457 11849 5491 11883
rect 6377 11849 6411 11883
rect 6837 11849 6871 11883
rect 7205 11849 7239 11883
rect 9321 11849 9355 11883
rect 9781 11849 9815 11883
rect 10149 11849 10183 11883
rect 10609 11849 10643 11883
rect 11529 11849 11563 11883
rect 18981 11849 19015 11883
rect 20913 11849 20947 11883
rect 4169 11781 4203 11815
rect 10517 11781 10551 11815
rect 11345 11781 11379 11815
rect 13676 11781 13710 11815
rect 4445 11713 4479 11747
rect 6193 11713 6227 11747
rect 6745 11713 6779 11747
rect 8033 11713 8067 11747
rect 9689 11713 9723 11747
rect 11897 11713 11931 11747
rect 17765 11713 17799 11747
rect 20462 11713 20496 11747
rect 20729 11713 20763 11747
rect 5181 11645 5215 11679
rect 6009 11645 6043 11679
rect 7021 11645 7055 11679
rect 7757 11645 7791 11679
rect 7941 11645 7975 11679
rect 9965 11645 9999 11679
rect 10793 11645 10827 11679
rect 11989 11645 12023 11679
rect 12173 11645 12207 11679
rect 12357 11645 12391 11679
rect 13921 11645 13955 11679
rect 17509 11645 17543 11679
rect 8401 11577 8435 11611
rect 12541 11577 12575 11611
rect 8585 11509 8619 11543
rect 11161 11509 11195 11543
rect 14013 11509 14047 11543
rect 16405 11509 16439 11543
rect 16773 11509 16807 11543
rect 18889 11509 18923 11543
rect 19349 11509 19383 11543
rect 1961 11305 1995 11339
rect 5365 11305 5399 11339
rect 6193 11305 6227 11339
rect 7021 11305 7055 11339
rect 7389 11305 7423 11339
rect 10057 11305 10091 11339
rect 11161 11305 11195 11339
rect 11345 11305 11379 11339
rect 14933 11305 14967 11339
rect 21189 11305 21223 11339
rect 2329 11237 2363 11271
rect 8953 11237 8987 11271
rect 12909 11237 12943 11271
rect 13645 11237 13679 11271
rect 16405 11237 16439 11271
rect 19625 11237 19659 11271
rect 4813 11169 4847 11203
rect 5641 11169 5675 11203
rect 6469 11169 6503 11203
rect 9597 11169 9631 11203
rect 10517 11169 10551 11203
rect 10609 11169 10643 11203
rect 11529 11169 11563 11203
rect 17785 11169 17819 11203
rect 21005 11169 21039 11203
rect 2145 11101 2179 11135
rect 2513 11101 2547 11135
rect 16313 11101 16347 11135
rect 17877 11101 17911 11135
rect 4261 11033 4295 11067
rect 4905 11033 4939 11067
rect 4997 11033 5031 11067
rect 5825 11033 5859 11067
rect 7113 11033 7147 11067
rect 9321 11033 9355 11067
rect 11069 11033 11103 11067
rect 11796 11033 11830 11067
rect 13093 11033 13127 11067
rect 16068 11033 16102 11067
rect 17518 11033 17552 11067
rect 18153 11033 18187 11067
rect 20738 11033 20772 11067
rect 4537 10965 4571 10999
rect 5733 10965 5767 10999
rect 6561 10965 6595 10999
rect 6653 10965 6687 10999
rect 8585 10965 8619 10999
rect 9413 10965 9447 10999
rect 9873 10965 9907 10999
rect 10425 10965 10459 10999
rect 13277 10965 13311 10999
rect 13369 10965 13403 10999
rect 3801 10761 3835 10795
rect 4721 10761 4755 10795
rect 5089 10761 5123 10795
rect 5917 10761 5951 10795
rect 7113 10761 7147 10795
rect 8217 10761 8251 10795
rect 8677 10761 8711 10795
rect 9045 10761 9079 10795
rect 9137 10761 9171 10795
rect 10333 10761 10367 10795
rect 16497 10761 16531 10795
rect 21005 10761 21039 10795
rect 6745 10693 6779 10727
rect 9597 10693 9631 10727
rect 12664 10693 12698 10727
rect 14473 10693 14507 10727
rect 14657 10693 14691 10727
rect 15384 10693 15418 10727
rect 5549 10625 5583 10659
rect 6009 10625 6043 10659
rect 7849 10625 7883 10659
rect 9505 10625 9539 10659
rect 10241 10625 10275 10659
rect 10701 10625 10735 10659
rect 12909 10625 12943 10659
rect 13001 10625 13035 10659
rect 13268 10625 13302 10659
rect 15117 10625 15151 10659
rect 16681 10625 16715 10659
rect 16937 10625 16971 10659
rect 20554 10625 20588 10659
rect 20821 10625 20855 10659
rect 2973 10557 3007 10591
rect 4261 10557 4295 10591
rect 4445 10557 4479 10591
rect 4629 10557 4663 10591
rect 5365 10557 5399 10591
rect 5457 10557 5491 10591
rect 6561 10557 6595 10591
rect 6653 10557 6687 10591
rect 7573 10557 7607 10591
rect 7757 10557 7791 10591
rect 8493 10557 8527 10591
rect 8585 10557 8619 10591
rect 9781 10557 9815 10591
rect 10793 10557 10827 10591
rect 10885 10557 10919 10591
rect 11253 10557 11287 10591
rect 18153 10557 18187 10591
rect 18337 10557 18371 10591
rect 3985 10421 4019 10455
rect 7297 10421 7331 10455
rect 11529 10421 11563 10455
rect 14381 10421 14415 10455
rect 18061 10421 18095 10455
rect 19441 10421 19475 10455
rect 1869 10217 1903 10251
rect 2145 10217 2179 10251
rect 3157 10217 3191 10251
rect 4629 10217 4663 10251
rect 5641 10217 5675 10251
rect 7297 10217 7331 10251
rect 8953 10217 8987 10251
rect 10149 10217 10183 10251
rect 19533 10217 19567 10251
rect 21005 10217 21039 10251
rect 4537 10149 4571 10183
rect 7205 10149 7239 10183
rect 13553 10149 13587 10183
rect 2605 10081 2639 10115
rect 3985 10081 4019 10115
rect 4997 10081 5031 10115
rect 5549 10081 5583 10115
rect 6193 10081 6227 10115
rect 6653 10081 6687 10115
rect 7849 10081 7883 10115
rect 8125 10081 8159 10115
rect 9413 10081 9447 10115
rect 9597 10081 9631 10115
rect 18797 10081 18831 10115
rect 20913 10081 20947 10115
rect 2329 10013 2363 10047
rect 2789 10013 2823 10047
rect 5273 10013 5307 10047
rect 6837 10013 6871 10047
rect 8401 10013 8435 10047
rect 11989 10013 12023 10047
rect 13461 10013 13495 10047
rect 14197 10013 14231 10047
rect 14464 10013 14498 10047
rect 17049 10013 17083 10047
rect 17141 10013 17175 10047
rect 3617 9945 3651 9979
rect 4169 9945 4203 9979
rect 6009 9945 6043 9979
rect 6745 9945 6779 9979
rect 8769 9945 8803 9979
rect 9321 9945 9355 9979
rect 10333 9945 10367 9979
rect 11744 9945 11778 9979
rect 13216 9945 13250 9979
rect 16782 9945 16816 9979
rect 17386 9945 17420 9979
rect 20646 9945 20680 9979
rect 2697 9877 2731 9911
rect 3249 9877 3283 9911
rect 4077 9877 4111 9911
rect 6101 9877 6135 9911
rect 7665 9877 7699 9911
rect 7757 9877 7791 9911
rect 9781 9877 9815 9911
rect 10609 9877 10643 9911
rect 12081 9877 12115 9911
rect 13829 9877 13863 9911
rect 15577 9877 15611 9911
rect 15669 9877 15703 9911
rect 18521 9877 18555 9911
rect 18705 9877 18739 9911
rect 18981 9877 19015 9911
rect 3341 9673 3375 9707
rect 8769 9673 8803 9707
rect 12081 9673 12115 9707
rect 13645 9673 13679 9707
rect 19533 9673 19567 9707
rect 6745 9605 6779 9639
rect 9321 9605 9355 9639
rect 16230 9605 16264 9639
rect 1777 9537 1811 9571
rect 2145 9537 2179 9571
rect 2789 9537 2823 9571
rect 2881 9537 2915 9571
rect 3709 9537 3743 9571
rect 4813 9537 4847 9571
rect 4905 9537 4939 9571
rect 5457 9537 5491 9571
rect 6101 9537 6135 9571
rect 6653 9537 6687 9571
rect 10333 9537 10367 9571
rect 10425 9537 10459 9571
rect 11069 9537 11103 9571
rect 13286 9537 13320 9571
rect 14758 9537 14792 9571
rect 15025 9537 15059 9571
rect 16497 9537 16531 9571
rect 17794 9537 17828 9571
rect 18409 9537 18443 9571
rect 19881 9537 19915 9571
rect 2513 9469 2547 9503
rect 3801 9469 3835 9503
rect 4261 9469 4295 9503
rect 4629 9469 4663 9503
rect 6469 9469 6503 9503
rect 9137 9469 9171 9503
rect 9229 9469 9263 9503
rect 10609 9469 10643 9503
rect 10793 9469 10827 9503
rect 13553 9469 13587 9503
rect 18061 9469 18095 9503
rect 18153 9469 18187 9503
rect 19625 9469 19659 9503
rect 1593 9401 1627 9435
rect 1961 9401 1995 9435
rect 3065 9401 3099 9435
rect 5273 9401 5307 9435
rect 5917 9401 5951 9435
rect 7113 9401 7147 9435
rect 9689 9401 9723 9435
rect 9873 9401 9907 9435
rect 11345 9401 11379 9435
rect 3985 9333 4019 9367
rect 4353 9333 4387 9367
rect 5733 9333 5767 9367
rect 7205 9333 7239 9367
rect 8217 9333 8251 9367
rect 8585 9333 8619 9367
rect 9965 9333 9999 9367
rect 12173 9333 12207 9367
rect 15117 9333 15151 9367
rect 16681 9333 16715 9367
rect 21005 9333 21039 9367
rect 21189 9333 21223 9367
rect 21281 9333 21315 9367
rect 1685 9129 1719 9163
rect 2973 9129 3007 9163
rect 6101 9129 6135 9163
rect 9505 9129 9539 9163
rect 9689 9129 9723 9163
rect 15669 9129 15703 9163
rect 15853 9129 15887 9163
rect 16037 9129 16071 9163
rect 16221 9129 16255 9163
rect 17877 9129 17911 9163
rect 18245 9129 18279 9163
rect 1961 9061 1995 9095
rect 5273 9061 5307 9095
rect 7021 9061 7055 9095
rect 12265 9061 12299 9095
rect 2421 8993 2455 9027
rect 3249 8993 3283 9027
rect 4629 8993 4663 9027
rect 5457 8993 5491 9027
rect 5641 8993 5675 9027
rect 6837 8993 6871 9027
rect 7665 8993 7699 9027
rect 8401 8993 8435 9027
rect 10149 8993 10183 9027
rect 10333 8993 10367 9027
rect 10701 8993 10735 9027
rect 11989 8993 12023 9027
rect 13645 8993 13679 9027
rect 13829 8993 13863 9027
rect 14105 8993 14139 9027
rect 16313 8993 16347 9027
rect 2145 8925 2179 8959
rect 2605 8925 2639 8959
rect 3525 8925 3559 8959
rect 4353 8925 4387 8959
rect 4905 8925 4939 8959
rect 10793 8925 10827 8959
rect 20637 8925 20671 8959
rect 1593 8857 1627 8891
rect 2513 8857 2547 8891
rect 4077 8857 4111 8891
rect 5733 8857 5767 8891
rect 7389 8857 7423 8891
rect 11713 8857 11747 8891
rect 13378 8857 13412 8891
rect 14350 8857 14384 8891
rect 16580 8857 16614 8891
rect 20370 8857 20404 8891
rect 4813 8789 4847 8823
rect 6193 8789 6227 8823
rect 6561 8789 6595 8823
rect 6653 8789 6687 8823
rect 7481 8789 7515 8823
rect 7849 8789 7883 8823
rect 8217 8789 8251 8823
rect 8309 8789 8343 8823
rect 8677 8789 8711 8823
rect 10057 8789 10091 8823
rect 10885 8789 10919 8823
rect 11253 8789 11287 8823
rect 11345 8789 11379 8823
rect 11805 8789 11839 8823
rect 15485 8789 15519 8823
rect 17693 8789 17727 8823
rect 19257 8789 19291 8823
rect 20821 8789 20855 8823
rect 2237 8585 2271 8619
rect 2605 8585 2639 8619
rect 4813 8585 4847 8619
rect 6193 8585 6227 8619
rect 8953 8585 8987 8619
rect 9965 8585 9999 8619
rect 10517 8585 10551 8619
rect 10977 8585 11011 8619
rect 13829 8585 13863 8619
rect 15761 8585 15795 8619
rect 20821 8585 20855 8619
rect 2881 8517 2915 8551
rect 3249 8517 3283 8551
rect 8033 8517 8067 8551
rect 8125 8517 8159 8551
rect 9413 8517 9447 8551
rect 19686 8517 19720 8551
rect 3157 8449 3191 8483
rect 3525 8449 3559 8483
rect 3985 8449 4019 8483
rect 4353 8449 4387 8483
rect 4445 8449 4479 8483
rect 4905 8449 4939 8483
rect 5825 8449 5859 8483
rect 6653 8449 6687 8483
rect 7297 8449 7331 8483
rect 10057 8449 10091 8483
rect 10885 8449 10919 8483
rect 11529 8449 11563 8483
rect 15402 8449 15436 8483
rect 15669 8449 15703 8483
rect 19082 8449 19116 8483
rect 2053 8381 2087 8415
rect 2145 8381 2179 8415
rect 3709 8381 3743 8415
rect 4261 8381 4295 8415
rect 5549 8381 5583 8415
rect 5733 8381 5767 8415
rect 7389 8381 7423 8415
rect 7573 8381 7607 8415
rect 7941 8381 7975 8415
rect 9045 8381 9079 8415
rect 9229 8381 9263 8415
rect 9873 8381 9907 8415
rect 11069 8381 11103 8415
rect 19349 8381 19383 8415
rect 19441 8381 19475 8415
rect 1501 8313 1535 8347
rect 1685 8313 1719 8347
rect 6929 8313 6963 8347
rect 8493 8313 8527 8347
rect 14289 8313 14323 8347
rect 5273 8245 5307 8279
rect 6377 8245 6411 8279
rect 6837 8245 6871 8279
rect 8585 8245 8619 8279
rect 10425 8245 10459 8279
rect 17969 8245 18003 8279
rect 21005 8245 21039 8279
rect 1501 8041 1535 8075
rect 3249 8041 3283 8075
rect 6469 8041 6503 8075
rect 7849 8041 7883 8075
rect 14381 8041 14415 8075
rect 14841 8041 14875 8075
rect 15761 8041 15795 8075
rect 19901 8041 19935 8075
rect 11897 7973 11931 8007
rect 17877 7973 17911 8007
rect 1961 7905 1995 7939
rect 2053 7905 2087 7939
rect 2881 7905 2915 7939
rect 4905 7905 4939 7939
rect 5549 7905 5583 7939
rect 7113 7905 7147 7939
rect 8401 7905 8435 7939
rect 9321 7905 9355 7939
rect 11253 7905 11287 7939
rect 12541 7905 12575 7939
rect 16681 7905 16715 7939
rect 18521 7905 18555 7939
rect 21281 7905 21315 7939
rect 21373 7905 21407 7939
rect 3065 7837 3099 7871
rect 5825 7837 5859 7871
rect 6377 7837 6411 7871
rect 6929 7837 6963 7871
rect 9413 7837 9447 7871
rect 16405 7837 16439 7871
rect 18337 7837 18371 7871
rect 19533 7837 19567 7871
rect 3341 7769 3375 7803
rect 5181 7769 5215 7803
rect 6101 7769 6135 7803
rect 8217 7769 8251 7803
rect 9505 7769 9539 7803
rect 9965 7769 9999 7803
rect 10425 7769 10459 7803
rect 10701 7769 10735 7803
rect 10977 7769 11011 7803
rect 11437 7769 11471 7803
rect 21014 7769 21048 7803
rect 2145 7701 2179 7735
rect 2513 7701 2547 7735
rect 4997 7701 5031 7735
rect 6837 7701 6871 7735
rect 7297 7701 7331 7735
rect 7573 7701 7607 7735
rect 8309 7701 8343 7735
rect 8677 7701 8711 7735
rect 9873 7701 9907 7735
rect 11345 7701 11379 7735
rect 11805 7701 11839 7735
rect 12265 7701 12299 7735
rect 12357 7701 12391 7735
rect 14289 7701 14323 7735
rect 15853 7701 15887 7735
rect 16037 7701 16071 7735
rect 16497 7701 16531 7735
rect 17509 7701 17543 7735
rect 17693 7701 17727 7735
rect 18245 7701 18279 7735
rect 1685 7497 1719 7531
rect 4261 7497 4295 7531
rect 4905 7497 4939 7531
rect 6193 7497 6227 7531
rect 7573 7497 7607 7531
rect 9137 7497 9171 7531
rect 9597 7497 9631 7531
rect 10517 7497 10551 7531
rect 12081 7497 12115 7531
rect 13461 7497 13495 7531
rect 14657 7497 14691 7531
rect 15117 7497 15151 7531
rect 15577 7497 15611 7531
rect 19349 7497 19383 7531
rect 20913 7497 20947 7531
rect 1501 7429 1535 7463
rect 9505 7429 9539 7463
rect 14749 7429 14783 7463
rect 4537 7361 4571 7395
rect 4997 7361 5031 7395
rect 5825 7361 5859 7395
rect 6837 7361 6871 7395
rect 7297 7361 7331 7395
rect 7941 7361 7975 7395
rect 8033 7361 8067 7395
rect 10885 7361 10919 7395
rect 11529 7361 11563 7395
rect 12449 7361 12483 7395
rect 12909 7361 12943 7395
rect 13829 7361 13863 7395
rect 15485 7361 15519 7395
rect 20462 7361 20496 7395
rect 20729 7361 20763 7395
rect 4813 7293 4847 7327
rect 5549 7293 5583 7327
rect 5733 7293 5767 7327
rect 6929 7293 6963 7327
rect 7113 7293 7147 7327
rect 8217 7293 8251 7327
rect 9689 7293 9723 7327
rect 10977 7293 11011 7327
rect 11069 7293 11103 7327
rect 12541 7293 12575 7327
rect 12725 7293 12759 7327
rect 13921 7293 13955 7327
rect 14105 7293 14139 7327
rect 14933 7293 14967 7327
rect 15761 7293 15795 7327
rect 6469 7225 6503 7259
rect 14289 7225 14323 7259
rect 5365 7157 5399 7191
rect 9965 7157 9999 7191
rect 10333 7157 10367 7191
rect 11897 7157 11931 7191
rect 6469 6953 6503 6987
rect 7389 6953 7423 6987
rect 8401 6953 8435 6987
rect 9321 6953 9355 6987
rect 14105 6953 14139 6987
rect 3985 6817 4019 6851
rect 4169 6817 4203 6851
rect 7021 6817 7055 6851
rect 7757 6817 7791 6851
rect 8585 6817 8619 6851
rect 9873 6817 9907 6851
rect 10241 6817 10275 6851
rect 11989 6817 12023 6851
rect 14565 6817 14599 6851
rect 14657 6817 14691 6851
rect 14933 6817 14967 6851
rect 3433 6749 3467 6783
rect 4261 6749 4295 6783
rect 6837 6749 6871 6783
rect 8953 6749 8987 6783
rect 9689 6749 9723 6783
rect 12081 6749 12115 6783
rect 3617 6681 3651 6715
rect 10517 6681 10551 6715
rect 4629 6613 4663 6647
rect 4813 6613 4847 6647
rect 5549 6613 5583 6647
rect 5733 6613 5767 6647
rect 5917 6613 5951 6647
rect 6101 6613 6135 6647
rect 6377 6613 6411 6647
rect 6929 6613 6963 6647
rect 7481 6613 7515 6647
rect 7941 6613 7975 6647
rect 8033 6613 8067 6647
rect 9137 6613 9171 6647
rect 9781 6613 9815 6647
rect 10425 6613 10459 6647
rect 10885 6613 10919 6647
rect 11621 6613 11655 6647
rect 12173 6613 12207 6647
rect 12541 6613 12575 6647
rect 13829 6613 13863 6647
rect 14473 6613 14507 6647
rect 2421 6409 2455 6443
rect 5181 6409 5215 6443
rect 5641 6409 5675 6443
rect 7113 6409 7147 6443
rect 7481 6409 7515 6443
rect 7941 6409 7975 6443
rect 8401 6409 8435 6443
rect 8769 6409 8803 6443
rect 9229 6409 9263 6443
rect 9965 6409 9999 6443
rect 12265 6409 12299 6443
rect 12725 6409 12759 6443
rect 14197 6409 14231 6443
rect 14289 6409 14323 6443
rect 3985 6341 4019 6375
rect 4353 6341 4387 6375
rect 4445 6341 4479 6375
rect 5733 6341 5767 6375
rect 2053 6273 2087 6307
rect 5273 6273 5307 6307
rect 6193 6273 6227 6307
rect 7021 6273 7055 6307
rect 8309 6273 8343 6307
rect 9137 6273 9171 6307
rect 10057 6273 10091 6307
rect 10977 6273 11011 6307
rect 12633 6273 12667 6307
rect 1869 6205 1903 6239
rect 1961 6205 1995 6239
rect 4169 6205 4203 6239
rect 5089 6205 5123 6239
rect 7573 6205 7607 6239
rect 7757 6205 7791 6239
rect 8585 6205 8619 6239
rect 9413 6205 9447 6239
rect 9873 6205 9907 6239
rect 10701 6205 10735 6239
rect 10885 6205 10919 6239
rect 11529 6205 11563 6239
rect 11713 6205 11747 6239
rect 12817 6205 12851 6239
rect 14105 6205 14139 6239
rect 4813 6137 4847 6171
rect 10425 6137 10459 6171
rect 11345 6137 11379 6171
rect 1501 6069 1535 6103
rect 6377 6069 6411 6103
rect 12081 6069 12115 6103
rect 14657 6069 14691 6103
rect 1501 5865 1535 5899
rect 5365 5865 5399 5899
rect 7205 5865 7239 5899
rect 7757 5865 7791 5899
rect 8769 5865 8803 5899
rect 11161 5865 11195 5899
rect 13277 5865 13311 5899
rect 7665 5797 7699 5831
rect 8953 5797 8987 5831
rect 9137 5797 9171 5831
rect 17325 5797 17359 5831
rect 5733 5729 5767 5763
rect 6561 5729 6595 5763
rect 8217 5729 8251 5763
rect 9689 5729 9723 5763
rect 10609 5729 10643 5763
rect 11621 5729 11655 5763
rect 12725 5729 12759 5763
rect 16681 5729 16715 5763
rect 17601 5729 17635 5763
rect 20177 5729 20211 5763
rect 5917 5661 5951 5695
rect 11805 5661 11839 5695
rect 13369 5661 13403 5695
rect 16865 5661 16899 5695
rect 6837 5593 6871 5627
rect 8309 5593 8343 5627
rect 9597 5593 9631 5627
rect 13645 5593 13679 5627
rect 17693 5593 17727 5627
rect 20361 5593 20395 5627
rect 4997 5525 5031 5559
rect 5181 5525 5215 5559
rect 5457 5525 5491 5559
rect 6009 5525 6043 5559
rect 6377 5525 6411 5559
rect 6745 5525 6779 5559
rect 8401 5525 8435 5559
rect 9505 5525 9539 5559
rect 10701 5525 10735 5559
rect 10793 5525 10827 5559
rect 11713 5525 11747 5559
rect 12173 5525 12207 5559
rect 12817 5525 12851 5559
rect 12909 5525 12943 5559
rect 16957 5525 16991 5559
rect 17785 5525 17819 5559
rect 18153 5525 18187 5559
rect 20269 5525 20303 5559
rect 20729 5525 20763 5559
rect 1777 5321 1811 5355
rect 2145 5321 2179 5355
rect 4721 5321 4755 5355
rect 5089 5321 5123 5355
rect 6653 5321 6687 5355
rect 7113 5321 7147 5355
rect 7941 5321 7975 5355
rect 8401 5321 8435 5355
rect 9045 5321 9079 5355
rect 9689 5321 9723 5355
rect 10149 5321 10183 5355
rect 10977 5321 11011 5355
rect 11897 5321 11931 5355
rect 13185 5321 13219 5355
rect 13829 5321 13863 5355
rect 17233 5321 17267 5355
rect 5549 5253 5583 5287
rect 11989 5253 12023 5287
rect 2237 5185 2271 5219
rect 2697 5185 2731 5219
rect 4629 5185 4663 5219
rect 6745 5185 6779 5219
rect 8309 5185 8343 5219
rect 8769 5185 8803 5219
rect 9781 5185 9815 5219
rect 10609 5185 10643 5219
rect 12817 5185 12851 5219
rect 13277 5185 13311 5219
rect 15393 5185 15427 5219
rect 15853 5185 15887 5219
rect 20637 5185 20671 5219
rect 2053 5117 2087 5151
rect 3801 5117 3835 5151
rect 4537 5117 4571 5151
rect 5273 5117 5307 5151
rect 5457 5117 5491 5151
rect 6009 5117 6043 5151
rect 6561 5117 6595 5151
rect 8493 5117 8527 5151
rect 9505 5117 9539 5151
rect 10333 5117 10367 5151
rect 10517 5117 10551 5151
rect 11805 5117 11839 5151
rect 12541 5117 12575 5151
rect 12725 5117 12759 5151
rect 13461 5117 13495 5151
rect 15485 5117 15519 5151
rect 15577 5117 15611 5151
rect 16129 5117 16163 5151
rect 20913 5117 20947 5151
rect 2605 5049 2639 5083
rect 5917 5049 5951 5083
rect 7757 5049 7791 5083
rect 11161 5049 11195 5083
rect 12357 5049 12391 5083
rect 4077 4981 4111 5015
rect 4169 4981 4203 5015
rect 9321 4981 9355 5015
rect 15025 4981 15059 5015
rect 4721 4777 4755 4811
rect 5825 4777 5859 4811
rect 6285 4777 6319 4811
rect 7113 4777 7147 4811
rect 8677 4777 8711 4811
rect 9781 4777 9815 4811
rect 10609 4777 10643 4811
rect 12265 4777 12299 4811
rect 15485 4777 15519 4811
rect 16957 4777 16991 4811
rect 18061 4777 18095 4811
rect 7573 4709 7607 4743
rect 8493 4709 8527 4743
rect 11437 4709 11471 4743
rect 5273 4641 5307 4675
rect 5917 4641 5951 4675
rect 6745 4641 6779 4675
rect 6929 4641 6963 4675
rect 7941 4641 7975 4675
rect 8033 4641 8067 4675
rect 9689 4641 9723 4675
rect 10241 4641 10275 4675
rect 10425 4641 10459 4675
rect 14841 4641 14875 4675
rect 15025 4641 15059 4675
rect 16037 4641 16071 4675
rect 16405 4641 16439 4675
rect 17509 4641 17543 4675
rect 5365 4573 5399 4607
rect 5457 4573 5491 4607
rect 9413 4573 9447 4607
rect 12173 4573 12207 4607
rect 14749 4573 14783 4607
rect 15853 4573 15887 4607
rect 16865 4573 16899 4607
rect 19257 4573 19291 4607
rect 4813 4505 4847 4539
rect 7389 4505 7423 4539
rect 8125 4505 8159 4539
rect 10149 4505 10183 4539
rect 19533 4505 19567 4539
rect 6101 4437 6135 4471
rect 6653 4437 6687 4471
rect 14381 4437 14415 4471
rect 15945 4437 15979 4471
rect 16681 4437 16715 4471
rect 17233 4437 17267 4471
rect 17601 4437 17635 4471
rect 17693 4437 17727 4471
rect 8953 4233 8987 4267
rect 9505 4233 9539 4267
rect 10517 4233 10551 4267
rect 10885 4233 10919 4267
rect 11897 4233 11931 4267
rect 12449 4233 12483 4267
rect 17601 4233 17635 4267
rect 5825 4165 5859 4199
rect 6377 4165 6411 4199
rect 7205 4165 7239 4199
rect 7665 4165 7699 4199
rect 8493 4165 8527 4199
rect 10057 4165 10091 4199
rect 17141 4165 17175 4199
rect 17969 4165 18003 4199
rect 7757 4097 7791 4131
rect 8585 4097 8619 4131
rect 10149 4097 10183 4131
rect 11989 4097 12023 4131
rect 14381 4097 14415 4131
rect 16405 4097 16439 4131
rect 17049 4097 17083 4131
rect 18061 4097 18095 4131
rect 5549 4029 5583 4063
rect 5733 4029 5767 4063
rect 7573 4029 7607 4063
rect 8401 4029 8435 4063
rect 10333 4029 10367 4063
rect 10977 4029 11011 4063
rect 11069 4029 11103 4063
rect 12081 4029 12115 4063
rect 14657 4029 14691 4063
rect 16221 4029 16255 4063
rect 17325 4029 17359 4063
rect 18153 4029 18187 4063
rect 8125 3961 8159 3995
rect 9689 3961 9723 3995
rect 11529 3961 11563 3995
rect 16681 3961 16715 3995
rect 6193 3893 6227 3927
rect 7021 3893 7055 3927
rect 9137 3893 9171 3927
rect 6101 3689 6135 3723
rect 10885 3689 10919 3723
rect 12357 3689 12391 3723
rect 17417 3689 17451 3723
rect 4537 3621 4571 3655
rect 7113 3621 7147 3655
rect 8033 3621 8067 3655
rect 10977 3621 11011 3655
rect 18613 3621 18647 3655
rect 5457 3553 5491 3587
rect 5917 3553 5951 3587
rect 6377 3553 6411 3587
rect 6561 3553 6595 3587
rect 9137 3553 9171 3587
rect 10333 3553 10367 3587
rect 10425 3553 10459 3587
rect 11529 3553 11563 3587
rect 13185 3553 13219 3587
rect 5273 3485 5307 3519
rect 5733 3485 5767 3519
rect 9321 3485 9355 3519
rect 13369 3485 13403 3519
rect 17325 3485 17359 3519
rect 5365 3417 5399 3451
rect 9229 3417 9263 3451
rect 11805 3417 11839 3451
rect 13277 3417 13311 3451
rect 4721 3349 4755 3383
rect 4905 3349 4939 3383
rect 6653 3349 6687 3383
rect 7021 3349 7055 3383
rect 9689 3349 9723 3383
rect 9965 3349 9999 3383
rect 10517 3349 10551 3383
rect 11161 3349 11195 3383
rect 11713 3349 11747 3383
rect 12173 3349 12207 3383
rect 13737 3349 13771 3383
rect 16589 3349 16623 3383
rect 5089 3145 5123 3179
rect 5457 3145 5491 3179
rect 6745 3145 6779 3179
rect 7113 3145 7147 3179
rect 10057 3145 10091 3179
rect 10517 3145 10551 3179
rect 10977 3145 11011 3179
rect 11345 3145 11379 3179
rect 11805 3145 11839 3179
rect 12081 3145 12115 3179
rect 15945 3145 15979 3179
rect 16313 3145 16347 3179
rect 18613 3145 18647 3179
rect 19349 3145 19383 3179
rect 20729 3145 20763 3179
rect 7665 3077 7699 3111
rect 8585 3077 8619 3111
rect 9229 3077 9263 3111
rect 10149 3077 10183 3111
rect 11529 3077 11563 3111
rect 12725 3077 12759 3111
rect 8769 3009 8803 3043
rect 9321 3009 9355 3043
rect 11897 3009 11931 3043
rect 12633 3009 12667 3043
rect 13461 3009 13495 3043
rect 13553 3009 13587 3043
rect 13737 3009 13771 3043
rect 14289 3009 14323 3043
rect 14657 3009 14691 3043
rect 15025 3009 15059 3043
rect 15393 3009 15427 3043
rect 15761 3009 15795 3043
rect 16129 3009 16163 3043
rect 16681 3009 16715 3043
rect 17049 3009 17083 3043
rect 17969 3009 18003 3043
rect 18061 3009 18095 3043
rect 18429 3009 18463 3043
rect 18797 3009 18831 3043
rect 19165 3009 19199 3043
rect 19717 3009 19751 3043
rect 19901 3009 19935 3043
rect 20269 3009 20303 3043
rect 20913 3009 20947 3043
rect 4813 2941 4847 2975
rect 4997 2941 5031 2975
rect 6561 2941 6595 2975
rect 6653 2941 6687 2975
rect 7757 2941 7791 2975
rect 7849 2941 7883 2975
rect 8125 2941 8159 2975
rect 9137 2941 9171 2975
rect 9873 2941 9907 2975
rect 10701 2941 10735 2975
rect 10885 2941 10919 2975
rect 12909 2941 12943 2975
rect 13921 2941 13955 2975
rect 7297 2873 7331 2907
rect 9689 2873 9723 2907
rect 12265 2873 12299 2907
rect 15577 2873 15611 2907
rect 16865 2873 16899 2907
rect 18245 2873 18279 2907
rect 18981 2873 19015 2907
rect 20085 2873 20119 2907
rect 13277 2805 13311 2839
rect 14473 2805 14507 2839
rect 14841 2805 14875 2839
rect 15209 2805 15243 2839
rect 17233 2805 17267 2839
rect 19533 2805 19567 2839
rect 20453 2805 20487 2839
rect 4997 2601 5031 2635
rect 5825 2601 5859 2635
rect 8953 2601 8987 2635
rect 9873 2601 9907 2635
rect 10609 2601 10643 2635
rect 10885 2601 10919 2635
rect 11805 2601 11839 2635
rect 14565 2601 14599 2635
rect 14933 2601 14967 2635
rect 15669 2601 15703 2635
rect 15945 2601 15979 2635
rect 18429 2601 18463 2635
rect 10057 2533 10091 2567
rect 18797 2533 18831 2567
rect 5641 2465 5675 2499
rect 9413 2465 9447 2499
rect 9597 2465 9631 2499
rect 7113 2397 7147 2431
rect 8677 2397 8711 2431
rect 14105 2397 14139 2431
rect 18613 2397 18647 2431
rect 4813 2329 4847 2363
rect 5457 2329 5491 2363
rect 8493 2329 8527 2363
rect 9321 2329 9355 2363
rect 18337 2329 18371 2363
rect 4629 2261 4663 2295
rect 5365 2261 5399 2295
rect 6929 2261 6963 2295
rect 14289 2261 14323 2295
<< metal1 >>
rect 11238 20952 11244 21004
rect 11296 20992 11302 21004
rect 11698 20992 11704 21004
rect 11296 20964 11704 20992
rect 11296 20952 11302 20964
rect 11698 20952 11704 20964
rect 11756 20952 11762 21004
rect 1104 20698 22056 20720
rect 1104 20646 6148 20698
rect 6200 20646 6212 20698
rect 6264 20646 6276 20698
rect 6328 20646 6340 20698
rect 6392 20646 6404 20698
rect 6456 20646 11346 20698
rect 11398 20646 11410 20698
rect 11462 20646 11474 20698
rect 11526 20646 11538 20698
rect 11590 20646 11602 20698
rect 11654 20646 16544 20698
rect 16596 20646 16608 20698
rect 16660 20646 16672 20698
rect 16724 20646 16736 20698
rect 16788 20646 16800 20698
rect 16852 20646 21742 20698
rect 21794 20646 21806 20698
rect 21858 20646 21870 20698
rect 21922 20646 21934 20698
rect 21986 20646 21998 20698
rect 22050 20646 22056 20698
rect 1104 20624 22056 20646
rect 7742 20544 7748 20596
rect 7800 20584 7806 20596
rect 15838 20584 15844 20596
rect 7800 20556 15844 20584
rect 7800 20544 7806 20556
rect 15838 20544 15844 20556
rect 15896 20544 15902 20596
rect 11054 20476 11060 20528
rect 11112 20516 11118 20528
rect 13998 20516 14004 20528
rect 11112 20488 14004 20516
rect 11112 20476 11118 20488
rect 13998 20476 14004 20488
rect 14056 20476 14062 20528
rect 9401 20451 9459 20457
rect 9401 20417 9413 20451
rect 9447 20448 9459 20451
rect 9953 20451 10011 20457
rect 9447 20420 9628 20448
rect 9447 20417 9459 20420
rect 9401 20411 9459 20417
rect 9214 20312 9220 20324
rect 9175 20284 9220 20312
rect 9214 20272 9220 20284
rect 9272 20272 9278 20324
rect 9600 20321 9628 20420
rect 9953 20417 9965 20451
rect 9999 20448 10011 20451
rect 10686 20448 10692 20460
rect 9999 20420 10692 20448
rect 9999 20417 10011 20420
rect 9953 20411 10011 20417
rect 10686 20408 10692 20420
rect 10744 20408 10750 20460
rect 20349 20451 20407 20457
rect 20349 20417 20361 20451
rect 20395 20448 20407 20451
rect 20625 20451 20683 20457
rect 20625 20448 20637 20451
rect 20395 20420 20637 20448
rect 20395 20417 20407 20420
rect 20349 20411 20407 20417
rect 20625 20417 20637 20420
rect 20671 20448 20683 20451
rect 22278 20448 22284 20460
rect 20671 20420 22284 20448
rect 20671 20417 20683 20420
rect 20625 20411 20683 20417
rect 22278 20408 22284 20420
rect 22336 20408 22342 20460
rect 9674 20340 9680 20392
rect 9732 20380 9738 20392
rect 14458 20380 14464 20392
rect 9732 20352 14464 20380
rect 9732 20340 9738 20352
rect 14458 20340 14464 20352
rect 14516 20340 14522 20392
rect 21269 20383 21327 20389
rect 21269 20349 21281 20383
rect 21315 20380 21327 20383
rect 21542 20380 21548 20392
rect 21315 20352 21548 20380
rect 21315 20349 21327 20352
rect 21269 20343 21327 20349
rect 21542 20340 21548 20352
rect 21600 20340 21606 20392
rect 9585 20315 9643 20321
rect 9585 20281 9597 20315
rect 9631 20312 9643 20315
rect 11146 20312 11152 20324
rect 9631 20284 11152 20312
rect 9631 20281 9643 20284
rect 9585 20275 9643 20281
rect 11146 20272 11152 20284
rect 11204 20272 11210 20324
rect 12526 20272 12532 20324
rect 12584 20312 12590 20324
rect 17218 20312 17224 20324
rect 12584 20284 17224 20312
rect 12584 20272 12590 20284
rect 17218 20272 17224 20284
rect 17276 20272 17282 20324
rect 8110 20204 8116 20256
rect 8168 20244 8174 20256
rect 8297 20247 8355 20253
rect 8297 20244 8309 20247
rect 8168 20216 8309 20244
rect 8168 20204 8174 20216
rect 8297 20213 8309 20216
rect 8343 20213 8355 20247
rect 8297 20207 8355 20213
rect 9769 20247 9827 20253
rect 9769 20213 9781 20247
rect 9815 20244 9827 20247
rect 20438 20244 20444 20256
rect 9815 20216 20444 20244
rect 9815 20213 9827 20216
rect 9769 20207 9827 20213
rect 20438 20204 20444 20216
rect 20496 20204 20502 20256
rect 1104 20154 21896 20176
rect 1104 20102 3549 20154
rect 3601 20102 3613 20154
rect 3665 20102 3677 20154
rect 3729 20102 3741 20154
rect 3793 20102 3805 20154
rect 3857 20102 8747 20154
rect 8799 20102 8811 20154
rect 8863 20102 8875 20154
rect 8927 20102 8939 20154
rect 8991 20102 9003 20154
rect 9055 20102 13945 20154
rect 13997 20102 14009 20154
rect 14061 20102 14073 20154
rect 14125 20102 14137 20154
rect 14189 20102 14201 20154
rect 14253 20102 19143 20154
rect 19195 20102 19207 20154
rect 19259 20102 19271 20154
rect 19323 20102 19335 20154
rect 19387 20102 19399 20154
rect 19451 20102 21896 20154
rect 1104 20080 21896 20102
rect 2774 20000 2780 20052
rect 2832 20040 2838 20052
rect 7742 20040 7748 20052
rect 2832 20012 2877 20040
rect 7703 20012 7748 20040
rect 2832 20000 2838 20012
rect 7742 20000 7748 20012
rect 7800 20000 7806 20052
rect 8665 20043 8723 20049
rect 8665 20009 8677 20043
rect 8711 20040 8723 20043
rect 9674 20040 9680 20052
rect 8711 20012 9680 20040
rect 8711 20009 8723 20012
rect 8665 20003 8723 20009
rect 9674 20000 9680 20012
rect 9732 20000 9738 20052
rect 10781 20043 10839 20049
rect 10781 20009 10793 20043
rect 10827 20040 10839 20043
rect 13538 20040 13544 20052
rect 10827 20012 13544 20040
rect 10827 20009 10839 20012
rect 10781 20003 10839 20009
rect 13538 20000 13544 20012
rect 13596 20000 13602 20052
rect 14461 20043 14519 20049
rect 14461 20009 14473 20043
rect 14507 20040 14519 20043
rect 19058 20040 19064 20052
rect 14507 20012 19064 20040
rect 14507 20009 14519 20012
rect 14461 20003 14519 20009
rect 19058 20000 19064 20012
rect 19116 20000 19122 20052
rect 21358 20040 21364 20052
rect 19168 20012 21364 20040
rect 9217 19975 9275 19981
rect 9217 19941 9229 19975
rect 9263 19941 9275 19975
rect 9217 19935 9275 19941
rect 9585 19975 9643 19981
rect 9585 19941 9597 19975
rect 9631 19972 9643 19975
rect 13725 19975 13783 19981
rect 9631 19944 12020 19972
rect 9631 19941 9643 19944
rect 9585 19935 9643 19941
rect 8113 19907 8171 19913
rect 8113 19904 8125 19907
rect 2976 19876 8125 19904
rect 2976 19845 3004 19876
rect 8113 19873 8125 19876
rect 8159 19873 8171 19907
rect 9232 19904 9260 19935
rect 11054 19904 11060 19916
rect 9232 19876 11060 19904
rect 8113 19867 8171 19873
rect 11054 19864 11060 19876
rect 11112 19864 11118 19916
rect 2961 19839 3019 19845
rect 2961 19805 2973 19839
rect 3007 19805 3019 19839
rect 7193 19839 7251 19845
rect 7193 19836 7205 19839
rect 2961 19799 3019 19805
rect 6932 19808 7205 19836
rect 6730 19660 6736 19712
rect 6788 19700 6794 19712
rect 6932 19709 6960 19808
rect 7193 19805 7205 19808
rect 7239 19805 7251 19839
rect 7193 19799 7251 19805
rect 7561 19839 7619 19845
rect 7561 19805 7573 19839
rect 7607 19836 7619 19839
rect 7650 19836 7656 19848
rect 7607 19808 7656 19836
rect 7607 19805 7619 19808
rect 7561 19799 7619 19805
rect 7101 19771 7159 19777
rect 7101 19737 7113 19771
rect 7147 19768 7159 19771
rect 7576 19768 7604 19799
rect 7650 19796 7656 19808
rect 7708 19796 7714 19848
rect 8386 19836 8392 19848
rect 8347 19808 8392 19836
rect 8386 19796 8392 19808
rect 8444 19796 8450 19848
rect 8481 19839 8539 19845
rect 8481 19805 8493 19839
rect 8527 19805 8539 19839
rect 9398 19836 9404 19848
rect 9359 19808 9404 19836
rect 8481 19799 8539 19805
rect 7147 19740 7604 19768
rect 7147 19737 7159 19740
rect 7101 19731 7159 19737
rect 8110 19728 8116 19780
rect 8168 19768 8174 19780
rect 8496 19768 8524 19799
rect 9398 19796 9404 19808
rect 9456 19796 9462 19848
rect 9766 19836 9772 19848
rect 9727 19808 9772 19836
rect 9766 19796 9772 19808
rect 9824 19796 9830 19848
rect 9861 19839 9919 19845
rect 9861 19805 9873 19839
rect 9907 19836 9919 19839
rect 9950 19836 9956 19848
rect 9907 19808 9956 19836
rect 9907 19805 9919 19808
rect 9861 19799 9919 19805
rect 8168 19740 8524 19768
rect 9033 19771 9091 19777
rect 8168 19728 8174 19740
rect 9033 19737 9045 19771
rect 9079 19768 9091 19771
rect 9876 19768 9904 19799
rect 9950 19796 9956 19808
rect 10008 19796 10014 19848
rect 10042 19796 10048 19848
rect 10100 19836 10106 19848
rect 10229 19839 10287 19845
rect 10229 19836 10241 19839
rect 10100 19808 10241 19836
rect 10100 19796 10106 19808
rect 10229 19805 10241 19808
rect 10275 19805 10287 19839
rect 10594 19836 10600 19848
rect 10555 19808 10600 19836
rect 10229 19799 10287 19805
rect 10594 19796 10600 19808
rect 10652 19796 10658 19848
rect 11992 19836 12020 19944
rect 13725 19941 13737 19975
rect 13771 19972 13783 19975
rect 19168 19972 19196 20012
rect 21358 20000 21364 20012
rect 21416 20000 21422 20052
rect 13771 19944 19196 19972
rect 13771 19941 13783 19944
rect 13725 19935 13783 19941
rect 21542 19904 21548 19916
rect 21503 19876 21548 19904
rect 21542 19864 21548 19876
rect 21600 19864 21606 19916
rect 12894 19836 12900 19848
rect 11992 19808 12900 19836
rect 12894 19796 12900 19808
rect 12952 19796 12958 19848
rect 12989 19839 13047 19845
rect 12989 19805 13001 19839
rect 13035 19836 13047 19839
rect 13078 19836 13084 19848
rect 13035 19808 13084 19836
rect 13035 19805 13047 19808
rect 12989 19799 13047 19805
rect 13078 19796 13084 19808
rect 13136 19796 13142 19848
rect 13541 19839 13599 19845
rect 13541 19805 13553 19839
rect 13587 19836 13599 19839
rect 13630 19836 13636 19848
rect 13587 19808 13636 19836
rect 13587 19805 13599 19808
rect 13541 19799 13599 19805
rect 13630 19796 13636 19808
rect 13688 19836 13694 19848
rect 14093 19839 14151 19845
rect 14093 19836 14105 19839
rect 13688 19808 14105 19836
rect 13688 19796 13694 19808
rect 14093 19805 14105 19808
rect 14139 19805 14151 19839
rect 14093 19799 14151 19805
rect 14277 19839 14335 19845
rect 14277 19805 14289 19839
rect 14323 19836 14335 19839
rect 14645 19839 14703 19845
rect 14645 19836 14657 19839
rect 14323 19808 14657 19836
rect 14323 19805 14335 19808
rect 14277 19799 14335 19805
rect 14645 19805 14657 19808
rect 14691 19836 14703 19839
rect 14826 19836 14832 19848
rect 14691 19808 14832 19836
rect 14691 19805 14703 19808
rect 14645 19799 14703 19805
rect 14826 19796 14832 19808
rect 14884 19796 14890 19848
rect 16301 19839 16359 19845
rect 16301 19805 16313 19839
rect 16347 19805 16359 19839
rect 16301 19799 16359 19805
rect 9079 19740 9904 19768
rect 9079 19737 9091 19740
rect 9033 19731 9091 19737
rect 12434 19728 12440 19780
rect 12492 19768 12498 19780
rect 12722 19771 12780 19777
rect 12722 19768 12734 19771
rect 12492 19740 12734 19768
rect 12492 19728 12498 19740
rect 12722 19737 12734 19740
rect 12768 19737 12780 19771
rect 14366 19768 14372 19780
rect 12722 19731 12780 19737
rect 12912 19740 14372 19768
rect 6917 19703 6975 19709
rect 6917 19700 6929 19703
rect 6788 19672 6929 19700
rect 6788 19660 6794 19672
rect 6917 19669 6929 19672
rect 6963 19669 6975 19703
rect 7374 19700 7380 19712
rect 7335 19672 7380 19700
rect 6917 19663 6975 19669
rect 7374 19660 7380 19672
rect 7432 19660 7438 19712
rect 10045 19703 10103 19709
rect 10045 19669 10057 19703
rect 10091 19700 10103 19703
rect 10134 19700 10140 19712
rect 10091 19672 10140 19700
rect 10091 19669 10103 19672
rect 10045 19663 10103 19669
rect 10134 19660 10140 19672
rect 10192 19660 10198 19712
rect 10410 19700 10416 19712
rect 10371 19672 10416 19700
rect 10410 19660 10416 19672
rect 10468 19660 10474 19712
rect 11054 19660 11060 19712
rect 11112 19700 11118 19712
rect 11609 19703 11667 19709
rect 11609 19700 11621 19703
rect 11112 19672 11621 19700
rect 11112 19660 11118 19672
rect 11609 19669 11621 19672
rect 11655 19669 11667 19703
rect 11609 19663 11667 19669
rect 11882 19660 11888 19712
rect 11940 19700 11946 19712
rect 12912 19700 12940 19740
rect 14366 19728 14372 19740
rect 14424 19728 14430 19780
rect 14458 19728 14464 19780
rect 14516 19768 14522 19780
rect 16117 19771 16175 19777
rect 16117 19768 16129 19771
rect 14516 19740 16129 19768
rect 14516 19728 14522 19740
rect 16117 19737 16129 19740
rect 16163 19768 16175 19771
rect 16316 19768 16344 19799
rect 16163 19740 16344 19768
rect 16163 19737 16175 19740
rect 16117 19731 16175 19737
rect 21082 19728 21088 19780
rect 21140 19768 21146 19780
rect 21278 19771 21336 19777
rect 21278 19768 21290 19771
rect 21140 19740 21290 19768
rect 21140 19728 21146 19740
rect 21278 19737 21290 19740
rect 21324 19737 21336 19771
rect 21278 19731 21336 19737
rect 13078 19700 13084 19712
rect 11940 19672 12940 19700
rect 13039 19672 13084 19700
rect 11940 19660 11946 19672
rect 13078 19660 13084 19672
rect 13136 19700 13142 19712
rect 13265 19703 13323 19709
rect 13265 19700 13277 19703
rect 13136 19672 13277 19700
rect 13136 19660 13142 19672
rect 13265 19669 13277 19672
rect 13311 19669 13323 19703
rect 13265 19663 13323 19669
rect 16485 19703 16543 19709
rect 16485 19669 16497 19703
rect 16531 19700 16543 19703
rect 16942 19700 16948 19712
rect 16531 19672 16948 19700
rect 16531 19669 16543 19672
rect 16485 19663 16543 19669
rect 16942 19660 16948 19672
rect 17000 19660 17006 19712
rect 20162 19700 20168 19712
rect 20123 19672 20168 19700
rect 20162 19660 20168 19672
rect 20220 19660 20226 19712
rect 1104 19610 22056 19632
rect 1104 19558 6148 19610
rect 6200 19558 6212 19610
rect 6264 19558 6276 19610
rect 6328 19558 6340 19610
rect 6392 19558 6404 19610
rect 6456 19558 11346 19610
rect 11398 19558 11410 19610
rect 11462 19558 11474 19610
rect 11526 19558 11538 19610
rect 11590 19558 11602 19610
rect 11654 19558 16544 19610
rect 16596 19558 16608 19610
rect 16660 19558 16672 19610
rect 16724 19558 16736 19610
rect 16788 19558 16800 19610
rect 16852 19558 21742 19610
rect 21794 19558 21806 19610
rect 21858 19558 21870 19610
rect 21922 19558 21934 19610
rect 21986 19558 21998 19610
rect 22050 19558 22056 19610
rect 1104 19536 22056 19558
rect 8294 19496 8300 19508
rect 8255 19468 8300 19496
rect 8294 19456 8300 19468
rect 8352 19456 8358 19508
rect 9401 19499 9459 19505
rect 9401 19465 9413 19499
rect 9447 19465 9459 19499
rect 9401 19459 9459 19465
rect 9861 19499 9919 19505
rect 9861 19465 9873 19499
rect 9907 19465 9919 19499
rect 9861 19459 9919 19465
rect 11517 19499 11575 19505
rect 11517 19465 11529 19499
rect 11563 19496 11575 19499
rect 11882 19496 11888 19508
rect 11563 19468 11888 19496
rect 11563 19465 11575 19468
rect 11517 19459 11575 19465
rect 9416 19428 9444 19459
rect 9876 19428 9904 19459
rect 11882 19456 11888 19468
rect 11940 19456 11946 19508
rect 12434 19456 12440 19508
rect 12492 19496 12498 19508
rect 12989 19499 13047 19505
rect 12989 19496 13001 19499
rect 12492 19468 13001 19496
rect 12492 19456 12498 19468
rect 12989 19465 13001 19468
rect 13035 19465 13047 19499
rect 12989 19459 13047 19465
rect 19337 19499 19395 19505
rect 19337 19465 19349 19499
rect 19383 19496 19395 19499
rect 19610 19496 19616 19508
rect 19383 19468 19616 19496
rect 19383 19465 19395 19468
rect 19337 19459 19395 19465
rect 19610 19456 19616 19468
rect 19668 19456 19674 19508
rect 20901 19499 20959 19505
rect 20901 19465 20913 19499
rect 20947 19496 20959 19499
rect 21542 19496 21548 19508
rect 20947 19468 21548 19496
rect 20947 19465 20959 19468
rect 20901 19459 20959 19465
rect 12526 19428 12532 19440
rect 9416 19400 9812 19428
rect 9876 19400 12532 19428
rect 8113 19363 8171 19369
rect 8113 19329 8125 19363
rect 8159 19360 8171 19363
rect 8159 19332 8294 19360
rect 8159 19329 8171 19332
rect 8113 19323 8171 19329
rect 8266 19292 8294 19332
rect 8662 19320 8668 19372
rect 8720 19360 8726 19372
rect 8757 19363 8815 19369
rect 8757 19360 8769 19363
rect 8720 19332 8769 19360
rect 8720 19320 8726 19332
rect 8757 19329 8769 19332
rect 8803 19329 8815 19363
rect 8757 19323 8815 19329
rect 9217 19363 9275 19369
rect 9217 19329 9229 19363
rect 9263 19329 9275 19363
rect 9217 19323 9275 19329
rect 9677 19363 9735 19369
rect 9677 19329 9689 19363
rect 9723 19329 9735 19363
rect 9677 19323 9735 19329
rect 8941 19295 8999 19301
rect 8941 19292 8953 19295
rect 8266 19264 8953 19292
rect 8941 19261 8953 19264
rect 8987 19292 8999 19295
rect 9122 19292 9128 19304
rect 8987 19264 9128 19292
rect 8987 19261 8999 19264
rect 8941 19255 8999 19261
rect 9122 19252 9128 19264
rect 9180 19252 9186 19304
rect 8570 19156 8576 19168
rect 8531 19128 8576 19156
rect 8570 19116 8576 19128
rect 8628 19116 8634 19168
rect 9125 19159 9183 19165
rect 9125 19125 9137 19159
rect 9171 19156 9183 19159
rect 9232 19156 9260 19323
rect 9692 19224 9720 19323
rect 9784 19292 9812 19400
rect 12526 19388 12532 19400
rect 12584 19388 12590 19440
rect 12630 19431 12688 19437
rect 12630 19397 12642 19431
rect 12676 19428 12688 19431
rect 12802 19428 12808 19440
rect 12676 19400 12808 19428
rect 12676 19397 12688 19400
rect 12630 19391 12688 19397
rect 12802 19388 12808 19400
rect 12860 19388 12866 19440
rect 14461 19431 14519 19437
rect 14461 19428 14473 19431
rect 13740 19400 14473 19428
rect 10042 19360 10048 19372
rect 10003 19332 10048 19360
rect 10042 19320 10048 19332
rect 10100 19320 10106 19372
rect 12897 19363 12955 19369
rect 11900 19332 12839 19360
rect 11900 19292 11928 19332
rect 9784 19264 11928 19292
rect 12811 19292 12839 19332
rect 12897 19329 12909 19363
rect 12943 19360 12955 19363
rect 13078 19360 13084 19372
rect 12943 19332 13084 19360
rect 12943 19329 12955 19332
rect 12897 19323 12955 19329
rect 13078 19320 13084 19332
rect 13136 19360 13142 19372
rect 13740 19360 13768 19400
rect 13136 19332 13768 19360
rect 13136 19320 13142 19332
rect 13814 19320 13820 19372
rect 13872 19360 13878 19372
rect 14102 19363 14160 19369
rect 14102 19360 14114 19363
rect 13872 19332 14114 19360
rect 13872 19320 13878 19332
rect 14102 19329 14114 19332
rect 14148 19329 14160 19363
rect 14102 19323 14160 19329
rect 14384 19301 14412 19400
rect 14461 19397 14473 19400
rect 14507 19397 14519 19431
rect 14461 19391 14519 19397
rect 20461 19363 20519 19369
rect 20461 19329 20473 19363
rect 20507 19360 20519 19363
rect 20717 19363 20775 19369
rect 20507 19332 20668 19360
rect 20507 19329 20519 19332
rect 20461 19323 20519 19329
rect 14369 19295 14427 19301
rect 12811 19264 13216 19292
rect 9692 19196 9812 19224
rect 9490 19156 9496 19168
rect 9171 19128 9496 19156
rect 9171 19125 9183 19128
rect 9125 19119 9183 19125
rect 9490 19116 9496 19128
rect 9548 19116 9554 19168
rect 9784 19156 9812 19196
rect 10134 19184 10140 19236
rect 10192 19224 10198 19236
rect 10192 19196 11652 19224
rect 10192 19184 10198 19196
rect 10321 19159 10379 19165
rect 10321 19156 10333 19159
rect 9784 19128 10333 19156
rect 10321 19125 10333 19128
rect 10367 19156 10379 19159
rect 10870 19156 10876 19168
rect 10367 19128 10876 19156
rect 10367 19125 10379 19128
rect 10321 19119 10379 19125
rect 10870 19116 10876 19128
rect 10928 19116 10934 19168
rect 11624 19156 11652 19196
rect 12894 19156 12900 19168
rect 11624 19128 12900 19156
rect 12894 19116 12900 19128
rect 12952 19116 12958 19168
rect 13188 19156 13216 19264
rect 14369 19261 14381 19295
rect 14415 19261 14427 19295
rect 14369 19255 14427 19261
rect 14642 19252 14648 19304
rect 14700 19292 14706 19304
rect 17034 19292 17040 19304
rect 14700 19264 17040 19292
rect 14700 19252 14706 19264
rect 17034 19252 17040 19264
rect 17092 19252 17098 19304
rect 20640 19292 20668 19332
rect 20717 19329 20729 19363
rect 20763 19360 20775 19363
rect 20916 19360 20944 19459
rect 21542 19456 21548 19468
rect 21600 19456 21606 19508
rect 20990 19360 20996 19372
rect 20763 19332 20996 19360
rect 20763 19329 20775 19332
rect 20717 19323 20775 19329
rect 20990 19320 20996 19332
rect 21048 19320 21054 19372
rect 20898 19292 20904 19304
rect 20640 19264 20904 19292
rect 20898 19252 20904 19264
rect 20956 19252 20962 19304
rect 16298 19224 16304 19236
rect 14384 19196 16304 19224
rect 14384 19156 14412 19196
rect 16298 19184 16304 19196
rect 16356 19184 16362 19236
rect 16942 19184 16948 19236
rect 17000 19224 17006 19236
rect 17000 19196 19472 19224
rect 17000 19184 17006 19196
rect 13188 19128 14412 19156
rect 14734 19116 14740 19168
rect 14792 19156 14798 19168
rect 18138 19156 18144 19168
rect 14792 19128 18144 19156
rect 14792 19116 14798 19128
rect 18138 19116 18144 19128
rect 18196 19116 18202 19168
rect 19444 19156 19472 19196
rect 21634 19156 21640 19168
rect 19444 19128 21640 19156
rect 21634 19116 21640 19128
rect 21692 19116 21698 19168
rect 1104 19066 21896 19088
rect 1104 19014 3549 19066
rect 3601 19014 3613 19066
rect 3665 19014 3677 19066
rect 3729 19014 3741 19066
rect 3793 19014 3805 19066
rect 3857 19014 8747 19066
rect 8799 19014 8811 19066
rect 8863 19014 8875 19066
rect 8927 19014 8939 19066
rect 8991 19014 9003 19066
rect 9055 19014 13945 19066
rect 13997 19014 14009 19066
rect 14061 19014 14073 19066
rect 14125 19014 14137 19066
rect 14189 19014 14201 19066
rect 14253 19014 19143 19066
rect 19195 19014 19207 19066
rect 19259 19014 19271 19066
rect 19323 19014 19335 19066
rect 19387 19014 19399 19066
rect 19451 19014 21896 19066
rect 1104 18992 21896 19014
rect 8938 18912 8944 18964
rect 8996 18952 9002 18964
rect 9950 18952 9956 18964
rect 8996 18924 9956 18952
rect 8996 18912 9002 18924
rect 9950 18912 9956 18924
rect 10008 18912 10014 18964
rect 10410 18912 10416 18964
rect 10468 18952 10474 18964
rect 10468 18924 12848 18952
rect 10468 18912 10474 18924
rect 9858 18844 9864 18896
rect 9916 18884 9922 18896
rect 10042 18884 10048 18896
rect 9916 18856 10048 18884
rect 9916 18844 9922 18856
rect 10042 18844 10048 18856
rect 10100 18844 10106 18896
rect 12820 18884 12848 18924
rect 12894 18912 12900 18964
rect 12952 18952 12958 18964
rect 17494 18952 17500 18964
rect 12952 18924 17500 18952
rect 12952 18912 12958 18924
rect 17494 18912 17500 18924
rect 17552 18912 17558 18964
rect 20990 18952 20996 18964
rect 20951 18924 20996 18952
rect 20990 18912 20996 18924
rect 21048 18912 21054 18964
rect 14734 18884 14740 18896
rect 12820 18856 14740 18884
rect 14734 18844 14740 18856
rect 14792 18844 14798 18896
rect 8941 18819 8999 18825
rect 8941 18816 8953 18819
rect 8588 18788 8953 18816
rect 8588 18760 8616 18788
rect 8941 18785 8953 18788
rect 8987 18785 8999 18819
rect 9398 18816 9404 18828
rect 9359 18788 9404 18816
rect 8941 18779 8999 18785
rect 9398 18776 9404 18788
rect 9456 18776 9462 18828
rect 9766 18776 9772 18828
rect 9824 18816 9830 18828
rect 10502 18816 10508 18828
rect 9824 18788 10508 18816
rect 9824 18776 9830 18788
rect 10502 18776 10508 18788
rect 10560 18776 10566 18828
rect 13354 18776 13360 18828
rect 13412 18816 13418 18828
rect 13541 18819 13599 18825
rect 13541 18816 13553 18819
rect 13412 18788 13553 18816
rect 13412 18776 13418 18788
rect 13541 18785 13553 18788
rect 13587 18785 13599 18819
rect 13541 18779 13599 18785
rect 14182 18776 14188 18828
rect 14240 18816 14246 18828
rect 14550 18816 14556 18828
rect 14240 18788 14556 18816
rect 14240 18776 14246 18788
rect 14550 18776 14556 18788
rect 14608 18776 14614 18828
rect 20901 18819 20959 18825
rect 20901 18785 20913 18819
rect 20947 18816 20959 18819
rect 21008 18816 21036 18912
rect 20947 18788 21036 18816
rect 20947 18785 20959 18788
rect 20901 18779 20959 18785
rect 8113 18751 8171 18757
rect 8113 18717 8125 18751
rect 8159 18748 8171 18751
rect 8570 18748 8576 18760
rect 8159 18720 8576 18748
rect 8159 18717 8171 18720
rect 8113 18711 8171 18717
rect 8570 18708 8576 18720
rect 8628 18708 8634 18760
rect 8757 18751 8815 18757
rect 8757 18717 8769 18751
rect 8803 18748 8815 18751
rect 9122 18748 9128 18760
rect 8803 18720 9128 18748
rect 8803 18717 8815 18720
rect 8757 18711 8815 18717
rect 9122 18708 9128 18720
rect 9180 18708 9186 18760
rect 9214 18708 9220 18760
rect 9272 18748 9278 18760
rect 10045 18751 10103 18757
rect 9272 18720 9317 18748
rect 9272 18708 9278 18720
rect 10045 18717 10057 18751
rect 10091 18748 10103 18751
rect 10962 18748 10968 18760
rect 10091 18720 10968 18748
rect 10091 18717 10103 18720
rect 10045 18711 10103 18717
rect 10962 18708 10968 18720
rect 11020 18708 11026 18760
rect 11054 18708 11060 18760
rect 11112 18748 11118 18760
rect 11526 18751 11584 18757
rect 11526 18748 11538 18751
rect 11112 18720 11538 18748
rect 11112 18708 11118 18720
rect 11526 18717 11538 18720
rect 11572 18717 11584 18751
rect 11526 18711 11584 18717
rect 11793 18751 11851 18757
rect 11793 18717 11805 18751
rect 11839 18748 11851 18751
rect 11885 18751 11943 18757
rect 11885 18748 11897 18751
rect 11839 18720 11897 18748
rect 11839 18717 11851 18720
rect 11793 18711 11851 18717
rect 11885 18717 11897 18720
rect 11931 18748 11943 18751
rect 13170 18748 13176 18760
rect 11931 18720 13176 18748
rect 11931 18717 11943 18720
rect 11885 18711 11943 18717
rect 13170 18708 13176 18720
rect 13228 18748 13234 18760
rect 13449 18751 13507 18757
rect 13449 18748 13461 18751
rect 13228 18720 13461 18748
rect 13228 18708 13234 18720
rect 13449 18717 13461 18720
rect 13495 18748 13507 18751
rect 13722 18748 13728 18760
rect 13495 18720 13728 18748
rect 13495 18717 13507 18720
rect 13449 18711 13507 18717
rect 13722 18708 13728 18720
rect 13780 18748 13786 18760
rect 13817 18751 13875 18757
rect 13817 18748 13829 18751
rect 13780 18720 13829 18748
rect 13780 18708 13786 18720
rect 13817 18717 13829 18720
rect 13863 18748 13875 18751
rect 14642 18748 14648 18760
rect 13863 18720 14648 18748
rect 13863 18717 13875 18720
rect 13817 18711 13875 18717
rect 14642 18708 14648 18720
rect 14700 18748 14706 18760
rect 14737 18751 14795 18757
rect 14737 18748 14749 18751
rect 14700 18720 14749 18748
rect 14700 18708 14706 18720
rect 14737 18717 14749 18720
rect 14783 18748 14795 18751
rect 16301 18751 16359 18757
rect 16301 18748 16313 18751
rect 14783 18720 16313 18748
rect 14783 18717 14795 18720
rect 14737 18711 14795 18717
rect 16301 18717 16313 18720
rect 16347 18748 16359 18751
rect 16390 18748 16396 18760
rect 16347 18720 16396 18748
rect 16347 18717 16359 18720
rect 16301 18711 16359 18717
rect 16390 18708 16396 18720
rect 16448 18748 16454 18760
rect 16669 18751 16727 18757
rect 16669 18748 16681 18751
rect 16448 18720 16681 18748
rect 16448 18708 16454 18720
rect 16669 18717 16681 18720
rect 16715 18748 16727 18751
rect 18141 18751 18199 18757
rect 18141 18748 18153 18751
rect 16715 18720 18153 18748
rect 16715 18717 16727 18720
rect 16669 18711 16727 18717
rect 18141 18717 18153 18720
rect 18187 18748 18199 18751
rect 18187 18720 18276 18748
rect 18187 18717 18199 18720
rect 18141 18711 18199 18717
rect 10134 18680 10140 18692
rect 8588 18652 10140 18680
rect 198 18572 204 18624
rect 256 18612 262 18624
rect 4614 18612 4620 18624
rect 256 18584 4620 18612
rect 256 18572 262 18584
rect 4614 18572 4620 18584
rect 4672 18572 4678 18624
rect 8294 18612 8300 18624
rect 8255 18584 8300 18612
rect 8294 18572 8300 18584
rect 8352 18572 8358 18624
rect 8588 18621 8616 18652
rect 10134 18640 10140 18652
rect 10192 18640 10198 18692
rect 10244 18652 11376 18680
rect 10244 18621 10272 18652
rect 8573 18615 8631 18621
rect 8573 18581 8585 18615
rect 8619 18581 8631 18615
rect 8573 18575 8631 18581
rect 10229 18615 10287 18621
rect 10229 18581 10241 18615
rect 10275 18581 10287 18615
rect 10410 18612 10416 18624
rect 10371 18584 10416 18612
rect 10229 18575 10287 18581
rect 10410 18572 10416 18584
rect 10468 18572 10474 18624
rect 11348 18612 11376 18652
rect 11974 18640 11980 18692
rect 12032 18680 12038 18692
rect 12130 18683 12188 18689
rect 12130 18680 12142 18683
rect 12032 18652 12142 18680
rect 12032 18640 12038 18652
rect 12130 18649 12142 18652
rect 12176 18649 12188 18683
rect 14274 18680 14280 18692
rect 12130 18643 12188 18649
rect 12406 18652 14280 18680
rect 12406 18612 12434 18652
rect 14274 18640 14280 18652
rect 14332 18640 14338 18692
rect 14366 18640 14372 18692
rect 14424 18680 14430 18692
rect 14982 18683 15040 18689
rect 14982 18680 14994 18683
rect 14424 18652 14994 18680
rect 14424 18640 14430 18652
rect 14982 18649 14994 18652
rect 15028 18649 15040 18683
rect 14982 18643 15040 18649
rect 17862 18640 17868 18692
rect 17920 18689 17926 18692
rect 17920 18680 17932 18689
rect 17920 18652 17965 18680
rect 17920 18643 17932 18652
rect 17920 18640 17926 18643
rect 18248 18624 18276 18720
rect 19702 18708 19708 18760
rect 19760 18748 19766 18760
rect 22738 18748 22744 18760
rect 19760 18720 22744 18748
rect 19760 18708 19766 18720
rect 22738 18708 22744 18720
rect 22796 18708 22802 18760
rect 20346 18640 20352 18692
rect 20404 18680 20410 18692
rect 20634 18683 20692 18689
rect 20634 18680 20646 18683
rect 20404 18652 20646 18680
rect 20404 18640 20410 18652
rect 20634 18649 20646 18652
rect 20680 18649 20692 18683
rect 20634 18643 20692 18649
rect 11348 18584 12434 18612
rect 12526 18572 12532 18624
rect 12584 18612 12590 18624
rect 13265 18615 13323 18621
rect 13265 18612 13277 18615
rect 12584 18584 13277 18612
rect 12584 18572 12590 18584
rect 13265 18581 13277 18584
rect 13311 18612 13323 18615
rect 13538 18612 13544 18624
rect 13311 18584 13544 18612
rect 13311 18581 13323 18584
rect 13265 18575 13323 18581
rect 13538 18572 13544 18584
rect 13596 18572 13602 18624
rect 16114 18612 16120 18624
rect 16075 18584 16120 18612
rect 16114 18572 16120 18584
rect 16172 18572 16178 18624
rect 16761 18615 16819 18621
rect 16761 18581 16773 18615
rect 16807 18612 16819 18615
rect 16942 18612 16948 18624
rect 16807 18584 16948 18612
rect 16807 18581 16819 18584
rect 16761 18575 16819 18581
rect 16942 18572 16948 18584
rect 17000 18572 17006 18624
rect 18230 18612 18236 18624
rect 18191 18584 18236 18612
rect 18230 18572 18236 18584
rect 18288 18572 18294 18624
rect 19521 18615 19579 18621
rect 19521 18581 19533 18615
rect 19567 18612 19579 18615
rect 19886 18612 19892 18624
rect 19567 18584 19892 18612
rect 19567 18581 19579 18584
rect 19521 18575 19579 18581
rect 19886 18572 19892 18584
rect 19944 18572 19950 18624
rect 1104 18522 22056 18544
rect 1104 18470 6148 18522
rect 6200 18470 6212 18522
rect 6264 18470 6276 18522
rect 6328 18470 6340 18522
rect 6392 18470 6404 18522
rect 6456 18470 11346 18522
rect 11398 18470 11410 18522
rect 11462 18470 11474 18522
rect 11526 18470 11538 18522
rect 11590 18470 11602 18522
rect 11654 18470 16544 18522
rect 16596 18470 16608 18522
rect 16660 18470 16672 18522
rect 16724 18470 16736 18522
rect 16788 18470 16800 18522
rect 16852 18470 21742 18522
rect 21794 18470 21806 18522
rect 21858 18470 21870 18522
rect 21922 18470 21934 18522
rect 21986 18470 21998 18522
rect 22050 18470 22056 18522
rect 1104 18448 22056 18470
rect 2133 18411 2191 18417
rect 2133 18377 2145 18411
rect 2179 18408 2191 18411
rect 2866 18408 2872 18420
rect 2179 18380 2872 18408
rect 2179 18377 2191 18380
rect 2133 18371 2191 18377
rect 2866 18368 2872 18380
rect 2924 18368 2930 18420
rect 4338 18368 4344 18420
rect 4396 18408 4402 18420
rect 8021 18411 8079 18417
rect 8021 18408 8033 18411
rect 4396 18380 8033 18408
rect 4396 18368 4402 18380
rect 8021 18377 8033 18380
rect 8067 18408 8079 18411
rect 8665 18411 8723 18417
rect 8665 18408 8677 18411
rect 8067 18380 8677 18408
rect 8067 18377 8079 18380
rect 8021 18371 8079 18377
rect 8665 18377 8677 18380
rect 8711 18377 8723 18411
rect 8665 18371 8723 18377
rect 9030 18368 9036 18420
rect 9088 18408 9094 18420
rect 9088 18380 10088 18408
rect 9088 18368 9094 18380
rect 2498 18300 2504 18352
rect 2556 18340 2562 18352
rect 4430 18340 4436 18352
rect 2556 18312 4436 18340
rect 2556 18300 2562 18312
rect 4430 18300 4436 18312
rect 4488 18340 4494 18352
rect 4801 18343 4859 18349
rect 4801 18340 4813 18343
rect 4488 18312 4813 18340
rect 4488 18300 4494 18312
rect 4801 18309 4813 18312
rect 4847 18340 4859 18343
rect 5537 18343 5595 18349
rect 5537 18340 5549 18343
rect 4847 18312 5549 18340
rect 4847 18309 4859 18312
rect 4801 18303 4859 18309
rect 5537 18309 5549 18312
rect 5583 18309 5595 18343
rect 5537 18303 5595 18309
rect 2317 18275 2375 18281
rect 2317 18241 2329 18275
rect 2363 18272 2375 18275
rect 3142 18272 3148 18284
rect 2363 18244 3148 18272
rect 2363 18241 2375 18244
rect 2317 18235 2375 18241
rect 3142 18232 3148 18244
rect 3200 18232 3206 18284
rect 3878 18232 3884 18284
rect 3936 18272 3942 18284
rect 5074 18272 5080 18284
rect 3936 18244 5080 18272
rect 3936 18232 3942 18244
rect 5074 18232 5080 18244
rect 5132 18232 5138 18284
rect 8018 18232 8024 18284
rect 8076 18272 8082 18284
rect 8573 18275 8631 18281
rect 8573 18272 8585 18275
rect 8076 18244 8585 18272
rect 8076 18232 8082 18244
rect 8573 18241 8585 18244
rect 8619 18241 8631 18275
rect 9030 18272 9036 18284
rect 8573 18235 8631 18241
rect 8680 18244 9036 18272
rect 2038 18164 2044 18216
rect 2096 18204 2102 18216
rect 4338 18204 4344 18216
rect 2096 18176 4344 18204
rect 2096 18164 2102 18176
rect 4338 18164 4344 18176
rect 4396 18204 4402 18216
rect 4985 18207 5043 18213
rect 4985 18204 4997 18207
rect 4396 18176 4997 18204
rect 4396 18164 4402 18176
rect 4985 18173 4997 18176
rect 5031 18204 5043 18207
rect 5629 18207 5687 18213
rect 5629 18204 5641 18207
rect 5031 18176 5641 18204
rect 5031 18173 5043 18176
rect 4985 18167 5043 18173
rect 5629 18173 5641 18176
rect 5675 18173 5687 18207
rect 5629 18167 5687 18173
rect 5813 18207 5871 18213
rect 5813 18173 5825 18207
rect 5859 18204 5871 18207
rect 6086 18204 6092 18216
rect 5859 18176 6092 18204
rect 5859 18173 5871 18176
rect 5813 18167 5871 18173
rect 6086 18164 6092 18176
rect 6144 18204 6150 18216
rect 8680 18204 8708 18244
rect 9030 18232 9036 18244
rect 9088 18232 9094 18284
rect 9628 18232 9634 18284
rect 9686 18281 9692 18284
rect 9686 18275 9704 18281
rect 9692 18241 9704 18275
rect 9686 18235 9704 18241
rect 9769 18275 9827 18281
rect 9769 18241 9781 18275
rect 9815 18272 9827 18275
rect 10060 18272 10088 18380
rect 10134 18368 10140 18420
rect 10192 18408 10198 18420
rect 14182 18408 14188 18420
rect 10192 18380 14188 18408
rect 10192 18368 10198 18380
rect 14182 18368 14188 18380
rect 14240 18368 14246 18420
rect 14642 18408 14648 18420
rect 14476 18380 14648 18408
rect 10226 18300 10232 18352
rect 10284 18340 10290 18352
rect 10410 18340 10416 18352
rect 10284 18312 10416 18340
rect 10284 18300 10290 18312
rect 10410 18300 10416 18312
rect 10468 18300 10474 18352
rect 13354 18340 13360 18352
rect 12645 18312 13360 18340
rect 12645 18281 12673 18312
rect 13354 18300 13360 18312
rect 13412 18340 13418 18352
rect 14366 18340 14372 18352
rect 13412 18312 14372 18340
rect 13412 18300 13418 18312
rect 14366 18300 14372 18312
rect 14424 18300 14430 18352
rect 12630 18275 12688 18281
rect 12630 18272 12642 18275
rect 9815 18244 9904 18272
rect 10060 18244 12642 18272
rect 9815 18241 9827 18244
rect 9769 18235 9827 18241
rect 9686 18232 9692 18235
rect 8846 18204 8852 18216
rect 6144 18176 8708 18204
rect 8807 18176 8852 18204
rect 6144 18164 6150 18176
rect 8846 18164 8852 18176
rect 8904 18164 8910 18216
rect 9398 18204 9404 18216
rect 9359 18176 9404 18204
rect 9398 18164 9404 18176
rect 9456 18164 9462 18216
rect 9876 18204 9904 18244
rect 12630 18241 12642 18244
rect 12676 18241 12688 18275
rect 12630 18235 12688 18241
rect 12897 18275 12955 18281
rect 12897 18241 12909 18275
rect 12943 18272 12955 18275
rect 13722 18272 13728 18284
rect 12943 18244 13728 18272
rect 12943 18241 12955 18244
rect 12897 18235 12955 18241
rect 13722 18232 13728 18244
rect 13780 18232 13786 18284
rect 14182 18232 14188 18284
rect 14240 18281 14246 18284
rect 14476 18281 14504 18380
rect 14642 18368 14648 18380
rect 14700 18368 14706 18420
rect 15105 18411 15163 18417
rect 15105 18377 15117 18411
rect 15151 18377 15163 18411
rect 16669 18411 16727 18417
rect 16669 18408 16681 18411
rect 15105 18371 15163 18377
rect 16316 18380 16681 18408
rect 15120 18340 15148 18371
rect 14568 18312 15148 18340
rect 14240 18272 14252 18281
rect 14461 18275 14519 18281
rect 14240 18244 14412 18272
rect 14240 18235 14252 18244
rect 14240 18232 14246 18235
rect 9508 18176 9904 18204
rect 10045 18207 10103 18213
rect 1578 18096 1584 18148
rect 1636 18136 1642 18148
rect 4154 18136 4160 18148
rect 1636 18108 4160 18136
rect 1636 18096 1642 18108
rect 4154 18096 4160 18108
rect 4212 18096 4218 18148
rect 4798 18096 4804 18148
rect 4856 18136 4862 18148
rect 6822 18136 6828 18148
rect 4856 18108 6828 18136
rect 4856 18096 4862 18108
rect 6822 18096 6828 18108
rect 6880 18096 6886 18148
rect 7006 18096 7012 18148
rect 7064 18136 7070 18148
rect 8938 18136 8944 18148
rect 7064 18108 8944 18136
rect 7064 18096 7070 18108
rect 8938 18096 8944 18108
rect 8996 18096 9002 18148
rect 1118 18028 1124 18080
rect 1176 18068 1182 18080
rect 3878 18068 3884 18080
rect 1176 18040 3884 18068
rect 1176 18028 1182 18040
rect 3878 18028 3884 18040
rect 3936 18028 3942 18080
rect 5169 18071 5227 18077
rect 5169 18037 5181 18071
rect 5215 18068 5227 18071
rect 5350 18068 5356 18080
rect 5215 18040 5356 18068
rect 5215 18037 5227 18040
rect 5169 18031 5227 18037
rect 5350 18028 5356 18040
rect 5408 18028 5414 18080
rect 6086 18068 6092 18080
rect 6047 18040 6092 18068
rect 6086 18028 6092 18040
rect 6144 18028 6150 18080
rect 7929 18071 7987 18077
rect 7929 18037 7941 18071
rect 7975 18068 7987 18071
rect 8018 18068 8024 18080
rect 7975 18040 8024 18068
rect 7975 18037 7987 18040
rect 7929 18031 7987 18037
rect 8018 18028 8024 18040
rect 8076 18028 8082 18080
rect 8202 18068 8208 18080
rect 8163 18040 8208 18068
rect 8202 18028 8208 18040
rect 8260 18028 8266 18080
rect 8478 18028 8484 18080
rect 8536 18068 8542 18080
rect 9508 18068 9536 18176
rect 10045 18173 10057 18207
rect 10091 18204 10103 18207
rect 10502 18204 10508 18216
rect 10091 18176 10508 18204
rect 10091 18173 10103 18176
rect 10045 18167 10103 18173
rect 10502 18164 10508 18176
rect 10560 18164 10566 18216
rect 14384 18204 14412 18244
rect 14461 18241 14473 18275
rect 14507 18241 14519 18275
rect 14461 18235 14519 18241
rect 14568 18204 14596 18312
rect 16218 18275 16276 18281
rect 16218 18272 16230 18275
rect 14384 18176 14596 18204
rect 15028 18244 16230 18272
rect 9950 18096 9956 18148
rect 10008 18136 10014 18148
rect 11517 18139 11575 18145
rect 11517 18136 11529 18139
rect 10008 18108 11529 18136
rect 10008 18096 10014 18108
rect 11517 18105 11529 18108
rect 11563 18105 11575 18139
rect 11517 18099 11575 18105
rect 11330 18068 11336 18080
rect 8536 18040 9536 18068
rect 11291 18040 11336 18068
rect 8536 18028 8542 18040
rect 11330 18028 11336 18040
rect 11388 18028 11394 18080
rect 11532 18068 11560 18099
rect 11974 18068 11980 18080
rect 11532 18040 11980 18068
rect 11974 18028 11980 18040
rect 12032 18028 12038 18080
rect 13078 18068 13084 18080
rect 13039 18040 13084 18068
rect 13078 18028 13084 18040
rect 13136 18028 13142 18080
rect 13170 18028 13176 18080
rect 13228 18068 13234 18080
rect 15028 18068 15056 18244
rect 16218 18241 16230 18244
rect 16264 18272 16276 18275
rect 16316 18272 16344 18380
rect 16669 18377 16681 18380
rect 16715 18377 16727 18411
rect 16669 18371 16727 18377
rect 17862 18368 17868 18420
rect 17920 18408 17926 18420
rect 18141 18411 18199 18417
rect 18141 18408 18153 18411
rect 17920 18380 18153 18408
rect 17920 18368 17926 18380
rect 18141 18377 18153 18380
rect 18187 18377 18199 18411
rect 18141 18371 18199 18377
rect 20990 18368 20996 18420
rect 21048 18408 21054 18420
rect 21085 18411 21143 18417
rect 21085 18408 21097 18411
rect 21048 18380 21097 18408
rect 21048 18368 21054 18380
rect 21085 18377 21097 18380
rect 21131 18377 21143 18411
rect 21085 18371 21143 18377
rect 18230 18340 18236 18352
rect 18064 18312 18236 18340
rect 16264 18244 16344 18272
rect 16264 18241 16276 18244
rect 16218 18235 16276 18241
rect 16390 18232 16396 18284
rect 16448 18272 16454 18284
rect 16485 18275 16543 18281
rect 16485 18272 16497 18275
rect 16448 18244 16497 18272
rect 16448 18232 16454 18244
rect 16485 18241 16497 18244
rect 16531 18241 16543 18275
rect 16485 18235 16543 18241
rect 17770 18232 17776 18284
rect 17828 18281 17834 18284
rect 18064 18281 18092 18312
rect 18230 18300 18236 18312
rect 18288 18340 18294 18352
rect 21008 18340 21036 18368
rect 18288 18312 21036 18340
rect 18288 18300 18294 18312
rect 17828 18272 17840 18281
rect 18049 18275 18107 18281
rect 17828 18244 17873 18272
rect 17828 18235 17840 18244
rect 18049 18241 18061 18275
rect 18095 18241 18107 18275
rect 18049 18235 18107 18241
rect 17828 18232 17834 18235
rect 18966 18232 18972 18284
rect 19024 18272 19030 18284
rect 19628 18281 19656 18312
rect 19254 18275 19312 18281
rect 19254 18272 19266 18275
rect 19024 18244 19266 18272
rect 19024 18232 19030 18244
rect 19254 18241 19266 18244
rect 19300 18241 19312 18275
rect 19254 18235 19312 18241
rect 19521 18275 19579 18281
rect 19521 18241 19533 18275
rect 19567 18272 19579 18275
rect 19613 18275 19671 18281
rect 19613 18272 19625 18275
rect 19567 18244 19625 18272
rect 19567 18241 19579 18244
rect 19521 18235 19579 18241
rect 19613 18241 19625 18244
rect 19659 18241 19671 18275
rect 19869 18275 19927 18281
rect 19869 18272 19881 18275
rect 19613 18235 19671 18241
rect 19720 18244 19881 18272
rect 19720 18204 19748 18244
rect 19869 18241 19881 18244
rect 19915 18241 19927 18275
rect 19869 18235 19927 18241
rect 19628 18176 19748 18204
rect 18064 18108 18644 18136
rect 13228 18040 15056 18068
rect 13228 18028 13234 18040
rect 16114 18028 16120 18080
rect 16172 18068 16178 18080
rect 18064 18068 18092 18108
rect 16172 18040 18092 18068
rect 18616 18068 18644 18108
rect 19628 18068 19656 18176
rect 20898 18096 20904 18148
rect 20956 18136 20962 18148
rect 20993 18139 21051 18145
rect 20993 18136 21005 18139
rect 20956 18108 21005 18136
rect 20956 18096 20962 18108
rect 20993 18105 21005 18108
rect 21039 18105 21051 18139
rect 20993 18099 21051 18105
rect 18616 18040 19656 18068
rect 16172 18028 16178 18040
rect 1104 17978 21896 18000
rect 1104 17926 3549 17978
rect 3601 17926 3613 17978
rect 3665 17926 3677 17978
rect 3729 17926 3741 17978
rect 3793 17926 3805 17978
rect 3857 17926 8747 17978
rect 8799 17926 8811 17978
rect 8863 17926 8875 17978
rect 8927 17926 8939 17978
rect 8991 17926 9003 17978
rect 9055 17926 13945 17978
rect 13997 17926 14009 17978
rect 14061 17926 14073 17978
rect 14125 17926 14137 17978
rect 14189 17926 14201 17978
rect 14253 17926 19143 17978
rect 19195 17926 19207 17978
rect 19259 17926 19271 17978
rect 19323 17926 19335 17978
rect 19387 17926 19399 17978
rect 19451 17926 21896 17978
rect 1104 17904 21896 17926
rect 2777 17867 2835 17873
rect 2777 17833 2789 17867
rect 2823 17864 2835 17867
rect 3050 17864 3056 17876
rect 2823 17836 3056 17864
rect 2823 17833 2835 17836
rect 2777 17827 2835 17833
rect 3050 17824 3056 17836
rect 3108 17824 3114 17876
rect 3418 17824 3424 17876
rect 3476 17864 3482 17876
rect 3789 17867 3847 17873
rect 3789 17864 3801 17867
rect 3476 17836 3801 17864
rect 3476 17824 3482 17836
rect 3789 17833 3801 17836
rect 3835 17864 3847 17867
rect 4522 17864 4528 17876
rect 3835 17836 4528 17864
rect 3835 17833 3847 17836
rect 3789 17827 3847 17833
rect 4522 17824 4528 17836
rect 4580 17824 4586 17876
rect 7006 17864 7012 17876
rect 5184 17836 7012 17864
rect 5184 17740 5212 17836
rect 7006 17824 7012 17836
rect 7064 17824 7070 17876
rect 8573 17867 8631 17873
rect 8573 17833 8585 17867
rect 8619 17864 8631 17867
rect 9214 17864 9220 17876
rect 8619 17836 9220 17864
rect 8619 17833 8631 17836
rect 8573 17827 8631 17833
rect 9214 17824 9220 17836
rect 9272 17824 9278 17876
rect 9950 17824 9956 17876
rect 10008 17864 10014 17876
rect 10962 17864 10968 17876
rect 10008 17836 10968 17864
rect 10008 17824 10014 17836
rect 10962 17824 10968 17836
rect 11020 17824 11026 17876
rect 11330 17824 11336 17876
rect 11388 17864 11394 17876
rect 11388 17836 13216 17864
rect 11388 17824 11394 17836
rect 6914 17756 6920 17808
rect 6972 17796 6978 17808
rect 11606 17796 11612 17808
rect 6972 17768 11612 17796
rect 6972 17756 6978 17768
rect 11606 17756 11612 17768
rect 11664 17756 11670 17808
rect 5166 17728 5172 17740
rect 5079 17700 5172 17728
rect 5166 17688 5172 17700
rect 5224 17688 5230 17740
rect 5350 17728 5356 17740
rect 5311 17700 5356 17728
rect 5350 17688 5356 17700
rect 5408 17688 5414 17740
rect 6086 17728 6092 17740
rect 5644 17700 6092 17728
rect 2961 17663 3019 17669
rect 2961 17629 2973 17663
rect 3007 17660 3019 17663
rect 3418 17660 3424 17672
rect 3007 17632 3424 17660
rect 3007 17629 3019 17632
rect 2961 17623 3019 17629
rect 3418 17620 3424 17632
rect 3476 17620 3482 17672
rect 4982 17620 4988 17672
rect 5040 17660 5046 17672
rect 5644 17660 5672 17700
rect 6086 17688 6092 17700
rect 6144 17728 6150 17740
rect 11716 17737 11744 17836
rect 13188 17805 13216 17836
rect 13446 17824 13452 17876
rect 13504 17864 13510 17876
rect 16850 17864 16856 17876
rect 13504 17836 16856 17864
rect 13504 17824 13510 17836
rect 16850 17824 16856 17836
rect 16908 17824 16914 17876
rect 18049 17867 18107 17873
rect 18049 17833 18061 17867
rect 18095 17864 18107 17867
rect 18233 17867 18291 17873
rect 18233 17864 18245 17867
rect 18095 17836 18245 17864
rect 18095 17833 18107 17836
rect 18049 17827 18107 17833
rect 18233 17833 18245 17836
rect 18279 17864 18291 17867
rect 19705 17867 19763 17873
rect 19705 17864 19717 17867
rect 18279 17836 19717 17864
rect 18279 17833 18291 17836
rect 18233 17827 18291 17833
rect 19705 17833 19717 17836
rect 19751 17864 19763 17867
rect 20990 17864 20996 17876
rect 19751 17836 20996 17864
rect 19751 17833 19763 17836
rect 19705 17827 19763 17833
rect 13173 17799 13231 17805
rect 13173 17765 13185 17799
rect 13219 17796 13231 17799
rect 13219 17768 13492 17796
rect 13219 17765 13231 17768
rect 13173 17759 13231 17765
rect 6457 17731 6515 17737
rect 6457 17728 6469 17731
rect 6144 17700 6469 17728
rect 6144 17688 6150 17700
rect 6457 17697 6469 17700
rect 6503 17728 6515 17731
rect 6733 17731 6791 17737
rect 6733 17728 6745 17731
rect 6503 17700 6745 17728
rect 6503 17697 6515 17700
rect 6457 17691 6515 17697
rect 6733 17697 6745 17700
rect 6779 17697 6791 17731
rect 6733 17691 6791 17697
rect 8021 17731 8079 17737
rect 8021 17697 8033 17731
rect 8067 17728 8079 17731
rect 11701 17731 11759 17737
rect 8067 17700 11652 17728
rect 8067 17697 8079 17700
rect 8021 17691 8079 17697
rect 5040 17632 5672 17660
rect 5040 17620 5046 17632
rect 5718 17620 5724 17672
rect 5776 17660 5782 17672
rect 6638 17660 6644 17672
rect 5776 17632 6644 17660
rect 5776 17620 5782 17632
rect 6638 17620 6644 17632
rect 6696 17620 6702 17672
rect 7466 17620 7472 17672
rect 7524 17660 7530 17672
rect 8205 17663 8263 17669
rect 8205 17660 8217 17663
rect 7524 17632 8217 17660
rect 7524 17620 7530 17632
rect 8205 17629 8217 17632
rect 8251 17629 8263 17663
rect 8205 17623 8263 17629
rect 9122 17620 9128 17672
rect 9180 17660 9186 17672
rect 9493 17663 9551 17669
rect 9493 17660 9505 17663
rect 9180 17632 9505 17660
rect 9180 17620 9186 17632
rect 9493 17629 9505 17632
rect 9539 17629 9551 17663
rect 9493 17623 9551 17629
rect 9769 17663 9827 17669
rect 9769 17629 9781 17663
rect 9815 17660 9827 17663
rect 9858 17660 9864 17672
rect 9815 17632 9864 17660
rect 9815 17629 9827 17632
rect 9769 17623 9827 17629
rect 9858 17620 9864 17632
rect 9916 17620 9922 17672
rect 11624 17660 11652 17700
rect 11701 17697 11713 17731
rect 11747 17697 11759 17731
rect 11701 17691 11759 17697
rect 12802 17688 12808 17740
rect 12860 17728 12866 17740
rect 13262 17728 13268 17740
rect 12860 17700 13268 17728
rect 12860 17688 12866 17700
rect 13262 17688 13268 17700
rect 13320 17688 13326 17740
rect 13464 17728 13492 17768
rect 13538 17756 13544 17808
rect 13596 17796 13602 17808
rect 13596 17768 14044 17796
rect 13596 17756 13602 17768
rect 13633 17731 13691 17737
rect 13633 17728 13645 17731
rect 13464 17700 13645 17728
rect 13633 17697 13645 17700
rect 13679 17728 13691 17731
rect 13722 17728 13728 17740
rect 13679 17700 13728 17728
rect 13679 17697 13691 17700
rect 13633 17691 13691 17697
rect 13722 17688 13728 17700
rect 13780 17688 13786 17740
rect 11624 17632 12480 17660
rect 3510 17552 3516 17604
rect 3568 17592 3574 17604
rect 4893 17595 4951 17601
rect 4893 17592 4905 17595
rect 3568 17564 4905 17592
rect 3568 17552 3574 17564
rect 4893 17561 4905 17564
rect 4939 17592 4951 17595
rect 6273 17595 6331 17601
rect 6273 17592 6285 17595
rect 4939 17564 6285 17592
rect 4939 17561 4951 17564
rect 4893 17555 4951 17561
rect 6273 17561 6285 17564
rect 6319 17561 6331 17595
rect 6273 17555 6331 17561
rect 7374 17552 7380 17604
rect 7432 17592 7438 17604
rect 8113 17595 8171 17601
rect 8113 17592 8125 17595
rect 7432 17564 8125 17592
rect 7432 17552 7438 17564
rect 8113 17561 8125 17564
rect 8159 17561 8171 17595
rect 8113 17555 8171 17561
rect 9214 17552 9220 17604
rect 9272 17592 9278 17604
rect 11968 17595 12026 17601
rect 9272 17564 11928 17592
rect 9272 17552 9278 17564
rect 4982 17484 4988 17536
rect 5040 17524 5046 17536
rect 5445 17527 5503 17533
rect 5445 17524 5457 17527
rect 5040 17496 5457 17524
rect 5040 17484 5046 17496
rect 5445 17493 5457 17496
rect 5491 17493 5503 17527
rect 5445 17487 5503 17493
rect 5718 17484 5724 17536
rect 5776 17524 5782 17536
rect 5813 17527 5871 17533
rect 5813 17524 5825 17527
rect 5776 17496 5825 17524
rect 5776 17484 5782 17496
rect 5813 17493 5825 17496
rect 5859 17493 5871 17527
rect 5813 17487 5871 17493
rect 5902 17484 5908 17536
rect 5960 17524 5966 17536
rect 6365 17527 6423 17533
rect 5960 17496 6005 17524
rect 5960 17484 5966 17496
rect 6365 17493 6377 17527
rect 6411 17524 6423 17527
rect 6546 17524 6552 17536
rect 6411 17496 6552 17524
rect 6411 17493 6423 17496
rect 6365 17487 6423 17493
rect 6546 17484 6552 17496
rect 6604 17484 6610 17536
rect 7745 17527 7803 17533
rect 7745 17493 7757 17527
rect 7791 17524 7803 17527
rect 7926 17524 7932 17536
rect 7791 17496 7932 17524
rect 7791 17493 7803 17496
rect 7745 17487 7803 17493
rect 7926 17484 7932 17496
rect 7984 17484 7990 17536
rect 9122 17484 9128 17536
rect 9180 17524 9186 17536
rect 9861 17527 9919 17533
rect 9861 17524 9873 17527
rect 9180 17496 9873 17524
rect 9180 17484 9186 17496
rect 9861 17493 9873 17496
rect 9907 17493 9919 17527
rect 11900 17524 11928 17564
rect 11968 17561 11980 17595
rect 12014 17592 12026 17595
rect 12342 17592 12348 17604
rect 12014 17564 12348 17592
rect 12014 17561 12026 17564
rect 11968 17555 12026 17561
rect 12342 17552 12348 17564
rect 12400 17552 12406 17604
rect 12452 17592 12480 17632
rect 12526 17620 12532 17672
rect 12584 17660 12590 17672
rect 14016 17660 14044 17768
rect 14366 17688 14372 17740
rect 14424 17728 14430 17740
rect 15102 17728 15108 17740
rect 14424 17700 15108 17728
rect 14424 17688 14430 17700
rect 15102 17688 15108 17700
rect 15160 17688 15166 17740
rect 16390 17688 16396 17740
rect 16448 17728 16454 17740
rect 19812 17737 19840 17836
rect 20990 17824 20996 17836
rect 21048 17864 21054 17876
rect 21269 17867 21327 17873
rect 21269 17864 21281 17867
rect 21048 17836 21281 17864
rect 21048 17824 21054 17836
rect 21269 17833 21281 17836
rect 21315 17833 21327 17867
rect 21269 17827 21327 17833
rect 16485 17731 16543 17737
rect 16485 17728 16497 17731
rect 16448 17700 16497 17728
rect 16448 17688 16454 17700
rect 16485 17697 16497 17700
rect 16531 17697 16543 17731
rect 16485 17691 16543 17697
rect 19797 17731 19855 17737
rect 19797 17697 19809 17731
rect 19843 17697 19855 17731
rect 19797 17691 19855 17697
rect 16741 17663 16799 17669
rect 16741 17660 16753 17663
rect 12584 17632 13584 17660
rect 14016 17632 16753 17660
rect 12584 17620 12590 17632
rect 13556 17592 13584 17632
rect 16741 17629 16753 17632
rect 16787 17629 16799 17663
rect 16741 17623 16799 17629
rect 19886 17620 19892 17672
rect 19944 17660 19950 17672
rect 20053 17663 20111 17669
rect 20053 17660 20065 17663
rect 19944 17632 20065 17660
rect 19944 17620 19950 17632
rect 20053 17629 20065 17632
rect 20099 17629 20111 17663
rect 20053 17623 20111 17629
rect 19702 17592 19708 17604
rect 12452 17564 12756 17592
rect 12526 17524 12532 17536
rect 11900 17496 12532 17524
rect 9861 17487 9919 17493
rect 12526 17484 12532 17496
rect 12584 17484 12590 17536
rect 12728 17524 12756 17564
rect 12912 17564 13492 17592
rect 13556 17564 19708 17592
rect 12912 17524 12940 17564
rect 12728 17496 12940 17524
rect 12986 17484 12992 17536
rect 13044 17524 13050 17536
rect 13081 17527 13139 17533
rect 13081 17524 13093 17527
rect 13044 17496 13093 17524
rect 13044 17484 13050 17496
rect 13081 17493 13093 17496
rect 13127 17493 13139 17527
rect 13464 17524 13492 17564
rect 19702 17552 19708 17564
rect 19760 17552 19766 17604
rect 17865 17527 17923 17533
rect 17865 17524 17877 17527
rect 13464 17496 17877 17524
rect 13081 17487 13139 17493
rect 17865 17493 17877 17496
rect 17911 17524 17923 17527
rect 18966 17524 18972 17536
rect 17911 17496 18972 17524
rect 17911 17493 17923 17496
rect 17865 17487 17923 17493
rect 18966 17484 18972 17496
rect 19024 17484 19030 17536
rect 21082 17484 21088 17536
rect 21140 17524 21146 17536
rect 21177 17527 21235 17533
rect 21177 17524 21189 17527
rect 21140 17496 21189 17524
rect 21140 17484 21146 17496
rect 21177 17493 21189 17496
rect 21223 17493 21235 17527
rect 21177 17487 21235 17493
rect 1104 17434 22056 17456
rect 1104 17382 6148 17434
rect 6200 17382 6212 17434
rect 6264 17382 6276 17434
rect 6328 17382 6340 17434
rect 6392 17382 6404 17434
rect 6456 17382 11346 17434
rect 11398 17382 11410 17434
rect 11462 17382 11474 17434
rect 11526 17382 11538 17434
rect 11590 17382 11602 17434
rect 11654 17382 16544 17434
rect 16596 17382 16608 17434
rect 16660 17382 16672 17434
rect 16724 17382 16736 17434
rect 16788 17382 16800 17434
rect 16852 17382 21742 17434
rect 21794 17382 21806 17434
rect 21858 17382 21870 17434
rect 21922 17382 21934 17434
rect 21986 17382 21998 17434
rect 22050 17382 22056 17434
rect 1104 17360 22056 17382
rect 2225 17323 2283 17329
rect 2225 17289 2237 17323
rect 2271 17320 2283 17323
rect 2958 17320 2964 17332
rect 2271 17292 2964 17320
rect 2271 17289 2283 17292
rect 2225 17283 2283 17289
rect 2958 17280 2964 17292
rect 3016 17280 3022 17332
rect 3326 17280 3332 17332
rect 3384 17320 3390 17332
rect 3973 17323 4031 17329
rect 3973 17320 3985 17323
rect 3384 17292 3985 17320
rect 3384 17280 3390 17292
rect 3973 17289 3985 17292
rect 4019 17320 4031 17323
rect 4062 17320 4068 17332
rect 4019 17292 4068 17320
rect 4019 17289 4031 17292
rect 3973 17283 4031 17289
rect 4062 17280 4068 17292
rect 4120 17320 4126 17332
rect 4433 17323 4491 17329
rect 4433 17320 4445 17323
rect 4120 17292 4445 17320
rect 4120 17280 4126 17292
rect 4433 17289 4445 17292
rect 4479 17289 4491 17323
rect 4433 17283 4491 17289
rect 4522 17280 4528 17332
rect 4580 17320 4586 17332
rect 4893 17323 4951 17329
rect 4580 17292 4625 17320
rect 4580 17280 4586 17292
rect 4893 17289 4905 17323
rect 4939 17320 4951 17323
rect 4982 17320 4988 17332
rect 4939 17292 4988 17320
rect 4939 17289 4951 17292
rect 4893 17283 4951 17289
rect 4982 17280 4988 17292
rect 5040 17280 5046 17332
rect 5445 17323 5503 17329
rect 5445 17289 5457 17323
rect 5491 17320 5503 17323
rect 5810 17320 5816 17332
rect 5491 17292 5816 17320
rect 5491 17289 5503 17292
rect 5445 17283 5503 17289
rect 5810 17280 5816 17292
rect 5868 17280 5874 17332
rect 5905 17323 5963 17329
rect 5905 17289 5917 17323
rect 5951 17320 5963 17323
rect 6917 17323 6975 17329
rect 6917 17320 6929 17323
rect 5951 17292 6929 17320
rect 5951 17289 5963 17292
rect 5905 17283 5963 17289
rect 6917 17289 6929 17292
rect 6963 17289 6975 17323
rect 7374 17320 7380 17332
rect 7335 17292 7380 17320
rect 6917 17283 6975 17289
rect 7374 17280 7380 17292
rect 7432 17280 7438 17332
rect 7926 17320 7932 17332
rect 7887 17292 7932 17320
rect 7926 17280 7932 17292
rect 7984 17280 7990 17332
rect 8297 17323 8355 17329
rect 8297 17289 8309 17323
rect 8343 17320 8355 17323
rect 8386 17320 8392 17332
rect 8343 17292 8392 17320
rect 8343 17289 8355 17292
rect 8297 17283 8355 17289
rect 8386 17280 8392 17292
rect 8444 17280 8450 17332
rect 9122 17320 9128 17332
rect 9083 17292 9128 17320
rect 9122 17280 9128 17292
rect 9180 17280 9186 17332
rect 9217 17323 9275 17329
rect 9217 17289 9229 17323
rect 9263 17320 9275 17323
rect 9585 17323 9643 17329
rect 9585 17320 9597 17323
rect 9263 17292 9597 17320
rect 9263 17289 9275 17292
rect 9217 17283 9275 17289
rect 9585 17289 9597 17292
rect 9631 17289 9643 17323
rect 13170 17320 13176 17332
rect 9585 17283 9643 17289
rect 10152 17292 13176 17320
rect 3418 17252 3424 17264
rect 3379 17224 3424 17252
rect 3418 17212 3424 17224
rect 3476 17212 3482 17264
rect 3881 17255 3939 17261
rect 3881 17221 3893 17255
rect 3927 17252 3939 17255
rect 4154 17252 4160 17264
rect 3927 17224 4160 17252
rect 3927 17221 3939 17224
rect 3881 17215 3939 17221
rect 4154 17212 4160 17224
rect 4212 17212 4218 17264
rect 5718 17212 5724 17264
rect 5776 17252 5782 17264
rect 7009 17255 7067 17261
rect 7009 17252 7021 17255
rect 5776 17224 7021 17252
rect 5776 17212 5782 17224
rect 7009 17221 7021 17224
rect 7055 17221 7067 17255
rect 7009 17215 7067 17221
rect 7837 17255 7895 17261
rect 7837 17221 7849 17255
rect 7883 17252 7895 17255
rect 8202 17252 8208 17264
rect 7883 17224 8208 17252
rect 7883 17221 7895 17224
rect 7837 17215 7895 17221
rect 8202 17212 8208 17224
rect 8260 17212 8266 17264
rect 8665 17255 8723 17261
rect 8665 17221 8677 17255
rect 8711 17252 8723 17255
rect 9306 17252 9312 17264
rect 8711 17224 9312 17252
rect 8711 17221 8723 17224
rect 8665 17215 8723 17221
rect 9306 17212 9312 17224
rect 9364 17252 9370 17264
rect 10045 17255 10103 17261
rect 10045 17252 10057 17255
rect 9364 17224 10057 17252
rect 9364 17212 9370 17224
rect 10045 17221 10057 17224
rect 10091 17221 10103 17255
rect 10045 17215 10103 17221
rect 2409 17187 2467 17193
rect 2409 17153 2421 17187
rect 2455 17153 2467 17187
rect 2409 17147 2467 17153
rect 2777 17187 2835 17193
rect 2777 17153 2789 17187
rect 2823 17184 2835 17187
rect 2958 17184 2964 17196
rect 2823 17156 2964 17184
rect 2823 17153 2835 17156
rect 2777 17147 2835 17153
rect 2424 17048 2452 17147
rect 2958 17144 2964 17156
rect 3016 17144 3022 17196
rect 3142 17184 3148 17196
rect 3103 17156 3148 17184
rect 3142 17144 3148 17156
rect 3200 17144 3206 17196
rect 3697 17187 3755 17193
rect 3697 17153 3709 17187
rect 3743 17153 3755 17187
rect 5534 17184 5540 17196
rect 5495 17156 5540 17184
rect 3697 17147 3755 17153
rect 2774 17048 2780 17060
rect 2424 17020 2780 17048
rect 2774 17008 2780 17020
rect 2832 17008 2838 17060
rect 2961 17051 3019 17057
rect 2961 17017 2973 17051
rect 3007 17048 3019 17051
rect 3234 17048 3240 17060
rect 3007 17020 3240 17048
rect 3007 17017 3019 17020
rect 2961 17011 3019 17017
rect 3234 17008 3240 17020
rect 3292 17008 3298 17060
rect 3712 17048 3740 17147
rect 5534 17144 5540 17156
rect 5592 17144 5598 17196
rect 8386 17144 8392 17196
rect 8444 17184 8450 17196
rect 9953 17187 10011 17193
rect 9953 17184 9965 17187
rect 8444 17156 9965 17184
rect 8444 17144 8450 17156
rect 9953 17153 9965 17156
rect 9999 17153 10011 17187
rect 9953 17147 10011 17153
rect 4341 17119 4399 17125
rect 4341 17085 4353 17119
rect 4387 17116 4399 17119
rect 4890 17116 4896 17128
rect 4387 17088 4896 17116
rect 4387 17085 4399 17088
rect 4341 17079 4399 17085
rect 4890 17076 4896 17088
rect 4948 17116 4954 17128
rect 4985 17119 5043 17125
rect 4985 17116 4997 17119
rect 4948 17088 4997 17116
rect 4948 17076 4954 17088
rect 4985 17085 4997 17088
rect 5031 17085 5043 17119
rect 4985 17079 5043 17085
rect 5166 17076 5172 17128
rect 5224 17116 5230 17128
rect 5261 17119 5319 17125
rect 5261 17116 5273 17119
rect 5224 17088 5273 17116
rect 5224 17076 5230 17088
rect 5261 17085 5273 17088
rect 5307 17116 5319 17119
rect 5442 17116 5448 17128
rect 5307 17088 5448 17116
rect 5307 17085 5319 17088
rect 5261 17079 5319 17085
rect 5442 17076 5448 17088
rect 5500 17076 5506 17128
rect 6825 17119 6883 17125
rect 6825 17085 6837 17119
rect 6871 17116 6883 17119
rect 6914 17116 6920 17128
rect 6871 17088 6920 17116
rect 6871 17085 6883 17088
rect 6825 17079 6883 17085
rect 6914 17076 6920 17088
rect 6972 17116 6978 17128
rect 7190 17116 7196 17128
rect 6972 17088 7196 17116
rect 6972 17076 6978 17088
rect 7190 17076 7196 17088
rect 7248 17076 7254 17128
rect 7742 17116 7748 17128
rect 7703 17088 7748 17116
rect 7742 17076 7748 17088
rect 7800 17076 7806 17128
rect 9401 17119 9459 17125
rect 9401 17085 9413 17119
rect 9447 17116 9459 17119
rect 10152 17116 10180 17292
rect 13170 17280 13176 17292
rect 13228 17280 13234 17332
rect 13354 17280 13360 17332
rect 13412 17320 13418 17332
rect 20162 17320 20168 17332
rect 13412 17292 16804 17320
rect 13412 17280 13418 17292
rect 10686 17252 10692 17264
rect 10647 17224 10692 17252
rect 10686 17212 10692 17224
rect 10744 17212 10750 17264
rect 10962 17212 10968 17264
rect 11020 17252 11026 17264
rect 12652 17255 12710 17261
rect 12652 17252 12664 17255
rect 11020 17224 12664 17252
rect 11020 17212 11026 17224
rect 12652 17221 12664 17224
rect 12698 17252 12710 17255
rect 12802 17252 12808 17264
rect 12698 17224 12808 17252
rect 12698 17221 12710 17224
rect 12652 17215 12710 17221
rect 12802 17212 12808 17224
rect 12860 17212 12866 17264
rect 14461 17255 14519 17261
rect 14461 17252 14473 17255
rect 13004 17224 14473 17252
rect 10410 17184 10416 17196
rect 10371 17156 10416 17184
rect 10410 17144 10416 17156
rect 10468 17144 10474 17196
rect 13004 17125 13032 17224
rect 14461 17221 14473 17224
rect 14507 17252 14519 17255
rect 15838 17252 15844 17264
rect 14507 17224 15844 17252
rect 14507 17221 14519 17224
rect 14461 17215 14519 17221
rect 15838 17212 15844 17224
rect 15896 17252 15902 17264
rect 16390 17252 16396 17264
rect 15896 17224 16396 17252
rect 15896 17212 15902 17224
rect 16390 17212 16396 17224
rect 16448 17252 16454 17264
rect 16448 17224 16528 17252
rect 16448 17212 16454 17224
rect 13256 17187 13314 17193
rect 13256 17153 13268 17187
rect 13302 17184 13314 17187
rect 14366 17184 14372 17196
rect 13302 17156 14372 17184
rect 13302 17153 13314 17156
rect 13256 17147 13314 17153
rect 14366 17144 14372 17156
rect 14424 17144 14430 17196
rect 16206 17144 16212 17196
rect 16264 17193 16270 17196
rect 16500 17193 16528 17224
rect 16264 17184 16276 17193
rect 16485 17187 16543 17193
rect 16264 17156 16309 17184
rect 16264 17147 16276 17156
rect 16485 17153 16497 17187
rect 16531 17153 16543 17187
rect 16776 17184 16804 17292
rect 17972 17292 20168 17320
rect 17782 17187 17840 17193
rect 17782 17184 17794 17187
rect 16776 17156 17794 17184
rect 16485 17147 16543 17153
rect 17782 17153 17794 17156
rect 17828 17184 17840 17187
rect 17972 17184 18000 17292
rect 20162 17280 20168 17292
rect 20220 17280 20226 17332
rect 20533 17323 20591 17329
rect 20533 17289 20545 17323
rect 20579 17320 20591 17323
rect 20990 17320 20996 17332
rect 20579 17292 20996 17320
rect 20579 17289 20591 17292
rect 20533 17283 20591 17289
rect 20548 17252 20576 17283
rect 20990 17280 20996 17292
rect 21048 17280 21054 17332
rect 17828 17156 18000 17184
rect 18984 17224 20576 17252
rect 17828 17153 17840 17156
rect 17782 17147 17840 17153
rect 16264 17144 16270 17147
rect 9447 17088 10180 17116
rect 10229 17119 10287 17125
rect 9447 17085 9459 17088
rect 9401 17079 9459 17085
rect 10229 17085 10241 17119
rect 10275 17116 10287 17119
rect 12897 17119 12955 17125
rect 10275 17088 11928 17116
rect 10275 17085 10287 17088
rect 10229 17079 10287 17085
rect 8757 17051 8815 17057
rect 8757 17048 8769 17051
rect 3712 17020 8769 17048
rect 8757 17017 8769 17020
rect 8803 17017 8815 17051
rect 8757 17011 8815 17017
rect 2593 16983 2651 16989
rect 2593 16949 2605 16983
rect 2639 16980 2651 16983
rect 2866 16980 2872 16992
rect 2639 16952 2872 16980
rect 2639 16949 2651 16952
rect 2593 16943 2651 16949
rect 2866 16940 2872 16952
rect 2924 16940 2930 16992
rect 4614 16940 4620 16992
rect 4672 16980 4678 16992
rect 5997 16983 6055 16989
rect 5997 16980 6009 16983
rect 4672 16952 6009 16980
rect 4672 16940 4678 16952
rect 5997 16949 6009 16952
rect 6043 16980 6055 16983
rect 6546 16980 6552 16992
rect 6043 16952 6552 16980
rect 6043 16949 6055 16952
rect 5997 16943 6055 16949
rect 6546 16940 6552 16952
rect 6604 16940 6610 16992
rect 8386 16980 8392 16992
rect 8347 16952 8392 16980
rect 8386 16940 8392 16952
rect 8444 16940 8450 16992
rect 9122 16940 9128 16992
rect 9180 16980 9186 16992
rect 9766 16980 9772 16992
rect 9180 16952 9772 16980
rect 9180 16940 9186 16952
rect 9766 16940 9772 16952
rect 9824 16940 9830 16992
rect 10686 16940 10692 16992
rect 10744 16980 10750 16992
rect 10962 16980 10968 16992
rect 10744 16952 10968 16980
rect 10744 16940 10750 16952
rect 10962 16940 10968 16952
rect 11020 16940 11026 16992
rect 11514 16980 11520 16992
rect 11475 16952 11520 16980
rect 11514 16940 11520 16952
rect 11572 16940 11578 16992
rect 11900 16980 11928 17088
rect 12897 17085 12909 17119
rect 12943 17116 12955 17119
rect 12989 17119 13047 17125
rect 12989 17116 13001 17119
rect 12943 17088 13001 17116
rect 12943 17085 12955 17088
rect 12897 17079 12955 17085
rect 12989 17085 13001 17088
rect 13035 17085 13047 17119
rect 18046 17116 18052 17128
rect 12989 17079 13047 17085
rect 14292 17088 15240 17116
rect 18007 17088 18052 17116
rect 14292 16980 14320 17088
rect 15102 17048 15108 17060
rect 15063 17020 15108 17048
rect 15102 17008 15108 17020
rect 15160 17008 15166 17060
rect 15212 17048 15240 17088
rect 18046 17076 18052 17088
rect 18104 17116 18110 17128
rect 18984 17125 19012 17224
rect 19058 17144 19064 17196
rect 19116 17184 19122 17196
rect 19225 17187 19283 17193
rect 19225 17184 19237 17187
rect 19116 17156 19237 17184
rect 19116 17144 19122 17156
rect 19225 17153 19237 17156
rect 19271 17153 19283 17187
rect 19225 17147 19283 17153
rect 18141 17119 18199 17125
rect 18141 17116 18153 17119
rect 18104 17088 18153 17116
rect 18104 17076 18110 17088
rect 18141 17085 18153 17088
rect 18187 17116 18199 17119
rect 18969 17119 19027 17125
rect 18969 17116 18981 17119
rect 18187 17088 18981 17116
rect 18187 17085 18199 17088
rect 18141 17079 18199 17085
rect 18969 17085 18981 17088
rect 19015 17085 19027 17119
rect 18969 17079 19027 17085
rect 15212 17020 15608 17048
rect 11900 16952 14320 16980
rect 14369 16983 14427 16989
rect 14369 16949 14381 16983
rect 14415 16980 14427 16983
rect 15470 16980 15476 16992
rect 14415 16952 15476 16980
rect 14415 16949 14427 16952
rect 14369 16943 14427 16949
rect 15470 16940 15476 16952
rect 15528 16940 15534 16992
rect 15580 16980 15608 17020
rect 16669 16983 16727 16989
rect 16669 16980 16681 16983
rect 15580 16952 16681 16980
rect 16669 16949 16681 16952
rect 16715 16980 16727 16983
rect 17770 16980 17776 16992
rect 16715 16952 17776 16980
rect 16715 16949 16727 16952
rect 16669 16943 16727 16949
rect 17770 16940 17776 16952
rect 17828 16940 17834 16992
rect 20346 16980 20352 16992
rect 20307 16952 20352 16980
rect 20346 16940 20352 16952
rect 20404 16940 20410 16992
rect 1104 16890 21896 16912
rect 1104 16838 3549 16890
rect 3601 16838 3613 16890
rect 3665 16838 3677 16890
rect 3729 16838 3741 16890
rect 3793 16838 3805 16890
rect 3857 16838 8747 16890
rect 8799 16838 8811 16890
rect 8863 16838 8875 16890
rect 8927 16838 8939 16890
rect 8991 16838 9003 16890
rect 9055 16838 13945 16890
rect 13997 16838 14009 16890
rect 14061 16838 14073 16890
rect 14125 16838 14137 16890
rect 14189 16838 14201 16890
rect 14253 16838 19143 16890
rect 19195 16838 19207 16890
rect 19259 16838 19271 16890
rect 19323 16838 19335 16890
rect 19387 16838 19399 16890
rect 19451 16838 21896 16890
rect 1104 16816 21896 16838
rect 3878 16776 3884 16788
rect 3839 16748 3884 16776
rect 3878 16736 3884 16748
rect 3936 16736 3942 16788
rect 4338 16736 4344 16788
rect 4396 16776 4402 16788
rect 6546 16776 6552 16788
rect 4396 16748 6552 16776
rect 4396 16736 4402 16748
rect 6546 16736 6552 16748
rect 6604 16736 6610 16788
rect 12526 16776 12532 16788
rect 10980 16748 12532 16776
rect 658 16668 664 16720
rect 716 16708 722 16720
rect 3418 16708 3424 16720
rect 716 16680 3424 16708
rect 716 16668 722 16680
rect 3418 16668 3424 16680
rect 3476 16668 3482 16720
rect 9122 16708 9128 16720
rect 7760 16680 9128 16708
rect 2958 16600 2964 16652
rect 3016 16640 3022 16652
rect 3329 16643 3387 16649
rect 3329 16640 3341 16643
rect 3016 16612 3341 16640
rect 3016 16600 3022 16612
rect 3329 16609 3341 16612
rect 3375 16609 3387 16643
rect 3329 16603 3387 16609
rect 4157 16643 4215 16649
rect 4157 16609 4169 16643
rect 4203 16640 4215 16643
rect 4890 16640 4896 16652
rect 4203 16612 4896 16640
rect 4203 16609 4215 16612
rect 4157 16603 4215 16609
rect 4890 16600 4896 16612
rect 4948 16600 4954 16652
rect 6178 16640 6184 16652
rect 5460 16612 5672 16640
rect 6139 16612 6184 16640
rect 2774 16532 2780 16584
rect 2832 16572 2838 16584
rect 3053 16575 3111 16581
rect 2832 16544 2877 16572
rect 2832 16532 2838 16544
rect 3053 16541 3065 16575
rect 3099 16541 3111 16575
rect 3602 16572 3608 16584
rect 3563 16544 3608 16572
rect 3053 16535 3111 16541
rect 3068 16504 3096 16535
rect 3602 16532 3608 16544
rect 3660 16532 3666 16584
rect 5460 16572 5488 16612
rect 3712 16544 5488 16572
rect 3712 16504 3740 16544
rect 5534 16532 5540 16584
rect 5592 16532 5598 16584
rect 3068 16476 3740 16504
rect 4154 16464 4160 16516
rect 4212 16504 4218 16516
rect 4341 16507 4399 16513
rect 4341 16504 4353 16507
rect 4212 16476 4353 16504
rect 4212 16464 4218 16476
rect 4341 16473 4353 16476
rect 4387 16473 4399 16507
rect 5552 16504 5580 16532
rect 4341 16467 4399 16473
rect 4724 16476 5580 16504
rect 5644 16504 5672 16612
rect 6178 16600 6184 16612
rect 6236 16600 6242 16652
rect 7558 16640 7564 16652
rect 7519 16612 7564 16640
rect 7558 16600 7564 16612
rect 7616 16600 7622 16652
rect 7760 16649 7788 16680
rect 9122 16668 9128 16680
rect 9180 16668 9186 16720
rect 10686 16708 10692 16720
rect 9692 16680 10692 16708
rect 7745 16643 7803 16649
rect 7745 16609 7757 16643
rect 7791 16609 7803 16643
rect 8110 16640 8116 16652
rect 8071 16612 8116 16640
rect 7745 16603 7803 16609
rect 8110 16600 8116 16612
rect 8168 16600 8174 16652
rect 9692 16649 9720 16680
rect 10686 16668 10692 16680
rect 10744 16668 10750 16720
rect 10980 16649 11008 16748
rect 12526 16736 12532 16748
rect 12584 16736 12590 16788
rect 13814 16736 13820 16788
rect 13872 16776 13878 16788
rect 14369 16779 14427 16785
rect 14369 16776 14381 16779
rect 13872 16748 14381 16776
rect 13872 16736 13878 16748
rect 14369 16745 14381 16748
rect 14415 16745 14427 16779
rect 15838 16776 15844 16788
rect 15799 16748 15844 16776
rect 14369 16739 14427 16745
rect 15838 16736 15844 16748
rect 15896 16776 15902 16788
rect 16577 16779 16635 16785
rect 16577 16776 16589 16779
rect 15896 16748 16589 16776
rect 15896 16736 15902 16748
rect 16577 16745 16589 16748
rect 16623 16776 16635 16779
rect 18046 16776 18052 16788
rect 16623 16748 18052 16776
rect 16623 16745 16635 16748
rect 16577 16739 16635 16745
rect 18046 16736 18052 16748
rect 18104 16776 18110 16788
rect 18325 16779 18383 16785
rect 18325 16776 18337 16779
rect 18104 16748 18337 16776
rect 18104 16736 18110 16748
rect 9677 16643 9735 16649
rect 9677 16609 9689 16643
rect 9723 16609 9735 16643
rect 9861 16643 9919 16649
rect 9861 16640 9873 16643
rect 9677 16603 9735 16609
rect 9784 16612 9873 16640
rect 5718 16532 5724 16584
rect 5776 16572 5782 16584
rect 6365 16575 6423 16581
rect 6365 16572 6377 16575
rect 5776 16544 6377 16572
rect 5776 16532 5782 16544
rect 6365 16541 6377 16544
rect 6411 16541 6423 16575
rect 6365 16535 6423 16541
rect 8662 16532 8668 16584
rect 8720 16572 8726 16584
rect 9217 16575 9275 16581
rect 9217 16572 9229 16575
rect 8720 16544 9229 16572
rect 8720 16532 8726 16544
rect 9217 16541 9229 16544
rect 9263 16541 9275 16575
rect 9490 16572 9496 16584
rect 9451 16544 9496 16572
rect 9217 16535 9275 16541
rect 9490 16532 9496 16544
rect 9548 16532 9554 16584
rect 9784 16572 9812 16612
rect 9861 16609 9873 16612
rect 9907 16609 9919 16643
rect 9861 16603 9919 16609
rect 10965 16643 11023 16649
rect 10965 16609 10977 16643
rect 11011 16609 11023 16643
rect 10965 16603 11023 16609
rect 11609 16643 11667 16649
rect 11609 16609 11621 16643
rect 11655 16640 11667 16643
rect 12250 16640 12256 16652
rect 11655 16612 12256 16640
rect 11655 16609 11667 16612
rect 11609 16603 11667 16609
rect 9600 16544 9812 16572
rect 9953 16575 10011 16581
rect 7009 16507 7067 16513
rect 5644 16476 6684 16504
rect 3878 16396 3884 16448
rect 3936 16436 3942 16448
rect 4724 16445 4752 16476
rect 4249 16439 4307 16445
rect 4249 16436 4261 16439
rect 3936 16408 4261 16436
rect 3936 16396 3942 16408
rect 4249 16405 4261 16408
rect 4295 16405 4307 16439
rect 4249 16399 4307 16405
rect 4709 16439 4767 16445
rect 4709 16405 4721 16439
rect 4755 16405 4767 16439
rect 4709 16399 4767 16405
rect 4890 16396 4896 16448
rect 4948 16436 4954 16448
rect 5350 16436 5356 16448
rect 4948 16408 5356 16436
rect 4948 16396 4954 16408
rect 5350 16396 5356 16408
rect 5408 16396 5414 16448
rect 5534 16436 5540 16448
rect 5495 16408 5540 16436
rect 5534 16396 5540 16408
rect 5592 16396 5598 16448
rect 5902 16436 5908 16448
rect 5863 16408 5908 16436
rect 5902 16396 5908 16408
rect 5960 16396 5966 16448
rect 5994 16396 6000 16448
rect 6052 16436 6058 16448
rect 6656 16436 6684 16476
rect 7009 16473 7021 16507
rect 7055 16504 7067 16507
rect 7469 16507 7527 16513
rect 7469 16504 7481 16507
rect 7055 16476 7481 16504
rect 7055 16473 7067 16476
rect 7009 16467 7067 16473
rect 7469 16473 7481 16476
rect 7515 16473 7527 16507
rect 8294 16504 8300 16516
rect 8255 16476 8300 16504
rect 7469 16467 7527 16473
rect 8294 16464 8300 16476
rect 8352 16464 8358 16516
rect 9122 16504 9128 16516
rect 8588 16476 9128 16504
rect 7101 16439 7159 16445
rect 7101 16436 7113 16439
rect 6052 16408 6097 16436
rect 6656 16408 7113 16436
rect 6052 16396 6058 16408
rect 7101 16405 7113 16408
rect 7147 16405 7159 16439
rect 7101 16399 7159 16405
rect 8205 16439 8263 16445
rect 8205 16405 8217 16439
rect 8251 16436 8263 16439
rect 8588 16436 8616 16476
rect 9122 16464 9128 16476
rect 9180 16464 9186 16516
rect 9306 16464 9312 16516
rect 9364 16504 9370 16516
rect 9600 16504 9628 16544
rect 9953 16541 9965 16575
rect 9999 16572 10011 16575
rect 11146 16572 11152 16584
rect 9999 16544 11152 16572
rect 9999 16541 10011 16544
rect 9953 16535 10011 16541
rect 11146 16532 11152 16544
rect 11204 16572 11210 16584
rect 11624 16572 11652 16603
rect 12250 16600 12256 16612
rect 12308 16600 12314 16652
rect 13541 16643 13599 16649
rect 13541 16640 13553 16643
rect 13208 16612 13553 16640
rect 11204 16544 11652 16572
rect 11204 16532 11210 16544
rect 9364 16476 9628 16504
rect 9364 16464 9370 16476
rect 9766 16464 9772 16516
rect 9824 16504 9830 16516
rect 10781 16507 10839 16513
rect 9824 16476 10456 16504
rect 9824 16464 9830 16476
rect 8251 16408 8616 16436
rect 8665 16439 8723 16445
rect 8251 16405 8263 16408
rect 8205 16399 8263 16405
rect 8665 16405 8677 16439
rect 8711 16436 8723 16439
rect 9398 16436 9404 16448
rect 8711 16408 9404 16436
rect 8711 16405 8723 16408
rect 8665 16399 8723 16405
rect 9398 16396 9404 16408
rect 9456 16396 9462 16448
rect 10318 16436 10324 16448
rect 10279 16408 10324 16436
rect 10318 16396 10324 16408
rect 10376 16396 10382 16448
rect 10428 16445 10456 16476
rect 10781 16473 10793 16507
rect 10827 16504 10839 16507
rect 11241 16507 11299 16513
rect 11241 16504 11253 16507
rect 10827 16476 11253 16504
rect 10827 16473 10839 16476
rect 10781 16467 10839 16473
rect 11241 16473 11253 16476
rect 11287 16473 11299 16507
rect 11241 16467 11299 16473
rect 12986 16464 12992 16516
rect 13044 16513 13050 16516
rect 13044 16504 13056 16513
rect 13208 16504 13236 16612
rect 13541 16609 13553 16612
rect 13587 16640 13599 16643
rect 14734 16640 14740 16652
rect 13587 16612 14740 16640
rect 13587 16609 13599 16612
rect 13541 16603 13599 16609
rect 14734 16600 14740 16612
rect 14792 16600 14798 16652
rect 15749 16643 15807 16649
rect 15749 16609 15761 16643
rect 15795 16640 15807 16643
rect 15856 16640 15884 16736
rect 18248 16649 18276 16748
rect 18325 16745 18337 16748
rect 18371 16745 18383 16779
rect 18325 16739 18383 16745
rect 20809 16779 20867 16785
rect 20809 16745 20821 16779
rect 20855 16776 20867 16779
rect 20990 16776 20996 16788
rect 20855 16748 20996 16776
rect 20855 16745 20867 16748
rect 20809 16739 20867 16745
rect 15795 16612 15884 16640
rect 18233 16643 18291 16649
rect 15795 16609 15807 16612
rect 15749 16603 15807 16609
rect 18233 16609 18245 16643
rect 18279 16609 18291 16643
rect 18233 16603 18291 16609
rect 20625 16643 20683 16649
rect 20625 16609 20637 16643
rect 20671 16640 20683 16643
rect 20824 16640 20852 16739
rect 20990 16736 20996 16748
rect 21048 16776 21054 16788
rect 21269 16779 21327 16785
rect 21269 16776 21281 16779
rect 21048 16748 21281 16776
rect 21048 16736 21054 16748
rect 21269 16745 21281 16748
rect 21315 16776 21327 16779
rect 21450 16776 21456 16788
rect 21315 16748 21456 16776
rect 21315 16745 21327 16748
rect 21269 16739 21327 16745
rect 21450 16736 21456 16748
rect 21508 16736 21514 16788
rect 20671 16612 20852 16640
rect 20671 16609 20683 16612
rect 20625 16603 20683 16609
rect 13265 16575 13323 16581
rect 13265 16541 13277 16575
rect 13311 16541 13323 16575
rect 13265 16535 13323 16541
rect 13044 16476 13236 16504
rect 13280 16504 13308 16535
rect 13354 16532 13360 16584
rect 13412 16572 13418 16584
rect 20358 16575 20416 16581
rect 20358 16572 20370 16575
rect 13412 16544 20370 16572
rect 13412 16532 13418 16544
rect 20358 16541 20370 16544
rect 20404 16541 20416 16575
rect 20358 16535 20416 16541
rect 13449 16507 13507 16513
rect 13449 16504 13461 16507
rect 13280 16476 13461 16504
rect 13044 16467 13056 16476
rect 13449 16473 13461 16476
rect 13495 16504 13507 16507
rect 13722 16504 13728 16516
rect 13495 16476 13728 16504
rect 13495 16473 13507 16476
rect 13449 16467 13507 16473
rect 13044 16464 13050 16467
rect 13722 16464 13728 16476
rect 13780 16504 13786 16516
rect 15194 16504 15200 16516
rect 13780 16476 15200 16504
rect 13780 16464 13786 16476
rect 15194 16464 15200 16476
rect 15252 16464 15258 16516
rect 15378 16464 15384 16516
rect 15436 16504 15442 16516
rect 15482 16507 15540 16513
rect 15482 16504 15494 16507
rect 15436 16476 15494 16504
rect 15436 16464 15442 16476
rect 15482 16473 15494 16476
rect 15528 16504 15540 16507
rect 16025 16507 16083 16513
rect 16025 16504 16037 16507
rect 15528 16476 16037 16504
rect 15528 16473 15540 16476
rect 15482 16467 15540 16473
rect 16025 16473 16037 16476
rect 16071 16504 16083 16507
rect 16390 16504 16396 16516
rect 16071 16476 16396 16504
rect 16071 16473 16083 16476
rect 16025 16467 16083 16473
rect 16390 16464 16396 16476
rect 16448 16464 16454 16516
rect 17954 16464 17960 16516
rect 18012 16513 18018 16516
rect 18012 16504 18024 16513
rect 18012 16476 18057 16504
rect 18012 16467 18024 16476
rect 18012 16464 18018 16467
rect 10413 16439 10471 16445
rect 10413 16405 10425 16439
rect 10459 16405 10471 16439
rect 10413 16399 10471 16405
rect 10873 16439 10931 16445
rect 10873 16405 10885 16439
rect 10919 16436 10931 16439
rect 11054 16436 11060 16448
rect 10919 16408 11060 16436
rect 10919 16405 10931 16408
rect 10873 16399 10931 16405
rect 11054 16396 11060 16408
rect 11112 16396 11118 16448
rect 11885 16439 11943 16445
rect 11885 16405 11897 16439
rect 11931 16436 11943 16439
rect 11974 16436 11980 16448
rect 11931 16408 11980 16436
rect 11931 16405 11943 16408
rect 11885 16399 11943 16405
rect 11974 16396 11980 16408
rect 12032 16396 12038 16448
rect 12066 16396 12072 16448
rect 12124 16436 12130 16448
rect 13814 16436 13820 16448
rect 12124 16408 13820 16436
rect 12124 16396 12130 16408
rect 13814 16396 13820 16408
rect 13872 16396 13878 16448
rect 14734 16396 14740 16448
rect 14792 16436 14798 16448
rect 16853 16439 16911 16445
rect 16853 16436 16865 16439
rect 14792 16408 16865 16436
rect 14792 16396 14798 16408
rect 16853 16405 16865 16408
rect 16899 16405 16911 16439
rect 16853 16399 16911 16405
rect 18966 16396 18972 16448
rect 19024 16436 19030 16448
rect 19245 16439 19303 16445
rect 19245 16436 19257 16439
rect 19024 16408 19257 16436
rect 19024 16396 19030 16408
rect 19245 16405 19257 16408
rect 19291 16405 19303 16439
rect 19245 16399 19303 16405
rect 21358 16396 21364 16448
rect 21416 16436 21422 16448
rect 21453 16439 21511 16445
rect 21453 16436 21465 16439
rect 21416 16408 21465 16436
rect 21416 16396 21422 16408
rect 21453 16405 21465 16408
rect 21499 16405 21511 16439
rect 21453 16399 21511 16405
rect 1104 16346 22056 16368
rect 1104 16294 6148 16346
rect 6200 16294 6212 16346
rect 6264 16294 6276 16346
rect 6328 16294 6340 16346
rect 6392 16294 6404 16346
rect 6456 16294 11346 16346
rect 11398 16294 11410 16346
rect 11462 16294 11474 16346
rect 11526 16294 11538 16346
rect 11590 16294 11602 16346
rect 11654 16294 16544 16346
rect 16596 16294 16608 16346
rect 16660 16294 16672 16346
rect 16724 16294 16736 16346
rect 16788 16294 16800 16346
rect 16852 16294 21742 16346
rect 21794 16294 21806 16346
rect 21858 16294 21870 16346
rect 21922 16294 21934 16346
rect 21986 16294 21998 16346
rect 22050 16294 22056 16346
rect 1104 16272 22056 16294
rect 4062 16232 4068 16244
rect 4023 16204 4068 16232
rect 4062 16192 4068 16204
rect 4120 16192 4126 16244
rect 4338 16232 4344 16244
rect 4299 16204 4344 16232
rect 4338 16192 4344 16204
rect 4396 16192 4402 16244
rect 5261 16235 5319 16241
rect 5261 16201 5273 16235
rect 5307 16232 5319 16235
rect 5902 16232 5908 16244
rect 5307 16204 5908 16232
rect 5307 16201 5319 16204
rect 5261 16195 5319 16201
rect 5902 16192 5908 16204
rect 5960 16192 5966 16244
rect 6089 16235 6147 16241
rect 6089 16201 6101 16235
rect 6135 16232 6147 16235
rect 7745 16235 7803 16241
rect 7745 16232 7757 16235
rect 6135 16204 7757 16232
rect 6135 16201 6147 16204
rect 6089 16195 6147 16201
rect 7745 16201 7757 16204
rect 7791 16201 7803 16235
rect 7745 16195 7803 16201
rect 9306 16192 9312 16244
rect 9364 16232 9370 16244
rect 10597 16235 10655 16241
rect 9364 16204 10088 16232
rect 9364 16192 9370 16204
rect 3050 16164 3056 16176
rect 3011 16136 3056 16164
rect 3050 16124 3056 16136
rect 3108 16124 3114 16176
rect 3142 16124 3148 16176
rect 3200 16164 3206 16176
rect 3605 16167 3663 16173
rect 3605 16164 3617 16167
rect 3200 16136 3617 16164
rect 3200 16124 3206 16136
rect 3605 16133 3617 16136
rect 3651 16133 3663 16167
rect 5534 16164 5540 16176
rect 3605 16127 3663 16133
rect 3804 16136 5540 16164
rect 3329 16099 3387 16105
rect 3329 16065 3341 16099
rect 3375 16096 3387 16099
rect 3804 16096 3832 16136
rect 5534 16124 5540 16136
rect 5592 16124 5598 16176
rect 6546 16124 6552 16176
rect 6604 16164 6610 16176
rect 6917 16167 6975 16173
rect 6917 16164 6929 16167
rect 6604 16136 6929 16164
rect 6604 16124 6610 16136
rect 6917 16133 6929 16136
rect 6963 16133 6975 16167
rect 6917 16127 6975 16133
rect 9769 16167 9827 16173
rect 9769 16133 9781 16167
rect 9815 16164 9827 16167
rect 9950 16164 9956 16176
rect 9815 16136 9956 16164
rect 9815 16133 9827 16136
rect 9769 16127 9827 16133
rect 9950 16124 9956 16136
rect 10008 16124 10014 16176
rect 10060 16164 10088 16204
rect 10597 16201 10609 16235
rect 10643 16232 10655 16235
rect 10778 16232 10784 16244
rect 10643 16204 10784 16232
rect 10643 16201 10655 16204
rect 10597 16195 10655 16201
rect 10778 16192 10784 16204
rect 10836 16192 10842 16244
rect 11054 16232 11060 16244
rect 11015 16204 11060 16232
rect 11054 16192 11060 16204
rect 11112 16192 11118 16244
rect 11146 16192 11152 16244
rect 11204 16232 11210 16244
rect 14826 16232 14832 16244
rect 11204 16204 14832 16232
rect 11204 16192 11210 16204
rect 14826 16192 14832 16204
rect 14884 16192 14890 16244
rect 10796 16164 10824 16192
rect 11517 16167 11575 16173
rect 11517 16164 11529 16167
rect 10060 16136 10732 16164
rect 10796 16136 11529 16164
rect 3375 16068 3832 16096
rect 3375 16065 3387 16068
rect 3329 16059 3387 16065
rect 3878 16056 3884 16108
rect 3936 16096 3942 16108
rect 3936 16068 3981 16096
rect 3936 16056 3942 16068
rect 5166 16056 5172 16108
rect 5224 16096 5230 16108
rect 5721 16099 5779 16105
rect 5721 16096 5733 16099
rect 5224 16068 5733 16096
rect 5224 16056 5230 16068
rect 5721 16065 5733 16068
rect 5767 16065 5779 16099
rect 5721 16059 5779 16065
rect 6362 16056 6368 16108
rect 6420 16096 6426 16108
rect 6825 16099 6883 16105
rect 6825 16096 6837 16099
rect 6420 16068 6837 16096
rect 6420 16056 6426 16068
rect 6825 16065 6837 16068
rect 6871 16065 6883 16099
rect 7834 16096 7840 16108
rect 7795 16068 7840 16096
rect 6825 16059 6883 16065
rect 7834 16056 7840 16068
rect 7892 16056 7898 16108
rect 10042 16096 10048 16108
rect 10003 16068 10048 16096
rect 10042 16056 10048 16068
rect 10100 16056 10106 16108
rect 10704 16105 10732 16136
rect 11517 16133 11529 16136
rect 11563 16133 11575 16167
rect 11517 16127 11575 16133
rect 11606 16124 11612 16176
rect 11664 16164 11670 16176
rect 15378 16164 15384 16176
rect 11664 16136 15384 16164
rect 11664 16124 11670 16136
rect 15378 16124 15384 16136
rect 15436 16124 15442 16176
rect 19429 16167 19487 16173
rect 19429 16164 19441 16167
rect 19260 16136 19441 16164
rect 10689 16099 10747 16105
rect 10689 16065 10701 16099
rect 10735 16065 10747 16099
rect 12066 16096 12072 16108
rect 10689 16059 10747 16065
rect 10980 16068 12072 16096
rect 3970 15988 3976 16040
rect 4028 16028 4034 16040
rect 4893 16031 4951 16037
rect 4893 16028 4905 16031
rect 4028 16000 4905 16028
rect 4028 15988 4034 16000
rect 4893 15997 4905 16000
rect 4939 16028 4951 16031
rect 5258 16028 5264 16040
rect 4939 16000 5264 16028
rect 4939 15997 4951 16000
rect 4893 15991 4951 15997
rect 5258 15988 5264 16000
rect 5316 15988 5322 16040
rect 5537 16031 5595 16037
rect 5537 15997 5549 16031
rect 5583 15997 5595 16031
rect 5537 15991 5595 15997
rect 5629 16031 5687 16037
rect 5629 15997 5641 16031
rect 5675 16028 5687 16031
rect 5994 16028 6000 16040
rect 5675 16000 6000 16028
rect 5675 15997 5687 16000
rect 5629 15991 5687 15997
rect 5552 15960 5580 15991
rect 5994 15988 6000 16000
rect 6052 15988 6058 16040
rect 6733 16031 6791 16037
rect 6733 15997 6745 16031
rect 6779 15997 6791 16031
rect 6733 15991 6791 15997
rect 7653 16031 7711 16037
rect 7653 15997 7665 16031
rect 7699 16028 7711 16031
rect 10502 16028 10508 16040
rect 7699 16000 9674 16028
rect 10463 16000 10508 16028
rect 7699 15997 7711 16000
rect 7653 15991 7711 15997
rect 5810 15960 5816 15972
rect 5552 15932 5816 15960
rect 5810 15920 5816 15932
rect 5868 15920 5874 15972
rect 6748 15960 6776 15991
rect 6914 15960 6920 15972
rect 6748 15932 6920 15960
rect 6914 15920 6920 15932
rect 6972 15920 6978 15972
rect 7285 15963 7343 15969
rect 7285 15929 7297 15963
rect 7331 15960 7343 15963
rect 8662 15960 8668 15972
rect 7331 15932 8668 15960
rect 7331 15929 7343 15932
rect 7285 15923 7343 15929
rect 8662 15920 8668 15932
rect 8720 15920 8726 15972
rect 8849 15963 8907 15969
rect 8849 15929 8861 15963
rect 8895 15960 8907 15963
rect 9122 15960 9128 15972
rect 8895 15932 9128 15960
rect 8895 15929 8907 15932
rect 8849 15923 8907 15929
rect 9122 15920 9128 15932
rect 9180 15920 9186 15972
rect 9646 15960 9674 16000
rect 10502 15988 10508 16000
rect 10560 15988 10566 16040
rect 10980 16028 11008 16068
rect 12066 16056 12072 16068
rect 12124 16056 12130 16108
rect 12526 16056 12532 16108
rect 12584 16096 12590 16108
rect 13274 16099 13332 16105
rect 13274 16096 13286 16099
rect 12584 16068 13286 16096
rect 12584 16056 12590 16068
rect 13274 16065 13286 16068
rect 13320 16065 13332 16099
rect 13274 16059 13332 16065
rect 14941 16099 14999 16105
rect 14941 16065 14953 16099
rect 14987 16096 14999 16099
rect 15102 16096 15108 16108
rect 14987 16068 15108 16096
rect 14987 16065 14999 16068
rect 14941 16059 14999 16065
rect 15102 16056 15108 16068
rect 15160 16096 15166 16108
rect 15473 16099 15531 16105
rect 15473 16096 15485 16099
rect 15160 16068 15485 16096
rect 15160 16056 15166 16068
rect 15473 16065 15485 16068
rect 15519 16065 15531 16099
rect 15473 16059 15531 16065
rect 18966 16056 18972 16108
rect 19024 16105 19030 16108
rect 19260 16105 19288 16136
rect 19429 16133 19441 16136
rect 19475 16164 19487 16167
rect 19475 16136 21496 16164
rect 19475 16133 19487 16136
rect 19429 16127 19487 16133
rect 21468 16108 21496 16136
rect 19024 16096 19036 16105
rect 19245 16099 19303 16105
rect 19024 16068 19069 16096
rect 19024 16059 19036 16068
rect 19245 16065 19257 16099
rect 19291 16065 19303 16099
rect 19245 16059 19303 16065
rect 19024 16056 19030 16059
rect 21174 16056 21180 16108
rect 21232 16105 21238 16108
rect 21232 16096 21244 16105
rect 21450 16096 21456 16108
rect 21232 16068 21277 16096
rect 21411 16068 21456 16096
rect 21232 16059 21244 16068
rect 21232 16056 21238 16059
rect 21450 16056 21456 16068
rect 21508 16056 21514 16108
rect 11146 16028 11152 16040
rect 10612 16000 11008 16028
rect 11107 16000 11152 16028
rect 9766 15960 9772 15972
rect 9646 15932 9772 15960
rect 9766 15920 9772 15932
rect 9824 15960 9830 15972
rect 10612 15960 10640 16000
rect 11146 15988 11152 16000
rect 11204 15988 11210 16040
rect 13541 16031 13599 16037
rect 13541 15997 13553 16031
rect 13587 16028 13599 16031
rect 15194 16028 15200 16040
rect 13587 16000 13768 16028
rect 15155 16000 15200 16028
rect 13587 15997 13599 16000
rect 13541 15991 13599 15997
rect 9824 15932 10640 15960
rect 9824 15920 9830 15932
rect 10778 15920 10784 15972
rect 10836 15960 10842 15972
rect 12161 15963 12219 15969
rect 12161 15960 12173 15963
rect 10836 15932 12173 15960
rect 10836 15920 10842 15932
rect 12161 15929 12173 15932
rect 12207 15960 12219 15963
rect 12342 15960 12348 15972
rect 12207 15932 12348 15960
rect 12207 15929 12219 15932
rect 12161 15923 12219 15929
rect 12342 15920 12348 15932
rect 12400 15920 12406 15972
rect 13740 15904 13768 16000
rect 15194 15988 15200 16000
rect 15252 16028 15258 16040
rect 15289 16031 15347 16037
rect 15289 16028 15301 16031
rect 15252 16000 15301 16028
rect 15252 15988 15258 16000
rect 15289 15997 15301 16000
rect 15335 15997 15347 16031
rect 15289 15991 15347 15997
rect 3878 15852 3884 15904
rect 3936 15892 3942 15904
rect 4982 15892 4988 15904
rect 3936 15864 4988 15892
rect 3936 15852 3942 15864
rect 4982 15852 4988 15864
rect 5040 15852 5046 15904
rect 6362 15892 6368 15904
rect 6323 15864 6368 15892
rect 6362 15852 6368 15864
rect 6420 15852 6426 15904
rect 7926 15852 7932 15904
rect 7984 15892 7990 15904
rect 8205 15895 8263 15901
rect 8205 15892 8217 15895
rect 7984 15864 8217 15892
rect 7984 15852 7990 15864
rect 8205 15861 8217 15864
rect 8251 15861 8263 15895
rect 8205 15855 8263 15861
rect 8294 15852 8300 15904
rect 8352 15892 8358 15904
rect 9214 15892 9220 15904
rect 8352 15864 8397 15892
rect 9175 15864 9220 15892
rect 8352 15852 8358 15864
rect 9214 15852 9220 15864
rect 9272 15852 9278 15904
rect 9306 15852 9312 15904
rect 9364 15892 9370 15904
rect 9401 15895 9459 15901
rect 9401 15892 9413 15895
rect 9364 15864 9413 15892
rect 9364 15852 9370 15864
rect 9401 15861 9413 15864
rect 9447 15861 9459 15895
rect 9401 15855 9459 15861
rect 9950 15852 9956 15904
rect 10008 15892 10014 15904
rect 10137 15895 10195 15901
rect 10137 15892 10149 15895
rect 10008 15864 10149 15892
rect 10008 15852 10014 15864
rect 10137 15861 10149 15864
rect 10183 15892 10195 15895
rect 11606 15892 11612 15904
rect 10183 15864 11612 15892
rect 10183 15861 10195 15864
rect 10137 15855 10195 15861
rect 11606 15852 11612 15864
rect 11664 15852 11670 15904
rect 13722 15892 13728 15904
rect 13683 15864 13728 15892
rect 13722 15852 13728 15864
rect 13780 15852 13786 15904
rect 13817 15895 13875 15901
rect 13817 15861 13829 15895
rect 13863 15892 13875 15895
rect 14826 15892 14832 15904
rect 13863 15864 14832 15892
rect 13863 15861 13875 15864
rect 13817 15855 13875 15861
rect 14826 15852 14832 15864
rect 14884 15852 14890 15904
rect 15838 15852 15844 15904
rect 15896 15892 15902 15904
rect 17865 15895 17923 15901
rect 17865 15892 17877 15895
rect 15896 15864 17877 15892
rect 15896 15852 15902 15864
rect 17865 15861 17877 15864
rect 17911 15861 17923 15895
rect 20070 15892 20076 15904
rect 20031 15864 20076 15892
rect 17865 15855 17923 15861
rect 20070 15852 20076 15864
rect 20128 15852 20134 15904
rect 1104 15802 21896 15824
rect 1104 15750 3549 15802
rect 3601 15750 3613 15802
rect 3665 15750 3677 15802
rect 3729 15750 3741 15802
rect 3793 15750 3805 15802
rect 3857 15750 8747 15802
rect 8799 15750 8811 15802
rect 8863 15750 8875 15802
rect 8927 15750 8939 15802
rect 8991 15750 9003 15802
rect 9055 15750 13945 15802
rect 13997 15750 14009 15802
rect 14061 15750 14073 15802
rect 14125 15750 14137 15802
rect 14189 15750 14201 15802
rect 14253 15750 19143 15802
rect 19195 15750 19207 15802
rect 19259 15750 19271 15802
rect 19323 15750 19335 15802
rect 19387 15750 19399 15802
rect 19451 15750 21896 15802
rect 1104 15728 21896 15750
rect 1946 15688 1952 15700
rect 1907 15660 1952 15688
rect 1946 15648 1952 15660
rect 2004 15648 2010 15700
rect 2314 15688 2320 15700
rect 2275 15660 2320 15688
rect 2314 15648 2320 15660
rect 2372 15648 2378 15700
rect 2682 15688 2688 15700
rect 2643 15660 2688 15688
rect 2682 15648 2688 15660
rect 2740 15648 2746 15700
rect 3326 15648 3332 15700
rect 3384 15688 3390 15700
rect 3605 15691 3663 15697
rect 3605 15688 3617 15691
rect 3384 15660 3617 15688
rect 3384 15648 3390 15660
rect 3605 15657 3617 15660
rect 3651 15688 3663 15691
rect 4062 15688 4068 15700
rect 3651 15660 4068 15688
rect 3651 15657 3663 15660
rect 3605 15651 3663 15657
rect 4062 15648 4068 15660
rect 4120 15688 4126 15700
rect 4798 15688 4804 15700
rect 4120 15660 4804 15688
rect 4120 15648 4126 15660
rect 4798 15648 4804 15660
rect 4856 15648 4862 15700
rect 5166 15688 5172 15700
rect 5127 15660 5172 15688
rect 5166 15648 5172 15660
rect 5224 15648 5230 15700
rect 5994 15688 6000 15700
rect 5955 15660 6000 15688
rect 5994 15648 6000 15660
rect 6052 15648 6058 15700
rect 6086 15648 6092 15700
rect 6144 15688 6150 15700
rect 6144 15660 6189 15688
rect 6144 15648 6150 15660
rect 7834 15648 7840 15700
rect 7892 15688 7898 15700
rect 8941 15691 8999 15697
rect 8941 15688 8953 15691
rect 7892 15660 8953 15688
rect 7892 15648 7898 15660
rect 8941 15657 8953 15660
rect 8987 15657 8999 15691
rect 8941 15651 8999 15657
rect 9122 15648 9128 15700
rect 9180 15688 9186 15700
rect 9953 15691 10011 15697
rect 9953 15688 9965 15691
rect 9180 15660 9965 15688
rect 9180 15648 9186 15660
rect 9953 15657 9965 15660
rect 9999 15657 10011 15691
rect 10226 15688 10232 15700
rect 10187 15660 10232 15688
rect 9953 15651 10011 15657
rect 10226 15648 10232 15660
rect 10284 15648 10290 15700
rect 19886 15688 19892 15700
rect 12406 15660 13492 15688
rect 3878 15620 3884 15632
rect 2516 15592 3884 15620
rect 2516 15493 2544 15592
rect 3878 15580 3884 15592
rect 3936 15580 3942 15632
rect 8110 15620 8116 15632
rect 4632 15592 8116 15620
rect 4246 15552 4252 15564
rect 2746 15524 4252 15552
rect 2133 15487 2191 15493
rect 2133 15453 2145 15487
rect 2179 15453 2191 15487
rect 2133 15447 2191 15453
rect 2501 15487 2559 15493
rect 2501 15453 2513 15487
rect 2547 15453 2559 15487
rect 2501 15447 2559 15453
rect 2148 15416 2176 15447
rect 2746 15416 2774 15524
rect 4246 15512 4252 15524
rect 4304 15512 4310 15564
rect 4632 15561 4660 15592
rect 5460 15561 5488 15592
rect 8110 15580 8116 15592
rect 8168 15580 8174 15632
rect 8389 15623 8447 15629
rect 8389 15589 8401 15623
rect 8435 15620 8447 15623
rect 8478 15620 8484 15632
rect 8435 15592 8484 15620
rect 8435 15589 8447 15592
rect 8389 15583 8447 15589
rect 8478 15580 8484 15592
rect 8536 15580 8542 15632
rect 12406 15620 12434 15660
rect 10888 15592 12434 15620
rect 13464 15620 13492 15660
rect 14568 15660 19892 15688
rect 14568 15620 14596 15660
rect 19886 15648 19892 15660
rect 19944 15648 19950 15700
rect 15838 15620 15844 15632
rect 13464 15592 14596 15620
rect 15799 15592 15844 15620
rect 4341 15555 4399 15561
rect 4341 15521 4353 15555
rect 4387 15552 4399 15555
rect 4617 15555 4675 15561
rect 4387 15524 4568 15552
rect 4387 15521 4399 15524
rect 4341 15515 4399 15521
rect 2869 15487 2927 15493
rect 2869 15453 2881 15487
rect 2915 15484 2927 15487
rect 4540 15484 4568 15524
rect 4617 15521 4629 15555
rect 4663 15521 4675 15555
rect 4617 15515 4675 15521
rect 5445 15555 5503 15561
rect 5445 15521 5457 15555
rect 5491 15521 5503 15555
rect 5445 15515 5503 15521
rect 5626 15512 5632 15564
rect 5684 15552 5690 15564
rect 6549 15555 6607 15561
rect 6549 15552 6561 15555
rect 5684 15524 6561 15552
rect 5684 15512 5690 15524
rect 6549 15521 6561 15524
rect 6595 15521 6607 15555
rect 6549 15515 6607 15521
rect 6733 15555 6791 15561
rect 6733 15521 6745 15555
rect 6779 15552 6791 15555
rect 6914 15552 6920 15564
rect 6779 15524 6920 15552
rect 6779 15521 6791 15524
rect 6733 15515 6791 15521
rect 6914 15512 6920 15524
rect 6972 15512 6978 15564
rect 7742 15552 7748 15564
rect 7703 15524 7748 15552
rect 7742 15512 7748 15524
rect 7800 15512 7806 15564
rect 7926 15552 7932 15564
rect 7887 15524 7932 15552
rect 7926 15512 7932 15524
rect 7984 15512 7990 15564
rect 9398 15552 9404 15564
rect 9359 15524 9404 15552
rect 9398 15512 9404 15524
rect 9456 15512 9462 15564
rect 9493 15555 9551 15561
rect 9493 15521 9505 15555
rect 9539 15552 9551 15555
rect 9950 15552 9956 15564
rect 9539 15524 9956 15552
rect 9539 15521 9551 15524
rect 9493 15515 9551 15521
rect 4706 15484 4712 15496
rect 2915 15456 4476 15484
rect 4540 15456 4712 15484
rect 2915 15453 2927 15456
rect 2869 15447 2927 15453
rect 2148 15388 2774 15416
rect 3234 15376 3240 15428
rect 3292 15416 3298 15428
rect 3881 15419 3939 15425
rect 3881 15416 3893 15419
rect 3292 15388 3893 15416
rect 3292 15376 3298 15388
rect 3881 15385 3893 15388
rect 3927 15385 3939 15419
rect 4448 15416 4476 15456
rect 4706 15444 4712 15456
rect 4764 15444 4770 15496
rect 4798 15444 4804 15496
rect 4856 15484 4862 15496
rect 4856 15456 4901 15484
rect 4856 15444 4862 15456
rect 5534 15444 5540 15496
rect 5592 15484 5598 15496
rect 6457 15487 6515 15493
rect 6457 15484 6469 15487
rect 5592 15456 6469 15484
rect 5592 15444 5598 15456
rect 6457 15453 6469 15456
rect 6503 15453 6515 15487
rect 9508 15484 9536 15515
rect 9950 15512 9956 15524
rect 10008 15512 10014 15564
rect 10686 15552 10692 15564
rect 10520 15524 10692 15552
rect 6457 15447 6515 15453
rect 7484 15456 9536 15484
rect 4614 15416 4620 15428
rect 4448 15388 4620 15416
rect 3881 15379 3939 15385
rect 4614 15376 4620 15388
rect 4672 15376 4678 15428
rect 4724 15416 4752 15444
rect 4724 15388 5212 15416
rect 3418 15348 3424 15360
rect 3379 15320 3424 15348
rect 3418 15308 3424 15320
rect 3476 15308 3482 15360
rect 4062 15308 4068 15360
rect 4120 15348 4126 15360
rect 4157 15351 4215 15357
rect 4157 15348 4169 15351
rect 4120 15320 4169 15348
rect 4120 15308 4126 15320
rect 4157 15317 4169 15320
rect 4203 15317 4215 15351
rect 4157 15311 4215 15317
rect 4338 15308 4344 15360
rect 4396 15348 4402 15360
rect 4709 15351 4767 15357
rect 4709 15348 4721 15351
rect 4396 15320 4721 15348
rect 4396 15308 4402 15320
rect 4709 15317 4721 15320
rect 4755 15317 4767 15351
rect 5184 15348 5212 15388
rect 5258 15376 5264 15428
rect 5316 15416 5322 15428
rect 5629 15419 5687 15425
rect 5629 15416 5641 15419
rect 5316 15388 5641 15416
rect 5316 15376 5322 15388
rect 5629 15385 5641 15388
rect 5675 15385 5687 15419
rect 5629 15379 5687 15385
rect 5810 15376 5816 15428
rect 5868 15416 5874 15428
rect 7484 15416 7512 15456
rect 5868 15388 7512 15416
rect 7561 15419 7619 15425
rect 5868 15376 5874 15388
rect 7561 15385 7573 15419
rect 7607 15416 7619 15419
rect 8202 15416 8208 15428
rect 7607 15388 8208 15416
rect 7607 15385 7619 15388
rect 7561 15379 7619 15385
rect 8202 15376 8208 15388
rect 8260 15376 8266 15428
rect 8754 15376 8760 15428
rect 8812 15416 8818 15428
rect 9769 15419 9827 15425
rect 9769 15416 9781 15419
rect 8812 15388 9781 15416
rect 8812 15376 8818 15388
rect 9769 15385 9781 15388
rect 9815 15416 9827 15419
rect 10520 15416 10548 15524
rect 10686 15512 10692 15524
rect 10744 15512 10750 15564
rect 10888 15561 10916 15592
rect 15838 15580 15844 15592
rect 15896 15580 15902 15632
rect 10873 15555 10931 15561
rect 10873 15521 10885 15555
rect 10919 15521 10931 15555
rect 15856 15552 15884 15580
rect 10873 15515 10931 15521
rect 15387 15524 15884 15552
rect 10597 15487 10655 15493
rect 10597 15453 10609 15487
rect 10643 15484 10655 15487
rect 11146 15484 11152 15496
rect 10643 15456 11152 15484
rect 10643 15453 10655 15456
rect 10597 15447 10655 15453
rect 11146 15444 11152 15456
rect 11204 15444 11210 15496
rect 13357 15487 13415 15493
rect 13357 15453 13369 15487
rect 13403 15484 13415 15487
rect 13722 15484 13728 15496
rect 13403 15456 13728 15484
rect 13403 15453 13415 15456
rect 13357 15447 13415 15453
rect 13722 15444 13728 15456
rect 13780 15444 13786 15496
rect 14918 15444 14924 15496
rect 14976 15484 14982 15496
rect 15217 15487 15275 15493
rect 15217 15484 15229 15487
rect 14976 15456 15229 15484
rect 14976 15444 14982 15456
rect 15217 15453 15229 15456
rect 15263 15484 15275 15487
rect 15387 15484 15415 15524
rect 15263 15456 15415 15484
rect 15473 15487 15531 15493
rect 15263 15453 15275 15456
rect 15217 15447 15275 15453
rect 15473 15453 15485 15487
rect 15519 15484 15531 15487
rect 15657 15487 15715 15493
rect 15657 15484 15669 15487
rect 15519 15456 15669 15484
rect 15519 15453 15531 15456
rect 15473 15447 15531 15453
rect 15657 15453 15669 15456
rect 15703 15484 15715 15487
rect 16117 15487 16175 15493
rect 16117 15484 16129 15487
rect 15703 15456 16129 15484
rect 15703 15453 15715 15456
rect 15657 15447 15715 15453
rect 16117 15453 16129 15456
rect 16163 15484 16175 15487
rect 17589 15487 17647 15493
rect 17589 15484 17601 15487
rect 16163 15456 17601 15484
rect 16163 15453 16175 15456
rect 16117 15447 16175 15453
rect 17589 15453 17601 15456
rect 17635 15453 17647 15487
rect 17589 15447 17647 15453
rect 19889 15487 19947 15493
rect 19889 15453 19901 15487
rect 19935 15484 19947 15487
rect 20073 15487 20131 15493
rect 20073 15484 20085 15487
rect 19935 15456 20085 15484
rect 19935 15453 19947 15456
rect 19889 15447 19947 15453
rect 20073 15453 20085 15456
rect 20119 15484 20131 15487
rect 20714 15484 20720 15496
rect 20119 15456 20720 15484
rect 20119 15453 20131 15456
rect 20073 15447 20131 15453
rect 9815 15388 10548 15416
rect 13112 15419 13170 15425
rect 9815 15385 9827 15388
rect 9769 15379 9827 15385
rect 13112 15385 13124 15419
rect 13158 15416 13170 15419
rect 14642 15416 14648 15428
rect 13158 15388 14648 15416
rect 13158 15385 13170 15388
rect 13112 15379 13170 15385
rect 14642 15376 14648 15388
rect 14700 15376 14706 15428
rect 15378 15376 15384 15428
rect 15436 15416 15442 15428
rect 15488 15416 15516 15447
rect 20714 15444 20720 15456
rect 20772 15484 20778 15496
rect 21450 15484 21456 15496
rect 20772 15456 21456 15484
rect 20772 15444 20778 15456
rect 21450 15444 21456 15456
rect 21508 15484 21514 15496
rect 21545 15487 21603 15493
rect 21545 15484 21557 15487
rect 21508 15456 21557 15484
rect 21508 15444 21514 15456
rect 21545 15453 21557 15456
rect 21591 15453 21603 15487
rect 21545 15447 21603 15453
rect 15436 15388 15516 15416
rect 15436 15376 15442 15388
rect 15562 15376 15568 15428
rect 15620 15416 15626 15428
rect 16362 15419 16420 15425
rect 16362 15416 16374 15419
rect 15620 15388 16374 15416
rect 15620 15376 15626 15388
rect 16362 15385 16374 15388
rect 16408 15385 16420 15419
rect 21266 15416 21272 15428
rect 21324 15425 21330 15428
rect 21236 15388 21272 15416
rect 16362 15379 16420 15385
rect 21266 15376 21272 15388
rect 21324 15379 21336 15425
rect 21324 15376 21330 15379
rect 5537 15351 5595 15357
rect 5537 15348 5549 15351
rect 5184 15320 5549 15348
rect 4709 15311 4767 15317
rect 5537 15317 5549 15320
rect 5583 15348 5595 15351
rect 6362 15348 6368 15360
rect 5583 15320 6368 15348
rect 5583 15317 5595 15320
rect 5537 15311 5595 15317
rect 6362 15308 6368 15320
rect 6420 15308 6426 15360
rect 7006 15308 7012 15360
rect 7064 15348 7070 15360
rect 8021 15351 8079 15357
rect 8021 15348 8033 15351
rect 7064 15320 8033 15348
rect 7064 15308 7070 15320
rect 8021 15317 8033 15320
rect 8067 15317 8079 15351
rect 8021 15311 8079 15317
rect 9309 15351 9367 15357
rect 9309 15317 9321 15351
rect 9355 15348 9367 15351
rect 9398 15348 9404 15360
rect 9355 15320 9404 15348
rect 9355 15317 9367 15320
rect 9309 15311 9367 15317
rect 9398 15308 9404 15320
rect 9456 15308 9462 15360
rect 10686 15308 10692 15360
rect 10744 15348 10750 15360
rect 11054 15348 11060 15360
rect 10744 15320 10789 15348
rect 11015 15320 11060 15348
rect 10744 15308 10750 15320
rect 11054 15308 11060 15320
rect 11112 15308 11118 15360
rect 11977 15351 12035 15357
rect 11977 15317 11989 15351
rect 12023 15348 12035 15351
rect 12526 15348 12532 15360
rect 12023 15320 12532 15348
rect 12023 15317 12035 15320
rect 11977 15311 12035 15317
rect 12526 15308 12532 15320
rect 12584 15308 12590 15360
rect 13541 15351 13599 15357
rect 13541 15317 13553 15351
rect 13587 15348 13599 15351
rect 13722 15348 13728 15360
rect 13587 15320 13728 15348
rect 13587 15317 13599 15320
rect 13541 15311 13599 15317
rect 13722 15308 13728 15320
rect 13780 15308 13786 15360
rect 13814 15308 13820 15360
rect 13872 15348 13878 15360
rect 14093 15351 14151 15357
rect 14093 15348 14105 15351
rect 13872 15320 14105 15348
rect 13872 15308 13878 15320
rect 14093 15317 14105 15320
rect 14139 15317 14151 15351
rect 14093 15311 14151 15317
rect 14734 15308 14740 15360
rect 14792 15348 14798 15360
rect 15580 15348 15608 15376
rect 17494 15348 17500 15360
rect 14792 15320 15608 15348
rect 17455 15320 17500 15348
rect 14792 15308 14798 15320
rect 17494 15308 17500 15320
rect 17552 15308 17558 15360
rect 20165 15351 20223 15357
rect 20165 15317 20177 15351
rect 20211 15348 20223 15351
rect 20530 15348 20536 15360
rect 20211 15320 20536 15348
rect 20211 15317 20223 15320
rect 20165 15311 20223 15317
rect 20530 15308 20536 15320
rect 20588 15308 20594 15360
rect 1104 15258 22056 15280
rect 1104 15206 6148 15258
rect 6200 15206 6212 15258
rect 6264 15206 6276 15258
rect 6328 15206 6340 15258
rect 6392 15206 6404 15258
rect 6456 15206 11346 15258
rect 11398 15206 11410 15258
rect 11462 15206 11474 15258
rect 11526 15206 11538 15258
rect 11590 15206 11602 15258
rect 11654 15206 16544 15258
rect 16596 15206 16608 15258
rect 16660 15206 16672 15258
rect 16724 15206 16736 15258
rect 16788 15206 16800 15258
rect 16852 15206 21742 15258
rect 21794 15206 21806 15258
rect 21858 15206 21870 15258
rect 21922 15206 21934 15258
rect 21986 15206 21998 15258
rect 22050 15206 22056 15258
rect 1104 15184 22056 15206
rect 1854 15104 1860 15156
rect 1912 15144 1918 15156
rect 1949 15147 2007 15153
rect 1949 15144 1961 15147
rect 1912 15116 1961 15144
rect 1912 15104 1918 15116
rect 1949 15113 1961 15116
rect 1995 15113 2007 15147
rect 1949 15107 2007 15113
rect 2590 15104 2596 15156
rect 2648 15144 2654 15156
rect 2685 15147 2743 15153
rect 2685 15144 2697 15147
rect 2648 15116 2697 15144
rect 2648 15104 2654 15116
rect 2685 15113 2697 15116
rect 2731 15113 2743 15147
rect 3326 15144 3332 15156
rect 3287 15116 3332 15144
rect 2685 15107 2743 15113
rect 3326 15104 3332 15116
rect 3384 15104 3390 15156
rect 3418 15104 3424 15156
rect 3476 15144 3482 15156
rect 4065 15147 4123 15153
rect 4065 15144 4077 15147
rect 3476 15116 4077 15144
rect 3476 15104 3482 15116
rect 4065 15113 4077 15116
rect 4111 15113 4123 15147
rect 4065 15107 4123 15113
rect 4157 15147 4215 15153
rect 4157 15113 4169 15147
rect 4203 15144 4215 15147
rect 4430 15144 4436 15156
rect 4203 15116 4436 15144
rect 4203 15113 4215 15116
rect 4157 15107 4215 15113
rect 4430 15104 4436 15116
rect 4488 15104 4494 15156
rect 4816 15116 5028 15144
rect 2501 15079 2559 15085
rect 2501 15045 2513 15079
rect 2547 15076 2559 15079
rect 4338 15076 4344 15088
rect 2547 15048 2774 15076
rect 2547 15045 2559 15048
rect 2501 15039 2559 15045
rect 2130 15008 2136 15020
rect 2091 14980 2136 15008
rect 2130 14968 2136 14980
rect 2188 14968 2194 15020
rect 2746 14940 2774 15048
rect 2884 15048 4344 15076
rect 2884 15017 2912 15048
rect 4338 15036 4344 15048
rect 4396 15036 4402 15088
rect 2869 15011 2927 15017
rect 2869 14977 2881 15011
rect 2915 14977 2927 15011
rect 3237 15011 3295 15017
rect 3237 15008 3249 15011
rect 2869 14971 2927 14977
rect 2976 14980 3249 15008
rect 2976 14940 3004 14980
rect 3237 14977 3249 14980
rect 3283 15008 3295 15011
rect 3970 15008 3976 15020
rect 3283 14980 3976 15008
rect 3283 14977 3295 14980
rect 3237 14971 3295 14977
rect 3970 14968 3976 14980
rect 4028 14968 4034 15020
rect 4062 14968 4068 15020
rect 4120 15008 4126 15020
rect 4448 15008 4476 15104
rect 4816 15076 4844 15116
rect 4724 15048 4844 15076
rect 4893 15079 4951 15085
rect 4724 15008 4752 15048
rect 4893 15045 4905 15079
rect 4939 15045 4951 15079
rect 5000 15076 5028 15116
rect 5626 15104 5632 15156
rect 5684 15144 5690 15156
rect 5905 15147 5963 15153
rect 5905 15144 5917 15147
rect 5684 15116 5917 15144
rect 5684 15104 5690 15116
rect 5905 15113 5917 15116
rect 5951 15113 5963 15147
rect 5905 15107 5963 15113
rect 7098 15104 7104 15156
rect 7156 15104 7162 15156
rect 7466 15144 7472 15156
rect 7427 15116 7472 15144
rect 7466 15104 7472 15116
rect 7524 15104 7530 15156
rect 7558 15104 7564 15156
rect 7616 15144 7622 15156
rect 7837 15147 7895 15153
rect 7837 15144 7849 15147
rect 7616 15116 7849 15144
rect 7616 15104 7622 15116
rect 7837 15113 7849 15116
rect 7883 15113 7895 15147
rect 8202 15144 8208 15156
rect 8163 15116 8208 15144
rect 7837 15107 7895 15113
rect 8202 15104 8208 15116
rect 8260 15104 8266 15156
rect 8662 15104 8668 15156
rect 8720 15144 8726 15156
rect 8941 15147 8999 15153
rect 8941 15144 8953 15147
rect 8720 15116 8953 15144
rect 8720 15104 8726 15116
rect 8941 15113 8953 15116
rect 8987 15113 8999 15147
rect 8941 15107 8999 15113
rect 9033 15147 9091 15153
rect 9033 15113 9045 15147
rect 9079 15144 9091 15147
rect 9122 15144 9128 15156
rect 9079 15116 9128 15144
rect 9079 15113 9091 15116
rect 9033 15107 9091 15113
rect 7116 15076 7144 15104
rect 7653 15079 7711 15085
rect 7653 15076 7665 15079
rect 5000 15048 5488 15076
rect 7116 15048 7665 15076
rect 4893 15039 4951 15045
rect 4120 14980 4476 15008
rect 4632 14980 4752 15008
rect 4120 14968 4126 14980
rect 2746 14912 3004 14940
rect 3145 14943 3203 14949
rect 3145 14909 3157 14943
rect 3191 14909 3203 14943
rect 3878 14940 3884 14952
rect 3839 14912 3884 14940
rect 3145 14903 3203 14909
rect 3160 14872 3188 14903
rect 3878 14900 3884 14912
rect 3936 14940 3942 14952
rect 4632 14940 4660 14980
rect 4798 14968 4804 15020
rect 4856 15008 4862 15020
rect 4908 15008 4936 15039
rect 4856 14980 4936 15008
rect 4985 15011 5043 15017
rect 4856 14968 4862 14980
rect 4985 14977 4997 15011
rect 5031 14977 5043 15011
rect 5460 15008 5488 15048
rect 7653 15045 7665 15048
rect 7699 15076 7711 15079
rect 8297 15079 8355 15085
rect 8297 15076 8309 15079
rect 7699 15048 8309 15076
rect 7699 15045 7711 15048
rect 7653 15039 7711 15045
rect 8297 15045 8309 15048
rect 8343 15045 8355 15079
rect 8297 15039 8355 15045
rect 8386 15036 8392 15088
rect 8444 15076 8450 15088
rect 9048 15076 9076 15107
rect 9122 15104 9128 15116
rect 9180 15104 9186 15156
rect 9493 15147 9551 15153
rect 9493 15113 9505 15147
rect 9539 15144 9551 15147
rect 9674 15144 9680 15156
rect 9539 15116 9680 15144
rect 9539 15113 9551 15116
rect 9493 15107 9551 15113
rect 9674 15104 9680 15116
rect 9732 15104 9738 15156
rect 10597 15147 10655 15153
rect 10597 15113 10609 15147
rect 10643 15144 10655 15147
rect 10686 15144 10692 15156
rect 10643 15116 10692 15144
rect 10643 15113 10655 15116
rect 10597 15107 10655 15113
rect 10686 15104 10692 15116
rect 10744 15104 10750 15156
rect 10962 15144 10968 15156
rect 10796 15116 10968 15144
rect 10796 15076 10824 15116
rect 10962 15104 10968 15116
rect 11020 15104 11026 15156
rect 11057 15147 11115 15153
rect 11057 15113 11069 15147
rect 11103 15144 11115 15147
rect 11609 15147 11667 15153
rect 11609 15144 11621 15147
rect 11103 15116 11621 15144
rect 11103 15113 11115 15116
rect 11057 15107 11115 15113
rect 11609 15113 11621 15116
rect 11655 15144 11667 15147
rect 12618 15144 12624 15156
rect 11655 15116 12624 15144
rect 11655 15113 11667 15116
rect 11609 15107 11667 15113
rect 12618 15104 12624 15116
rect 12676 15104 12682 15156
rect 13909 15147 13967 15153
rect 13909 15113 13921 15147
rect 13955 15144 13967 15147
rect 14550 15144 14556 15156
rect 13955 15116 14556 15144
rect 13955 15113 13967 15116
rect 13909 15107 13967 15113
rect 14550 15104 14556 15116
rect 14608 15104 14614 15156
rect 16390 15104 16396 15156
rect 16448 15144 16454 15156
rect 16669 15147 16727 15153
rect 16669 15144 16681 15147
rect 16448 15116 16681 15144
rect 16448 15104 16454 15116
rect 16669 15113 16681 15116
rect 16715 15113 16727 15147
rect 20070 15144 20076 15156
rect 16669 15107 16727 15113
rect 17880 15116 20076 15144
rect 12894 15076 12900 15088
rect 8444 15048 9076 15076
rect 9692 15048 10824 15076
rect 10888 15048 12900 15076
rect 8444 15036 8450 15048
rect 5460 14980 5672 15008
rect 4985 14971 5043 14977
rect 3936 14912 4660 14940
rect 4709 14943 4767 14949
rect 3936 14900 3942 14912
rect 4709 14909 4721 14943
rect 4755 14909 4767 14943
rect 4709 14903 4767 14909
rect 4525 14875 4583 14881
rect 3160 14844 3280 14872
rect 3252 14816 3280 14844
rect 4525 14841 4537 14875
rect 4571 14872 4583 14875
rect 4614 14872 4620 14884
rect 4571 14844 4620 14872
rect 4571 14841 4583 14844
rect 4525 14835 4583 14841
rect 4614 14832 4620 14844
rect 4672 14832 4678 14884
rect 4724 14872 4752 14903
rect 4798 14872 4804 14884
rect 4724 14844 4804 14872
rect 4798 14832 4804 14844
rect 4856 14832 4862 14884
rect 3234 14764 3240 14816
rect 3292 14764 3298 14816
rect 3697 14807 3755 14813
rect 3697 14773 3709 14807
rect 3743 14804 3755 14807
rect 4062 14804 4068 14816
rect 3743 14776 4068 14804
rect 3743 14773 3755 14776
rect 3697 14767 3755 14773
rect 4062 14764 4068 14776
rect 4120 14764 4126 14816
rect 4430 14764 4436 14816
rect 4488 14804 4494 14816
rect 5000 14804 5028 14971
rect 5350 14900 5356 14952
rect 5408 14940 5414 14952
rect 5445 14943 5503 14949
rect 5445 14940 5457 14943
rect 5408 14912 5457 14940
rect 5408 14900 5414 14912
rect 5445 14909 5457 14912
rect 5491 14909 5503 14943
rect 5644 14940 5672 14980
rect 5718 14968 5724 15020
rect 5776 15008 5782 15020
rect 7101 15011 7159 15017
rect 7101 15008 7113 15011
rect 5776 14980 7113 15008
rect 5776 14968 5782 14980
rect 7101 14977 7113 14980
rect 7147 14977 7159 15011
rect 9692 15008 9720 15048
rect 9858 15008 9864 15020
rect 7101 14971 7159 14977
rect 8312 14980 9720 15008
rect 9819 14980 9864 15008
rect 6089 14943 6147 14949
rect 6089 14940 6101 14943
rect 5644 14912 6101 14940
rect 5445 14903 5503 14909
rect 6089 14909 6101 14912
rect 6135 14909 6147 14943
rect 6089 14903 6147 14909
rect 6917 14943 6975 14949
rect 6917 14909 6929 14943
rect 6963 14909 6975 14943
rect 6917 14903 6975 14909
rect 7009 14943 7067 14949
rect 7009 14909 7021 14943
rect 7055 14940 7067 14943
rect 7282 14940 7288 14952
rect 7055 14912 7288 14940
rect 7055 14909 7067 14912
rect 7009 14903 7067 14909
rect 5534 14832 5540 14884
rect 5592 14872 5598 14884
rect 5721 14875 5779 14881
rect 5721 14872 5733 14875
rect 5592 14844 5733 14872
rect 5592 14832 5598 14844
rect 5721 14841 5733 14844
rect 5767 14841 5779 14875
rect 5721 14835 5779 14841
rect 4488 14776 5028 14804
rect 5353 14807 5411 14813
rect 4488 14764 4494 14776
rect 5353 14773 5365 14807
rect 5399 14804 5411 14807
rect 5626 14804 5632 14816
rect 5399 14776 5632 14804
rect 5399 14773 5411 14776
rect 5353 14767 5411 14773
rect 5626 14764 5632 14776
rect 5684 14764 5690 14816
rect 6104 14804 6132 14903
rect 6932 14872 6960 14903
rect 7282 14900 7288 14912
rect 7340 14900 7346 14952
rect 7742 14900 7748 14952
rect 7800 14940 7806 14952
rect 8312 14940 8340 14980
rect 9858 14968 9864 14980
rect 9916 14968 9922 15020
rect 7800 14912 8340 14940
rect 8389 14943 8447 14949
rect 7800 14900 7806 14912
rect 8389 14909 8401 14943
rect 8435 14909 8447 14943
rect 8389 14903 8447 14909
rect 7190 14872 7196 14884
rect 6932 14844 7196 14872
rect 7190 14832 7196 14844
rect 7248 14832 7254 14884
rect 8202 14832 8208 14884
rect 8260 14872 8266 14884
rect 8404 14872 8432 14903
rect 8662 14900 8668 14952
rect 8720 14940 8726 14952
rect 8757 14943 8815 14949
rect 8757 14940 8769 14943
rect 8720 14912 8769 14940
rect 8720 14900 8726 14912
rect 8757 14909 8769 14912
rect 8803 14909 8815 14943
rect 8757 14903 8815 14909
rect 9122 14900 9128 14952
rect 9180 14940 9186 14952
rect 9953 14943 10011 14949
rect 9953 14940 9965 14943
rect 9180 14912 9965 14940
rect 9180 14900 9186 14912
rect 9953 14909 9965 14912
rect 9999 14909 10011 14943
rect 9953 14903 10011 14909
rect 10137 14943 10195 14949
rect 10137 14909 10149 14943
rect 10183 14940 10195 14943
rect 10888 14940 10916 15048
rect 12894 15036 12900 15048
rect 12952 15036 12958 15088
rect 13538 15076 13544 15088
rect 13096 15048 13544 15076
rect 10965 15011 11023 15017
rect 10965 14977 10977 15011
rect 11011 14977 11023 15011
rect 13096 15008 13124 15048
rect 13538 15036 13544 15048
rect 13596 15036 13602 15088
rect 10965 14971 11023 14977
rect 11256 14980 13124 15008
rect 13193 15011 13251 15017
rect 10183 14912 10916 14940
rect 10183 14909 10195 14912
rect 10137 14903 10195 14909
rect 10502 14872 10508 14884
rect 8260 14844 8432 14872
rect 9232 14844 10508 14872
rect 8260 14832 8266 14844
rect 9232 14804 9260 14844
rect 10502 14832 10508 14844
rect 10560 14832 10566 14884
rect 9398 14804 9404 14816
rect 6104 14776 9260 14804
rect 9359 14776 9404 14804
rect 9398 14764 9404 14776
rect 9456 14764 9462 14816
rect 10226 14764 10232 14816
rect 10284 14804 10290 14816
rect 10413 14807 10471 14813
rect 10413 14804 10425 14807
rect 10284 14776 10425 14804
rect 10284 14764 10290 14776
rect 10413 14773 10425 14776
rect 10459 14804 10471 14807
rect 10980 14804 11008 14971
rect 11256 14949 11284 14980
rect 13193 14977 13205 15011
rect 13239 15008 13251 15011
rect 13354 15008 13360 15020
rect 13239 14980 13360 15008
rect 13239 14977 13251 14980
rect 13193 14971 13251 14977
rect 13354 14968 13360 14980
rect 13412 14968 13418 15020
rect 13449 15011 13507 15017
rect 13449 14977 13461 15011
rect 13495 15008 13507 15011
rect 13495 14980 13676 15008
rect 13495 14977 13507 14980
rect 13449 14971 13507 14977
rect 13648 14949 13676 14980
rect 15010 14968 15016 15020
rect 15068 15017 15074 15020
rect 15068 15008 15080 15017
rect 15068 14980 15113 15008
rect 15068 14971 15080 14980
rect 15068 14968 15074 14971
rect 15194 14968 15200 15020
rect 15252 15008 15258 15020
rect 15289 15011 15347 15017
rect 15289 15008 15301 15011
rect 15252 14980 15301 15008
rect 15252 14968 15258 14980
rect 15289 14977 15301 14980
rect 15335 15008 15347 15011
rect 15381 15011 15439 15017
rect 15381 15008 15393 15011
rect 15335 14980 15393 15008
rect 15335 14977 15347 14980
rect 15289 14971 15347 14977
rect 15381 14977 15393 14980
rect 15427 14977 15439 15011
rect 17782 15011 17840 15017
rect 17782 15008 17794 15011
rect 15381 14971 15439 14977
rect 16040 14980 17794 15008
rect 11241 14943 11299 14949
rect 11241 14909 11253 14943
rect 11287 14909 11299 14943
rect 11241 14903 11299 14909
rect 13633 14943 13691 14949
rect 13633 14909 13645 14943
rect 13679 14940 13691 14943
rect 13722 14940 13728 14952
rect 13679 14912 13728 14940
rect 13679 14909 13691 14912
rect 13633 14903 13691 14909
rect 13722 14900 13728 14912
rect 13780 14900 13786 14952
rect 13446 14832 13452 14884
rect 13504 14872 13510 14884
rect 13504 14844 14412 14872
rect 13504 14832 13510 14844
rect 12066 14804 12072 14816
rect 10459 14776 11008 14804
rect 12027 14776 12072 14804
rect 10459 14773 10471 14776
rect 10413 14767 10471 14773
rect 12066 14764 12072 14776
rect 12124 14764 12130 14816
rect 12526 14764 12532 14816
rect 12584 14804 12590 14816
rect 13630 14804 13636 14816
rect 12584 14776 13636 14804
rect 12584 14764 12590 14776
rect 13630 14764 13636 14776
rect 13688 14764 13694 14816
rect 14384 14804 14412 14844
rect 16040 14804 16068 14980
rect 17782 14977 17794 14980
rect 17828 15008 17840 15011
rect 17880 15008 17908 15116
rect 20070 15104 20076 15116
rect 20128 15104 20134 15156
rect 17828 14980 17908 15008
rect 18156 15048 20116 15076
rect 17828 14977 17840 14980
rect 17782 14971 17840 14977
rect 18046 14940 18052 14952
rect 18007 14912 18052 14940
rect 18046 14900 18052 14912
rect 18104 14940 18110 14952
rect 18156 14949 18184 15048
rect 19794 14968 19800 15020
rect 19852 15017 19858 15020
rect 20088 15017 20116 15048
rect 20162 15036 20168 15088
rect 20220 15076 20226 15088
rect 21278 15079 21336 15085
rect 21278 15076 21290 15079
rect 20220 15048 21290 15076
rect 20220 15036 20226 15048
rect 21278 15045 21290 15048
rect 21324 15045 21336 15079
rect 21278 15039 21336 15045
rect 19852 15008 19864 15017
rect 20073 15011 20131 15017
rect 19852 14980 19897 15008
rect 19852 14971 19864 14980
rect 20073 14977 20085 15011
rect 20119 15008 20131 15011
rect 20714 15008 20720 15020
rect 20119 14980 20720 15008
rect 20119 14977 20131 14980
rect 20073 14971 20131 14977
rect 19852 14968 19858 14971
rect 20714 14968 20720 14980
rect 20772 15008 20778 15020
rect 21545 15011 21603 15017
rect 21545 15008 21557 15011
rect 20772 14980 21557 15008
rect 20772 14968 20778 14980
rect 21545 14977 21557 14980
rect 21591 14977 21603 15011
rect 21545 14971 21603 14977
rect 18141 14943 18199 14949
rect 18141 14940 18153 14943
rect 18104 14912 18153 14940
rect 18104 14900 18110 14912
rect 18141 14909 18153 14912
rect 18187 14909 18199 14943
rect 18141 14903 18199 14909
rect 16206 14872 16212 14884
rect 16119 14844 16212 14872
rect 16206 14832 16212 14844
rect 16264 14872 16270 14884
rect 16264 14844 16804 14872
rect 16264 14832 16270 14844
rect 14384 14776 16068 14804
rect 16776 14804 16804 14844
rect 18064 14844 18828 14872
rect 18064 14804 18092 14844
rect 18690 14804 18696 14816
rect 16776 14776 18092 14804
rect 18651 14776 18696 14804
rect 18690 14764 18696 14776
rect 18748 14764 18754 14816
rect 18800 14804 18828 14844
rect 20165 14807 20223 14813
rect 20165 14804 20177 14807
rect 18800 14776 20177 14804
rect 20165 14773 20177 14776
rect 20211 14773 20223 14807
rect 20165 14767 20223 14773
rect 1104 14714 21896 14736
rect 1104 14662 3549 14714
rect 3601 14662 3613 14714
rect 3665 14662 3677 14714
rect 3729 14662 3741 14714
rect 3793 14662 3805 14714
rect 3857 14662 8747 14714
rect 8799 14662 8811 14714
rect 8863 14662 8875 14714
rect 8927 14662 8939 14714
rect 8991 14662 9003 14714
rect 9055 14662 13945 14714
rect 13997 14662 14009 14714
rect 14061 14662 14073 14714
rect 14125 14662 14137 14714
rect 14189 14662 14201 14714
rect 14253 14662 19143 14714
rect 19195 14662 19207 14714
rect 19259 14662 19271 14714
rect 19323 14662 19335 14714
rect 19387 14662 19399 14714
rect 19451 14662 21896 14714
rect 1104 14640 21896 14662
rect 3421 14603 3479 14609
rect 3421 14569 3433 14603
rect 3467 14600 3479 14603
rect 4154 14600 4160 14612
rect 3467 14572 4160 14600
rect 3467 14569 3479 14572
rect 3421 14563 3479 14569
rect 4154 14560 4160 14572
rect 4212 14560 4218 14612
rect 4617 14603 4675 14609
rect 4617 14569 4629 14603
rect 4663 14600 4675 14603
rect 4890 14600 4896 14612
rect 4663 14572 4896 14600
rect 4663 14569 4675 14572
rect 4617 14563 4675 14569
rect 4890 14560 4896 14572
rect 4948 14560 4954 14612
rect 6641 14603 6699 14609
rect 5000 14572 6592 14600
rect 3237 14535 3295 14541
rect 3237 14501 3249 14535
rect 3283 14532 3295 14535
rect 4430 14532 4436 14544
rect 3283 14504 4436 14532
rect 3283 14501 3295 14504
rect 3237 14495 3295 14501
rect 4430 14492 4436 14504
rect 4488 14492 4494 14544
rect 3418 14424 3424 14476
rect 3476 14464 3482 14476
rect 3605 14467 3663 14473
rect 3605 14464 3617 14467
rect 3476 14436 3617 14464
rect 3476 14424 3482 14436
rect 3605 14433 3617 14436
rect 3651 14433 3663 14467
rect 3605 14427 3663 14433
rect 4065 14467 4123 14473
rect 4065 14433 4077 14467
rect 4111 14464 4123 14467
rect 5000 14464 5028 14572
rect 5626 14492 5632 14544
rect 5684 14532 5690 14544
rect 6564 14532 6592 14572
rect 6641 14569 6653 14603
rect 6687 14600 6699 14603
rect 9122 14600 9128 14612
rect 6687 14572 9128 14600
rect 6687 14569 6699 14572
rect 6641 14563 6699 14569
rect 9122 14560 9128 14572
rect 9180 14560 9186 14612
rect 9861 14603 9919 14609
rect 9861 14569 9873 14603
rect 9907 14600 9919 14603
rect 10042 14600 10048 14612
rect 9907 14572 10048 14600
rect 9907 14569 9919 14572
rect 9861 14563 9919 14569
rect 10042 14560 10048 14572
rect 10100 14560 10106 14612
rect 10502 14560 10508 14612
rect 10560 14600 10566 14612
rect 10560 14572 10824 14600
rect 10560 14560 10566 14572
rect 7742 14532 7748 14544
rect 5684 14504 6224 14532
rect 6564 14504 7748 14532
rect 5684 14492 5690 14504
rect 4111 14436 5028 14464
rect 5077 14467 5135 14473
rect 4111 14433 4123 14436
rect 4065 14427 4123 14433
rect 5077 14433 5089 14467
rect 5123 14464 5135 14467
rect 5258 14464 5264 14476
rect 5123 14436 5264 14464
rect 5123 14433 5135 14436
rect 5077 14427 5135 14433
rect 3620 14260 3648 14427
rect 5258 14424 5264 14436
rect 5316 14424 5322 14476
rect 6196 14473 6224 14504
rect 7742 14492 7748 14504
rect 7800 14492 7806 14544
rect 8386 14532 8392 14544
rect 8036 14504 8392 14532
rect 6089 14467 6147 14473
rect 6089 14433 6101 14467
rect 6135 14433 6147 14467
rect 6089 14427 6147 14433
rect 6181 14467 6239 14473
rect 6181 14433 6193 14467
rect 6227 14433 6239 14467
rect 7374 14464 7380 14476
rect 6181 14427 6239 14433
rect 6288 14436 7380 14464
rect 4154 14356 4160 14408
rect 4212 14396 4218 14408
rect 4249 14399 4307 14405
rect 4249 14396 4261 14399
rect 4212 14368 4261 14396
rect 4212 14356 4218 14368
rect 4249 14365 4261 14368
rect 4295 14396 4307 14399
rect 4709 14399 4767 14405
rect 4709 14396 4721 14399
rect 4295 14368 4721 14396
rect 4295 14365 4307 14368
rect 4249 14359 4307 14365
rect 4709 14365 4721 14368
rect 4755 14396 4767 14399
rect 5169 14399 5227 14405
rect 5169 14396 5181 14399
rect 4755 14368 5181 14396
rect 4755 14365 4767 14368
rect 4709 14359 4767 14365
rect 5169 14365 5181 14368
rect 5215 14365 5227 14399
rect 6104 14396 6132 14427
rect 6288 14396 6316 14436
rect 7374 14424 7380 14436
rect 7432 14424 7438 14476
rect 7469 14467 7527 14473
rect 7469 14433 7481 14467
rect 7515 14464 7527 14467
rect 7650 14464 7656 14476
rect 7515 14436 7656 14464
rect 7515 14433 7527 14436
rect 7469 14427 7527 14433
rect 7650 14424 7656 14436
rect 7708 14464 7714 14476
rect 7834 14464 7840 14476
rect 7708 14436 7840 14464
rect 7708 14424 7714 14436
rect 7834 14424 7840 14436
rect 7892 14424 7898 14476
rect 8036 14473 8064 14504
rect 8386 14492 8392 14504
rect 8444 14492 8450 14544
rect 10796 14532 10824 14572
rect 11054 14560 11060 14612
rect 11112 14600 11118 14612
rect 12526 14600 12532 14612
rect 11112 14572 12532 14600
rect 11112 14560 11118 14572
rect 12526 14560 12532 14572
rect 12584 14560 12590 14612
rect 14918 14600 14924 14612
rect 12636 14572 14924 14600
rect 11238 14532 11244 14544
rect 8496 14504 10732 14532
rect 10796 14504 11244 14532
rect 8021 14467 8079 14473
rect 8021 14433 8033 14467
rect 8067 14433 8079 14467
rect 8202 14464 8208 14476
rect 8163 14436 8208 14464
rect 8021 14427 8079 14433
rect 8202 14424 8208 14436
rect 8260 14424 8266 14476
rect 8294 14424 8300 14476
rect 8352 14464 8358 14476
rect 8496 14464 8524 14504
rect 8352 14436 8524 14464
rect 8352 14424 8358 14436
rect 9122 14424 9128 14476
rect 9180 14464 9186 14476
rect 9217 14467 9275 14473
rect 9217 14464 9229 14467
rect 9180 14436 9229 14464
rect 9180 14424 9186 14436
rect 9217 14433 9229 14436
rect 9263 14433 9275 14467
rect 9217 14427 9275 14433
rect 9398 14424 9404 14476
rect 9456 14464 9462 14476
rect 10597 14467 10655 14473
rect 9456 14436 10180 14464
rect 9456 14424 9462 14436
rect 6104 14368 6316 14396
rect 5169 14359 5227 14365
rect 7098 14356 7104 14408
rect 7156 14396 7162 14408
rect 9493 14399 9551 14405
rect 9493 14396 9505 14399
rect 7156 14368 9505 14396
rect 7156 14356 7162 14368
rect 9493 14365 9505 14368
rect 9539 14365 9551 14399
rect 9493 14359 9551 14365
rect 4522 14288 4528 14340
rect 4580 14328 4586 14340
rect 5261 14331 5319 14337
rect 5261 14328 5273 14331
rect 4580 14300 5273 14328
rect 4580 14288 4586 14300
rect 5261 14297 5273 14300
rect 5307 14297 5319 14331
rect 7466 14328 7472 14340
rect 5261 14291 5319 14297
rect 5644 14300 7472 14328
rect 5644 14269 5672 14300
rect 7466 14288 7472 14300
rect 7524 14288 7530 14340
rect 9401 14331 9459 14337
rect 9401 14297 9413 14331
rect 9447 14328 9459 14331
rect 10152 14328 10180 14436
rect 10597 14433 10609 14467
rect 10643 14433 10655 14467
rect 10704 14464 10732 14504
rect 11238 14492 11244 14504
rect 11296 14532 11302 14544
rect 12636 14532 12664 14572
rect 14918 14560 14924 14572
rect 14976 14560 14982 14612
rect 15194 14560 15200 14612
rect 15252 14600 15258 14612
rect 15933 14603 15991 14609
rect 15933 14600 15945 14603
rect 15252 14572 15945 14600
rect 15252 14560 15258 14572
rect 11296 14504 12664 14532
rect 11296 14492 11302 14504
rect 13630 14492 13636 14544
rect 13688 14532 13694 14544
rect 13688 14504 14872 14532
rect 13688 14492 13694 14504
rect 13541 14467 13599 14473
rect 10704 14436 12434 14464
rect 10597 14427 10655 14433
rect 10318 14396 10324 14408
rect 10279 14368 10324 14396
rect 10318 14356 10324 14368
rect 10376 14356 10382 14408
rect 10502 14356 10508 14408
rect 10560 14396 10566 14408
rect 10612 14396 10640 14427
rect 11790 14396 11796 14408
rect 10560 14368 11796 14396
rect 10560 14356 10566 14368
rect 11790 14356 11796 14368
rect 11848 14356 11854 14408
rect 10413 14331 10471 14337
rect 10413 14328 10425 14331
rect 9447 14300 9996 14328
rect 10152 14300 10425 14328
rect 9447 14297 9459 14300
rect 9401 14291 9459 14297
rect 4157 14263 4215 14269
rect 4157 14260 4169 14263
rect 3620 14232 4169 14260
rect 4157 14229 4169 14232
rect 4203 14229 4215 14263
rect 4157 14223 4215 14229
rect 5629 14263 5687 14269
rect 5629 14229 5641 14263
rect 5675 14229 5687 14263
rect 5629 14223 5687 14229
rect 6273 14263 6331 14269
rect 6273 14229 6285 14263
rect 6319 14260 6331 14263
rect 6546 14260 6552 14272
rect 6319 14232 6552 14260
rect 6319 14229 6331 14232
rect 6273 14223 6331 14229
rect 6546 14220 6552 14232
rect 6604 14220 6610 14272
rect 7561 14263 7619 14269
rect 7561 14229 7573 14263
rect 7607 14260 7619 14263
rect 7742 14260 7748 14272
rect 7607 14232 7748 14260
rect 7607 14229 7619 14232
rect 7561 14223 7619 14229
rect 7742 14220 7748 14232
rect 7800 14220 7806 14272
rect 7834 14220 7840 14272
rect 7892 14260 7898 14272
rect 7929 14263 7987 14269
rect 7929 14260 7941 14263
rect 7892 14232 7941 14260
rect 7892 14220 7898 14232
rect 7929 14229 7941 14232
rect 7975 14229 7987 14263
rect 7929 14223 7987 14229
rect 8018 14220 8024 14272
rect 8076 14260 8082 14272
rect 8202 14260 8208 14272
rect 8076 14232 8208 14260
rect 8076 14220 8082 14232
rect 8202 14220 8208 14232
rect 8260 14260 8266 14272
rect 8573 14263 8631 14269
rect 8573 14260 8585 14263
rect 8260 14232 8585 14260
rect 8260 14220 8266 14232
rect 8573 14229 8585 14232
rect 8619 14229 8631 14263
rect 8573 14223 8631 14229
rect 9122 14220 9128 14272
rect 9180 14260 9186 14272
rect 9582 14260 9588 14272
rect 9180 14232 9588 14260
rect 9180 14220 9186 14232
rect 9582 14220 9588 14232
rect 9640 14220 9646 14272
rect 9968 14269 9996 14300
rect 10413 14297 10425 14300
rect 10459 14297 10471 14331
rect 12406 14328 12434 14436
rect 13541 14433 13553 14467
rect 13587 14464 13599 14467
rect 13722 14464 13728 14476
rect 13587 14436 13728 14464
rect 13587 14433 13599 14436
rect 13541 14427 13599 14433
rect 13722 14424 13728 14436
rect 13780 14424 13786 14476
rect 12526 14356 12532 14408
rect 12584 14396 12590 14408
rect 13274 14399 13332 14405
rect 13274 14396 13286 14399
rect 12584 14368 13286 14396
rect 12584 14356 12590 14368
rect 13274 14365 13286 14368
rect 13320 14396 13332 14399
rect 13814 14396 13820 14408
rect 13320 14368 13820 14396
rect 13320 14365 13332 14368
rect 13274 14359 13332 14365
rect 13814 14356 13820 14368
rect 13872 14356 13878 14408
rect 13446 14328 13452 14340
rect 12406 14300 13452 14328
rect 10413 14291 10471 14297
rect 13446 14288 13452 14300
rect 13504 14288 13510 14340
rect 13538 14288 13544 14340
rect 13596 14328 13602 14340
rect 14844 14328 14872 14504
rect 15856 14473 15884 14572
rect 15933 14569 15945 14572
rect 15979 14569 15991 14603
rect 17681 14603 17739 14609
rect 17681 14600 17693 14603
rect 15933 14563 15991 14569
rect 16408 14572 17693 14600
rect 16408 14476 16436 14572
rect 15841 14467 15899 14473
rect 15841 14433 15853 14467
rect 15887 14464 15899 14467
rect 16390 14464 16396 14476
rect 15887 14436 16396 14464
rect 15887 14433 15899 14436
rect 15841 14427 15899 14433
rect 16390 14424 16396 14436
rect 16448 14424 16454 14476
rect 17604 14473 17632 14572
rect 17681 14569 17693 14572
rect 17727 14600 17739 14603
rect 18046 14600 18052 14612
rect 17727 14572 18052 14600
rect 17727 14569 17739 14572
rect 17681 14563 17739 14569
rect 18046 14560 18052 14572
rect 18104 14560 18110 14612
rect 20714 14560 20720 14612
rect 20772 14600 20778 14612
rect 21177 14603 21235 14609
rect 21177 14600 21189 14603
rect 20772 14572 21189 14600
rect 20772 14560 20778 14572
rect 21100 14473 21128 14572
rect 21177 14569 21189 14572
rect 21223 14600 21235 14603
rect 21450 14600 21456 14612
rect 21223 14572 21456 14600
rect 21223 14569 21235 14572
rect 21177 14563 21235 14569
rect 21450 14560 21456 14572
rect 21508 14560 21514 14612
rect 17589 14467 17647 14473
rect 17589 14433 17601 14467
rect 17635 14433 17647 14467
rect 17589 14427 17647 14433
rect 21085 14467 21143 14473
rect 21085 14433 21097 14467
rect 21131 14433 21143 14467
rect 21085 14427 21143 14433
rect 15562 14396 15568 14408
rect 15620 14405 15626 14408
rect 15620 14399 15643 14405
rect 15495 14368 15568 14396
rect 15562 14356 15568 14368
rect 15631 14396 15643 14399
rect 16206 14396 16212 14408
rect 15631 14368 16212 14396
rect 15631 14365 15643 14368
rect 15620 14359 15643 14365
rect 15620 14356 15626 14359
rect 16206 14356 16212 14368
rect 16264 14356 16270 14408
rect 20346 14396 20352 14408
rect 17144 14368 20352 14396
rect 17144 14328 17172 14368
rect 20346 14356 20352 14368
rect 20404 14356 20410 14408
rect 13596 14300 14504 14328
rect 14844 14300 17172 14328
rect 13596 14288 13602 14300
rect 9953 14263 10011 14269
rect 9953 14229 9965 14263
rect 9999 14229 10011 14263
rect 9953 14223 10011 14229
rect 10042 14220 10048 14272
rect 10100 14260 10106 14272
rect 10318 14260 10324 14272
rect 10100 14232 10324 14260
rect 10100 14220 10106 14232
rect 10318 14220 10324 14232
rect 10376 14220 10382 14272
rect 11882 14220 11888 14272
rect 11940 14260 11946 14272
rect 12161 14263 12219 14269
rect 12161 14260 12173 14263
rect 11940 14232 12173 14260
rect 11940 14220 11946 14232
rect 12161 14229 12173 14232
rect 12207 14260 12219 14263
rect 12342 14260 12348 14272
rect 12207 14232 12348 14260
rect 12207 14229 12219 14232
rect 12161 14223 12219 14229
rect 12342 14220 12348 14232
rect 12400 14220 12406 14272
rect 12710 14220 12716 14272
rect 12768 14260 12774 14272
rect 13170 14260 13176 14272
rect 12768 14232 13176 14260
rect 12768 14220 12774 14232
rect 13170 14220 13176 14232
rect 13228 14220 13234 14272
rect 13630 14260 13636 14272
rect 13591 14232 13636 14260
rect 13630 14220 13636 14232
rect 13688 14220 13694 14272
rect 14476 14269 14504 14300
rect 17218 14288 17224 14340
rect 17276 14328 17282 14340
rect 17322 14331 17380 14337
rect 17322 14328 17334 14331
rect 17276 14300 17334 14328
rect 17276 14288 17282 14300
rect 17322 14297 17334 14300
rect 17368 14297 17380 14331
rect 17322 14291 17380 14297
rect 20806 14288 20812 14340
rect 20864 14337 20870 14340
rect 20864 14328 20876 14337
rect 20864 14300 20909 14328
rect 20864 14291 20876 14300
rect 20864 14288 20870 14291
rect 14461 14263 14519 14269
rect 14461 14229 14473 14263
rect 14507 14229 14519 14263
rect 16206 14260 16212 14272
rect 16119 14232 16212 14260
rect 14461 14223 14519 14229
rect 16206 14220 16212 14232
rect 16264 14260 16270 14272
rect 19058 14260 19064 14272
rect 16264 14232 19064 14260
rect 16264 14220 16270 14232
rect 19058 14220 19064 14232
rect 19116 14220 19122 14272
rect 19705 14263 19763 14269
rect 19705 14229 19717 14263
rect 19751 14260 19763 14263
rect 19794 14260 19800 14272
rect 19751 14232 19800 14260
rect 19751 14229 19763 14232
rect 19705 14223 19763 14229
rect 19794 14220 19800 14232
rect 19852 14220 19858 14272
rect 1104 14170 22056 14192
rect 1104 14118 6148 14170
rect 6200 14118 6212 14170
rect 6264 14118 6276 14170
rect 6328 14118 6340 14170
rect 6392 14118 6404 14170
rect 6456 14118 11346 14170
rect 11398 14118 11410 14170
rect 11462 14118 11474 14170
rect 11526 14118 11538 14170
rect 11590 14118 11602 14170
rect 11654 14118 16544 14170
rect 16596 14118 16608 14170
rect 16660 14118 16672 14170
rect 16724 14118 16736 14170
rect 16788 14118 16800 14170
rect 16852 14118 21742 14170
rect 21794 14118 21806 14170
rect 21858 14118 21870 14170
rect 21922 14118 21934 14170
rect 21986 14118 21998 14170
rect 22050 14118 22056 14170
rect 1104 14096 22056 14118
rect 2130 14016 2136 14068
rect 2188 14056 2194 14068
rect 4154 14056 4160 14068
rect 2188 14028 4160 14056
rect 2188 14016 2194 14028
rect 4154 14016 4160 14028
rect 4212 14016 4218 14068
rect 4522 14056 4528 14068
rect 4483 14028 4528 14056
rect 4522 14016 4528 14028
rect 4580 14016 4586 14068
rect 5350 14056 5356 14068
rect 5311 14028 5356 14056
rect 5350 14016 5356 14028
rect 5408 14016 5414 14068
rect 5718 14056 5724 14068
rect 5679 14028 5724 14056
rect 5718 14016 5724 14028
rect 5776 14016 5782 14068
rect 6365 14059 6423 14065
rect 6365 14025 6377 14059
rect 6411 14056 6423 14059
rect 6546 14056 6552 14068
rect 6411 14028 6552 14056
rect 6411 14025 6423 14028
rect 6365 14019 6423 14025
rect 6546 14016 6552 14028
rect 6604 14016 6610 14068
rect 7282 14056 7288 14068
rect 7243 14028 7288 14056
rect 7282 14016 7288 14028
rect 7340 14016 7346 14068
rect 7742 14056 7748 14068
rect 7703 14028 7748 14056
rect 7742 14016 7748 14028
rect 7800 14016 7806 14068
rect 9766 14056 9772 14068
rect 8772 14028 9772 14056
rect 4540 13988 4568 14016
rect 5905 13991 5963 13997
rect 5905 13988 5917 13991
rect 4540 13960 5917 13988
rect 5905 13957 5917 13960
rect 5951 13988 5963 13991
rect 6825 13991 6883 13997
rect 6825 13988 6837 13991
rect 5951 13960 6837 13988
rect 5951 13957 5963 13960
rect 5905 13951 5963 13957
rect 6825 13957 6837 13960
rect 6871 13957 6883 13991
rect 6825 13951 6883 13957
rect 7190 13948 7196 14000
rect 7248 13988 7254 14000
rect 8662 13988 8668 14000
rect 7248 13960 8668 13988
rect 7248 13948 7254 13960
rect 8662 13948 8668 13960
rect 8720 13948 8726 14000
rect 6730 13920 6736 13932
rect 6643 13892 6736 13920
rect 6730 13880 6736 13892
rect 6788 13880 6794 13932
rect 7650 13920 7656 13932
rect 6840 13892 7052 13920
rect 7611 13892 7656 13920
rect 5077 13855 5135 13861
rect 5077 13821 5089 13855
rect 5123 13821 5135 13855
rect 5077 13815 5135 13821
rect 5092 13784 5120 13815
rect 5166 13812 5172 13864
rect 5224 13852 5230 13864
rect 5261 13855 5319 13861
rect 5261 13852 5273 13855
rect 5224 13824 5273 13852
rect 5224 13812 5230 13824
rect 5261 13821 5273 13824
rect 5307 13821 5319 13855
rect 6086 13852 6092 13864
rect 6047 13824 6092 13852
rect 5261 13815 5319 13821
rect 6086 13812 6092 13824
rect 6144 13852 6150 13864
rect 6748 13852 6776 13880
rect 6144 13824 6776 13852
rect 6144 13812 6150 13824
rect 5442 13784 5448 13796
rect 5092 13756 5448 13784
rect 5442 13744 5448 13756
rect 5500 13784 5506 13796
rect 6840 13784 6868 13892
rect 6917 13855 6975 13861
rect 6917 13821 6929 13855
rect 6963 13821 6975 13855
rect 6917 13815 6975 13821
rect 5500 13756 6868 13784
rect 5500 13744 5506 13756
rect 4798 13676 4804 13728
rect 4856 13716 4862 13728
rect 6932 13716 6960 13815
rect 7024 13784 7052 13892
rect 7650 13880 7656 13892
rect 7708 13880 7714 13932
rect 8772 13920 8800 14028
rect 9766 14016 9772 14028
rect 9824 14016 9830 14068
rect 10410 14056 10416 14068
rect 10152 14028 10416 14056
rect 9217 13991 9275 13997
rect 9217 13957 9229 13991
rect 9263 13988 9275 13991
rect 10152 13988 10180 14028
rect 10410 14016 10416 14028
rect 10468 14016 10474 14068
rect 10505 14059 10563 14065
rect 10505 14025 10517 14059
rect 10551 14056 10563 14059
rect 11054 14056 11060 14068
rect 10551 14028 11060 14056
rect 10551 14025 10563 14028
rect 10505 14019 10563 14025
rect 11054 14016 11060 14028
rect 11112 14016 11118 14068
rect 11238 14056 11244 14068
rect 11199 14028 11244 14056
rect 11238 14016 11244 14028
rect 11296 14016 11302 14068
rect 12526 14056 12532 14068
rect 12268 14028 12532 14056
rect 9263 13960 10180 13988
rect 9263 13957 9275 13960
rect 9217 13951 9275 13957
rect 10318 13948 10324 14000
rect 10376 13988 10382 14000
rect 11256 13988 11284 14016
rect 10376 13960 11284 13988
rect 10376 13948 10382 13960
rect 7760 13892 8800 13920
rect 9677 13923 9735 13929
rect 7374 13812 7380 13864
rect 7432 13852 7438 13864
rect 7760 13852 7788 13892
rect 9677 13889 9689 13923
rect 9723 13920 9735 13923
rect 9766 13920 9772 13932
rect 9723 13892 9772 13920
rect 9723 13889 9735 13892
rect 9677 13883 9735 13889
rect 9766 13880 9772 13892
rect 9824 13880 9830 13932
rect 12268 13929 12296 14028
rect 12526 14016 12532 14028
rect 12584 14056 12590 14068
rect 13630 14056 13636 14068
rect 12584 14028 13636 14056
rect 12584 14016 12590 14028
rect 13630 14016 13636 14028
rect 13688 14016 13694 14068
rect 15102 14056 15108 14068
rect 15063 14028 15108 14056
rect 15102 14016 15108 14028
rect 15160 14016 15166 14068
rect 17218 14016 17224 14068
rect 17276 14056 17282 14068
rect 18141 14059 18199 14065
rect 18141 14056 18153 14059
rect 17276 14028 18153 14056
rect 17276 14016 17282 14028
rect 18141 14025 18153 14028
rect 18187 14025 18199 14059
rect 18141 14019 18199 14025
rect 19705 14059 19763 14065
rect 19705 14025 19717 14059
rect 19751 14056 19763 14059
rect 20714 14056 20720 14068
rect 19751 14028 20720 14056
rect 19751 14025 19763 14028
rect 19705 14019 19763 14025
rect 12342 13948 12348 14000
rect 12400 13988 12406 14000
rect 16218 13991 16276 13997
rect 16218 13988 16230 13991
rect 12400 13960 16230 13988
rect 12400 13948 12406 13960
rect 16218 13957 16230 13960
rect 16264 13957 16276 13991
rect 16914 13991 16972 13997
rect 16914 13988 16926 13991
rect 16218 13951 16276 13957
rect 16316 13960 16926 13988
rect 12253 13923 12311 13929
rect 12253 13889 12265 13923
rect 12299 13889 12311 13923
rect 12509 13923 12567 13929
rect 12509 13920 12521 13923
rect 12253 13883 12311 13889
rect 12360 13892 12521 13920
rect 7432 13824 7788 13852
rect 7837 13855 7895 13861
rect 7432 13812 7438 13824
rect 7837 13821 7849 13855
rect 7883 13821 7895 13855
rect 7837 13815 7895 13821
rect 9493 13855 9551 13861
rect 9493 13821 9505 13855
rect 9539 13821 9551 13855
rect 9493 13815 9551 13821
rect 9585 13855 9643 13861
rect 9585 13821 9597 13855
rect 9631 13852 9643 13855
rect 10226 13852 10232 13864
rect 9631 13824 9720 13852
rect 10187 13824 10232 13852
rect 9631 13821 9643 13824
rect 9585 13815 9643 13821
rect 7852 13784 7880 13815
rect 7024 13756 7880 13784
rect 7282 13716 7288 13728
rect 4856 13688 7288 13716
rect 4856 13676 4862 13688
rect 7282 13676 7288 13688
rect 7340 13716 7346 13728
rect 7558 13716 7564 13728
rect 7340 13688 7564 13716
rect 7340 13676 7346 13688
rect 7558 13676 7564 13688
rect 7616 13676 7622 13728
rect 9508 13716 9536 13815
rect 9692 13796 9720 13824
rect 10226 13812 10232 13824
rect 10284 13812 10290 13864
rect 10413 13855 10471 13861
rect 10413 13821 10425 13855
rect 10459 13852 10471 13855
rect 10502 13852 10508 13864
rect 10459 13824 10508 13852
rect 10459 13821 10471 13824
rect 10413 13815 10471 13821
rect 10502 13812 10508 13824
rect 10560 13852 10566 13864
rect 10870 13852 10876 13864
rect 10560 13824 10876 13852
rect 10560 13812 10566 13824
rect 10870 13812 10876 13824
rect 10928 13812 10934 13864
rect 11790 13812 11796 13864
rect 11848 13852 11854 13864
rect 11974 13852 11980 13864
rect 11848 13824 11980 13852
rect 11848 13812 11854 13824
rect 11974 13812 11980 13824
rect 12032 13852 12038 13864
rect 12360 13852 12388 13892
rect 12509 13889 12521 13892
rect 12555 13889 12567 13923
rect 12509 13883 12567 13889
rect 13538 13880 13544 13932
rect 13596 13920 13602 13932
rect 16316 13920 16344 13960
rect 16914 13957 16926 13960
rect 16960 13957 16972 13991
rect 16914 13951 16972 13957
rect 18690 13948 18696 14000
rect 18748 13988 18754 14000
rect 18966 13988 18972 14000
rect 18748 13960 18972 13988
rect 18748 13948 18754 13960
rect 18966 13948 18972 13960
rect 19024 13988 19030 14000
rect 19254 13991 19312 13997
rect 19254 13988 19266 13991
rect 19024 13960 19266 13988
rect 19024 13948 19030 13960
rect 19254 13957 19266 13960
rect 19300 13957 19312 13991
rect 19254 13951 19312 13957
rect 13596 13892 16344 13920
rect 13596 13880 13602 13892
rect 16390 13880 16396 13932
rect 16448 13920 16454 13932
rect 16485 13923 16543 13929
rect 16485 13920 16497 13923
rect 16448 13892 16497 13920
rect 16448 13880 16454 13892
rect 16485 13889 16497 13892
rect 16531 13920 16543 13923
rect 16669 13923 16727 13929
rect 16669 13920 16681 13923
rect 16531 13892 16681 13920
rect 16531 13889 16543 13892
rect 16485 13883 16543 13889
rect 16669 13889 16681 13892
rect 16715 13889 16727 13923
rect 16669 13883 16727 13889
rect 19521 13923 19579 13929
rect 19521 13889 19533 13923
rect 19567 13920 19579 13923
rect 19720 13920 19748 14019
rect 20180 13929 20208 14028
rect 20714 14016 20720 14028
rect 20772 14016 20778 14068
rect 21266 14016 21272 14068
rect 21324 14056 21330 14068
rect 21542 14056 21548 14068
rect 21324 14028 21548 14056
rect 21324 14016 21330 14028
rect 21542 14016 21548 14028
rect 21600 14016 21606 14068
rect 19567 13892 19748 13920
rect 20165 13923 20223 13929
rect 19567 13889 19579 13892
rect 19521 13883 19579 13889
rect 20165 13889 20177 13923
rect 20211 13889 20223 13923
rect 20165 13883 20223 13889
rect 20254 13880 20260 13932
rect 20312 13920 20318 13932
rect 20421 13923 20479 13929
rect 20421 13920 20433 13923
rect 20312 13892 20433 13920
rect 20312 13880 20318 13892
rect 20421 13889 20433 13892
rect 20467 13889 20479 13923
rect 20421 13883 20479 13889
rect 12032 13824 12388 13852
rect 12032 13812 12038 13824
rect 13354 13812 13360 13864
rect 13412 13852 13418 13864
rect 13412 13824 13676 13852
rect 13412 13812 13418 13824
rect 9674 13744 9680 13796
rect 9732 13744 9738 13796
rect 10042 13784 10048 13796
rect 10003 13756 10048 13784
rect 10042 13744 10048 13756
rect 10100 13744 10106 13796
rect 13648 13793 13676 13824
rect 17954 13812 17960 13864
rect 18012 13852 18018 13864
rect 18012 13824 18092 13852
rect 18012 13812 18018 13824
rect 18064 13793 18092 13824
rect 13633 13787 13691 13793
rect 13633 13753 13645 13787
rect 13679 13753 13691 13787
rect 13633 13747 13691 13753
rect 18049 13787 18107 13793
rect 18049 13753 18061 13787
rect 18095 13753 18107 13787
rect 18049 13747 18107 13753
rect 10594 13716 10600 13728
rect 9508 13688 10600 13716
rect 10594 13676 10600 13688
rect 10652 13676 10658 13728
rect 10870 13716 10876 13728
rect 10831 13688 10876 13716
rect 10870 13676 10876 13688
rect 10928 13676 10934 13728
rect 12250 13676 12256 13728
rect 12308 13716 12314 13728
rect 13538 13716 13544 13728
rect 12308 13688 13544 13716
rect 12308 13676 12314 13688
rect 13538 13676 13544 13688
rect 13596 13676 13602 13728
rect 13817 13719 13875 13725
rect 13817 13685 13829 13719
rect 13863 13716 13875 13719
rect 14274 13716 14280 13728
rect 13863 13688 14280 13716
rect 13863 13685 13875 13688
rect 13817 13679 13875 13685
rect 14274 13676 14280 13688
rect 14332 13676 14338 13728
rect 1104 13626 21896 13648
rect 1104 13574 3549 13626
rect 3601 13574 3613 13626
rect 3665 13574 3677 13626
rect 3729 13574 3741 13626
rect 3793 13574 3805 13626
rect 3857 13574 8747 13626
rect 8799 13574 8811 13626
rect 8863 13574 8875 13626
rect 8927 13574 8939 13626
rect 8991 13574 9003 13626
rect 9055 13574 13945 13626
rect 13997 13574 14009 13626
rect 14061 13574 14073 13626
rect 14125 13574 14137 13626
rect 14189 13574 14201 13626
rect 14253 13574 19143 13626
rect 19195 13574 19207 13626
rect 19259 13574 19271 13626
rect 19323 13574 19335 13626
rect 19387 13574 19399 13626
rect 19451 13574 21896 13626
rect 1104 13552 21896 13574
rect 4798 13472 4804 13524
rect 4856 13512 4862 13524
rect 5534 13512 5540 13524
rect 4856 13484 5540 13512
rect 4856 13472 4862 13484
rect 5534 13472 5540 13484
rect 5592 13472 5598 13524
rect 6089 13515 6147 13521
rect 6089 13481 6101 13515
rect 6135 13512 6147 13515
rect 6822 13512 6828 13524
rect 6135 13484 6828 13512
rect 6135 13481 6147 13484
rect 6089 13475 6147 13481
rect 6822 13472 6828 13484
rect 6880 13472 6886 13524
rect 7098 13512 7104 13524
rect 7059 13484 7104 13512
rect 7098 13472 7104 13484
rect 7156 13472 7162 13524
rect 7929 13515 7987 13521
rect 7929 13481 7941 13515
rect 7975 13512 7987 13515
rect 9674 13512 9680 13524
rect 7975 13484 9680 13512
rect 7975 13481 7987 13484
rect 7929 13475 7987 13481
rect 9674 13472 9680 13484
rect 9732 13472 9738 13524
rect 9784 13484 13768 13512
rect 5074 13404 5080 13456
rect 5132 13444 5138 13456
rect 5442 13444 5448 13456
rect 5132 13416 5448 13444
rect 5132 13404 5138 13416
rect 5442 13404 5448 13416
rect 5500 13444 5506 13456
rect 6181 13447 6239 13453
rect 6181 13444 6193 13447
rect 5500 13416 6193 13444
rect 5500 13404 5506 13416
rect 6181 13413 6193 13416
rect 6227 13413 6239 13447
rect 7742 13444 7748 13456
rect 6181 13407 6239 13413
rect 7300 13416 7748 13444
rect 4706 13376 4712 13388
rect 4667 13348 4712 13376
rect 4706 13336 4712 13348
rect 4764 13336 4770 13388
rect 6546 13376 6552 13388
rect 6507 13348 6552 13376
rect 6546 13336 6552 13348
rect 6604 13336 6610 13388
rect 7300 13385 7328 13416
rect 7742 13404 7748 13416
rect 7800 13404 7806 13456
rect 8021 13447 8079 13453
rect 8021 13413 8033 13447
rect 8067 13413 8079 13447
rect 8021 13407 8079 13413
rect 9401 13447 9459 13453
rect 9401 13413 9413 13447
rect 9447 13444 9459 13447
rect 9490 13444 9496 13456
rect 9447 13416 9496 13444
rect 9447 13413 9459 13416
rect 9401 13407 9459 13413
rect 7285 13379 7343 13385
rect 7285 13345 7297 13379
rect 7331 13345 7343 13379
rect 7466 13376 7472 13388
rect 7427 13348 7472 13376
rect 7285 13339 7343 13345
rect 7466 13336 7472 13348
rect 7524 13336 7530 13388
rect 2133 13311 2191 13317
rect 2133 13277 2145 13311
rect 2179 13308 2191 13311
rect 3326 13308 3332 13320
rect 2179 13280 3332 13308
rect 2179 13277 2191 13280
rect 2133 13271 2191 13277
rect 3326 13268 3332 13280
rect 3384 13268 3390 13320
rect 4985 13311 5043 13317
rect 4985 13277 4997 13311
rect 5031 13308 5043 13311
rect 8036 13308 8064 13407
rect 9490 13404 9496 13416
rect 9548 13404 9554 13456
rect 8662 13376 8668 13388
rect 8623 13348 8668 13376
rect 8662 13336 8668 13348
rect 8720 13336 8726 13388
rect 9784 13376 9812 13484
rect 11057 13447 11115 13453
rect 11057 13444 11069 13447
rect 9876 13416 11069 13444
rect 9876 13385 9904 13416
rect 11057 13413 11069 13416
rect 11103 13413 11115 13447
rect 12434 13444 12440 13456
rect 11057 13407 11115 13413
rect 11624 13416 12440 13444
rect 9646 13348 9812 13376
rect 9861 13379 9919 13385
rect 5031 13280 8064 13308
rect 5031 13277 5043 13280
rect 4985 13271 5043 13277
rect 8202 13268 8208 13320
rect 8260 13308 8266 13320
rect 9646 13308 9674 13348
rect 9861 13345 9873 13379
rect 9907 13345 9919 13379
rect 9861 13339 9919 13345
rect 10045 13379 10103 13385
rect 10045 13345 10057 13379
rect 10091 13376 10103 13379
rect 10873 13379 10931 13385
rect 10091 13348 10824 13376
rect 10091 13345 10103 13348
rect 10045 13339 10103 13345
rect 8260 13280 9674 13308
rect 10689 13311 10747 13317
rect 8260 13268 8266 13280
rect 10689 13277 10701 13311
rect 10735 13277 10747 13311
rect 10689 13271 10747 13277
rect 5350 13200 5356 13252
rect 5408 13240 5414 13252
rect 6641 13243 6699 13249
rect 6641 13240 6653 13243
rect 5408 13212 6653 13240
rect 5408 13200 5414 13212
rect 6641 13209 6653 13212
rect 6687 13209 6699 13243
rect 6641 13203 6699 13209
rect 6914 13200 6920 13252
rect 6972 13240 6978 13252
rect 10704 13240 10732 13271
rect 6972 13212 10732 13240
rect 10796 13240 10824 13348
rect 10873 13345 10885 13379
rect 10919 13376 10931 13379
rect 10962 13376 10968 13388
rect 10919 13348 10968 13376
rect 10919 13345 10931 13348
rect 10873 13339 10931 13345
rect 10962 13336 10968 13348
rect 11020 13376 11026 13388
rect 11624 13376 11652 13416
rect 12434 13404 12440 13416
rect 12492 13404 12498 13456
rect 13740 13444 13768 13484
rect 13814 13472 13820 13524
rect 13872 13512 13878 13524
rect 13909 13515 13967 13521
rect 13909 13512 13921 13515
rect 13872 13484 13921 13512
rect 13872 13472 13878 13484
rect 13909 13481 13921 13484
rect 13955 13512 13967 13515
rect 14366 13512 14372 13524
rect 13955 13484 14372 13512
rect 13955 13481 13967 13484
rect 13909 13475 13967 13481
rect 14366 13472 14372 13484
rect 14424 13472 14430 13524
rect 15010 13472 15016 13524
rect 15068 13512 15074 13524
rect 16117 13515 16175 13521
rect 16117 13512 16129 13515
rect 15068 13484 16129 13512
rect 15068 13472 15074 13484
rect 16117 13481 16129 13484
rect 16163 13481 16175 13515
rect 21450 13512 21456 13524
rect 21411 13484 21456 13512
rect 16117 13475 16175 13481
rect 21450 13472 21456 13484
rect 21508 13472 21514 13524
rect 15562 13444 15568 13456
rect 13740 13416 15568 13444
rect 15562 13404 15568 13416
rect 15620 13404 15626 13456
rect 11020 13348 11652 13376
rect 11701 13379 11759 13385
rect 11020 13336 11026 13348
rect 11701 13345 11713 13379
rect 11747 13376 11759 13379
rect 11974 13376 11980 13388
rect 11747 13348 11980 13376
rect 11747 13345 11759 13348
rect 11701 13339 11759 13345
rect 11974 13336 11980 13348
rect 12032 13336 12038 13388
rect 11514 13308 11520 13320
rect 11475 13280 11520 13308
rect 11514 13268 11520 13280
rect 11572 13268 11578 13320
rect 12526 13308 12532 13320
rect 12487 13280 12532 13308
rect 12526 13268 12532 13280
rect 12584 13268 12590 13320
rect 12728 13280 17273 13308
rect 12728 13240 12756 13280
rect 12802 13249 12808 13252
rect 10796 13212 12756 13240
rect 6972 13200 6978 13212
rect 12796 13203 12808 13249
rect 12860 13240 12866 13252
rect 17245 13249 17273 13280
rect 17402 13268 17408 13320
rect 17460 13308 17466 13320
rect 17497 13311 17555 13317
rect 17497 13308 17509 13311
rect 17460 13280 17509 13308
rect 17460 13268 17466 13280
rect 17497 13277 17509 13280
rect 17543 13277 17555 13311
rect 19702 13308 19708 13320
rect 17497 13271 17555 13277
rect 18156 13280 19708 13308
rect 17230 13243 17288 13249
rect 12860 13212 12896 13240
rect 12802 13200 12808 13203
rect 12860 13200 12866 13212
rect 17230 13209 17242 13243
rect 17276 13240 17288 13243
rect 18046 13240 18052 13252
rect 17276 13212 18052 13240
rect 17276 13209 17288 13212
rect 17230 13203 17288 13209
rect 18046 13200 18052 13212
rect 18104 13200 18110 13252
rect 18156 13184 18184 13280
rect 19702 13268 19708 13280
rect 19760 13308 19766 13320
rect 19889 13311 19947 13317
rect 19889 13308 19901 13311
rect 19760 13280 19901 13308
rect 19760 13268 19766 13280
rect 19889 13277 19901 13280
rect 19935 13308 19947 13311
rect 20714 13308 20720 13320
rect 19935 13280 20720 13308
rect 19935 13277 19947 13280
rect 19889 13271 19947 13277
rect 20714 13268 20720 13280
rect 20772 13268 20778 13320
rect 20156 13243 20214 13249
rect 20156 13209 20168 13243
rect 20202 13240 20214 13243
rect 20622 13240 20628 13252
rect 20202 13212 20628 13240
rect 20202 13209 20214 13212
rect 20156 13203 20214 13209
rect 20622 13200 20628 13212
rect 20680 13200 20686 13252
rect 1946 13172 1952 13184
rect 1907 13144 1952 13172
rect 1946 13132 1952 13144
rect 2004 13132 2010 13184
rect 6730 13172 6736 13184
rect 6691 13144 6736 13172
rect 6730 13132 6736 13144
rect 6788 13132 6794 13184
rect 7558 13132 7564 13184
rect 7616 13172 7622 13184
rect 8386 13172 8392 13184
rect 7616 13144 7661 13172
rect 8347 13144 8392 13172
rect 7616 13132 7622 13144
rect 8386 13132 8392 13144
rect 8444 13132 8450 13184
rect 8481 13175 8539 13181
rect 8481 13141 8493 13175
rect 8527 13172 8539 13175
rect 9306 13172 9312 13184
rect 8527 13144 9312 13172
rect 8527 13141 8539 13144
rect 8481 13135 8539 13141
rect 9306 13132 9312 13144
rect 9364 13132 9370 13184
rect 9398 13132 9404 13184
rect 9456 13172 9462 13184
rect 9582 13172 9588 13184
rect 9456 13144 9588 13172
rect 9456 13132 9462 13144
rect 9582 13132 9588 13144
rect 9640 13132 9646 13184
rect 9674 13132 9680 13184
rect 9732 13172 9738 13184
rect 9769 13175 9827 13181
rect 9769 13172 9781 13175
rect 9732 13144 9781 13172
rect 9732 13132 9738 13144
rect 9769 13141 9781 13144
rect 9815 13141 9827 13175
rect 9769 13135 9827 13141
rect 10229 13175 10287 13181
rect 10229 13141 10241 13175
rect 10275 13172 10287 13175
rect 10410 13172 10416 13184
rect 10275 13144 10416 13172
rect 10275 13141 10287 13144
rect 10229 13135 10287 13141
rect 10410 13132 10416 13144
rect 10468 13132 10474 13184
rect 10597 13175 10655 13181
rect 10597 13141 10609 13175
rect 10643 13172 10655 13175
rect 10870 13172 10876 13184
rect 10643 13144 10876 13172
rect 10643 13141 10655 13144
rect 10597 13135 10655 13141
rect 10870 13132 10876 13144
rect 10928 13132 10934 13184
rect 11238 13132 11244 13184
rect 11296 13172 11302 13184
rect 11425 13175 11483 13181
rect 11425 13172 11437 13175
rect 11296 13144 11437 13172
rect 11296 13132 11302 13144
rect 11425 13141 11437 13144
rect 11471 13141 11483 13175
rect 11425 13135 11483 13141
rect 11974 13132 11980 13184
rect 12032 13172 12038 13184
rect 14090 13172 14096 13184
rect 12032 13144 14096 13172
rect 12032 13132 12038 13144
rect 14090 13132 14096 13144
rect 14148 13132 14154 13184
rect 14185 13175 14243 13181
rect 14185 13141 14197 13175
rect 14231 13172 14243 13175
rect 14274 13172 14280 13184
rect 14231 13144 14280 13172
rect 14231 13141 14243 13144
rect 14185 13135 14243 13141
rect 14274 13132 14280 13144
rect 14332 13132 14338 13184
rect 15930 13172 15936 13184
rect 15891 13144 15936 13172
rect 15930 13132 15936 13144
rect 15988 13172 15994 13184
rect 17402 13172 17408 13184
rect 15988 13144 17408 13172
rect 15988 13132 15994 13144
rect 17402 13132 17408 13144
rect 17460 13172 17466 13184
rect 17589 13175 17647 13181
rect 17589 13172 17601 13175
rect 17460 13144 17601 13172
rect 17460 13132 17466 13144
rect 17589 13141 17601 13144
rect 17635 13172 17647 13175
rect 18138 13172 18144 13184
rect 17635 13144 18144 13172
rect 17635 13141 17647 13144
rect 17589 13135 17647 13141
rect 18138 13132 18144 13144
rect 18196 13132 18202 13184
rect 20898 13132 20904 13184
rect 20956 13172 20962 13184
rect 21174 13172 21180 13184
rect 20956 13144 21180 13172
rect 20956 13132 20962 13144
rect 21174 13132 21180 13144
rect 21232 13172 21238 13184
rect 21269 13175 21327 13181
rect 21269 13172 21281 13175
rect 21232 13144 21281 13172
rect 21232 13132 21238 13144
rect 21269 13141 21281 13144
rect 21315 13141 21327 13175
rect 21269 13135 21327 13141
rect 1104 13082 22056 13104
rect 1104 13030 6148 13082
rect 6200 13030 6212 13082
rect 6264 13030 6276 13082
rect 6328 13030 6340 13082
rect 6392 13030 6404 13082
rect 6456 13030 11346 13082
rect 11398 13030 11410 13082
rect 11462 13030 11474 13082
rect 11526 13030 11538 13082
rect 11590 13030 11602 13082
rect 11654 13030 16544 13082
rect 16596 13030 16608 13082
rect 16660 13030 16672 13082
rect 16724 13030 16736 13082
rect 16788 13030 16800 13082
rect 16852 13030 21742 13082
rect 21794 13030 21806 13082
rect 21858 13030 21870 13082
rect 21922 13030 21934 13082
rect 21986 13030 21998 13082
rect 22050 13030 22056 13082
rect 1104 13008 22056 13030
rect 5077 12971 5135 12977
rect 5077 12937 5089 12971
rect 5123 12968 5135 12971
rect 5445 12971 5503 12977
rect 5445 12968 5457 12971
rect 5123 12940 5457 12968
rect 5123 12937 5135 12940
rect 5077 12931 5135 12937
rect 5445 12937 5457 12940
rect 5491 12937 5503 12971
rect 5445 12931 5503 12937
rect 5905 12971 5963 12977
rect 5905 12937 5917 12971
rect 5951 12968 5963 12971
rect 6365 12971 6423 12977
rect 6365 12968 6377 12971
rect 5951 12940 6377 12968
rect 5951 12937 5963 12940
rect 5905 12931 5963 12937
rect 6365 12937 6377 12940
rect 6411 12937 6423 12971
rect 6365 12931 6423 12937
rect 6733 12971 6791 12977
rect 6733 12937 6745 12971
rect 6779 12968 6791 12971
rect 6822 12968 6828 12980
rect 6779 12940 6828 12968
rect 6779 12937 6791 12940
rect 6733 12931 6791 12937
rect 6822 12928 6828 12940
rect 6880 12928 6886 12980
rect 7285 12971 7343 12977
rect 7285 12937 7297 12971
rect 7331 12968 7343 12971
rect 8202 12968 8208 12980
rect 7331 12940 8208 12968
rect 7331 12937 7343 12940
rect 7285 12931 7343 12937
rect 3326 12900 3332 12912
rect 3287 12872 3332 12900
rect 3326 12860 3332 12872
rect 3384 12860 3390 12912
rect 4246 12900 4252 12912
rect 4207 12872 4252 12900
rect 4246 12860 4252 12872
rect 4304 12860 4310 12912
rect 3605 12835 3663 12841
rect 3605 12801 3617 12835
rect 3651 12801 3663 12835
rect 4522 12832 4528 12844
rect 4483 12804 4528 12832
rect 3605 12795 3663 12801
rect 3620 12696 3648 12795
rect 4522 12792 4528 12804
rect 4580 12792 4586 12844
rect 4985 12835 5043 12841
rect 4985 12801 4997 12835
rect 5031 12832 5043 12835
rect 5626 12832 5632 12844
rect 5031 12804 5632 12832
rect 5031 12801 5043 12804
rect 4985 12795 5043 12801
rect 5626 12792 5632 12804
rect 5684 12792 5690 12844
rect 5810 12832 5816 12844
rect 5771 12804 5816 12832
rect 5810 12792 5816 12804
rect 5868 12792 5874 12844
rect 6825 12835 6883 12841
rect 6825 12832 6837 12835
rect 5920 12804 6837 12832
rect 5258 12764 5264 12776
rect 5219 12736 5264 12764
rect 5258 12724 5264 12736
rect 5316 12724 5322 12776
rect 5442 12724 5448 12776
rect 5500 12764 5506 12776
rect 5920 12764 5948 12804
rect 6825 12801 6837 12804
rect 6871 12801 6883 12835
rect 6825 12795 6883 12801
rect 5500 12736 5948 12764
rect 6089 12767 6147 12773
rect 5500 12724 5506 12736
rect 6089 12733 6101 12767
rect 6135 12764 6147 12767
rect 6546 12764 6552 12776
rect 6135 12736 6552 12764
rect 6135 12733 6147 12736
rect 6089 12727 6147 12733
rect 6546 12724 6552 12736
rect 6604 12724 6610 12776
rect 7009 12767 7067 12773
rect 7009 12733 7021 12767
rect 7055 12764 7067 12767
rect 7098 12764 7104 12776
rect 7055 12736 7104 12764
rect 7055 12733 7067 12736
rect 7009 12727 7067 12733
rect 7098 12724 7104 12736
rect 7156 12764 7162 12776
rect 7300 12764 7328 12931
rect 8202 12928 8208 12940
rect 8260 12928 8266 12980
rect 8386 12928 8392 12980
rect 8444 12968 8450 12980
rect 8573 12971 8631 12977
rect 8573 12968 8585 12971
rect 8444 12940 8585 12968
rect 8444 12928 8450 12940
rect 8573 12937 8585 12940
rect 8619 12937 8631 12971
rect 9950 12968 9956 12980
rect 9911 12940 9956 12968
rect 8573 12931 8631 12937
rect 9950 12928 9956 12940
rect 10008 12928 10014 12980
rect 10410 12968 10416 12980
rect 10371 12940 10416 12968
rect 10410 12928 10416 12940
rect 10468 12928 10474 12980
rect 14090 12928 14096 12980
rect 14148 12968 14154 12980
rect 14826 12968 14832 12980
rect 14148 12940 14832 12968
rect 14148 12928 14154 12940
rect 14826 12928 14832 12940
rect 14884 12968 14890 12980
rect 18046 12968 18052 12980
rect 14884 12940 16620 12968
rect 18007 12940 18052 12968
rect 14884 12928 14890 12940
rect 10321 12903 10379 12909
rect 10321 12900 10333 12903
rect 8404 12872 10333 12900
rect 8404 12844 8432 12872
rect 10321 12869 10333 12872
rect 10367 12869 10379 12903
rect 10321 12863 10379 12869
rect 14274 12860 14280 12912
rect 14332 12900 14338 12912
rect 16592 12900 16620 12940
rect 18046 12928 18052 12940
rect 18104 12928 18110 12980
rect 19518 12968 19524 12980
rect 19479 12940 19524 12968
rect 19518 12928 19524 12940
rect 19576 12928 19582 12980
rect 20714 12928 20720 12980
rect 20772 12968 20778 12980
rect 21085 12971 21143 12977
rect 21085 12968 21097 12971
rect 20772 12940 21097 12968
rect 20772 12928 20778 12940
rect 16914 12903 16972 12909
rect 16914 12900 16926 12903
rect 14332 12872 15608 12900
rect 16592 12872 16926 12900
rect 14332 12860 14338 12872
rect 7561 12835 7619 12841
rect 7561 12801 7573 12835
rect 7607 12832 7619 12835
rect 8021 12835 8079 12841
rect 8021 12832 8033 12835
rect 7607 12804 8033 12832
rect 7607 12801 7619 12804
rect 7561 12795 7619 12801
rect 8021 12801 8033 12804
rect 8067 12801 8079 12835
rect 8021 12795 8079 12801
rect 8386 12792 8392 12844
rect 8444 12792 8450 12844
rect 8941 12835 8999 12841
rect 8941 12801 8953 12835
rect 8987 12832 8999 12835
rect 9582 12832 9588 12844
rect 8987 12804 9588 12832
rect 8987 12801 8999 12804
rect 8941 12795 8999 12801
rect 9582 12792 9588 12804
rect 9640 12792 9646 12844
rect 12066 12792 12072 12844
rect 12124 12832 12130 12844
rect 13826 12835 13884 12841
rect 13826 12832 13838 12835
rect 12124 12804 13838 12832
rect 12124 12792 12130 12804
rect 13826 12801 13838 12804
rect 13872 12801 13884 12835
rect 13826 12795 13884 12801
rect 14366 12792 14372 12844
rect 14424 12832 14430 12844
rect 15580 12841 15608 12872
rect 16914 12869 16926 12872
rect 16960 12869 16972 12903
rect 16914 12863 16972 12869
rect 15298 12835 15356 12841
rect 15298 12832 15310 12835
rect 14424 12804 15310 12832
rect 14424 12792 14430 12804
rect 15298 12801 15310 12804
rect 15344 12801 15356 12835
rect 15298 12795 15356 12801
rect 15565 12835 15623 12841
rect 15565 12801 15577 12835
rect 15611 12832 15623 12835
rect 15657 12835 15715 12841
rect 15657 12832 15669 12835
rect 15611 12804 15669 12832
rect 15611 12801 15623 12804
rect 15565 12795 15623 12801
rect 15657 12801 15669 12804
rect 15703 12832 15715 12835
rect 15930 12832 15936 12844
rect 15703 12804 15936 12832
rect 15703 12801 15715 12804
rect 15657 12795 15715 12801
rect 15930 12792 15936 12804
rect 15988 12832 15994 12844
rect 16666 12832 16672 12844
rect 15988 12804 16672 12832
rect 15988 12792 15994 12804
rect 16666 12792 16672 12804
rect 16724 12792 16730 12844
rect 17494 12792 17500 12844
rect 17552 12832 17558 12844
rect 18397 12835 18455 12841
rect 18397 12832 18409 12835
rect 17552 12804 18409 12832
rect 17552 12792 17558 12804
rect 7742 12764 7748 12776
rect 7156 12736 7328 12764
rect 7703 12736 7748 12764
rect 7156 12724 7162 12736
rect 7742 12724 7748 12736
rect 7800 12724 7806 12776
rect 7834 12724 7840 12776
rect 7892 12764 7898 12776
rect 7929 12767 7987 12773
rect 7929 12764 7941 12767
rect 7892 12736 7941 12764
rect 7892 12724 7898 12736
rect 7929 12733 7941 12736
rect 7975 12733 7987 12767
rect 7929 12727 7987 12733
rect 8294 12724 8300 12776
rect 8352 12764 8358 12776
rect 9033 12767 9091 12773
rect 9033 12764 9045 12767
rect 8352 12736 9045 12764
rect 8352 12724 8358 12736
rect 9033 12733 9045 12736
rect 9079 12733 9091 12767
rect 9033 12727 9091 12733
rect 9217 12767 9275 12773
rect 9217 12733 9229 12767
rect 9263 12764 9275 12767
rect 10597 12767 10655 12773
rect 9263 12736 10548 12764
rect 9263 12733 9275 12736
rect 9217 12727 9275 12733
rect 4617 12699 4675 12705
rect 4617 12696 4629 12699
rect 3620 12668 4629 12696
rect 4617 12665 4629 12668
rect 4663 12665 4675 12699
rect 4617 12659 4675 12665
rect 5534 12656 5540 12708
rect 5592 12696 5598 12708
rect 6730 12696 6736 12708
rect 5592 12668 6736 12696
rect 5592 12656 5598 12668
rect 6730 12656 6736 12668
rect 6788 12656 6794 12708
rect 8389 12699 8447 12705
rect 8389 12665 8401 12699
rect 8435 12696 8447 12699
rect 9766 12696 9772 12708
rect 8435 12668 9772 12696
rect 8435 12665 8447 12668
rect 8389 12659 8447 12665
rect 9766 12656 9772 12668
rect 9824 12656 9830 12708
rect 10520 12696 10548 12736
rect 10597 12733 10609 12767
rect 10643 12764 10655 12767
rect 11882 12764 11888 12776
rect 10643 12736 11888 12764
rect 10643 12733 10655 12736
rect 10597 12727 10655 12733
rect 11882 12724 11888 12736
rect 11940 12724 11946 12776
rect 14093 12767 14151 12773
rect 14093 12733 14105 12767
rect 14139 12764 14151 12767
rect 14274 12764 14280 12776
rect 14139 12736 14280 12764
rect 14139 12733 14151 12736
rect 14093 12727 14151 12733
rect 14274 12724 14280 12736
rect 14332 12724 14338 12776
rect 10870 12696 10876 12708
rect 10520 12668 10876 12696
rect 10870 12656 10876 12668
rect 10928 12696 10934 12708
rect 10928 12668 13216 12696
rect 10928 12656 10934 12668
rect 3326 12588 3332 12640
rect 3384 12628 3390 12640
rect 4246 12628 4252 12640
rect 3384 12600 4252 12628
rect 3384 12588 3390 12600
rect 4246 12588 4252 12600
rect 4304 12588 4310 12640
rect 6546 12588 6552 12640
rect 6604 12628 6610 12640
rect 12250 12628 12256 12640
rect 6604 12600 12256 12628
rect 6604 12588 6610 12600
rect 12250 12588 12256 12600
rect 12308 12588 12314 12640
rect 12526 12628 12532 12640
rect 12487 12600 12532 12628
rect 12526 12588 12532 12600
rect 12584 12588 12590 12640
rect 12710 12628 12716 12640
rect 12671 12600 12716 12628
rect 12710 12588 12716 12600
rect 12768 12588 12774 12640
rect 13188 12628 13216 12668
rect 14108 12668 14688 12696
rect 14108 12628 14136 12668
rect 13188 12600 14136 12628
rect 14185 12631 14243 12637
rect 14185 12597 14197 12631
rect 14231 12628 14243 12631
rect 14550 12628 14556 12640
rect 14231 12600 14556 12628
rect 14231 12597 14243 12600
rect 14185 12591 14243 12597
rect 14550 12588 14556 12600
rect 14608 12588 14614 12640
rect 14660 12628 14688 12668
rect 17696 12628 17724 12804
rect 18397 12801 18409 12804
rect 18443 12801 18455 12835
rect 18397 12795 18455 12801
rect 20737 12835 20795 12841
rect 20737 12801 20749 12835
rect 20783 12832 20795 12835
rect 20898 12832 20904 12844
rect 20783 12804 20904 12832
rect 20783 12801 20795 12804
rect 20737 12795 20795 12801
rect 20898 12792 20904 12804
rect 20956 12792 20962 12844
rect 21008 12841 21036 12940
rect 21085 12937 21097 12940
rect 21131 12968 21143 12971
rect 21266 12968 21272 12980
rect 21131 12940 21272 12968
rect 21131 12937 21143 12940
rect 21085 12931 21143 12937
rect 21266 12928 21272 12940
rect 21324 12968 21330 12980
rect 21361 12971 21419 12977
rect 21361 12968 21373 12971
rect 21324 12940 21373 12968
rect 21324 12928 21330 12940
rect 21361 12937 21373 12940
rect 21407 12937 21419 12971
rect 21361 12931 21419 12937
rect 20993 12835 21051 12841
rect 20993 12801 21005 12835
rect 21039 12801 21051 12835
rect 20993 12795 21051 12801
rect 18138 12764 18144 12776
rect 18099 12736 18144 12764
rect 18138 12724 18144 12736
rect 18196 12724 18202 12776
rect 14660 12600 17724 12628
rect 19610 12588 19616 12640
rect 19668 12628 19674 12640
rect 19668 12600 19713 12628
rect 19668 12588 19674 12600
rect 1104 12538 21896 12560
rect 1104 12486 3549 12538
rect 3601 12486 3613 12538
rect 3665 12486 3677 12538
rect 3729 12486 3741 12538
rect 3793 12486 3805 12538
rect 3857 12486 8747 12538
rect 8799 12486 8811 12538
rect 8863 12486 8875 12538
rect 8927 12486 8939 12538
rect 8991 12486 9003 12538
rect 9055 12486 13945 12538
rect 13997 12486 14009 12538
rect 14061 12486 14073 12538
rect 14125 12486 14137 12538
rect 14189 12486 14201 12538
rect 14253 12486 19143 12538
rect 19195 12486 19207 12538
rect 19259 12486 19271 12538
rect 19323 12486 19335 12538
rect 19387 12486 19399 12538
rect 19451 12486 21896 12538
rect 1104 12464 21896 12486
rect 1949 12427 2007 12433
rect 1949 12393 1961 12427
rect 1995 12424 2007 12427
rect 2866 12424 2872 12436
rect 1995 12396 2872 12424
rect 1995 12393 2007 12396
rect 1949 12387 2007 12393
rect 2866 12384 2872 12396
rect 2924 12384 2930 12436
rect 5626 12424 5632 12436
rect 5587 12396 5632 12424
rect 5626 12384 5632 12396
rect 5684 12384 5690 12436
rect 6822 12384 6828 12436
rect 6880 12424 6886 12436
rect 7282 12424 7288 12436
rect 6880 12396 7288 12424
rect 6880 12384 6886 12396
rect 7282 12384 7288 12396
rect 7340 12384 7346 12436
rect 7469 12427 7527 12433
rect 7469 12393 7481 12427
rect 7515 12424 7527 12427
rect 7650 12424 7656 12436
rect 7515 12396 7656 12424
rect 7515 12393 7527 12396
rect 7469 12387 7527 12393
rect 7650 12384 7656 12396
rect 7708 12384 7714 12436
rect 7742 12384 7748 12436
rect 7800 12424 7806 12436
rect 8294 12424 8300 12436
rect 7800 12396 8300 12424
rect 7800 12384 7806 12396
rect 8294 12384 8300 12396
rect 8352 12424 8358 12436
rect 8389 12427 8447 12433
rect 8389 12424 8401 12427
rect 8352 12396 8401 12424
rect 8352 12384 8358 12396
rect 8389 12393 8401 12396
rect 8435 12393 8447 12427
rect 8389 12387 8447 12393
rect 9306 12384 9312 12436
rect 9364 12424 9370 12436
rect 10229 12427 10287 12433
rect 10229 12424 10241 12427
rect 9364 12396 10241 12424
rect 9364 12384 9370 12396
rect 10229 12393 10241 12396
rect 10275 12393 10287 12427
rect 10229 12387 10287 12393
rect 10594 12384 10600 12436
rect 10652 12424 10658 12436
rect 18141 12427 18199 12433
rect 18141 12424 18153 12427
rect 10652 12396 18153 12424
rect 10652 12384 10658 12396
rect 18141 12393 18153 12396
rect 18187 12393 18199 12427
rect 18141 12387 18199 12393
rect 4522 12316 4528 12368
rect 4580 12356 4586 12368
rect 8941 12359 8999 12365
rect 8941 12356 8953 12359
rect 4580 12328 8953 12356
rect 4580 12316 4586 12328
rect 8941 12325 8953 12328
rect 8987 12325 8999 12359
rect 8941 12319 8999 12325
rect 10962 12316 10968 12368
rect 11020 12356 11026 12368
rect 11146 12356 11152 12368
rect 11020 12328 11152 12356
rect 11020 12316 11026 12328
rect 11146 12316 11152 12328
rect 11204 12316 11210 12368
rect 14642 12316 14648 12368
rect 14700 12356 14706 12368
rect 15289 12359 15347 12365
rect 15289 12356 15301 12359
rect 14700 12328 15301 12356
rect 14700 12316 14706 12328
rect 15289 12325 15301 12328
rect 15335 12325 15347 12359
rect 15289 12319 15347 12325
rect 4982 12248 4988 12300
rect 5040 12288 5046 12300
rect 5077 12291 5135 12297
rect 5077 12288 5089 12291
rect 5040 12260 5089 12288
rect 5040 12248 5046 12260
rect 5077 12257 5089 12260
rect 5123 12257 5135 12291
rect 5077 12251 5135 12257
rect 6273 12291 6331 12297
rect 6273 12257 6285 12291
rect 6319 12288 6331 12291
rect 6546 12288 6552 12300
rect 6319 12260 6552 12288
rect 6319 12257 6331 12260
rect 6273 12251 6331 12257
rect 6546 12248 6552 12260
rect 6604 12248 6610 12300
rect 6638 12248 6644 12300
rect 6696 12288 6702 12300
rect 8018 12288 8024 12300
rect 6696 12260 8024 12288
rect 6696 12248 6702 12260
rect 8018 12248 8024 12260
rect 8076 12288 8082 12300
rect 8573 12291 8631 12297
rect 8573 12288 8585 12291
rect 8076 12260 8585 12288
rect 8076 12248 8082 12260
rect 8573 12257 8585 12260
rect 8619 12257 8631 12291
rect 9490 12288 9496 12300
rect 9451 12260 9496 12288
rect 8573 12251 8631 12257
rect 9490 12248 9496 12260
rect 9548 12248 9554 12300
rect 9582 12248 9588 12300
rect 9640 12288 9646 12300
rect 9769 12291 9827 12297
rect 9769 12288 9781 12291
rect 9640 12260 9781 12288
rect 9640 12248 9646 12260
rect 9769 12257 9781 12260
rect 9815 12257 9827 12291
rect 10870 12288 10876 12300
rect 10831 12260 10876 12288
rect 9769 12251 9827 12257
rect 10870 12248 10876 12260
rect 10928 12248 10934 12300
rect 12437 12291 12495 12297
rect 12437 12257 12449 12291
rect 12483 12288 12495 12291
rect 12526 12288 12532 12300
rect 12483 12260 12532 12288
rect 12483 12257 12495 12260
rect 12437 12251 12495 12257
rect 12526 12248 12532 12260
rect 12584 12248 12590 12300
rect 16666 12288 16672 12300
rect 16627 12260 16672 12288
rect 16666 12248 16672 12260
rect 16724 12288 16730 12300
rect 16761 12291 16819 12297
rect 16761 12288 16773 12291
rect 16724 12260 16773 12288
rect 16724 12248 16730 12260
rect 16761 12257 16773 12260
rect 16807 12257 16819 12291
rect 18156 12288 18184 12387
rect 18230 12384 18236 12436
rect 18288 12424 18294 12436
rect 18417 12427 18475 12433
rect 18417 12424 18429 12427
rect 18288 12396 18429 12424
rect 18288 12384 18294 12396
rect 18417 12393 18429 12396
rect 18463 12393 18475 12427
rect 19702 12424 19708 12436
rect 19663 12396 19708 12424
rect 18417 12387 18475 12393
rect 19702 12384 19708 12396
rect 19760 12384 19766 12436
rect 21266 12424 21272 12436
rect 21227 12396 21272 12424
rect 21266 12384 21272 12396
rect 21324 12384 21330 12436
rect 21177 12291 21235 12297
rect 18156 12260 20024 12288
rect 16761 12251 16819 12257
rect 2133 12223 2191 12229
rect 2133 12189 2145 12223
rect 2179 12220 2191 12223
rect 4062 12220 4068 12232
rect 2179 12192 4068 12220
rect 2179 12189 2191 12192
rect 2133 12183 2191 12189
rect 4062 12180 4068 12192
rect 4120 12180 4126 12232
rect 5353 12223 5411 12229
rect 5353 12189 5365 12223
rect 5399 12220 5411 12223
rect 9306 12220 9312 12232
rect 5399 12192 9312 12220
rect 5399 12189 5411 12192
rect 5353 12183 5411 12189
rect 9306 12180 9312 12192
rect 9364 12180 9370 12232
rect 10597 12223 10655 12229
rect 10597 12189 10609 12223
rect 10643 12220 10655 12223
rect 11146 12220 11152 12232
rect 10643 12192 11152 12220
rect 10643 12189 10655 12192
rect 10597 12183 10655 12189
rect 11146 12180 11152 12192
rect 11204 12220 11210 12232
rect 11790 12220 11796 12232
rect 11204 12192 11796 12220
rect 11204 12180 11210 12192
rect 11790 12180 11796 12192
rect 11848 12180 11854 12232
rect 11882 12180 11888 12232
rect 11940 12220 11946 12232
rect 12170 12223 12228 12229
rect 12170 12220 12182 12223
rect 11940 12192 12182 12220
rect 11940 12180 11946 12192
rect 12170 12189 12182 12192
rect 12216 12189 12228 12223
rect 12170 12183 12228 12189
rect 13906 12180 13912 12232
rect 13964 12220 13970 12232
rect 14366 12220 14372 12232
rect 13964 12192 14372 12220
rect 13964 12180 13970 12192
rect 14366 12180 14372 12192
rect 14424 12180 14430 12232
rect 14918 12180 14924 12232
rect 14976 12220 14982 12232
rect 16402 12223 16460 12229
rect 16402 12220 16414 12223
rect 14976 12192 16414 12220
rect 14976 12180 14982 12192
rect 16402 12189 16414 12192
rect 16448 12189 16460 12223
rect 19996 12220 20024 12260
rect 21177 12257 21189 12291
rect 21223 12288 21235 12291
rect 21284 12288 21312 12384
rect 21223 12260 21312 12288
rect 21223 12257 21235 12260
rect 21177 12251 21235 12257
rect 20910 12223 20968 12229
rect 20910 12220 20922 12223
rect 19996 12192 20922 12220
rect 16402 12183 16460 12189
rect 20910 12189 20922 12192
rect 20956 12189 20968 12223
rect 20910 12183 20968 12189
rect 5442 12112 5448 12164
rect 5500 12152 5506 12164
rect 7190 12152 7196 12164
rect 5500 12124 7196 12152
rect 5500 12112 5506 12124
rect 7190 12112 7196 12124
rect 7248 12112 7254 12164
rect 7650 12112 7656 12164
rect 7708 12152 7714 12164
rect 10689 12155 10747 12161
rect 7708 12124 10640 12152
rect 7708 12112 7714 12124
rect 5994 12084 6000 12096
rect 5955 12056 6000 12084
rect 5994 12044 6000 12056
rect 6052 12044 6058 12096
rect 6089 12087 6147 12093
rect 6089 12053 6101 12087
rect 6135 12084 6147 12087
rect 6546 12084 6552 12096
rect 6135 12056 6552 12084
rect 6135 12053 6147 12056
rect 6089 12047 6147 12053
rect 6546 12044 6552 12056
rect 6604 12044 6610 12096
rect 7282 12084 7288 12096
rect 7243 12056 7288 12084
rect 7282 12044 7288 12056
rect 7340 12084 7346 12096
rect 7837 12087 7895 12093
rect 7837 12084 7849 12087
rect 7340 12056 7849 12084
rect 7340 12044 7346 12056
rect 7837 12053 7849 12056
rect 7883 12053 7895 12087
rect 7837 12047 7895 12053
rect 7929 12087 7987 12093
rect 7929 12053 7941 12087
rect 7975 12084 7987 12087
rect 8294 12084 8300 12096
rect 7975 12056 8300 12084
rect 7975 12053 7987 12056
rect 7929 12047 7987 12053
rect 8294 12044 8300 12056
rect 8352 12044 8358 12096
rect 9122 12044 9128 12096
rect 9180 12084 9186 12096
rect 9309 12087 9367 12093
rect 9309 12084 9321 12087
rect 9180 12056 9321 12084
rect 9180 12044 9186 12056
rect 9309 12053 9321 12056
rect 9355 12053 9367 12087
rect 9309 12047 9367 12053
rect 9401 12087 9459 12093
rect 9401 12053 9413 12087
rect 9447 12084 9459 12087
rect 10042 12084 10048 12096
rect 9447 12056 10048 12084
rect 9447 12053 9459 12056
rect 9401 12047 9459 12053
rect 10042 12044 10048 12056
rect 10100 12044 10106 12096
rect 10612 12084 10640 12124
rect 10689 12121 10701 12155
rect 10735 12152 10747 12155
rect 11698 12152 11704 12164
rect 10735 12124 11704 12152
rect 10735 12121 10747 12124
rect 10689 12115 10747 12121
rect 11698 12112 11704 12124
rect 11756 12112 11762 12164
rect 11974 12112 11980 12164
rect 12032 12152 12038 12164
rect 12250 12152 12256 12164
rect 12032 12124 12256 12152
rect 12032 12112 12038 12124
rect 12250 12112 12256 12124
rect 12308 12112 12314 12164
rect 12618 12112 12624 12164
rect 12676 12152 12682 12164
rect 12774 12155 12832 12161
rect 12774 12152 12786 12155
rect 12676 12124 12786 12152
rect 12676 12112 12682 12124
rect 12774 12121 12786 12124
rect 12820 12121 12832 12155
rect 14642 12152 14648 12164
rect 12774 12115 12832 12121
rect 13004 12124 14648 12152
rect 13004 12096 13032 12124
rect 14642 12112 14648 12124
rect 14700 12112 14706 12164
rect 16574 12112 16580 12164
rect 16632 12152 16638 12164
rect 17006 12155 17064 12161
rect 17006 12152 17018 12155
rect 16632 12124 17018 12152
rect 16632 12112 16638 12124
rect 17006 12121 17018 12124
rect 17052 12121 17064 12155
rect 17006 12115 17064 12121
rect 11057 12087 11115 12093
rect 11057 12084 11069 12087
rect 10612 12056 11069 12084
rect 11057 12053 11069 12056
rect 11103 12084 11115 12087
rect 12526 12084 12532 12096
rect 11103 12056 12532 12084
rect 11103 12053 11115 12056
rect 11057 12047 11115 12053
rect 12526 12044 12532 12056
rect 12584 12044 12590 12096
rect 12986 12044 12992 12096
rect 13044 12044 13050 12096
rect 13906 12084 13912 12096
rect 13867 12056 13912 12084
rect 13906 12044 13912 12056
rect 13964 12044 13970 12096
rect 14182 12084 14188 12096
rect 14143 12056 14188 12084
rect 14182 12044 14188 12056
rect 14240 12084 14246 12096
rect 14369 12087 14427 12093
rect 14369 12084 14381 12087
rect 14240 12056 14381 12084
rect 14240 12044 14246 12056
rect 14369 12053 14381 12056
rect 14415 12053 14427 12087
rect 14369 12047 14427 12053
rect 14734 12044 14740 12096
rect 14792 12084 14798 12096
rect 19797 12087 19855 12093
rect 19797 12084 19809 12087
rect 14792 12056 19809 12084
rect 14792 12044 14798 12056
rect 19797 12053 19809 12056
rect 19843 12053 19855 12087
rect 19797 12047 19855 12053
rect 1104 11994 22056 12016
rect 1104 11942 6148 11994
rect 6200 11942 6212 11994
rect 6264 11942 6276 11994
rect 6328 11942 6340 11994
rect 6392 11942 6404 11994
rect 6456 11942 11346 11994
rect 11398 11942 11410 11994
rect 11462 11942 11474 11994
rect 11526 11942 11538 11994
rect 11590 11942 11602 11994
rect 11654 11942 16544 11994
rect 16596 11942 16608 11994
rect 16660 11942 16672 11994
rect 16724 11942 16736 11994
rect 16788 11942 16800 11994
rect 16852 11942 21742 11994
rect 21794 11942 21806 11994
rect 21858 11942 21870 11994
rect 21922 11942 21934 11994
rect 21986 11942 21998 11994
rect 22050 11942 22056 11994
rect 1104 11920 22056 11942
rect 5442 11880 5448 11892
rect 5403 11852 5448 11880
rect 5442 11840 5448 11852
rect 5500 11840 5506 11892
rect 6365 11883 6423 11889
rect 6365 11849 6377 11883
rect 6411 11880 6423 11883
rect 6546 11880 6552 11892
rect 6411 11852 6552 11880
rect 6411 11849 6423 11852
rect 6365 11843 6423 11849
rect 6546 11840 6552 11852
rect 6604 11840 6610 11892
rect 6825 11883 6883 11889
rect 6825 11880 6837 11883
rect 6656 11852 6837 11880
rect 4154 11812 4160 11824
rect 4115 11784 4160 11812
rect 4154 11772 4160 11784
rect 4212 11772 4218 11824
rect 4430 11744 4436 11756
rect 4391 11716 4436 11744
rect 4430 11704 4436 11716
rect 4488 11704 4494 11756
rect 6181 11747 6239 11753
rect 6181 11713 6193 11747
rect 6227 11744 6239 11747
rect 6656 11744 6684 11852
rect 6825 11849 6837 11852
rect 6871 11880 6883 11883
rect 6914 11880 6920 11892
rect 6871 11852 6920 11880
rect 6871 11849 6883 11852
rect 6825 11843 6883 11849
rect 6914 11840 6920 11852
rect 6972 11840 6978 11892
rect 7098 11840 7104 11892
rect 7156 11880 7162 11892
rect 7193 11883 7251 11889
rect 7193 11880 7205 11883
rect 7156 11852 7205 11880
rect 7156 11840 7162 11852
rect 7193 11849 7205 11852
rect 7239 11849 7251 11883
rect 9306 11880 9312 11892
rect 9267 11852 9312 11880
rect 7193 11843 7251 11849
rect 9306 11840 9312 11852
rect 9364 11840 9370 11892
rect 9769 11883 9827 11889
rect 9769 11849 9781 11883
rect 9815 11880 9827 11883
rect 10137 11883 10195 11889
rect 10137 11880 10149 11883
rect 9815 11852 10149 11880
rect 9815 11849 9827 11852
rect 9769 11843 9827 11849
rect 10137 11849 10149 11852
rect 10183 11849 10195 11883
rect 10137 11843 10195 11849
rect 10597 11883 10655 11889
rect 10597 11849 10609 11883
rect 10643 11880 10655 11883
rect 10962 11880 10968 11892
rect 10643 11852 10968 11880
rect 10643 11849 10655 11852
rect 10597 11843 10655 11849
rect 10962 11840 10968 11852
rect 11020 11840 11026 11892
rect 11238 11840 11244 11892
rect 11296 11880 11302 11892
rect 11517 11883 11575 11889
rect 11517 11880 11529 11883
rect 11296 11852 11529 11880
rect 11296 11840 11302 11852
rect 11517 11849 11529 11852
rect 11563 11849 11575 11883
rect 13814 11880 13820 11892
rect 11517 11843 11575 11849
rect 11808 11852 13820 11880
rect 7926 11772 7932 11824
rect 7984 11812 7990 11824
rect 8202 11812 8208 11824
rect 7984 11784 8208 11812
rect 7984 11772 7990 11784
rect 8202 11772 8208 11784
rect 8260 11772 8266 11824
rect 10505 11815 10563 11821
rect 10505 11781 10517 11815
rect 10551 11812 10563 11815
rect 11054 11812 11060 11824
rect 10551 11784 11060 11812
rect 10551 11781 10563 11784
rect 10505 11775 10563 11781
rect 11054 11772 11060 11784
rect 11112 11772 11118 11824
rect 11333 11815 11391 11821
rect 11333 11781 11345 11815
rect 11379 11812 11391 11815
rect 11698 11812 11704 11824
rect 11379 11784 11704 11812
rect 11379 11781 11391 11784
rect 11333 11775 11391 11781
rect 11698 11772 11704 11784
rect 11756 11772 11762 11824
rect 6227 11716 6684 11744
rect 6733 11747 6791 11753
rect 6227 11713 6239 11716
rect 6181 11707 6239 11713
rect 6733 11713 6745 11747
rect 6779 11713 6791 11747
rect 8018 11744 8024 11756
rect 7979 11716 8024 11744
rect 6733 11707 6791 11713
rect 4982 11636 4988 11688
rect 5040 11676 5046 11688
rect 5169 11679 5227 11685
rect 5169 11676 5181 11679
rect 5040 11648 5181 11676
rect 5040 11636 5046 11648
rect 5169 11645 5181 11648
rect 5215 11645 5227 11679
rect 5169 11639 5227 11645
rect 5997 11679 6055 11685
rect 5997 11645 6009 11679
rect 6043 11676 6055 11679
rect 6638 11676 6644 11688
rect 6043 11648 6644 11676
rect 6043 11645 6055 11648
rect 5997 11639 6055 11645
rect 6638 11636 6644 11648
rect 6696 11676 6702 11688
rect 6748 11676 6776 11707
rect 8018 11704 8024 11716
rect 8076 11704 8082 11756
rect 9674 11744 9680 11756
rect 9635 11716 9680 11744
rect 9674 11704 9680 11716
rect 9732 11704 9738 11756
rect 10686 11704 10692 11756
rect 10744 11744 10750 11756
rect 11808 11744 11836 11852
rect 13814 11840 13820 11852
rect 13872 11840 13878 11892
rect 18230 11840 18236 11892
rect 18288 11880 18294 11892
rect 18969 11883 19027 11889
rect 18969 11880 18981 11883
rect 18288 11852 18981 11880
rect 18288 11840 18294 11852
rect 18969 11849 18981 11852
rect 19015 11849 19027 11883
rect 18969 11843 19027 11849
rect 20901 11883 20959 11889
rect 20901 11849 20913 11883
rect 20947 11880 20959 11883
rect 21266 11880 21272 11892
rect 20947 11852 21272 11880
rect 20947 11849 20959 11852
rect 20901 11843 20959 11849
rect 11974 11772 11980 11824
rect 12032 11812 12038 11824
rect 13664 11815 13722 11821
rect 13664 11812 13676 11815
rect 12032 11784 13676 11812
rect 12032 11772 12038 11784
rect 13664 11781 13676 11784
rect 13710 11812 13722 11815
rect 14550 11812 14556 11824
rect 13710 11784 14556 11812
rect 13710 11781 13722 11784
rect 13664 11775 13722 11781
rect 14550 11772 14556 11784
rect 14608 11772 14614 11824
rect 10744 11716 11836 11744
rect 10744 11704 10750 11716
rect 11882 11704 11888 11756
rect 11940 11744 11946 11756
rect 12710 11744 12716 11756
rect 11940 11716 12716 11744
rect 11940 11704 11946 11716
rect 12710 11704 12716 11716
rect 12768 11704 12774 11756
rect 15102 11744 15108 11756
rect 12912 11716 15108 11744
rect 6696 11648 6776 11676
rect 7009 11679 7067 11685
rect 6696 11636 6702 11648
rect 7009 11645 7021 11679
rect 7055 11676 7067 11679
rect 7098 11676 7104 11688
rect 7055 11648 7104 11676
rect 7055 11645 7067 11648
rect 7009 11639 7067 11645
rect 5626 11568 5632 11620
rect 5684 11608 5690 11620
rect 7024 11608 7052 11639
rect 7098 11636 7104 11648
rect 7156 11636 7162 11688
rect 7466 11636 7472 11688
rect 7524 11676 7530 11688
rect 7745 11679 7803 11685
rect 7745 11676 7757 11679
rect 7524 11648 7757 11676
rect 7524 11636 7530 11648
rect 7745 11645 7757 11648
rect 7791 11645 7803 11679
rect 7926 11676 7932 11688
rect 7887 11648 7932 11676
rect 7745 11639 7803 11645
rect 7926 11636 7932 11648
rect 7984 11636 7990 11688
rect 9950 11676 9956 11688
rect 9911 11648 9956 11676
rect 9950 11636 9956 11648
rect 10008 11636 10014 11688
rect 10778 11676 10784 11688
rect 10739 11648 10784 11676
rect 10778 11636 10784 11648
rect 10836 11636 10842 11688
rect 11330 11636 11336 11688
rect 11388 11676 11394 11688
rect 11977 11679 12035 11685
rect 11977 11676 11989 11679
rect 11388 11648 11989 11676
rect 11388 11636 11394 11648
rect 11977 11645 11989 11648
rect 12023 11645 12035 11679
rect 11977 11639 12035 11645
rect 12161 11679 12219 11685
rect 12161 11645 12173 11679
rect 12207 11676 12219 11679
rect 12250 11676 12256 11688
rect 12207 11648 12256 11676
rect 12207 11645 12219 11648
rect 12161 11639 12219 11645
rect 12250 11636 12256 11648
rect 12308 11676 12314 11688
rect 12345 11679 12403 11685
rect 12345 11676 12357 11679
rect 12308 11648 12357 11676
rect 12308 11636 12314 11648
rect 12345 11645 12357 11648
rect 12391 11676 12403 11679
rect 12912 11676 12940 11716
rect 15102 11704 15108 11716
rect 15160 11704 15166 11756
rect 16390 11704 16396 11756
rect 16448 11744 16454 11756
rect 17753 11747 17811 11753
rect 17753 11744 17765 11747
rect 16448 11716 17765 11744
rect 16448 11704 16454 11716
rect 17753 11713 17765 11716
rect 17799 11713 17811 11747
rect 17753 11707 17811 11713
rect 19886 11704 19892 11756
rect 19944 11744 19950 11756
rect 20450 11747 20508 11753
rect 20450 11744 20462 11747
rect 19944 11716 20462 11744
rect 19944 11704 19950 11716
rect 20450 11713 20462 11716
rect 20496 11713 20508 11747
rect 20450 11707 20508 11713
rect 20717 11747 20775 11753
rect 20717 11713 20729 11747
rect 20763 11744 20775 11747
rect 20916 11744 20944 11843
rect 21266 11840 21272 11852
rect 21324 11840 21330 11892
rect 20763 11716 20944 11744
rect 20763 11713 20775 11716
rect 20717 11707 20775 11713
rect 12391 11648 12940 11676
rect 13909 11679 13967 11685
rect 12391 11645 12403 11648
rect 12345 11639 12403 11645
rect 13909 11645 13921 11679
rect 13955 11676 13967 11679
rect 14182 11676 14188 11688
rect 13955 11648 14188 11676
rect 13955 11645 13967 11648
rect 13909 11639 13967 11645
rect 5684 11580 7052 11608
rect 8389 11611 8447 11617
rect 5684 11568 5690 11580
rect 8389 11577 8401 11611
rect 8435 11608 8447 11611
rect 9858 11608 9864 11620
rect 8435 11580 9864 11608
rect 8435 11577 8447 11580
rect 8389 11571 8447 11577
rect 9858 11568 9864 11580
rect 9916 11568 9922 11620
rect 10962 11568 10968 11620
rect 11020 11608 11026 11620
rect 11020 11580 11744 11608
rect 11020 11568 11026 11580
rect 6362 11500 6368 11552
rect 6420 11540 6426 11552
rect 7742 11540 7748 11552
rect 6420 11512 7748 11540
rect 6420 11500 6426 11512
rect 7742 11500 7748 11512
rect 7800 11500 7806 11552
rect 8294 11500 8300 11552
rect 8352 11540 8358 11552
rect 8573 11543 8631 11549
rect 8573 11540 8585 11543
rect 8352 11512 8585 11540
rect 8352 11500 8358 11512
rect 8573 11509 8585 11512
rect 8619 11540 8631 11543
rect 9030 11540 9036 11552
rect 8619 11512 9036 11540
rect 8619 11509 8631 11512
rect 8573 11503 8631 11509
rect 9030 11500 9036 11512
rect 9088 11540 9094 11552
rect 10226 11540 10232 11552
rect 9088 11512 10232 11540
rect 9088 11500 9094 11512
rect 10226 11500 10232 11512
rect 10284 11500 10290 11552
rect 11146 11540 11152 11552
rect 11107 11512 11152 11540
rect 11146 11500 11152 11512
rect 11204 11500 11210 11552
rect 11716 11540 11744 11580
rect 11790 11568 11796 11620
rect 11848 11608 11854 11620
rect 12529 11611 12587 11617
rect 12529 11608 12541 11611
rect 11848 11580 12541 11608
rect 11848 11568 11854 11580
rect 12529 11577 12541 11580
rect 12575 11577 12587 11611
rect 12529 11571 12587 11577
rect 12066 11540 12072 11552
rect 11716 11512 12072 11540
rect 12066 11500 12072 11512
rect 12124 11500 12130 11552
rect 13722 11500 13728 11552
rect 13780 11540 13786 11552
rect 13924 11540 13952 11639
rect 14182 11636 14188 11648
rect 14240 11636 14246 11688
rect 17497 11679 17555 11685
rect 17497 11676 17509 11679
rect 16776 11648 17509 11676
rect 14001 11543 14059 11549
rect 14001 11540 14013 11543
rect 13780 11512 14013 11540
rect 13780 11500 13786 11512
rect 14001 11509 14013 11512
rect 14047 11509 14059 11543
rect 14001 11503 14059 11509
rect 16298 11500 16304 11552
rect 16356 11540 16362 11552
rect 16776 11549 16804 11648
rect 17497 11645 17509 11648
rect 17543 11645 17555 11679
rect 17497 11639 17555 11645
rect 16393 11543 16451 11549
rect 16393 11540 16405 11543
rect 16356 11512 16405 11540
rect 16356 11500 16362 11512
rect 16393 11509 16405 11512
rect 16439 11540 16451 11543
rect 16761 11543 16819 11549
rect 16761 11540 16773 11543
rect 16439 11512 16773 11540
rect 16439 11509 16451 11512
rect 16393 11503 16451 11509
rect 16761 11509 16773 11512
rect 16807 11509 16819 11543
rect 18874 11540 18880 11552
rect 18835 11512 18880 11540
rect 16761 11503 16819 11509
rect 18874 11500 18880 11512
rect 18932 11500 18938 11552
rect 18966 11500 18972 11552
rect 19024 11540 19030 11552
rect 19337 11543 19395 11549
rect 19337 11540 19349 11543
rect 19024 11512 19349 11540
rect 19024 11500 19030 11512
rect 19337 11509 19349 11512
rect 19383 11509 19395 11543
rect 19337 11503 19395 11509
rect 1104 11450 21896 11472
rect 1104 11398 3549 11450
rect 3601 11398 3613 11450
rect 3665 11398 3677 11450
rect 3729 11398 3741 11450
rect 3793 11398 3805 11450
rect 3857 11398 8747 11450
rect 8799 11398 8811 11450
rect 8863 11398 8875 11450
rect 8927 11398 8939 11450
rect 8991 11398 9003 11450
rect 9055 11398 13945 11450
rect 13997 11398 14009 11450
rect 14061 11398 14073 11450
rect 14125 11398 14137 11450
rect 14189 11398 14201 11450
rect 14253 11398 19143 11450
rect 19195 11398 19207 11450
rect 19259 11398 19271 11450
rect 19323 11398 19335 11450
rect 19387 11398 19399 11450
rect 19451 11398 21896 11450
rect 1104 11376 21896 11398
rect 1949 11339 2007 11345
rect 1949 11305 1961 11339
rect 1995 11336 2007 11339
rect 2774 11336 2780 11348
rect 1995 11308 2780 11336
rect 1995 11305 2007 11308
rect 1949 11299 2007 11305
rect 2774 11296 2780 11308
rect 2832 11296 2838 11348
rect 5353 11339 5411 11345
rect 5353 11305 5365 11339
rect 5399 11336 5411 11339
rect 5534 11336 5540 11348
rect 5399 11308 5540 11336
rect 5399 11305 5411 11308
rect 5353 11299 5411 11305
rect 5534 11296 5540 11308
rect 5592 11296 5598 11348
rect 5994 11296 6000 11348
rect 6052 11336 6058 11348
rect 6181 11339 6239 11345
rect 6181 11336 6193 11339
rect 6052 11308 6193 11336
rect 6052 11296 6058 11308
rect 6181 11305 6193 11308
rect 6227 11305 6239 11339
rect 7006 11336 7012 11348
rect 6967 11308 7012 11336
rect 6181 11299 6239 11305
rect 7006 11296 7012 11308
rect 7064 11296 7070 11348
rect 7098 11296 7104 11348
rect 7156 11336 7162 11348
rect 7377 11339 7435 11345
rect 7377 11336 7389 11339
rect 7156 11308 7389 11336
rect 7156 11296 7162 11308
rect 7377 11305 7389 11308
rect 7423 11305 7435 11339
rect 10042 11336 10048 11348
rect 10003 11308 10048 11336
rect 7377 11299 7435 11305
rect 10042 11296 10048 11308
rect 10100 11296 10106 11348
rect 10962 11296 10968 11348
rect 11020 11336 11026 11348
rect 11149 11339 11207 11345
rect 11149 11336 11161 11339
rect 11020 11308 11161 11336
rect 11020 11296 11026 11308
rect 11149 11305 11161 11308
rect 11195 11305 11207 11339
rect 11330 11336 11336 11348
rect 11291 11308 11336 11336
rect 11149 11299 11207 11305
rect 11330 11296 11336 11308
rect 11388 11296 11394 11348
rect 12434 11336 12440 11348
rect 11532 11308 12440 11336
rect 2317 11271 2375 11277
rect 2317 11237 2329 11271
rect 2363 11268 2375 11271
rect 3050 11268 3056 11280
rect 2363 11240 3056 11268
rect 2363 11237 2375 11240
rect 2317 11231 2375 11237
rect 3050 11228 3056 11240
rect 3108 11228 3114 11280
rect 4430 11228 4436 11280
rect 4488 11268 4494 11280
rect 8941 11271 8999 11277
rect 8941 11268 8953 11271
rect 4488 11240 8953 11268
rect 4488 11228 4494 11240
rect 8941 11237 8953 11240
rect 8987 11237 8999 11271
rect 8941 11231 8999 11237
rect 9306 11228 9312 11280
rect 9364 11268 9370 11280
rect 10686 11268 10692 11280
rect 9364 11240 10692 11268
rect 9364 11228 9370 11240
rect 4338 11160 4344 11212
rect 4396 11200 4402 11212
rect 4801 11203 4859 11209
rect 4801 11200 4813 11203
rect 4396 11172 4813 11200
rect 4396 11160 4402 11172
rect 4801 11169 4813 11172
rect 4847 11200 4859 11203
rect 5442 11200 5448 11212
rect 4847 11172 5448 11200
rect 4847 11169 4859 11172
rect 4801 11163 4859 11169
rect 5442 11160 5448 11172
rect 5500 11160 5506 11212
rect 5626 11200 5632 11212
rect 5587 11172 5632 11200
rect 5626 11160 5632 11172
rect 5684 11200 5690 11212
rect 5994 11200 6000 11212
rect 5684 11172 6000 11200
rect 5684 11160 5690 11172
rect 5994 11160 6000 11172
rect 6052 11160 6058 11212
rect 6457 11203 6515 11209
rect 6457 11169 6469 11203
rect 6503 11200 6515 11203
rect 9398 11200 9404 11212
rect 6503 11172 9404 11200
rect 6503 11169 6515 11172
rect 6457 11163 6515 11169
rect 9398 11160 9404 11172
rect 9456 11160 9462 11212
rect 9585 11203 9643 11209
rect 9585 11169 9597 11203
rect 9631 11169 9643 11203
rect 10502 11200 10508 11212
rect 10463 11172 10508 11200
rect 9585 11163 9643 11169
rect 2133 11135 2191 11141
rect 2133 11101 2145 11135
rect 2179 11101 2191 11135
rect 2133 11095 2191 11101
rect 2501 11135 2559 11141
rect 2501 11101 2513 11135
rect 2547 11132 2559 11135
rect 3050 11132 3056 11144
rect 2547 11104 3056 11132
rect 2547 11101 2559 11104
rect 2501 11095 2559 11101
rect 2148 11064 2176 11095
rect 3050 11092 3056 11104
rect 3108 11092 3114 11144
rect 4430 11092 4436 11144
rect 4488 11132 4494 11144
rect 6546 11132 6552 11144
rect 4488 11104 6552 11132
rect 4488 11092 4494 11104
rect 6546 11092 6552 11104
rect 6604 11092 6610 11144
rect 6638 11092 6644 11144
rect 6696 11132 6702 11144
rect 8294 11132 8300 11144
rect 6696 11104 8300 11132
rect 6696 11092 6702 11104
rect 8294 11092 8300 11104
rect 8352 11132 8358 11144
rect 8570 11132 8576 11144
rect 8352 11104 8576 11132
rect 8352 11092 8358 11104
rect 8570 11092 8576 11104
rect 8628 11092 8634 11144
rect 9600 11132 9628 11163
rect 10502 11160 10508 11172
rect 10560 11160 10566 11212
rect 10612 11209 10640 11240
rect 10686 11228 10692 11240
rect 10744 11228 10750 11280
rect 11532 11209 11560 11308
rect 12434 11296 12440 11308
rect 12492 11296 12498 11348
rect 14274 11296 14280 11348
rect 14332 11336 14338 11348
rect 14921 11339 14979 11345
rect 14921 11336 14933 11339
rect 14332 11308 14933 11336
rect 14332 11296 14338 11308
rect 14921 11305 14933 11308
rect 14967 11336 14979 11339
rect 20254 11336 20260 11348
rect 14967 11308 20260 11336
rect 14967 11305 14979 11308
rect 14921 11299 14979 11305
rect 20254 11296 20260 11308
rect 20312 11296 20318 11348
rect 21177 11339 21235 11345
rect 21177 11305 21189 11339
rect 21223 11336 21235 11339
rect 21266 11336 21272 11348
rect 21223 11308 21272 11336
rect 21223 11305 21235 11308
rect 21177 11299 21235 11305
rect 12897 11271 12955 11277
rect 12897 11237 12909 11271
rect 12943 11268 12955 11271
rect 13170 11268 13176 11280
rect 12943 11240 13176 11268
rect 12943 11237 12955 11240
rect 12897 11231 12955 11237
rect 13170 11228 13176 11240
rect 13228 11228 13234 11280
rect 13538 11228 13544 11280
rect 13596 11268 13602 11280
rect 13633 11271 13691 11277
rect 13633 11268 13645 11271
rect 13596 11240 13645 11268
rect 13596 11228 13602 11240
rect 13633 11237 13645 11240
rect 13679 11268 13691 11271
rect 14734 11268 14740 11280
rect 13679 11240 14740 11268
rect 13679 11237 13691 11240
rect 13633 11231 13691 11237
rect 14734 11228 14740 11240
rect 14792 11228 14798 11280
rect 16393 11271 16451 11277
rect 16393 11237 16405 11271
rect 16439 11268 16451 11271
rect 16758 11268 16764 11280
rect 16439 11240 16764 11268
rect 16439 11237 16451 11240
rect 16393 11231 16451 11237
rect 16758 11228 16764 11240
rect 16816 11228 16822 11280
rect 19613 11271 19671 11277
rect 19613 11237 19625 11271
rect 19659 11237 19671 11271
rect 19613 11231 19671 11237
rect 10597 11203 10655 11209
rect 10597 11169 10609 11203
rect 10643 11169 10655 11203
rect 10597 11163 10655 11169
rect 11517 11203 11575 11209
rect 11517 11169 11529 11203
rect 11563 11169 11575 11203
rect 11517 11163 11575 11169
rect 12526 11160 12532 11212
rect 12584 11200 12590 11212
rect 14366 11200 14372 11212
rect 12584 11172 14372 11200
rect 12584 11160 12590 11172
rect 14366 11160 14372 11172
rect 14424 11160 14430 11212
rect 17773 11203 17831 11209
rect 17773 11169 17785 11203
rect 17819 11200 17831 11203
rect 19628 11200 19656 11231
rect 17819 11172 17853 11200
rect 19306 11172 19656 11200
rect 17819 11169 17831 11172
rect 17773 11163 17831 11169
rect 12802 11132 12808 11144
rect 9600 11104 12808 11132
rect 12802 11092 12808 11104
rect 12860 11092 12866 11144
rect 15102 11092 15108 11144
rect 15160 11132 15166 11144
rect 16298 11132 16304 11144
rect 15160 11104 16304 11132
rect 15160 11092 15166 11104
rect 16298 11092 16304 11104
rect 16356 11132 16362 11144
rect 17788 11132 17816 11163
rect 17865 11135 17923 11141
rect 17865 11132 17877 11135
rect 16356 11104 17877 11132
rect 16356 11092 16362 11104
rect 17865 11101 17877 11104
rect 17911 11101 17923 11135
rect 17865 11095 17923 11101
rect 3234 11064 3240 11076
rect 2148 11036 3240 11064
rect 3234 11024 3240 11036
rect 3292 11024 3298 11076
rect 4246 11064 4252 11076
rect 4207 11036 4252 11064
rect 4246 11024 4252 11036
rect 4304 11064 4310 11076
rect 4893 11067 4951 11073
rect 4893 11064 4905 11067
rect 4304 11036 4905 11064
rect 4304 11024 4310 11036
rect 4893 11033 4905 11036
rect 4939 11033 4951 11067
rect 4893 11027 4951 11033
rect 4982 11024 4988 11076
rect 5040 11064 5046 11076
rect 5813 11067 5871 11073
rect 5040 11036 5085 11064
rect 5040 11024 5046 11036
rect 5813 11033 5825 11067
rect 5859 11064 5871 11067
rect 7101 11067 7159 11073
rect 7101 11064 7113 11067
rect 5859 11036 7113 11064
rect 5859 11033 5871 11036
rect 5813 11027 5871 11033
rect 7101 11033 7113 11036
rect 7147 11033 7159 11067
rect 7101 11027 7159 11033
rect 9309 11067 9367 11073
rect 9309 11033 9321 11067
rect 9355 11064 9367 11067
rect 9766 11064 9772 11076
rect 9355 11036 9772 11064
rect 9355 11033 9367 11036
rect 9309 11027 9367 11033
rect 9766 11024 9772 11036
rect 9824 11024 9830 11076
rect 9950 11024 9956 11076
rect 10008 11064 10014 11076
rect 11054 11064 11060 11076
rect 10008 11036 10916 11064
rect 10967 11036 11060 11064
rect 10008 11024 10014 11036
rect 4525 10999 4583 11005
rect 4525 10965 4537 10999
rect 4571 10996 4583 10999
rect 4798 10996 4804 11008
rect 4571 10968 4804 10996
rect 4571 10965 4583 10968
rect 4525 10959 4583 10965
rect 4798 10956 4804 10968
rect 4856 10996 4862 11008
rect 5721 10999 5779 11005
rect 5721 10996 5733 10999
rect 4856 10968 5733 10996
rect 4856 10956 4862 10968
rect 5721 10965 5733 10968
rect 5767 10996 5779 10999
rect 6362 10996 6368 11008
rect 5767 10968 6368 10996
rect 5767 10965 5779 10968
rect 5721 10959 5779 10965
rect 6362 10956 6368 10968
rect 6420 10956 6426 11008
rect 6546 10996 6552 11008
rect 6507 10968 6552 10996
rect 6546 10956 6552 10968
rect 6604 10956 6610 11008
rect 6638 10956 6644 11008
rect 6696 10996 6702 11008
rect 8570 10996 8576 11008
rect 6696 10968 6741 10996
rect 8531 10968 8576 10996
rect 6696 10956 6702 10968
rect 8570 10956 8576 10968
rect 8628 10956 8634 11008
rect 9398 10956 9404 11008
rect 9456 10996 9462 11008
rect 9861 10999 9919 11005
rect 9456 10968 9501 10996
rect 9456 10956 9462 10968
rect 9861 10965 9873 10999
rect 9907 10996 9919 10999
rect 10226 10996 10232 11008
rect 9907 10968 10232 10996
rect 9907 10965 9919 10968
rect 9861 10959 9919 10965
rect 10226 10956 10232 10968
rect 10284 10996 10290 11008
rect 10413 10999 10471 11005
rect 10413 10996 10425 10999
rect 10284 10968 10425 10996
rect 10284 10956 10290 10968
rect 10413 10965 10425 10968
rect 10459 10965 10471 10999
rect 10888 10996 10916 11036
rect 11054 11024 11060 11036
rect 11112 11064 11118 11076
rect 11238 11064 11244 11076
rect 11112 11036 11244 11064
rect 11112 11024 11118 11036
rect 11238 11024 11244 11036
rect 11296 11024 11302 11076
rect 11784 11067 11842 11073
rect 11784 11033 11796 11067
rect 11830 11064 11842 11067
rect 12250 11064 12256 11076
rect 11830 11036 12256 11064
rect 11830 11033 11842 11036
rect 11784 11027 11842 11033
rect 12250 11024 12256 11036
rect 12308 11024 12314 11076
rect 12710 11024 12716 11076
rect 12768 11064 12774 11076
rect 13081 11067 13139 11073
rect 13081 11064 13093 11067
rect 12768 11036 13093 11064
rect 12768 11024 12774 11036
rect 13081 11033 13093 11036
rect 13127 11064 13139 11067
rect 14458 11064 14464 11076
rect 13127 11036 14464 11064
rect 13127 11033 13139 11036
rect 13081 11027 13139 11033
rect 14458 11024 14464 11036
rect 14516 11024 14522 11076
rect 16056 11067 16114 11073
rect 16056 11033 16068 11067
rect 16102 11033 16114 11067
rect 16056 11027 16114 11033
rect 17506 11067 17564 11073
rect 17506 11033 17518 11067
rect 17552 11064 17564 11067
rect 17678 11064 17684 11076
rect 17552 11036 17684 11064
rect 17552 11033 17564 11036
rect 17506 11027 17564 11033
rect 11974 10996 11980 11008
rect 10888 10968 11980 10996
rect 10413 10959 10471 10965
rect 11974 10956 11980 10968
rect 12032 10956 12038 11008
rect 12434 10956 12440 11008
rect 12492 10996 12498 11008
rect 13265 10999 13323 11005
rect 13265 10996 13277 10999
rect 12492 10968 13277 10996
rect 12492 10956 12498 10968
rect 13265 10965 13277 10968
rect 13311 10996 13323 10999
rect 13357 10999 13415 11005
rect 13357 10996 13369 10999
rect 13311 10968 13369 10996
rect 13311 10965 13323 10968
rect 13265 10959 13323 10965
rect 13357 10965 13369 10968
rect 13403 10965 13415 10999
rect 13357 10959 13415 10965
rect 15194 10956 15200 11008
rect 15252 10996 15258 11008
rect 16071 10996 16099 11027
rect 17678 11024 17684 11036
rect 17736 11024 17742 11076
rect 18138 11064 18144 11076
rect 18099 11036 18144 11064
rect 18138 11024 18144 11036
rect 18196 11024 18202 11076
rect 19306 10996 19334 11172
rect 20990 11160 20996 11212
rect 21048 11200 21054 11212
rect 21192 11200 21220 11299
rect 21266 11296 21272 11308
rect 21324 11296 21330 11348
rect 21048 11172 21220 11200
rect 21048 11160 21054 11172
rect 19518 11024 19524 11076
rect 19576 11064 19582 11076
rect 20726 11067 20784 11073
rect 20726 11064 20738 11067
rect 19576 11036 20738 11064
rect 19576 11024 19582 11036
rect 20726 11033 20738 11036
rect 20772 11033 20784 11067
rect 20726 11027 20784 11033
rect 15252 10968 19334 10996
rect 15252 10956 15258 10968
rect 1104 10906 22056 10928
rect 1104 10854 6148 10906
rect 6200 10854 6212 10906
rect 6264 10854 6276 10906
rect 6328 10854 6340 10906
rect 6392 10854 6404 10906
rect 6456 10854 11346 10906
rect 11398 10854 11410 10906
rect 11462 10854 11474 10906
rect 11526 10854 11538 10906
rect 11590 10854 11602 10906
rect 11654 10854 16544 10906
rect 16596 10854 16608 10906
rect 16660 10854 16672 10906
rect 16724 10854 16736 10906
rect 16788 10854 16800 10906
rect 16852 10854 21742 10906
rect 21794 10854 21806 10906
rect 21858 10854 21870 10906
rect 21922 10854 21934 10906
rect 21986 10854 21998 10906
rect 22050 10854 22056 10906
rect 1104 10832 22056 10854
rect 3418 10752 3424 10804
rect 3476 10792 3482 10804
rect 3789 10795 3847 10801
rect 3789 10792 3801 10795
rect 3476 10764 3801 10792
rect 3476 10752 3482 10764
rect 3789 10761 3801 10764
rect 3835 10792 3847 10795
rect 4709 10795 4767 10801
rect 4709 10792 4721 10795
rect 3835 10764 4721 10792
rect 3835 10761 3847 10764
rect 3789 10755 3847 10761
rect 4709 10761 4721 10764
rect 4755 10761 4767 10795
rect 4709 10755 4767 10761
rect 5077 10795 5135 10801
rect 5077 10761 5089 10795
rect 5123 10792 5135 10795
rect 5166 10792 5172 10804
rect 5123 10764 5172 10792
rect 5123 10761 5135 10764
rect 5077 10755 5135 10761
rect 5166 10752 5172 10764
rect 5224 10752 5230 10804
rect 5905 10795 5963 10801
rect 5905 10761 5917 10795
rect 5951 10792 5963 10795
rect 6638 10792 6644 10804
rect 5951 10764 6644 10792
rect 5951 10761 5963 10764
rect 5905 10755 5963 10761
rect 6638 10752 6644 10764
rect 6696 10752 6702 10804
rect 7101 10795 7159 10801
rect 7101 10761 7113 10795
rect 7147 10761 7159 10795
rect 7101 10755 7159 10761
rect 3326 10684 3332 10736
rect 3384 10724 3390 10736
rect 6733 10727 6791 10733
rect 6733 10724 6745 10727
rect 3384 10696 6745 10724
rect 3384 10684 3390 10696
rect 6733 10693 6745 10696
rect 6779 10693 6791 10727
rect 7116 10724 7144 10755
rect 7926 10752 7932 10804
rect 7984 10792 7990 10804
rect 8205 10795 8263 10801
rect 8205 10792 8217 10795
rect 7984 10764 8217 10792
rect 7984 10752 7990 10764
rect 8205 10761 8217 10764
rect 8251 10761 8263 10795
rect 8205 10755 8263 10761
rect 8478 10752 8484 10804
rect 8536 10752 8542 10804
rect 8570 10752 8576 10804
rect 8628 10792 8634 10804
rect 8665 10795 8723 10801
rect 8665 10792 8677 10795
rect 8628 10764 8677 10792
rect 8628 10752 8634 10764
rect 8665 10761 8677 10764
rect 8711 10761 8723 10795
rect 9030 10792 9036 10804
rect 8991 10764 9036 10792
rect 8665 10755 8723 10761
rect 9030 10752 9036 10764
rect 9088 10752 9094 10804
rect 9125 10795 9183 10801
rect 9125 10761 9137 10795
rect 9171 10792 9183 10795
rect 9398 10792 9404 10804
rect 9171 10764 9404 10792
rect 9171 10761 9183 10764
rect 9125 10755 9183 10761
rect 9398 10752 9404 10764
rect 9456 10752 9462 10804
rect 9674 10752 9680 10804
rect 9732 10792 9738 10804
rect 10321 10795 10379 10801
rect 10321 10792 10333 10795
rect 9732 10764 10333 10792
rect 9732 10752 9738 10764
rect 10321 10761 10333 10764
rect 10367 10761 10379 10795
rect 10321 10755 10379 10761
rect 10686 10752 10692 10804
rect 10744 10792 10750 10804
rect 16390 10792 16396 10804
rect 10744 10764 16396 10792
rect 10744 10752 10750 10764
rect 16390 10752 16396 10764
rect 16448 10792 16454 10804
rect 16485 10795 16543 10801
rect 16485 10792 16497 10795
rect 16448 10764 16497 10792
rect 16448 10752 16454 10764
rect 16485 10761 16497 10764
rect 16531 10761 16543 10795
rect 16942 10792 16948 10804
rect 16485 10755 16543 10761
rect 16684 10764 16948 10792
rect 8496 10724 8524 10752
rect 7116 10696 8524 10724
rect 9585 10727 9643 10733
rect 6733 10687 6791 10693
rect 9585 10693 9597 10727
rect 9631 10724 9643 10727
rect 10134 10724 10140 10736
rect 9631 10696 10140 10724
rect 9631 10693 9643 10696
rect 9585 10687 9643 10693
rect 10134 10684 10140 10696
rect 10192 10684 10198 10736
rect 10502 10684 10508 10736
rect 10560 10724 10566 10736
rect 10560 10696 11284 10724
rect 10560 10684 10566 10696
rect 5534 10656 5540 10668
rect 5495 10628 5540 10656
rect 5534 10616 5540 10628
rect 5592 10616 5598 10668
rect 5718 10616 5724 10668
rect 5776 10656 5782 10668
rect 5997 10659 6055 10665
rect 5997 10656 6009 10659
rect 5776 10628 6009 10656
rect 5776 10616 5782 10628
rect 5997 10625 6009 10628
rect 6043 10625 6055 10659
rect 6914 10656 6920 10668
rect 5997 10619 6055 10625
rect 6564 10628 6920 10656
rect 2774 10548 2780 10600
rect 2832 10588 2838 10600
rect 2961 10591 3019 10597
rect 2961 10588 2973 10591
rect 2832 10560 2973 10588
rect 2832 10548 2838 10560
rect 2961 10557 2973 10560
rect 3007 10557 3019 10591
rect 2961 10551 3019 10557
rect 4249 10591 4307 10597
rect 4249 10557 4261 10591
rect 4295 10588 4307 10591
rect 4430 10588 4436 10600
rect 4295 10560 4436 10588
rect 4295 10557 4307 10560
rect 4249 10551 4307 10557
rect 4430 10548 4436 10560
rect 4488 10548 4494 10600
rect 4617 10591 4675 10597
rect 4617 10557 4629 10591
rect 4663 10557 4675 10591
rect 4617 10551 4675 10557
rect 5353 10591 5411 10597
rect 5353 10557 5365 10591
rect 5399 10557 5411 10591
rect 5353 10551 5411 10557
rect 4632 10520 4660 10551
rect 3988 10492 4660 10520
rect 5368 10520 5396 10551
rect 5442 10548 5448 10600
rect 5500 10588 5506 10600
rect 5500 10560 5545 10588
rect 5500 10548 5506 10560
rect 5736 10520 5764 10616
rect 6564 10597 6592 10628
rect 6914 10616 6920 10628
rect 6972 10616 6978 10668
rect 7190 10616 7196 10668
rect 7248 10656 7254 10668
rect 7837 10659 7895 10665
rect 7837 10656 7849 10659
rect 7248 10628 7849 10656
rect 7248 10616 7254 10628
rect 7837 10625 7849 10628
rect 7883 10625 7895 10659
rect 9306 10656 9312 10668
rect 7837 10619 7895 10625
rect 8496 10628 9312 10656
rect 6549 10591 6607 10597
rect 6549 10557 6561 10591
rect 6595 10557 6607 10591
rect 6549 10551 6607 10557
rect 6641 10591 6699 10597
rect 6641 10557 6653 10591
rect 6687 10557 6699 10591
rect 6641 10551 6699 10557
rect 5368 10492 5764 10520
rect 3988 10464 4016 10492
rect 5902 10480 5908 10532
rect 5960 10520 5966 10532
rect 6656 10520 6684 10551
rect 6822 10548 6828 10600
rect 6880 10588 6886 10600
rect 7561 10591 7619 10597
rect 7561 10588 7573 10591
rect 6880 10560 7573 10588
rect 6880 10548 6886 10560
rect 7561 10557 7573 10560
rect 7607 10557 7619 10591
rect 7561 10551 7619 10557
rect 7745 10591 7803 10597
rect 7745 10557 7757 10591
rect 7791 10588 7803 10591
rect 8386 10588 8392 10600
rect 7791 10560 8392 10588
rect 7791 10557 7803 10560
rect 7745 10551 7803 10557
rect 5960 10492 6684 10520
rect 7576 10520 7604 10551
rect 8386 10548 8392 10560
rect 8444 10548 8450 10600
rect 8496 10597 8524 10628
rect 9306 10616 9312 10628
rect 9364 10616 9370 10668
rect 9493 10659 9551 10665
rect 9493 10625 9505 10659
rect 9539 10656 9551 10659
rect 10042 10656 10048 10668
rect 9539 10628 10048 10656
rect 9539 10625 9551 10628
rect 9493 10619 9551 10625
rect 10042 10616 10048 10628
rect 10100 10616 10106 10668
rect 10229 10659 10287 10665
rect 10229 10625 10241 10659
rect 10275 10656 10287 10659
rect 10689 10659 10747 10665
rect 10689 10656 10701 10659
rect 10275 10628 10701 10656
rect 10275 10625 10287 10628
rect 10229 10619 10287 10625
rect 10689 10625 10701 10628
rect 10735 10625 10747 10659
rect 10689 10619 10747 10625
rect 8481 10591 8539 10597
rect 8481 10557 8493 10591
rect 8527 10557 8539 10591
rect 8481 10551 8539 10557
rect 8570 10548 8576 10600
rect 8628 10588 8634 10600
rect 9582 10588 9588 10600
rect 8628 10560 8673 10588
rect 9048 10560 9588 10588
rect 8628 10548 8634 10560
rect 9048 10520 9076 10560
rect 9582 10548 9588 10560
rect 9640 10548 9646 10600
rect 9769 10591 9827 10597
rect 9769 10557 9781 10591
rect 9815 10557 9827 10591
rect 10778 10588 10784 10600
rect 10739 10560 10784 10588
rect 9769 10551 9827 10557
rect 7576 10492 9076 10520
rect 5960 10480 5966 10492
rect 9122 10480 9128 10532
rect 9180 10520 9186 10532
rect 9784 10520 9812 10551
rect 10778 10548 10784 10560
rect 10836 10548 10842 10600
rect 10870 10548 10876 10600
rect 10928 10588 10934 10600
rect 11256 10597 11284 10696
rect 12434 10684 12440 10736
rect 12492 10684 12498 10736
rect 12652 10727 12710 10733
rect 12652 10693 12664 10727
rect 12698 10724 12710 10727
rect 12802 10724 12808 10736
rect 12698 10696 12808 10724
rect 12698 10693 12710 10696
rect 12652 10687 12710 10693
rect 12802 10684 12808 10696
rect 12860 10684 12866 10736
rect 13722 10724 13728 10736
rect 13004 10696 13728 10724
rect 12452 10656 12480 10684
rect 13004 10665 13032 10696
rect 13722 10684 13728 10696
rect 13780 10724 13786 10736
rect 14458 10724 14464 10736
rect 13780 10696 14464 10724
rect 13780 10684 13786 10696
rect 14458 10684 14464 10696
rect 14516 10724 14522 10736
rect 14645 10727 14703 10733
rect 14645 10724 14657 10727
rect 14516 10696 14657 10724
rect 14516 10684 14522 10696
rect 14645 10693 14657 10696
rect 14691 10724 14703 10727
rect 15372 10727 15430 10733
rect 14691 10696 15148 10724
rect 14691 10693 14703 10696
rect 14645 10687 14703 10693
rect 15120 10668 15148 10696
rect 15372 10693 15384 10727
rect 15418 10724 15430 10727
rect 15562 10724 15568 10736
rect 15418 10696 15568 10724
rect 15418 10693 15430 10696
rect 15372 10687 15430 10693
rect 15562 10684 15568 10696
rect 15620 10684 15626 10736
rect 12897 10659 12955 10665
rect 12897 10656 12909 10659
rect 12452 10628 12909 10656
rect 12897 10625 12909 10628
rect 12943 10656 12955 10659
rect 12989 10659 13047 10665
rect 12989 10656 13001 10659
rect 12943 10628 13001 10656
rect 12943 10625 12955 10628
rect 12897 10619 12955 10625
rect 12989 10625 13001 10628
rect 13035 10625 13047 10659
rect 12989 10619 13047 10625
rect 13256 10659 13314 10665
rect 13256 10625 13268 10659
rect 13302 10656 13314 10659
rect 13630 10656 13636 10668
rect 13302 10628 13636 10656
rect 13302 10625 13314 10628
rect 13256 10619 13314 10625
rect 13630 10616 13636 10628
rect 13688 10616 13694 10668
rect 15102 10656 15108 10668
rect 15015 10628 15108 10656
rect 15102 10616 15108 10628
rect 15160 10616 15166 10668
rect 16298 10616 16304 10668
rect 16356 10656 16362 10668
rect 16684 10665 16712 10764
rect 16942 10752 16948 10764
rect 17000 10752 17006 10804
rect 20990 10792 20996 10804
rect 20951 10764 20996 10792
rect 20990 10752 20996 10764
rect 21048 10752 21054 10804
rect 16669 10659 16727 10665
rect 16669 10656 16681 10659
rect 16356 10628 16681 10656
rect 16356 10616 16362 10628
rect 16669 10625 16681 10628
rect 16715 10625 16727 10659
rect 16925 10659 16983 10665
rect 16925 10656 16937 10659
rect 16669 10619 16727 10625
rect 16776 10628 16937 10656
rect 11241 10591 11299 10597
rect 10928 10560 10973 10588
rect 10928 10548 10934 10560
rect 11241 10557 11253 10591
rect 11287 10588 11299 10591
rect 11698 10588 11704 10600
rect 11287 10560 11704 10588
rect 11287 10557 11299 10560
rect 11241 10551 11299 10557
rect 11698 10548 11704 10560
rect 11756 10548 11762 10600
rect 16776 10588 16804 10628
rect 16925 10625 16937 10628
rect 16971 10625 16983 10659
rect 16925 10619 16983 10625
rect 20070 10616 20076 10668
rect 20128 10656 20134 10668
rect 20542 10659 20600 10665
rect 20542 10656 20554 10659
rect 20128 10628 20554 10656
rect 20128 10616 20134 10628
rect 20542 10625 20554 10628
rect 20588 10625 20600 10659
rect 20542 10619 20600 10625
rect 20809 10659 20867 10665
rect 20809 10625 20821 10659
rect 20855 10656 20867 10659
rect 21008 10656 21036 10752
rect 20855 10628 21036 10656
rect 20855 10625 20867 10628
rect 20809 10619 20867 10625
rect 16132 10560 16804 10588
rect 9180 10492 11744 10520
rect 9180 10480 9186 10492
rect 3970 10452 3976 10464
rect 3931 10424 3976 10452
rect 3970 10412 3976 10424
rect 4028 10412 4034 10464
rect 7190 10412 7196 10464
rect 7248 10452 7254 10464
rect 7285 10455 7343 10461
rect 7285 10452 7297 10455
rect 7248 10424 7297 10452
rect 7248 10412 7254 10424
rect 7285 10421 7297 10424
rect 7331 10421 7343 10455
rect 7285 10415 7343 10421
rect 9306 10412 9312 10464
rect 9364 10452 9370 10464
rect 9858 10452 9864 10464
rect 9364 10424 9864 10452
rect 9364 10412 9370 10424
rect 9858 10412 9864 10424
rect 9916 10412 9922 10464
rect 11517 10455 11575 10461
rect 11517 10421 11529 10455
rect 11563 10452 11575 10455
rect 11606 10452 11612 10464
rect 11563 10424 11612 10452
rect 11563 10421 11575 10424
rect 11517 10415 11575 10421
rect 11606 10412 11612 10424
rect 11664 10412 11670 10464
rect 11716 10452 11744 10492
rect 13924 10492 14780 10520
rect 12986 10452 12992 10464
rect 11716 10424 12992 10452
rect 12986 10412 12992 10424
rect 13044 10412 13050 10464
rect 13722 10412 13728 10464
rect 13780 10452 13786 10464
rect 13924 10452 13952 10492
rect 13780 10424 13952 10452
rect 14369 10455 14427 10461
rect 13780 10412 13786 10424
rect 14369 10421 14381 10455
rect 14415 10452 14427 10455
rect 14642 10452 14648 10464
rect 14415 10424 14648 10452
rect 14415 10421 14427 10424
rect 14369 10415 14427 10421
rect 14642 10412 14648 10424
rect 14700 10412 14706 10464
rect 14752 10452 14780 10492
rect 16132 10452 16160 10560
rect 17954 10548 17960 10600
rect 18012 10588 18018 10600
rect 18141 10591 18199 10597
rect 18141 10588 18153 10591
rect 18012 10560 18153 10588
rect 18012 10548 18018 10560
rect 18141 10557 18153 10560
rect 18187 10588 18199 10591
rect 18325 10591 18383 10597
rect 18325 10588 18337 10591
rect 18187 10560 18337 10588
rect 18187 10557 18199 10560
rect 18141 10551 18199 10557
rect 18325 10557 18337 10560
rect 18371 10557 18383 10591
rect 18325 10551 18383 10557
rect 19702 10520 19708 10532
rect 18064 10492 19708 10520
rect 18064 10461 18092 10492
rect 19702 10480 19708 10492
rect 19760 10480 19766 10532
rect 14752 10424 16160 10452
rect 18049 10455 18107 10461
rect 18049 10421 18061 10455
rect 18095 10421 18107 10455
rect 18049 10415 18107 10421
rect 19429 10455 19487 10461
rect 19429 10421 19441 10455
rect 19475 10452 19487 10455
rect 19518 10452 19524 10464
rect 19475 10424 19524 10452
rect 19475 10421 19487 10424
rect 19429 10415 19487 10421
rect 19518 10412 19524 10424
rect 19576 10412 19582 10464
rect 1104 10362 21896 10384
rect 1104 10310 3549 10362
rect 3601 10310 3613 10362
rect 3665 10310 3677 10362
rect 3729 10310 3741 10362
rect 3793 10310 3805 10362
rect 3857 10310 8747 10362
rect 8799 10310 8811 10362
rect 8863 10310 8875 10362
rect 8927 10310 8939 10362
rect 8991 10310 9003 10362
rect 9055 10310 13945 10362
rect 13997 10310 14009 10362
rect 14061 10310 14073 10362
rect 14125 10310 14137 10362
rect 14189 10310 14201 10362
rect 14253 10310 19143 10362
rect 19195 10310 19207 10362
rect 19259 10310 19271 10362
rect 19323 10310 19335 10362
rect 19387 10310 19399 10362
rect 19451 10310 21896 10362
rect 1104 10288 21896 10310
rect 1762 10208 1768 10260
rect 1820 10248 1826 10260
rect 1857 10251 1915 10257
rect 1857 10248 1869 10251
rect 1820 10220 1869 10248
rect 1820 10208 1826 10220
rect 1857 10217 1869 10220
rect 1903 10217 1915 10251
rect 1857 10211 1915 10217
rect 2133 10251 2191 10257
rect 2133 10217 2145 10251
rect 2179 10248 2191 10251
rect 2958 10248 2964 10260
rect 2179 10220 2964 10248
rect 2179 10217 2191 10220
rect 2133 10211 2191 10217
rect 2958 10208 2964 10220
rect 3016 10208 3022 10260
rect 3145 10251 3203 10257
rect 3145 10217 3157 10251
rect 3191 10248 3203 10251
rect 3326 10248 3332 10260
rect 3191 10220 3332 10248
rect 3191 10217 3203 10220
rect 3145 10211 3203 10217
rect 3326 10208 3332 10220
rect 3384 10208 3390 10260
rect 4062 10208 4068 10260
rect 4120 10248 4126 10260
rect 4430 10248 4436 10260
rect 4120 10220 4436 10248
rect 4120 10208 4126 10220
rect 4430 10208 4436 10220
rect 4488 10248 4494 10260
rect 4617 10251 4675 10257
rect 4617 10248 4629 10251
rect 4488 10220 4629 10248
rect 4488 10208 4494 10220
rect 4617 10217 4629 10220
rect 4663 10248 4675 10251
rect 5442 10248 5448 10260
rect 4663 10220 5448 10248
rect 4663 10217 4675 10220
rect 4617 10211 4675 10217
rect 5442 10208 5448 10220
rect 5500 10208 5506 10260
rect 5629 10251 5687 10257
rect 5629 10217 5641 10251
rect 5675 10248 5687 10251
rect 5810 10248 5816 10260
rect 5675 10220 5816 10248
rect 5675 10217 5687 10220
rect 5629 10211 5687 10217
rect 5810 10208 5816 10220
rect 5868 10208 5874 10260
rect 6546 10208 6552 10260
rect 6604 10248 6610 10260
rect 7098 10248 7104 10260
rect 6604 10220 7104 10248
rect 6604 10208 6610 10220
rect 7098 10208 7104 10220
rect 7156 10208 7162 10260
rect 7285 10251 7343 10257
rect 7285 10217 7297 10251
rect 7331 10248 7343 10251
rect 7558 10248 7564 10260
rect 7331 10220 7564 10248
rect 7331 10217 7343 10220
rect 7285 10211 7343 10217
rect 7558 10208 7564 10220
rect 7616 10208 7622 10260
rect 8018 10208 8024 10260
rect 8076 10248 8082 10260
rect 8941 10251 8999 10257
rect 8941 10248 8953 10251
rect 8076 10220 8953 10248
rect 8076 10208 8082 10220
rect 8941 10217 8953 10220
rect 8987 10217 8999 10251
rect 10134 10248 10140 10260
rect 10095 10220 10140 10248
rect 8941 10211 8999 10217
rect 10134 10208 10140 10220
rect 10192 10208 10198 10260
rect 11606 10208 11612 10260
rect 11664 10248 11670 10260
rect 12526 10248 12532 10260
rect 11664 10220 12532 10248
rect 11664 10208 11670 10220
rect 12526 10208 12532 10220
rect 12584 10248 12590 10260
rect 13722 10248 13728 10260
rect 12584 10220 13728 10248
rect 12584 10208 12590 10220
rect 13722 10208 13728 10220
rect 13780 10208 13786 10260
rect 14458 10248 14464 10260
rect 14209 10220 14464 10248
rect 4525 10183 4583 10189
rect 4525 10149 4537 10183
rect 4571 10180 4583 10183
rect 7193 10183 7251 10189
rect 4571 10152 6408 10180
rect 4571 10149 4583 10152
rect 4525 10143 4583 10149
rect 2593 10115 2651 10121
rect 2593 10081 2605 10115
rect 2639 10112 2651 10115
rect 3786 10112 3792 10124
rect 2639 10084 3792 10112
rect 2639 10081 2651 10084
rect 2593 10075 2651 10081
rect 3786 10072 3792 10084
rect 3844 10072 3850 10124
rect 3973 10115 4031 10121
rect 3973 10081 3985 10115
rect 4019 10112 4031 10115
rect 4019 10084 4568 10112
rect 4019 10081 4031 10084
rect 3973 10075 4031 10081
rect 2317 10047 2375 10053
rect 2317 10013 2329 10047
rect 2363 10013 2375 10047
rect 2317 10007 2375 10013
rect 2332 9976 2360 10007
rect 2774 10004 2780 10056
rect 2832 10044 2838 10056
rect 2832 10016 2877 10044
rect 2832 10004 2838 10016
rect 3694 10004 3700 10056
rect 3752 10044 3758 10056
rect 3988 10044 4016 10075
rect 3752 10016 4016 10044
rect 4540 10044 4568 10084
rect 4614 10072 4620 10124
rect 4672 10112 4678 10124
rect 4985 10115 5043 10121
rect 4985 10112 4997 10115
rect 4672 10084 4997 10112
rect 4672 10072 4678 10084
rect 4985 10081 4997 10084
rect 5031 10081 5043 10115
rect 5534 10112 5540 10124
rect 5495 10084 5540 10112
rect 4985 10075 5043 10081
rect 5534 10072 5540 10084
rect 5592 10072 5598 10124
rect 5994 10072 6000 10124
rect 6052 10112 6058 10124
rect 6181 10115 6239 10121
rect 6181 10112 6193 10115
rect 6052 10084 6193 10112
rect 6052 10072 6058 10084
rect 6181 10081 6193 10084
rect 6227 10081 6239 10115
rect 6181 10075 6239 10081
rect 5074 10044 5080 10056
rect 4540 10016 5080 10044
rect 3752 10004 3758 10016
rect 5074 10004 5080 10016
rect 5132 10004 5138 10056
rect 5258 10044 5264 10056
rect 5219 10016 5264 10044
rect 5258 10004 5264 10016
rect 5316 10004 5322 10056
rect 6380 10044 6408 10152
rect 7193 10149 7205 10183
rect 7239 10180 7251 10183
rect 9306 10180 9312 10192
rect 7239 10152 9312 10180
rect 7239 10149 7251 10152
rect 7193 10143 7251 10149
rect 9306 10140 9312 10152
rect 9364 10140 9370 10192
rect 12158 10140 12164 10192
rect 12216 10180 12222 10192
rect 12342 10180 12348 10192
rect 12216 10152 12348 10180
rect 12216 10140 12222 10152
rect 12342 10140 12348 10152
rect 12400 10140 12406 10192
rect 13446 10140 13452 10192
rect 13504 10180 13510 10192
rect 13541 10183 13599 10189
rect 13541 10180 13553 10183
rect 13504 10152 13553 10180
rect 13504 10140 13510 10152
rect 13541 10149 13553 10152
rect 13587 10180 13599 10183
rect 13587 10152 13768 10180
rect 13587 10149 13599 10152
rect 13541 10143 13599 10149
rect 13740 10124 13768 10152
rect 6638 10112 6644 10124
rect 6599 10084 6644 10112
rect 6638 10072 6644 10084
rect 6696 10072 6702 10124
rect 6730 10072 6736 10124
rect 6788 10112 6794 10124
rect 7837 10115 7895 10121
rect 7837 10112 7849 10115
rect 6788 10084 7849 10112
rect 6788 10072 6794 10084
rect 7837 10081 7849 10084
rect 7883 10081 7895 10115
rect 8110 10112 8116 10124
rect 8071 10084 8116 10112
rect 7837 10075 7895 10081
rect 8110 10072 8116 10084
rect 8168 10112 8174 10124
rect 8570 10112 8576 10124
rect 8168 10084 8576 10112
rect 8168 10072 8174 10084
rect 8570 10072 8576 10084
rect 8628 10072 8634 10124
rect 9398 10112 9404 10124
rect 9359 10084 9404 10112
rect 9398 10072 9404 10084
rect 9456 10072 9462 10124
rect 9582 10112 9588 10124
rect 9543 10084 9588 10112
rect 9582 10072 9588 10084
rect 9640 10072 9646 10124
rect 13722 10072 13728 10124
rect 13780 10072 13786 10124
rect 6825 10047 6883 10053
rect 6825 10044 6837 10047
rect 6380 10016 6837 10044
rect 6825 10013 6837 10016
rect 6871 10013 6883 10047
rect 8386 10044 8392 10056
rect 8299 10016 8392 10044
rect 6825 10007 6883 10013
rect 8386 10004 8392 10016
rect 8444 10044 8450 10056
rect 10042 10044 10048 10056
rect 8444 10016 10048 10044
rect 8444 10004 8450 10016
rect 10042 10004 10048 10016
rect 10100 10004 10106 10056
rect 11977 10047 12035 10053
rect 11977 10013 11989 10047
rect 12023 10044 12035 10047
rect 12066 10044 12072 10056
rect 12023 10016 12072 10044
rect 12023 10013 12035 10016
rect 11977 10007 12035 10013
rect 12066 10004 12072 10016
rect 12124 10044 12130 10056
rect 12434 10044 12440 10056
rect 12124 10016 12440 10044
rect 12124 10004 12130 10016
rect 12434 10004 12440 10016
rect 12492 10004 12498 10056
rect 14209 10053 14237 10220
rect 14458 10208 14464 10220
rect 14516 10208 14522 10260
rect 14918 10208 14924 10260
rect 14976 10248 14982 10260
rect 19521 10251 19579 10257
rect 19521 10248 19533 10251
rect 14976 10220 19533 10248
rect 14976 10208 14982 10220
rect 19521 10217 19533 10220
rect 19567 10217 19579 10251
rect 20990 10248 20996 10260
rect 20951 10220 20996 10248
rect 19521 10211 19579 10217
rect 20990 10208 20996 10220
rect 21048 10208 21054 10260
rect 18785 10115 18843 10121
rect 18785 10112 18797 10115
rect 18156 10084 18797 10112
rect 14458 10053 14464 10056
rect 13449 10047 13507 10053
rect 13449 10013 13461 10047
rect 13495 10044 13507 10047
rect 14185 10047 14243 10053
rect 14185 10044 14197 10047
rect 13495 10016 14197 10044
rect 13495 10013 13507 10016
rect 13449 10007 13507 10013
rect 14185 10013 14197 10016
rect 14231 10013 14243 10047
rect 14185 10007 14243 10013
rect 14452 10007 14464 10053
rect 14516 10044 14522 10056
rect 14516 10016 14552 10044
rect 14458 10004 14464 10007
rect 14516 10004 14522 10016
rect 15286 10004 15292 10056
rect 15344 10044 15350 10056
rect 15344 10016 16896 10044
rect 15344 10004 15350 10016
rect 3418 9976 3424 9988
rect 2332 9948 3424 9976
rect 3418 9936 3424 9948
rect 3476 9936 3482 9988
rect 3605 9979 3663 9985
rect 3605 9945 3617 9979
rect 3651 9976 3663 9979
rect 4157 9979 4215 9985
rect 4157 9976 4169 9979
rect 3651 9948 4169 9976
rect 3651 9945 3663 9948
rect 3605 9939 3663 9945
rect 4157 9945 4169 9948
rect 4203 9945 4215 9979
rect 4157 9939 4215 9945
rect 4982 9936 4988 9988
rect 5040 9976 5046 9988
rect 5997 9979 6055 9985
rect 5997 9976 6009 9979
rect 5040 9948 6009 9976
rect 5040 9936 5046 9948
rect 5997 9945 6009 9948
rect 6043 9976 6055 9979
rect 6043 9948 6224 9976
rect 6043 9945 6055 9948
rect 5997 9939 6055 9945
rect 1762 9868 1768 9920
rect 1820 9908 1826 9920
rect 2685 9911 2743 9917
rect 2685 9908 2697 9911
rect 1820 9880 2697 9908
rect 1820 9868 1826 9880
rect 2685 9877 2697 9880
rect 2731 9877 2743 9911
rect 2685 9871 2743 9877
rect 2958 9868 2964 9920
rect 3016 9908 3022 9920
rect 3237 9911 3295 9917
rect 3237 9908 3249 9911
rect 3016 9880 3249 9908
rect 3016 9868 3022 9880
rect 3237 9877 3249 9880
rect 3283 9908 3295 9911
rect 4065 9911 4123 9917
rect 4065 9908 4077 9911
rect 3283 9880 4077 9908
rect 3283 9877 3295 9880
rect 3237 9871 3295 9877
rect 4065 9877 4077 9880
rect 4111 9877 4123 9911
rect 4065 9871 4123 9877
rect 5534 9868 5540 9920
rect 5592 9908 5598 9920
rect 6086 9908 6092 9920
rect 5592 9880 6092 9908
rect 5592 9868 5598 9880
rect 6086 9868 6092 9880
rect 6144 9868 6150 9920
rect 6196 9908 6224 9948
rect 6270 9936 6276 9988
rect 6328 9976 6334 9988
rect 6733 9979 6791 9985
rect 6733 9976 6745 9979
rect 6328 9948 6745 9976
rect 6328 9936 6334 9948
rect 6733 9945 6745 9948
rect 6779 9945 6791 9979
rect 8018 9976 8024 9988
rect 6733 9939 6791 9945
rect 6932 9948 8024 9976
rect 6932 9908 6960 9948
rect 8018 9936 8024 9948
rect 8076 9936 8082 9988
rect 8757 9979 8815 9985
rect 8757 9945 8769 9979
rect 8803 9976 8815 9979
rect 9309 9979 9367 9985
rect 9309 9976 9321 9979
rect 8803 9948 9321 9976
rect 8803 9945 8815 9948
rect 8757 9939 8815 9945
rect 9309 9945 9321 9948
rect 9355 9945 9367 9979
rect 10321 9979 10379 9985
rect 10321 9976 10333 9979
rect 9309 9939 9367 9945
rect 9508 9948 10333 9976
rect 6196 9880 6960 9908
rect 7006 9868 7012 9920
rect 7064 9908 7070 9920
rect 7653 9911 7711 9917
rect 7653 9908 7665 9911
rect 7064 9880 7665 9908
rect 7064 9868 7070 9880
rect 7653 9877 7665 9880
rect 7699 9877 7711 9911
rect 7653 9871 7711 9877
rect 7742 9868 7748 9920
rect 7800 9908 7806 9920
rect 7800 9880 7845 9908
rect 7800 9868 7806 9880
rect 8202 9868 8208 9920
rect 8260 9908 8266 9920
rect 9508 9908 9536 9948
rect 10321 9945 10333 9948
rect 10367 9976 10379 9979
rect 10778 9976 10784 9988
rect 10367 9948 10784 9976
rect 10367 9945 10379 9948
rect 10321 9939 10379 9945
rect 10778 9936 10784 9948
rect 10836 9936 10842 9988
rect 11732 9979 11790 9985
rect 11732 9945 11744 9979
rect 11778 9976 11790 9979
rect 13204 9979 13262 9985
rect 11778 9948 13124 9976
rect 11778 9945 11790 9948
rect 11732 9939 11790 9945
rect 9766 9908 9772 9920
rect 8260 9880 9536 9908
rect 9727 9880 9772 9908
rect 8260 9868 8266 9880
rect 9766 9868 9772 9880
rect 9824 9868 9830 9920
rect 10594 9908 10600 9920
rect 10555 9880 10600 9908
rect 10594 9868 10600 9880
rect 10652 9868 10658 9920
rect 12069 9911 12127 9917
rect 12069 9877 12081 9911
rect 12115 9908 12127 9911
rect 12710 9908 12716 9920
rect 12115 9880 12716 9908
rect 12115 9877 12127 9880
rect 12069 9871 12127 9877
rect 12710 9868 12716 9880
rect 12768 9868 12774 9920
rect 13096 9908 13124 9948
rect 13204 9945 13216 9979
rect 13250 9976 13262 9979
rect 13354 9976 13360 9988
rect 13250 9948 13360 9976
rect 13250 9945 13262 9948
rect 13204 9939 13262 9945
rect 13354 9936 13360 9948
rect 13412 9936 13418 9988
rect 16298 9936 16304 9988
rect 16356 9976 16362 9988
rect 16770 9979 16828 9985
rect 16770 9976 16782 9979
rect 16356 9948 16782 9976
rect 16356 9936 16362 9948
rect 16770 9945 16782 9948
rect 16816 9945 16828 9979
rect 16868 9976 16896 10016
rect 16942 10004 16948 10056
rect 17000 10044 17006 10056
rect 17037 10047 17095 10053
rect 17037 10044 17049 10047
rect 17000 10016 17049 10044
rect 17000 10004 17006 10016
rect 17037 10013 17049 10016
rect 17083 10044 17095 10047
rect 17129 10047 17187 10053
rect 17129 10044 17141 10047
rect 17083 10016 17141 10044
rect 17083 10013 17095 10016
rect 17037 10007 17095 10013
rect 17129 10013 17141 10016
rect 17175 10044 17187 10047
rect 17954 10044 17960 10056
rect 17175 10016 17960 10044
rect 17175 10013 17187 10016
rect 17129 10007 17187 10013
rect 17954 10004 17960 10016
rect 18012 10004 18018 10056
rect 18156 10044 18184 10084
rect 18785 10081 18797 10084
rect 18831 10112 18843 10115
rect 19610 10112 19616 10124
rect 18831 10084 19616 10112
rect 18831 10081 18843 10084
rect 18785 10075 18843 10081
rect 19610 10072 19616 10084
rect 19668 10072 19674 10124
rect 20901 10115 20959 10121
rect 20901 10081 20913 10115
rect 20947 10112 20959 10115
rect 21008 10112 21036 10208
rect 20947 10084 21036 10112
rect 20947 10081 20959 10084
rect 20901 10075 20959 10081
rect 19886 10044 19892 10056
rect 18064 10016 18184 10044
rect 18524 10016 19892 10044
rect 17374 9979 17432 9985
rect 17374 9976 17386 9979
rect 16868 9948 17386 9976
rect 16770 9939 16828 9945
rect 17374 9945 17386 9948
rect 17420 9945 17432 9979
rect 18064 9976 18092 10016
rect 17374 9939 17432 9945
rect 17512 9948 18092 9976
rect 13817 9911 13875 9917
rect 13817 9908 13829 9911
rect 13096 9880 13829 9908
rect 13817 9877 13829 9880
rect 13863 9908 13875 9911
rect 13906 9908 13912 9920
rect 13863 9880 13912 9908
rect 13863 9877 13875 9880
rect 13817 9871 13875 9877
rect 13906 9868 13912 9880
rect 13964 9868 13970 9920
rect 15562 9908 15568 9920
rect 15523 9880 15568 9908
rect 15562 9868 15568 9880
rect 15620 9868 15626 9920
rect 15654 9868 15660 9920
rect 15712 9908 15718 9920
rect 16776 9908 16804 9939
rect 17512 9908 17540 9948
rect 18524 9920 18552 10016
rect 19886 10004 19892 10016
rect 19944 10004 19950 10056
rect 19334 9936 19340 9988
rect 19392 9976 19398 9988
rect 20530 9976 20536 9988
rect 19392 9948 20536 9976
rect 19392 9936 19398 9948
rect 20530 9936 20536 9948
rect 20588 9976 20594 9988
rect 20634 9979 20692 9985
rect 20634 9976 20646 9979
rect 20588 9948 20646 9976
rect 20588 9936 20594 9948
rect 20634 9945 20646 9948
rect 20680 9945 20692 9979
rect 20634 9939 20692 9945
rect 18506 9908 18512 9920
rect 15712 9880 15757 9908
rect 16776 9880 17540 9908
rect 18467 9880 18512 9908
rect 15712 9868 15718 9880
rect 18506 9868 18512 9880
rect 18564 9868 18570 9920
rect 18693 9911 18751 9917
rect 18693 9877 18705 9911
rect 18739 9908 18751 9911
rect 18969 9911 19027 9917
rect 18969 9908 18981 9911
rect 18739 9880 18981 9908
rect 18739 9877 18751 9880
rect 18693 9871 18751 9877
rect 18969 9877 18981 9880
rect 19015 9908 19027 9911
rect 19150 9908 19156 9920
rect 19015 9880 19156 9908
rect 19015 9877 19027 9880
rect 18969 9871 19027 9877
rect 19150 9868 19156 9880
rect 19208 9868 19214 9920
rect 1104 9818 22056 9840
rect 1104 9766 6148 9818
rect 6200 9766 6212 9818
rect 6264 9766 6276 9818
rect 6328 9766 6340 9818
rect 6392 9766 6404 9818
rect 6456 9766 11346 9818
rect 11398 9766 11410 9818
rect 11462 9766 11474 9818
rect 11526 9766 11538 9818
rect 11590 9766 11602 9818
rect 11654 9766 16544 9818
rect 16596 9766 16608 9818
rect 16660 9766 16672 9818
rect 16724 9766 16736 9818
rect 16788 9766 16800 9818
rect 16852 9766 21742 9818
rect 21794 9766 21806 9818
rect 21858 9766 21870 9818
rect 21922 9766 21934 9818
rect 21986 9766 21998 9818
rect 22050 9766 22056 9818
rect 1104 9744 22056 9766
rect 2774 9664 2780 9716
rect 2832 9704 2838 9716
rect 3329 9707 3387 9713
rect 3329 9704 3341 9707
rect 2832 9676 3341 9704
rect 2832 9664 2838 9676
rect 3329 9673 3341 9676
rect 3375 9704 3387 9707
rect 3786 9704 3792 9716
rect 3375 9676 3792 9704
rect 3375 9673 3387 9676
rect 3329 9667 3387 9673
rect 3786 9664 3792 9676
rect 3844 9664 3850 9716
rect 3878 9664 3884 9716
rect 3936 9704 3942 9716
rect 8757 9707 8815 9713
rect 8757 9704 8769 9707
rect 3936 9676 8769 9704
rect 3936 9664 3942 9676
rect 8757 9673 8769 9676
rect 8803 9704 8815 9707
rect 9398 9704 9404 9716
rect 8803 9676 9404 9704
rect 8803 9673 8815 9676
rect 8757 9667 8815 9673
rect 9398 9664 9404 9676
rect 9456 9704 9462 9716
rect 9456 9676 9904 9704
rect 9456 9664 9462 9676
rect 6178 9636 6184 9648
rect 2792 9608 6184 9636
rect 1765 9571 1823 9577
rect 1765 9537 1777 9571
rect 1811 9537 1823 9571
rect 2130 9568 2136 9580
rect 2091 9540 2136 9568
rect 1765 9531 1823 9537
rect 1780 9500 1808 9531
rect 2130 9528 2136 9540
rect 2188 9528 2194 9580
rect 2792 9577 2820 9608
rect 6178 9596 6184 9608
rect 6236 9596 6242 9648
rect 6362 9596 6368 9648
rect 6420 9636 6426 9648
rect 6733 9639 6791 9645
rect 6733 9636 6745 9639
rect 6420 9608 6745 9636
rect 6420 9596 6426 9608
rect 6733 9605 6745 9608
rect 6779 9605 6791 9639
rect 6733 9599 6791 9605
rect 9309 9639 9367 9645
rect 9309 9605 9321 9639
rect 9355 9636 9367 9639
rect 9766 9636 9772 9648
rect 9355 9608 9772 9636
rect 9355 9605 9367 9608
rect 9309 9599 9367 9605
rect 9766 9596 9772 9608
rect 9824 9596 9830 9648
rect 9876 9636 9904 9676
rect 10778 9664 10784 9716
rect 10836 9704 10842 9716
rect 12066 9704 12072 9716
rect 10836 9676 11100 9704
rect 12027 9676 12072 9704
rect 10836 9664 10842 9676
rect 10962 9636 10968 9648
rect 9876 9608 10968 9636
rect 10962 9596 10968 9608
rect 11020 9596 11026 9648
rect 11072 9636 11100 9676
rect 12066 9664 12072 9676
rect 12124 9664 12130 9716
rect 13630 9704 13636 9716
rect 12406 9676 13636 9704
rect 12406 9636 12434 9676
rect 13630 9664 13636 9676
rect 13688 9664 13694 9716
rect 15010 9664 15016 9716
rect 15068 9704 15074 9716
rect 19334 9704 19340 9716
rect 15068 9676 19340 9704
rect 15068 9664 15074 9676
rect 19334 9664 19340 9676
rect 19392 9664 19398 9716
rect 19521 9707 19579 9713
rect 19521 9673 19533 9707
rect 19567 9673 19579 9707
rect 19521 9667 19579 9673
rect 11072 9608 12434 9636
rect 14642 9596 14648 9648
rect 14700 9636 14706 9648
rect 16218 9639 16276 9645
rect 16218 9636 16230 9639
rect 14700 9608 16230 9636
rect 14700 9596 14706 9608
rect 16218 9605 16230 9608
rect 16264 9605 16276 9639
rect 19536 9636 19564 9667
rect 19610 9636 19616 9648
rect 16218 9599 16276 9605
rect 16316 9608 18440 9636
rect 19536 9608 19616 9636
rect 2777 9571 2835 9577
rect 2777 9537 2789 9571
rect 2823 9537 2835 9571
rect 2777 9531 2835 9537
rect 2866 9528 2872 9580
rect 2924 9568 2930 9580
rect 3697 9571 3755 9577
rect 2924 9540 2969 9568
rect 2924 9528 2930 9540
rect 3697 9537 3709 9571
rect 3743 9568 3755 9571
rect 4154 9568 4160 9580
rect 3743 9540 4160 9568
rect 3743 9537 3755 9540
rect 3697 9531 3755 9537
rect 4154 9528 4160 9540
rect 4212 9568 4218 9580
rect 4801 9571 4859 9577
rect 4801 9568 4813 9571
rect 4212 9540 4813 9568
rect 4212 9528 4218 9540
rect 4801 9537 4813 9540
rect 4847 9537 4859 9571
rect 4801 9531 4859 9537
rect 4893 9571 4951 9577
rect 4893 9537 4905 9571
rect 4939 9537 4951 9571
rect 4893 9531 4951 9537
rect 2501 9503 2559 9509
rect 2501 9500 2513 9503
rect 1780 9472 2513 9500
rect 2501 9469 2513 9472
rect 2547 9469 2559 9503
rect 3786 9500 3792 9512
rect 3747 9472 3792 9500
rect 2501 9463 2559 9469
rect 3786 9460 3792 9472
rect 3844 9460 3850 9512
rect 4249 9503 4307 9509
rect 4249 9469 4261 9503
rect 4295 9500 4307 9503
rect 4338 9500 4344 9512
rect 4295 9472 4344 9500
rect 4295 9469 4307 9472
rect 4249 9463 4307 9469
rect 4338 9460 4344 9472
rect 4396 9500 4402 9512
rect 4617 9503 4675 9509
rect 4617 9500 4629 9503
rect 4396 9472 4629 9500
rect 4396 9460 4402 9472
rect 4617 9469 4629 9472
rect 4663 9469 4675 9503
rect 4617 9463 4675 9469
rect 1578 9432 1584 9444
rect 1539 9404 1584 9432
rect 1578 9392 1584 9404
rect 1636 9392 1642 9444
rect 1854 9392 1860 9444
rect 1912 9432 1918 9444
rect 1949 9435 2007 9441
rect 1949 9432 1961 9435
rect 1912 9404 1961 9432
rect 1912 9392 1918 9404
rect 1949 9401 1961 9404
rect 1995 9401 2007 9435
rect 1949 9395 2007 9401
rect 3053 9435 3111 9441
rect 3053 9401 3065 9435
rect 3099 9432 3111 9435
rect 3142 9432 3148 9444
rect 3099 9404 3148 9432
rect 3099 9401 3111 9404
rect 3053 9395 3111 9401
rect 3142 9392 3148 9404
rect 3200 9392 3206 9444
rect 3804 9432 3832 9460
rect 4430 9432 4436 9444
rect 3804 9404 4436 9432
rect 4430 9392 4436 9404
rect 4488 9432 4494 9444
rect 4908 9432 4936 9531
rect 5258 9528 5264 9580
rect 5316 9568 5322 9580
rect 5445 9571 5503 9577
rect 5445 9568 5457 9571
rect 5316 9540 5457 9568
rect 5316 9528 5322 9540
rect 5445 9537 5457 9540
rect 5491 9568 5503 9571
rect 5534 9568 5540 9580
rect 5491 9540 5540 9568
rect 5491 9537 5503 9540
rect 5445 9531 5503 9537
rect 5534 9528 5540 9540
rect 5592 9528 5598 9580
rect 6086 9568 6092 9580
rect 6047 9540 6092 9568
rect 6086 9528 6092 9540
rect 6144 9528 6150 9580
rect 6270 9528 6276 9580
rect 6328 9568 6334 9580
rect 6641 9571 6699 9577
rect 6641 9568 6653 9571
rect 6328 9540 6653 9568
rect 6328 9528 6334 9540
rect 6641 9537 6653 9540
rect 6687 9537 6699 9571
rect 6641 9531 6699 9537
rect 10321 9571 10379 9577
rect 10321 9537 10333 9571
rect 10367 9537 10379 9571
rect 10321 9531 10379 9537
rect 10413 9571 10471 9577
rect 10413 9537 10425 9571
rect 10459 9568 10471 9571
rect 11057 9571 11115 9577
rect 11057 9568 11069 9571
rect 10459 9540 11069 9568
rect 10459 9537 10471 9540
rect 10413 9531 10471 9537
rect 11057 9537 11069 9540
rect 11103 9568 11115 9571
rect 12434 9568 12440 9580
rect 11103 9540 12440 9568
rect 11103 9537 11115 9540
rect 11057 9531 11115 9537
rect 5626 9460 5632 9512
rect 5684 9500 5690 9512
rect 6457 9503 6515 9509
rect 6457 9500 6469 9503
rect 5684 9472 6469 9500
rect 5684 9460 5690 9472
rect 6457 9469 6469 9472
rect 6503 9469 6515 9503
rect 9122 9500 9128 9512
rect 9083 9472 9128 9500
rect 6457 9463 6515 9469
rect 4488 9404 4936 9432
rect 5261 9435 5319 9441
rect 4488 9392 4494 9404
rect 5261 9401 5273 9435
rect 5307 9432 5319 9435
rect 5350 9432 5356 9444
rect 5307 9404 5356 9432
rect 5307 9401 5319 9404
rect 5261 9395 5319 9401
rect 5350 9392 5356 9404
rect 5408 9392 5414 9444
rect 5810 9392 5816 9444
rect 5868 9432 5874 9444
rect 5905 9435 5963 9441
rect 5905 9432 5917 9435
rect 5868 9404 5917 9432
rect 5868 9392 5874 9404
rect 5905 9401 5917 9404
rect 5951 9432 5963 9435
rect 6362 9432 6368 9444
rect 5951 9404 6368 9432
rect 5951 9401 5963 9404
rect 5905 9395 5963 9401
rect 6362 9392 6368 9404
rect 6420 9392 6426 9444
rect 6472 9432 6500 9463
rect 9122 9460 9128 9472
rect 9180 9460 9186 9512
rect 9217 9503 9275 9509
rect 9217 9469 9229 9503
rect 9263 9469 9275 9503
rect 10336 9500 10364 9531
rect 12434 9528 12440 9540
rect 12492 9528 12498 9580
rect 12710 9528 12716 9580
rect 12768 9568 12774 9580
rect 13274 9571 13332 9577
rect 13274 9568 13286 9571
rect 12768 9540 13286 9568
rect 12768 9528 12774 9540
rect 13274 9537 13286 9540
rect 13320 9537 13332 9571
rect 13274 9531 13332 9537
rect 13630 9528 13636 9580
rect 13688 9568 13694 9580
rect 14746 9571 14804 9577
rect 14746 9568 14758 9571
rect 13688 9540 14758 9568
rect 13688 9528 13694 9540
rect 14746 9537 14758 9540
rect 14792 9537 14804 9571
rect 14746 9531 14804 9537
rect 15013 9571 15071 9577
rect 15013 9537 15025 9571
rect 15059 9568 15071 9571
rect 15102 9568 15108 9580
rect 15059 9540 15108 9568
rect 15059 9537 15071 9540
rect 15013 9531 15071 9537
rect 15102 9528 15108 9540
rect 15160 9528 15166 9580
rect 15654 9528 15660 9580
rect 15712 9568 15718 9580
rect 16316 9568 16344 9608
rect 16482 9568 16488 9580
rect 15712 9540 16344 9568
rect 16443 9540 16488 9568
rect 15712 9528 15718 9540
rect 16482 9528 16488 9540
rect 16540 9528 16546 9580
rect 17770 9528 17776 9580
rect 17828 9577 17834 9580
rect 18412 9577 18440 9608
rect 19610 9596 19616 9608
rect 19668 9636 19674 9648
rect 20162 9636 20168 9648
rect 19668 9608 20168 9636
rect 19668 9596 19674 9608
rect 20162 9596 20168 9608
rect 20220 9596 20226 9648
rect 17828 9568 17840 9577
rect 18397 9571 18455 9577
rect 17828 9540 17873 9568
rect 17828 9531 17840 9540
rect 18397 9537 18409 9571
rect 18443 9537 18455 9571
rect 18397 9531 18455 9537
rect 17828 9528 17834 9531
rect 18874 9528 18880 9580
rect 18932 9568 18938 9580
rect 19869 9571 19927 9577
rect 19869 9568 19881 9571
rect 18932 9540 19881 9568
rect 18932 9528 18938 9540
rect 19869 9537 19881 9540
rect 19915 9537 19927 9571
rect 19869 9531 19927 9537
rect 10597 9503 10655 9509
rect 10336 9472 10456 9500
rect 9217 9463 9275 9469
rect 6730 9432 6736 9444
rect 6472 9404 6736 9432
rect 6730 9392 6736 9404
rect 6788 9392 6794 9444
rect 7101 9435 7159 9441
rect 7101 9401 7113 9435
rect 7147 9432 7159 9435
rect 7834 9432 7840 9444
rect 7147 9404 7840 9432
rect 7147 9401 7159 9404
rect 7101 9395 7159 9401
rect 7834 9392 7840 9404
rect 7892 9392 7898 9444
rect 3694 9324 3700 9376
rect 3752 9364 3758 9376
rect 3878 9364 3884 9376
rect 3752 9336 3884 9364
rect 3752 9324 3758 9336
rect 3878 9324 3884 9336
rect 3936 9364 3942 9376
rect 3973 9367 4031 9373
rect 3973 9364 3985 9367
rect 3936 9336 3985 9364
rect 3936 9324 3942 9336
rect 3973 9333 3985 9336
rect 4019 9333 4031 9367
rect 3973 9327 4031 9333
rect 4341 9367 4399 9373
rect 4341 9333 4353 9367
rect 4387 9364 4399 9367
rect 4982 9364 4988 9376
rect 4387 9336 4988 9364
rect 4387 9333 4399 9336
rect 4341 9327 4399 9333
rect 4982 9324 4988 9336
rect 5040 9324 5046 9376
rect 5626 9324 5632 9376
rect 5684 9364 5690 9376
rect 5721 9367 5779 9373
rect 5721 9364 5733 9367
rect 5684 9336 5733 9364
rect 5684 9324 5690 9336
rect 5721 9333 5733 9336
rect 5767 9333 5779 9367
rect 5721 9327 5779 9333
rect 7006 9324 7012 9376
rect 7064 9364 7070 9376
rect 7193 9367 7251 9373
rect 7193 9364 7205 9367
rect 7064 9336 7205 9364
rect 7064 9324 7070 9336
rect 7193 9333 7205 9336
rect 7239 9333 7251 9367
rect 7193 9327 7251 9333
rect 7742 9324 7748 9376
rect 7800 9364 7806 9376
rect 8205 9367 8263 9373
rect 8205 9364 8217 9367
rect 7800 9336 8217 9364
rect 7800 9324 7806 9336
rect 8205 9333 8217 9336
rect 8251 9364 8263 9367
rect 8386 9364 8392 9376
rect 8251 9336 8392 9364
rect 8251 9333 8263 9336
rect 8205 9327 8263 9333
rect 8386 9324 8392 9336
rect 8444 9324 8450 9376
rect 8478 9324 8484 9376
rect 8536 9364 8542 9376
rect 8573 9367 8631 9373
rect 8573 9364 8585 9367
rect 8536 9336 8585 9364
rect 8536 9324 8542 9336
rect 8573 9333 8585 9336
rect 8619 9364 8631 9367
rect 9232 9364 9260 9463
rect 9674 9432 9680 9444
rect 9635 9404 9680 9432
rect 9674 9392 9680 9404
rect 9732 9392 9738 9444
rect 9861 9435 9919 9441
rect 9861 9401 9873 9435
rect 9907 9432 9919 9435
rect 10042 9432 10048 9444
rect 9907 9404 10048 9432
rect 9907 9401 9919 9404
rect 9861 9395 9919 9401
rect 10042 9392 10048 9404
rect 10100 9392 10106 9444
rect 8619 9336 9260 9364
rect 9953 9367 10011 9373
rect 8619 9333 8631 9336
rect 8573 9327 8631 9333
rect 9953 9333 9965 9367
rect 9999 9364 10011 9367
rect 10134 9364 10140 9376
rect 9999 9336 10140 9364
rect 9999 9333 10011 9336
rect 9953 9327 10011 9333
rect 10134 9324 10140 9336
rect 10192 9324 10198 9376
rect 10428 9364 10456 9472
rect 10597 9469 10609 9503
rect 10643 9469 10655 9503
rect 10597 9463 10655 9469
rect 10781 9503 10839 9509
rect 10781 9469 10793 9503
rect 10827 9500 10839 9503
rect 10870 9500 10876 9512
rect 10827 9472 10876 9500
rect 10827 9469 10839 9472
rect 10781 9463 10839 9469
rect 10612 9432 10640 9463
rect 10870 9460 10876 9472
rect 10928 9460 10934 9512
rect 13541 9503 13599 9509
rect 10980 9472 12388 9500
rect 10980 9432 11008 9472
rect 11054 9432 11060 9444
rect 10612 9404 11060 9432
rect 11054 9392 11060 9404
rect 11112 9392 11118 9444
rect 11333 9435 11391 9441
rect 11333 9401 11345 9435
rect 11379 9432 11391 9435
rect 11882 9432 11888 9444
rect 11379 9404 11888 9432
rect 11379 9401 11391 9404
rect 11333 9395 11391 9401
rect 11348 9364 11376 9395
rect 11882 9392 11888 9404
rect 11940 9432 11946 9444
rect 12250 9432 12256 9444
rect 11940 9404 12256 9432
rect 11940 9392 11946 9404
rect 12250 9392 12256 9404
rect 12308 9392 12314 9444
rect 10428 9336 11376 9364
rect 11606 9324 11612 9376
rect 11664 9364 11670 9376
rect 12158 9364 12164 9376
rect 11664 9336 12164 9364
rect 11664 9324 11670 9336
rect 12158 9324 12164 9336
rect 12216 9324 12222 9376
rect 12360 9364 12388 9472
rect 13541 9469 13553 9503
rect 13587 9500 13599 9503
rect 13814 9500 13820 9512
rect 13587 9472 13820 9500
rect 13587 9469 13599 9472
rect 13541 9463 13599 9469
rect 13814 9460 13820 9472
rect 13872 9460 13878 9512
rect 18046 9500 18052 9512
rect 18007 9472 18052 9500
rect 18046 9460 18052 9472
rect 18104 9500 18110 9512
rect 18141 9503 18199 9509
rect 18141 9500 18153 9503
rect 18104 9472 18153 9500
rect 18104 9460 18110 9472
rect 18141 9469 18153 9472
rect 18187 9469 18199 9503
rect 18141 9463 18199 9469
rect 19150 9460 19156 9512
rect 19208 9500 19214 9512
rect 19613 9503 19671 9509
rect 19613 9500 19625 9503
rect 19208 9472 19625 9500
rect 19208 9460 19214 9472
rect 19613 9469 19625 9472
rect 19659 9469 19671 9503
rect 19613 9463 19671 9469
rect 13998 9432 14004 9444
rect 13556 9404 14004 9432
rect 13556 9364 13584 9404
rect 13998 9392 14004 9404
rect 14056 9392 14062 9444
rect 12360 9336 13584 9364
rect 13906 9324 13912 9376
rect 13964 9364 13970 9376
rect 14826 9364 14832 9376
rect 13964 9336 14832 9364
rect 13964 9324 13970 9336
rect 14826 9324 14832 9336
rect 14884 9364 14890 9376
rect 15105 9367 15163 9373
rect 15105 9364 15117 9367
rect 14884 9336 15117 9364
rect 14884 9324 14890 9336
rect 15105 9333 15117 9336
rect 15151 9333 15163 9367
rect 15105 9327 15163 9333
rect 16669 9367 16727 9373
rect 16669 9333 16681 9367
rect 16715 9364 16727 9367
rect 16942 9364 16948 9376
rect 16715 9336 16948 9364
rect 16715 9333 16727 9336
rect 16669 9327 16727 9333
rect 16942 9324 16948 9336
rect 17000 9324 17006 9376
rect 19628 9364 19656 9463
rect 20548 9404 21220 9432
rect 20548 9364 20576 9404
rect 19628 9336 20576 9364
rect 20806 9324 20812 9376
rect 20864 9364 20870 9376
rect 21192 9373 21220 9404
rect 20993 9367 21051 9373
rect 20993 9364 21005 9367
rect 20864 9336 21005 9364
rect 20864 9324 20870 9336
rect 20993 9333 21005 9336
rect 21039 9333 21051 9367
rect 20993 9327 21051 9333
rect 21177 9367 21235 9373
rect 21177 9333 21189 9367
rect 21223 9364 21235 9367
rect 21266 9364 21272 9376
rect 21223 9336 21272 9364
rect 21223 9333 21235 9336
rect 21177 9327 21235 9333
rect 21266 9324 21272 9336
rect 21324 9324 21330 9376
rect 1104 9274 21896 9296
rect 1104 9222 3549 9274
rect 3601 9222 3613 9274
rect 3665 9222 3677 9274
rect 3729 9222 3741 9274
rect 3793 9222 3805 9274
rect 3857 9222 8747 9274
rect 8799 9222 8811 9274
rect 8863 9222 8875 9274
rect 8927 9222 8939 9274
rect 8991 9222 9003 9274
rect 9055 9222 13945 9274
rect 13997 9222 14009 9274
rect 14061 9222 14073 9274
rect 14125 9222 14137 9274
rect 14189 9222 14201 9274
rect 14253 9222 19143 9274
rect 19195 9222 19207 9274
rect 19259 9222 19271 9274
rect 19323 9222 19335 9274
rect 19387 9222 19399 9274
rect 19451 9222 21896 9274
rect 1104 9200 21896 9222
rect 1670 9160 1676 9172
rect 1631 9132 1676 9160
rect 1670 9120 1676 9132
rect 1728 9160 1734 9172
rect 2038 9160 2044 9172
rect 1728 9132 2044 9160
rect 1728 9120 1734 9132
rect 2038 9120 2044 9132
rect 2096 9160 2102 9172
rect 2961 9163 3019 9169
rect 2096 9132 2636 9160
rect 2096 9120 2102 9132
rect 1949 9095 2007 9101
rect 1949 9061 1961 9095
rect 1995 9092 2007 9095
rect 2222 9092 2228 9104
rect 1995 9064 2228 9092
rect 1995 9061 2007 9064
rect 1949 9055 2007 9061
rect 2222 9052 2228 9064
rect 2280 9052 2286 9104
rect 2409 9027 2467 9033
rect 2409 8993 2421 9027
rect 2455 9024 2467 9027
rect 2498 9024 2504 9036
rect 2455 8996 2504 9024
rect 2455 8993 2467 8996
rect 2409 8987 2467 8993
rect 2498 8984 2504 8996
rect 2556 8984 2562 9036
rect 1670 8916 1676 8968
rect 1728 8956 1734 8968
rect 2608 8965 2636 9132
rect 2961 9129 2973 9163
rect 3007 9160 3019 9163
rect 5902 9160 5908 9172
rect 3007 9132 5908 9160
rect 3007 9129 3019 9132
rect 2961 9123 3019 9129
rect 5902 9120 5908 9132
rect 5960 9120 5966 9172
rect 6089 9163 6147 9169
rect 6089 9129 6101 9163
rect 6135 9160 6147 9163
rect 6546 9160 6552 9172
rect 6135 9132 6552 9160
rect 6135 9129 6147 9132
rect 6089 9123 6147 9129
rect 6546 9120 6552 9132
rect 6604 9120 6610 9172
rect 8018 9120 8024 9172
rect 8076 9160 8082 9172
rect 9493 9163 9551 9169
rect 9493 9160 9505 9163
rect 8076 9132 9505 9160
rect 8076 9120 8082 9132
rect 9493 9129 9505 9132
rect 9539 9160 9551 9163
rect 9582 9160 9588 9172
rect 9539 9132 9588 9160
rect 9539 9129 9551 9132
rect 9493 9123 9551 9129
rect 9582 9120 9588 9132
rect 9640 9120 9646 9172
rect 9677 9163 9735 9169
rect 9677 9129 9689 9163
rect 9723 9160 9735 9163
rect 9858 9160 9864 9172
rect 9723 9132 9864 9160
rect 9723 9129 9735 9132
rect 9677 9123 9735 9129
rect 9858 9120 9864 9132
rect 9916 9120 9922 9172
rect 11790 9160 11796 9172
rect 9968 9132 11796 9160
rect 3528 9064 5028 9092
rect 3234 9024 3240 9036
rect 3195 8996 3240 9024
rect 3234 8984 3240 8996
rect 3292 8984 3298 9036
rect 3528 8965 3556 9064
rect 3970 8984 3976 9036
rect 4028 9024 4034 9036
rect 4614 9024 4620 9036
rect 4028 8996 4476 9024
rect 4575 8996 4620 9024
rect 4028 8984 4034 8996
rect 2133 8959 2191 8965
rect 2133 8956 2145 8959
rect 1728 8928 2145 8956
rect 1728 8916 1734 8928
rect 2133 8925 2145 8928
rect 2179 8925 2191 8959
rect 2133 8919 2191 8925
rect 2593 8959 2651 8965
rect 2593 8925 2605 8959
rect 2639 8925 2651 8959
rect 2593 8919 2651 8925
rect 3513 8959 3571 8965
rect 3513 8925 3525 8959
rect 3559 8925 3571 8959
rect 4338 8956 4344 8968
rect 4299 8928 4344 8956
rect 3513 8919 3571 8925
rect 4338 8916 4344 8928
rect 4396 8916 4402 8968
rect 4448 8956 4476 8996
rect 4614 8984 4620 8996
rect 4672 8984 4678 9036
rect 4893 8959 4951 8965
rect 4893 8956 4905 8959
rect 4448 8928 4905 8956
rect 4893 8925 4905 8928
rect 4939 8925 4951 8959
rect 5000 8956 5028 9064
rect 5074 9052 5080 9104
rect 5132 9092 5138 9104
rect 5261 9095 5319 9101
rect 5261 9092 5273 9095
rect 5132 9064 5273 9092
rect 5132 9052 5138 9064
rect 5261 9061 5273 9064
rect 5307 9061 5319 9095
rect 7009 9095 7067 9101
rect 7009 9092 7021 9095
rect 5261 9055 5319 9061
rect 5368 9064 7021 9092
rect 5368 8956 5396 9064
rect 7009 9061 7021 9064
rect 7055 9061 7067 9095
rect 7009 9055 7067 9061
rect 7834 9052 7840 9104
rect 7892 9092 7898 9104
rect 8202 9092 8208 9104
rect 7892 9064 8208 9092
rect 7892 9052 7898 9064
rect 8202 9052 8208 9064
rect 8260 9052 8266 9104
rect 9968 9092 9996 9132
rect 11790 9120 11796 9132
rect 11848 9120 11854 9172
rect 13630 9160 13636 9172
rect 12406 9132 13636 9160
rect 12253 9095 12311 9101
rect 12253 9092 12265 9095
rect 8404 9064 9996 9092
rect 11900 9064 12265 9092
rect 5445 9027 5503 9033
rect 5445 8993 5457 9027
rect 5491 8993 5503 9027
rect 5445 8987 5503 8993
rect 5629 9027 5687 9033
rect 5629 8993 5641 9027
rect 5675 9024 5687 9027
rect 6086 9024 6092 9036
rect 5675 8996 6092 9024
rect 5675 8993 5687 8996
rect 5629 8987 5687 8993
rect 5000 8928 5396 8956
rect 4893 8919 4951 8925
rect 1581 8891 1639 8897
rect 1581 8857 1593 8891
rect 1627 8888 1639 8891
rect 2501 8891 2559 8897
rect 2501 8888 2513 8891
rect 1627 8860 2513 8888
rect 1627 8857 1639 8860
rect 1581 8851 1639 8857
rect 2501 8857 2513 8860
rect 2547 8888 2559 8891
rect 3142 8888 3148 8900
rect 2547 8860 3148 8888
rect 2547 8857 2559 8860
rect 2501 8851 2559 8857
rect 3142 8848 3148 8860
rect 3200 8848 3206 8900
rect 3418 8848 3424 8900
rect 3476 8888 3482 8900
rect 4065 8891 4123 8897
rect 4065 8888 4077 8891
rect 3476 8860 4077 8888
rect 3476 8848 3482 8860
rect 4065 8857 4077 8860
rect 4111 8857 4123 8891
rect 4065 8851 4123 8857
rect 5074 8848 5080 8900
rect 5132 8888 5138 8900
rect 5460 8888 5488 8987
rect 6086 8984 6092 8996
rect 6144 8984 6150 9036
rect 6822 9024 6828 9036
rect 6783 8996 6828 9024
rect 6822 8984 6828 8996
rect 6880 8984 6886 9036
rect 7650 9024 7656 9036
rect 7611 8996 7656 9024
rect 7650 8984 7656 8996
rect 7708 8984 7714 9036
rect 8110 8984 8116 9036
rect 8168 9024 8174 9036
rect 8404 9033 8432 9064
rect 8389 9027 8447 9033
rect 8389 9024 8401 9027
rect 8168 8996 8401 9024
rect 8168 8984 8174 8996
rect 8389 8993 8401 8996
rect 8435 8993 8447 9027
rect 8389 8987 8447 8993
rect 9582 8984 9588 9036
rect 9640 9024 9646 9036
rect 9640 8996 10088 9024
rect 9640 8984 9646 8996
rect 7466 8916 7472 8968
rect 7524 8956 7530 8968
rect 9950 8956 9956 8968
rect 7524 8928 9956 8956
rect 7524 8916 7530 8928
rect 9950 8916 9956 8928
rect 10008 8916 10014 8968
rect 10060 8956 10088 8996
rect 10134 8984 10140 9036
rect 10192 9024 10198 9036
rect 10318 9024 10324 9036
rect 10192 8996 10237 9024
rect 10279 8996 10324 9024
rect 10192 8984 10198 8996
rect 10318 8984 10324 8996
rect 10376 8984 10382 9036
rect 10686 9024 10692 9036
rect 10647 8996 10692 9024
rect 10686 8984 10692 8996
rect 10744 8984 10750 9036
rect 11900 9024 11928 9064
rect 12253 9061 12265 9064
rect 12299 9092 12311 9095
rect 12406 9092 12434 9132
rect 13630 9120 13636 9132
rect 13688 9120 13694 9172
rect 15657 9163 15715 9169
rect 15657 9160 15669 9163
rect 14108 9132 15669 9160
rect 12299 9064 12434 9092
rect 12299 9061 12311 9064
rect 12253 9055 12311 9061
rect 10980 8996 11928 9024
rect 11977 9027 12035 9033
rect 10594 8956 10600 8968
rect 10060 8928 10600 8956
rect 10594 8916 10600 8928
rect 10652 8956 10658 8968
rect 10781 8959 10839 8965
rect 10781 8956 10793 8959
rect 10652 8928 10793 8956
rect 10652 8916 10658 8928
rect 10781 8925 10793 8928
rect 10827 8925 10839 8959
rect 10781 8919 10839 8925
rect 5718 8888 5724 8900
rect 5132 8860 5488 8888
rect 5679 8860 5724 8888
rect 5132 8848 5138 8860
rect 5718 8848 5724 8860
rect 5776 8848 5782 8900
rect 7282 8888 7288 8900
rect 6012 8860 7288 8888
rect 3694 8780 3700 8832
rect 3752 8820 3758 8832
rect 4801 8823 4859 8829
rect 4801 8820 4813 8823
rect 3752 8792 4813 8820
rect 3752 8780 3758 8792
rect 4801 8789 4813 8792
rect 4847 8820 4859 8823
rect 6012 8820 6040 8860
rect 7282 8848 7288 8860
rect 7340 8848 7346 8900
rect 7377 8891 7435 8897
rect 7377 8857 7389 8891
rect 7423 8888 7435 8891
rect 7423 8860 7880 8888
rect 7423 8857 7435 8860
rect 7377 8851 7435 8857
rect 6178 8820 6184 8832
rect 4847 8792 6040 8820
rect 6139 8792 6184 8820
rect 4847 8789 4859 8792
rect 4801 8783 4859 8789
rect 6178 8780 6184 8792
rect 6236 8780 6242 8832
rect 6546 8820 6552 8832
rect 6507 8792 6552 8820
rect 6546 8780 6552 8792
rect 6604 8780 6610 8832
rect 6638 8780 6644 8832
rect 6696 8820 6702 8832
rect 7466 8820 7472 8832
rect 6696 8792 6741 8820
rect 7427 8792 7472 8820
rect 6696 8780 6702 8792
rect 7466 8780 7472 8792
rect 7524 8780 7530 8832
rect 7852 8829 7880 8860
rect 9122 8848 9128 8900
rect 9180 8888 9186 8900
rect 9490 8888 9496 8900
rect 9180 8860 9496 8888
rect 9180 8848 9186 8860
rect 9490 8848 9496 8860
rect 9548 8848 9554 8900
rect 9582 8848 9588 8900
rect 9640 8888 9646 8900
rect 10980 8888 11008 8996
rect 11977 8993 11989 9027
rect 12023 8993 12035 9027
rect 11977 8987 12035 8993
rect 13633 9027 13691 9033
rect 13633 8993 13645 9027
rect 13679 9024 13691 9027
rect 13814 9024 13820 9036
rect 13679 8996 13820 9024
rect 13679 8993 13691 8996
rect 13633 8987 13691 8993
rect 11992 8956 12020 8987
rect 13814 8984 13820 8996
rect 13872 9024 13878 9036
rect 14108 9033 14136 9132
rect 15657 9129 15669 9132
rect 15703 9160 15715 9163
rect 15746 9160 15752 9172
rect 15703 9132 15752 9160
rect 15703 9129 15715 9132
rect 15657 9123 15715 9129
rect 15746 9120 15752 9132
rect 15804 9160 15810 9172
rect 15841 9163 15899 9169
rect 15841 9160 15853 9163
rect 15804 9132 15853 9160
rect 15804 9120 15810 9132
rect 15841 9129 15853 9132
rect 15887 9160 15899 9163
rect 16025 9163 16083 9169
rect 16025 9160 16037 9163
rect 15887 9132 16037 9160
rect 15887 9129 15899 9132
rect 15841 9123 15899 9129
rect 16025 9129 16037 9132
rect 16071 9160 16083 9163
rect 16209 9163 16267 9169
rect 16209 9160 16221 9163
rect 16071 9132 16221 9160
rect 16071 9129 16083 9132
rect 16025 9123 16083 9129
rect 16209 9129 16221 9132
rect 16255 9160 16267 9163
rect 16482 9160 16488 9172
rect 16255 9132 16488 9160
rect 16255 9129 16267 9132
rect 16209 9123 16267 9129
rect 16316 9033 16344 9132
rect 16482 9120 16488 9132
rect 16540 9160 16546 9172
rect 17865 9163 17923 9169
rect 17865 9160 17877 9163
rect 16540 9132 17877 9160
rect 16540 9120 16546 9132
rect 17865 9129 17877 9132
rect 17911 9160 17923 9163
rect 18046 9160 18052 9172
rect 17911 9132 18052 9160
rect 17911 9129 17923 9132
rect 17865 9123 17923 9129
rect 18046 9120 18052 9132
rect 18104 9160 18110 9172
rect 18233 9163 18291 9169
rect 18233 9160 18245 9163
rect 18104 9132 18245 9160
rect 18104 9120 18110 9132
rect 18233 9129 18245 9132
rect 18279 9160 18291 9163
rect 19058 9160 19064 9172
rect 18279 9132 19064 9160
rect 18279 9129 18291 9132
rect 18233 9123 18291 9129
rect 19058 9120 19064 9132
rect 19116 9120 19122 9172
rect 14093 9027 14151 9033
rect 14093 9024 14105 9027
rect 13872 8996 14105 9024
rect 13872 8984 13878 8996
rect 14093 8993 14105 8996
rect 14139 8993 14151 9027
rect 14093 8987 14151 8993
rect 16301 9027 16359 9033
rect 16301 8993 16313 9027
rect 16347 8993 16359 9027
rect 16301 8987 16359 8993
rect 18874 8956 18880 8968
rect 11992 8928 18880 8956
rect 18874 8916 18880 8928
rect 18932 8916 18938 8968
rect 20070 8956 20076 8968
rect 19628 8928 20076 8956
rect 11701 8891 11759 8897
rect 11701 8888 11713 8891
rect 9640 8860 11008 8888
rect 11256 8860 11713 8888
rect 9640 8848 9646 8860
rect 7837 8823 7895 8829
rect 7837 8789 7849 8823
rect 7883 8789 7895 8823
rect 8202 8820 8208 8832
rect 8163 8792 8208 8820
rect 7837 8783 7895 8789
rect 8202 8780 8208 8792
rect 8260 8780 8266 8832
rect 8297 8823 8355 8829
rect 8297 8789 8309 8823
rect 8343 8820 8355 8823
rect 8570 8820 8576 8832
rect 8343 8792 8576 8820
rect 8343 8789 8355 8792
rect 8297 8783 8355 8789
rect 8570 8780 8576 8792
rect 8628 8780 8634 8832
rect 8662 8780 8668 8832
rect 8720 8820 8726 8832
rect 10045 8823 10103 8829
rect 8720 8792 8765 8820
rect 8720 8780 8726 8792
rect 10045 8789 10057 8823
rect 10091 8820 10103 8823
rect 10502 8820 10508 8832
rect 10091 8792 10508 8820
rect 10091 8789 10103 8792
rect 10045 8783 10103 8789
rect 10502 8780 10508 8792
rect 10560 8780 10566 8832
rect 10870 8820 10876 8832
rect 10831 8792 10876 8820
rect 10870 8780 10876 8792
rect 10928 8780 10934 8832
rect 11256 8829 11284 8860
rect 11701 8857 11713 8860
rect 11747 8857 11759 8891
rect 11701 8851 11759 8857
rect 13262 8848 13268 8900
rect 13320 8888 13326 8900
rect 13366 8891 13424 8897
rect 13366 8888 13378 8891
rect 13320 8860 13378 8888
rect 13320 8848 13326 8860
rect 13366 8857 13378 8860
rect 13412 8857 13424 8891
rect 13366 8851 13424 8857
rect 13538 8848 13544 8900
rect 13596 8888 13602 8900
rect 14338 8891 14396 8897
rect 14338 8888 14350 8891
rect 13596 8860 14350 8888
rect 13596 8848 13602 8860
rect 14338 8857 14350 8860
rect 14384 8857 14396 8891
rect 16206 8888 16212 8900
rect 14338 8851 14396 8857
rect 15212 8860 16212 8888
rect 11241 8823 11299 8829
rect 11241 8789 11253 8823
rect 11287 8789 11299 8823
rect 11241 8783 11299 8789
rect 11330 8780 11336 8832
rect 11388 8820 11394 8832
rect 11790 8820 11796 8832
rect 11388 8792 11433 8820
rect 11751 8792 11796 8820
rect 11388 8780 11394 8792
rect 11790 8780 11796 8792
rect 11848 8780 11854 8832
rect 12434 8780 12440 8832
rect 12492 8820 12498 8832
rect 15212 8820 15240 8860
rect 16206 8848 16212 8860
rect 16264 8848 16270 8900
rect 16568 8891 16626 8897
rect 16568 8857 16580 8891
rect 16614 8857 16626 8891
rect 16568 8851 16626 8857
rect 12492 8792 15240 8820
rect 12492 8780 12498 8792
rect 15286 8780 15292 8832
rect 15344 8820 15350 8832
rect 15473 8823 15531 8829
rect 15473 8820 15485 8823
rect 15344 8792 15485 8820
rect 15344 8780 15350 8792
rect 15473 8789 15485 8792
rect 15519 8789 15531 8823
rect 16592 8820 16620 8851
rect 16942 8848 16948 8900
rect 17000 8888 17006 8900
rect 19628 8888 19656 8928
rect 20070 8916 20076 8928
rect 20128 8916 20134 8968
rect 20625 8959 20683 8965
rect 20625 8925 20637 8959
rect 20671 8956 20683 8959
rect 20671 8928 20852 8956
rect 20671 8925 20683 8928
rect 20625 8919 20683 8925
rect 17000 8860 19656 8888
rect 17000 8848 17006 8860
rect 19702 8848 19708 8900
rect 19760 8888 19766 8900
rect 20358 8891 20416 8897
rect 20358 8888 20370 8891
rect 19760 8860 20370 8888
rect 19760 8848 19766 8860
rect 20358 8857 20370 8860
rect 20404 8857 20416 8891
rect 20358 8851 20416 8857
rect 17034 8820 17040 8832
rect 16592 8792 17040 8820
rect 15473 8783 15531 8789
rect 17034 8780 17040 8792
rect 17092 8780 17098 8832
rect 17586 8780 17592 8832
rect 17644 8820 17650 8832
rect 17681 8823 17739 8829
rect 17681 8820 17693 8823
rect 17644 8792 17693 8820
rect 17644 8780 17650 8792
rect 17681 8789 17693 8792
rect 17727 8789 17739 8823
rect 17681 8783 17739 8789
rect 18874 8780 18880 8832
rect 18932 8820 18938 8832
rect 20824 8829 20852 8928
rect 19245 8823 19303 8829
rect 19245 8820 19257 8823
rect 18932 8792 19257 8820
rect 18932 8780 18938 8792
rect 19245 8789 19257 8792
rect 19291 8789 19303 8823
rect 19245 8783 19303 8789
rect 20809 8823 20867 8829
rect 20809 8789 20821 8823
rect 20855 8820 20867 8823
rect 21266 8820 21272 8832
rect 20855 8792 21272 8820
rect 20855 8789 20867 8792
rect 20809 8783 20867 8789
rect 21266 8780 21272 8792
rect 21324 8780 21330 8832
rect 1104 8730 22056 8752
rect 1104 8678 6148 8730
rect 6200 8678 6212 8730
rect 6264 8678 6276 8730
rect 6328 8678 6340 8730
rect 6392 8678 6404 8730
rect 6456 8678 11346 8730
rect 11398 8678 11410 8730
rect 11462 8678 11474 8730
rect 11526 8678 11538 8730
rect 11590 8678 11602 8730
rect 11654 8678 16544 8730
rect 16596 8678 16608 8730
rect 16660 8678 16672 8730
rect 16724 8678 16736 8730
rect 16788 8678 16800 8730
rect 16852 8678 21742 8730
rect 21794 8678 21806 8730
rect 21858 8678 21870 8730
rect 21922 8678 21934 8730
rect 21986 8678 21998 8730
rect 22050 8678 22056 8730
rect 1104 8656 22056 8678
rect 1486 8576 1492 8628
rect 1544 8616 1550 8628
rect 2225 8619 2283 8625
rect 2225 8616 2237 8619
rect 1544 8588 2237 8616
rect 1544 8576 1550 8588
rect 2225 8585 2237 8588
rect 2271 8585 2283 8619
rect 2225 8579 2283 8585
rect 2593 8619 2651 8625
rect 2593 8585 2605 8619
rect 2639 8616 2651 8619
rect 4801 8619 4859 8625
rect 2639 8588 4752 8616
rect 2639 8585 2651 8588
rect 2593 8579 2651 8585
rect 2130 8508 2136 8560
rect 2188 8548 2194 8560
rect 2869 8551 2927 8557
rect 2869 8548 2881 8551
rect 2188 8520 2881 8548
rect 2188 8508 2194 8520
rect 2869 8517 2881 8520
rect 2915 8517 2927 8551
rect 3237 8551 3295 8557
rect 3237 8548 3249 8551
rect 2869 8511 2927 8517
rect 3068 8520 3249 8548
rect 1504 8452 2176 8480
rect 1394 8304 1400 8356
rect 1452 8344 1458 8356
rect 1504 8353 1532 8452
rect 2148 8421 2176 8452
rect 2774 8440 2780 8492
rect 2832 8480 2838 8492
rect 3068 8480 3096 8520
rect 3237 8517 3249 8520
rect 3283 8517 3295 8551
rect 4724 8548 4752 8588
rect 4801 8585 4813 8619
rect 4847 8616 4859 8619
rect 6181 8619 6239 8625
rect 4847 8588 6132 8616
rect 4847 8585 4859 8588
rect 4801 8579 4859 8585
rect 5166 8548 5172 8560
rect 4724 8520 5172 8548
rect 3237 8511 3295 8517
rect 5166 8508 5172 8520
rect 5224 8508 5230 8560
rect 6104 8548 6132 8588
rect 6181 8585 6193 8619
rect 6227 8616 6239 8619
rect 6546 8616 6552 8628
rect 6227 8588 6552 8616
rect 6227 8585 6239 8588
rect 6181 8579 6239 8585
rect 6546 8576 6552 8588
rect 6604 8576 6610 8628
rect 6822 8576 6828 8628
rect 6880 8616 6886 8628
rect 7926 8616 7932 8628
rect 6880 8588 7932 8616
rect 6880 8576 6886 8588
rect 7926 8576 7932 8588
rect 7984 8616 7990 8628
rect 8662 8616 8668 8628
rect 7984 8588 8668 8616
rect 7984 8576 7990 8588
rect 8662 8576 8668 8588
rect 8720 8616 8726 8628
rect 8941 8619 8999 8625
rect 8941 8616 8953 8619
rect 8720 8588 8953 8616
rect 8720 8576 8726 8588
rect 8941 8585 8953 8588
rect 8987 8585 8999 8619
rect 9950 8616 9956 8628
rect 9911 8588 9956 8616
rect 8941 8579 8999 8585
rect 9950 8576 9956 8588
rect 10008 8576 10014 8628
rect 10502 8616 10508 8628
rect 10463 8588 10508 8616
rect 10502 8576 10508 8588
rect 10560 8576 10566 8628
rect 10594 8576 10600 8628
rect 10652 8616 10658 8628
rect 10965 8619 11023 8625
rect 10965 8616 10977 8619
rect 10652 8588 10977 8616
rect 10652 8576 10658 8588
rect 10965 8585 10977 8588
rect 11011 8585 11023 8619
rect 13814 8616 13820 8628
rect 13775 8588 13820 8616
rect 10965 8579 11023 8585
rect 13814 8576 13820 8588
rect 13872 8576 13878 8628
rect 14550 8576 14556 8628
rect 14608 8616 14614 8628
rect 15102 8616 15108 8628
rect 14608 8588 15108 8616
rect 14608 8576 14614 8588
rect 15102 8576 15108 8588
rect 15160 8576 15166 8628
rect 15746 8616 15752 8628
rect 15707 8588 15752 8616
rect 15746 8576 15752 8588
rect 15804 8576 15810 8628
rect 18874 8576 18880 8628
rect 18932 8616 18938 8628
rect 18932 8588 19104 8616
rect 18932 8576 18938 8588
rect 6104 8520 7420 8548
rect 2832 8452 3096 8480
rect 3145 8483 3203 8489
rect 2832 8440 2838 8452
rect 3145 8449 3157 8483
rect 3191 8449 3203 8483
rect 3145 8443 3203 8449
rect 2041 8415 2099 8421
rect 2041 8381 2053 8415
rect 2087 8381 2099 8415
rect 2041 8375 2099 8381
rect 2133 8415 2191 8421
rect 2133 8381 2145 8415
rect 2179 8381 2191 8415
rect 2133 8375 2191 8381
rect 1489 8347 1547 8353
rect 1489 8344 1501 8347
rect 1452 8316 1501 8344
rect 1452 8304 1458 8316
rect 1489 8313 1501 8316
rect 1535 8313 1547 8347
rect 1670 8344 1676 8356
rect 1631 8316 1676 8344
rect 1489 8307 1547 8313
rect 1670 8304 1676 8316
rect 1728 8304 1734 8356
rect 2056 8344 2084 8375
rect 2774 8344 2780 8356
rect 2056 8316 2780 8344
rect 2774 8304 2780 8316
rect 2832 8304 2838 8356
rect 3160 8344 3188 8443
rect 3326 8440 3332 8492
rect 3384 8480 3390 8492
rect 3513 8483 3571 8489
rect 3513 8480 3525 8483
rect 3384 8452 3525 8480
rect 3384 8440 3390 8452
rect 3513 8449 3525 8452
rect 3559 8480 3571 8483
rect 3970 8480 3976 8492
rect 3559 8452 3832 8480
rect 3931 8452 3976 8480
rect 3559 8449 3571 8452
rect 3513 8443 3571 8449
rect 3418 8372 3424 8424
rect 3476 8412 3482 8424
rect 3694 8412 3700 8424
rect 3476 8384 3700 8412
rect 3476 8372 3482 8384
rect 3694 8372 3700 8384
rect 3752 8372 3758 8424
rect 3804 8412 3832 8452
rect 3970 8440 3976 8452
rect 4028 8440 4034 8492
rect 4341 8483 4399 8489
rect 4341 8480 4353 8483
rect 4080 8452 4353 8480
rect 4080 8412 4108 8452
rect 4341 8449 4353 8452
rect 4387 8449 4399 8483
rect 4341 8443 4399 8449
rect 4433 8483 4491 8489
rect 4433 8449 4445 8483
rect 4479 8480 4491 8483
rect 4893 8483 4951 8489
rect 4893 8480 4905 8483
rect 4479 8452 4905 8480
rect 4479 8449 4491 8452
rect 4433 8443 4491 8449
rect 4893 8449 4905 8452
rect 4939 8449 4951 8483
rect 4893 8443 4951 8449
rect 5813 8483 5871 8489
rect 5813 8449 5825 8483
rect 5859 8480 5871 8483
rect 5994 8480 6000 8492
rect 5859 8452 6000 8480
rect 5859 8449 5871 8452
rect 5813 8443 5871 8449
rect 5994 8440 6000 8452
rect 6052 8440 6058 8492
rect 6641 8483 6699 8489
rect 6641 8449 6653 8483
rect 6687 8480 6699 8483
rect 6914 8480 6920 8492
rect 6687 8452 6920 8480
rect 6687 8449 6699 8452
rect 6641 8443 6699 8449
rect 6914 8440 6920 8452
rect 6972 8440 6978 8492
rect 7282 8480 7288 8492
rect 7243 8452 7288 8480
rect 7282 8440 7288 8452
rect 7340 8440 7346 8492
rect 7392 8480 7420 8520
rect 7650 8508 7656 8560
rect 7708 8548 7714 8560
rect 7834 8548 7840 8560
rect 7708 8520 7840 8548
rect 7708 8508 7714 8520
rect 7834 8508 7840 8520
rect 7892 8548 7898 8560
rect 8021 8551 8079 8557
rect 8021 8548 8033 8551
rect 7892 8520 8033 8548
rect 7892 8508 7898 8520
rect 8021 8517 8033 8520
rect 8067 8517 8079 8551
rect 8021 8511 8079 8517
rect 8113 8551 8171 8557
rect 8113 8517 8125 8551
rect 8159 8548 8171 8551
rect 9401 8551 9459 8557
rect 9401 8548 9413 8551
rect 8159 8520 9413 8548
rect 8159 8517 8171 8520
rect 8113 8511 8171 8517
rect 9401 8517 9413 8520
rect 9447 8517 9459 8551
rect 9401 8511 9459 8517
rect 10045 8483 10103 8489
rect 10045 8480 10057 8483
rect 7392 8452 10057 8480
rect 10045 8449 10057 8452
rect 10091 8449 10103 8483
rect 10045 8443 10103 8449
rect 10873 8483 10931 8489
rect 10873 8449 10885 8483
rect 10919 8480 10931 8483
rect 11517 8483 11575 8489
rect 11517 8480 11529 8483
rect 10919 8452 11529 8480
rect 10919 8449 10931 8452
rect 10873 8443 10931 8449
rect 11517 8449 11529 8452
rect 11563 8449 11575 8483
rect 11517 8443 11575 8449
rect 15378 8440 15384 8492
rect 15436 8489 15442 8492
rect 15436 8480 15448 8489
rect 15657 8483 15715 8489
rect 15436 8452 15481 8480
rect 15436 8443 15448 8452
rect 15657 8449 15669 8483
rect 15703 8480 15715 8483
rect 15764 8480 15792 8576
rect 18966 8508 18972 8560
rect 19024 8508 19030 8560
rect 19076 8548 19104 8588
rect 20622 8576 20628 8628
rect 20680 8616 20686 8628
rect 20809 8619 20867 8625
rect 20809 8616 20821 8619
rect 20680 8588 20821 8616
rect 20680 8576 20686 8588
rect 20809 8585 20821 8588
rect 20855 8585 20867 8619
rect 20809 8579 20867 8585
rect 19674 8551 19732 8557
rect 19674 8548 19686 8551
rect 19076 8520 19686 8548
rect 19674 8517 19686 8520
rect 19720 8517 19732 8551
rect 19674 8511 19732 8517
rect 15703 8452 15792 8480
rect 15703 8449 15715 8452
rect 15657 8443 15715 8449
rect 15436 8440 15442 8443
rect 17310 8440 17316 8492
rect 17368 8480 17374 8492
rect 18984 8480 19012 8508
rect 19070 8483 19128 8489
rect 19070 8480 19082 8483
rect 17368 8452 19082 8480
rect 17368 8440 17374 8452
rect 19070 8449 19082 8452
rect 19116 8449 19128 8483
rect 19070 8443 19128 8449
rect 3804 8384 4108 8412
rect 4249 8415 4307 8421
rect 4249 8381 4261 8415
rect 4295 8412 4307 8415
rect 4614 8412 4620 8424
rect 4295 8384 4620 8412
rect 4295 8381 4307 8384
rect 4249 8375 4307 8381
rect 4614 8372 4620 8384
rect 4672 8412 4678 8424
rect 5074 8412 5080 8424
rect 4672 8384 5080 8412
rect 4672 8372 4678 8384
rect 5074 8372 5080 8384
rect 5132 8372 5138 8424
rect 5442 8372 5448 8424
rect 5500 8412 5506 8424
rect 5537 8415 5595 8421
rect 5537 8412 5549 8415
rect 5500 8384 5549 8412
rect 5500 8372 5506 8384
rect 5537 8381 5549 8384
rect 5583 8381 5595 8415
rect 5718 8412 5724 8424
rect 5679 8384 5724 8412
rect 5537 8375 5595 8381
rect 5718 8372 5724 8384
rect 5776 8372 5782 8424
rect 7374 8412 7380 8424
rect 7335 8384 7380 8412
rect 7374 8372 7380 8384
rect 7432 8372 7438 8424
rect 7558 8412 7564 8424
rect 7519 8384 7564 8412
rect 7558 8372 7564 8384
rect 7616 8372 7622 8424
rect 7929 8415 7987 8421
rect 7929 8381 7941 8415
rect 7975 8412 7987 8415
rect 7975 8384 8616 8412
rect 7975 8381 7987 8384
rect 7929 8375 7987 8381
rect 6917 8347 6975 8353
rect 6917 8344 6929 8347
rect 3160 8316 6929 8344
rect 6917 8313 6929 8316
rect 6963 8313 6975 8347
rect 6917 8307 6975 8313
rect 5074 8236 5080 8288
rect 5132 8276 5138 8288
rect 5261 8279 5319 8285
rect 5261 8276 5273 8279
rect 5132 8248 5273 8276
rect 5132 8236 5138 8248
rect 5261 8245 5273 8248
rect 5307 8245 5319 8279
rect 5261 8239 5319 8245
rect 5810 8236 5816 8288
rect 5868 8276 5874 8288
rect 6365 8279 6423 8285
rect 6365 8276 6377 8279
rect 5868 8248 6377 8276
rect 5868 8236 5874 8248
rect 6365 8245 6377 8248
rect 6411 8245 6423 8279
rect 6822 8276 6828 8288
rect 6783 8248 6828 8276
rect 6365 8239 6423 8245
rect 6822 8236 6828 8248
rect 6880 8236 6886 8288
rect 7742 8236 7748 8288
rect 7800 8276 7806 8288
rect 7944 8276 7972 8375
rect 8202 8304 8208 8356
rect 8260 8344 8266 8356
rect 8481 8347 8539 8353
rect 8481 8344 8493 8347
rect 8260 8316 8493 8344
rect 8260 8304 8266 8316
rect 8481 8313 8493 8316
rect 8527 8313 8539 8347
rect 8588 8344 8616 8384
rect 8662 8372 8668 8424
rect 8720 8412 8726 8424
rect 9033 8415 9091 8421
rect 9033 8412 9045 8415
rect 8720 8384 9045 8412
rect 8720 8372 8726 8384
rect 9033 8381 9045 8384
rect 9079 8412 9091 8415
rect 9122 8412 9128 8424
rect 9079 8384 9128 8412
rect 9079 8381 9091 8384
rect 9033 8375 9091 8381
rect 9122 8372 9128 8384
rect 9180 8372 9186 8424
rect 9217 8415 9275 8421
rect 9217 8381 9229 8415
rect 9263 8412 9275 8415
rect 9766 8412 9772 8424
rect 9263 8384 9772 8412
rect 9263 8381 9275 8384
rect 9217 8375 9275 8381
rect 9232 8344 9260 8375
rect 9766 8372 9772 8384
rect 9824 8372 9830 8424
rect 9858 8372 9864 8424
rect 9916 8412 9922 8424
rect 11054 8412 11060 8424
rect 9916 8384 9961 8412
rect 11015 8384 11060 8412
rect 9916 8372 9922 8384
rect 11054 8372 11060 8384
rect 11112 8372 11118 8424
rect 14458 8412 14464 8424
rect 12452 8384 14464 8412
rect 8588 8316 9260 8344
rect 8481 8307 8539 8313
rect 8570 8276 8576 8288
rect 7800 8248 7972 8276
rect 8531 8248 8576 8276
rect 7800 8236 7806 8248
rect 8570 8236 8576 8248
rect 8628 8236 8634 8288
rect 9858 8236 9864 8288
rect 9916 8276 9922 8288
rect 10318 8276 10324 8288
rect 9916 8248 10324 8276
rect 9916 8236 9922 8248
rect 10318 8236 10324 8248
rect 10376 8236 10382 8288
rect 10413 8279 10471 8285
rect 10413 8245 10425 8279
rect 10459 8276 10471 8279
rect 12452 8276 12480 8384
rect 14458 8372 14464 8384
rect 14516 8372 14522 8424
rect 19337 8415 19395 8421
rect 19337 8381 19349 8415
rect 19383 8412 19395 8415
rect 19429 8415 19487 8421
rect 19429 8412 19441 8415
rect 19383 8384 19441 8412
rect 19383 8381 19395 8384
rect 19337 8375 19395 8381
rect 19429 8381 19441 8384
rect 19475 8381 19487 8415
rect 19429 8375 19487 8381
rect 13262 8304 13268 8356
rect 13320 8344 13326 8356
rect 14277 8347 14335 8353
rect 14277 8344 14289 8347
rect 13320 8316 14289 8344
rect 13320 8304 13326 8316
rect 14277 8313 14289 8316
rect 14323 8313 14335 8347
rect 14277 8307 14335 8313
rect 18138 8304 18144 8356
rect 18196 8304 18202 8356
rect 10459 8248 12480 8276
rect 10459 8245 10471 8248
rect 10413 8239 10471 8245
rect 12526 8236 12532 8288
rect 12584 8276 12590 8288
rect 12802 8276 12808 8288
rect 12584 8248 12808 8276
rect 12584 8236 12590 8248
rect 12802 8236 12808 8248
rect 12860 8236 12866 8288
rect 13446 8236 13452 8288
rect 13504 8276 13510 8288
rect 13722 8276 13728 8288
rect 13504 8248 13728 8276
rect 13504 8236 13510 8248
rect 13722 8236 13728 8248
rect 13780 8276 13786 8288
rect 16482 8276 16488 8288
rect 13780 8248 16488 8276
rect 13780 8236 13786 8248
rect 16482 8236 16488 8248
rect 16540 8236 16546 8288
rect 17402 8236 17408 8288
rect 17460 8276 17466 8288
rect 17957 8279 18015 8285
rect 17957 8276 17969 8279
rect 17460 8248 17969 8276
rect 17460 8236 17466 8248
rect 17957 8245 17969 8248
rect 18003 8276 18015 8279
rect 18156 8276 18184 8304
rect 18003 8248 18184 8276
rect 19444 8276 19472 8375
rect 20993 8279 21051 8285
rect 20993 8276 21005 8279
rect 19444 8248 21005 8276
rect 18003 8245 18015 8248
rect 17957 8239 18015 8245
rect 20993 8245 21005 8248
rect 21039 8276 21051 8279
rect 21266 8276 21272 8288
rect 21039 8248 21272 8276
rect 21039 8245 21051 8248
rect 20993 8239 21051 8245
rect 21266 8236 21272 8248
rect 21324 8236 21330 8288
rect 1104 8186 21896 8208
rect 1104 8134 3549 8186
rect 3601 8134 3613 8186
rect 3665 8134 3677 8186
rect 3729 8134 3741 8186
rect 3793 8134 3805 8186
rect 3857 8134 8747 8186
rect 8799 8134 8811 8186
rect 8863 8134 8875 8186
rect 8927 8134 8939 8186
rect 8991 8134 9003 8186
rect 9055 8134 13945 8186
rect 13997 8134 14009 8186
rect 14061 8134 14073 8186
rect 14125 8134 14137 8186
rect 14189 8134 14201 8186
rect 14253 8134 19143 8186
rect 19195 8134 19207 8186
rect 19259 8134 19271 8186
rect 19323 8134 19335 8186
rect 19387 8134 19399 8186
rect 19451 8134 21896 8186
rect 1104 8112 21896 8134
rect 1486 8072 1492 8084
rect 1447 8044 1492 8072
rect 1486 8032 1492 8044
rect 1544 8032 1550 8084
rect 2774 8032 2780 8084
rect 2832 8072 2838 8084
rect 3237 8075 3295 8081
rect 3237 8072 3249 8075
rect 2832 8044 3249 8072
rect 2832 8032 2838 8044
rect 3237 8041 3249 8044
rect 3283 8072 3295 8075
rect 3878 8072 3884 8084
rect 3283 8044 3884 8072
rect 3283 8041 3295 8044
rect 3237 8035 3295 8041
rect 3878 8032 3884 8044
rect 3936 8032 3942 8084
rect 4982 8032 4988 8084
rect 5040 8072 5046 8084
rect 5626 8072 5632 8084
rect 5040 8044 5632 8072
rect 5040 8032 5046 8044
rect 5626 8032 5632 8044
rect 5684 8032 5690 8084
rect 5718 8032 5724 8084
rect 5776 8072 5782 8084
rect 6457 8075 6515 8081
rect 6457 8072 6469 8075
rect 5776 8044 6469 8072
rect 5776 8032 5782 8044
rect 6457 8041 6469 8044
rect 6503 8041 6515 8075
rect 6457 8035 6515 8041
rect 7466 8032 7472 8084
rect 7524 8072 7530 8084
rect 7837 8075 7895 8081
rect 7837 8072 7849 8075
rect 7524 8044 7849 8072
rect 7524 8032 7530 8044
rect 7837 8041 7849 8044
rect 7883 8041 7895 8075
rect 7837 8035 7895 8041
rect 8202 8032 8208 8084
rect 8260 8072 8266 8084
rect 12618 8072 12624 8084
rect 8260 8044 12624 8072
rect 8260 8032 8266 8044
rect 12618 8032 12624 8044
rect 12676 8032 12682 8084
rect 13722 8032 13728 8084
rect 13780 8072 13786 8084
rect 14369 8075 14427 8081
rect 14369 8072 14381 8075
rect 13780 8044 14381 8072
rect 13780 8032 13786 8044
rect 14369 8041 14381 8044
rect 14415 8041 14427 8075
rect 14369 8035 14427 8041
rect 14829 8075 14887 8081
rect 14829 8041 14841 8075
rect 14875 8072 14887 8075
rect 15102 8072 15108 8084
rect 14875 8044 15108 8072
rect 14875 8041 14887 8044
rect 14829 8035 14887 8041
rect 15102 8032 15108 8044
rect 15160 8072 15166 8084
rect 15470 8072 15476 8084
rect 15160 8044 15476 8072
rect 15160 8032 15166 8044
rect 15470 8032 15476 8044
rect 15528 8032 15534 8084
rect 15749 8075 15807 8081
rect 15749 8041 15761 8075
rect 15795 8072 15807 8075
rect 16390 8072 16396 8084
rect 15795 8044 16396 8072
rect 15795 8041 15807 8044
rect 15749 8035 15807 8041
rect 16390 8032 16396 8044
rect 16448 8032 16454 8084
rect 16482 8032 16488 8084
rect 16540 8072 16546 8084
rect 19889 8075 19947 8081
rect 19889 8072 19901 8075
rect 16540 8044 19901 8072
rect 16540 8032 16546 8044
rect 19889 8041 19901 8044
rect 19935 8041 19947 8075
rect 21542 8072 21548 8084
rect 19889 8035 19947 8041
rect 19996 8044 21548 8072
rect 3050 7964 3056 8016
rect 3108 8004 3114 8016
rect 11885 8007 11943 8013
rect 11885 8004 11897 8007
rect 3108 7976 5580 8004
rect 3108 7964 3114 7976
rect 1949 7939 2007 7945
rect 1949 7905 1961 7939
rect 1995 7905 2007 7939
rect 1949 7899 2007 7905
rect 1964 7800 1992 7899
rect 2038 7896 2044 7948
rect 2096 7936 2102 7948
rect 2866 7936 2872 7948
rect 2096 7908 2141 7936
rect 2827 7908 2872 7936
rect 2096 7896 2102 7908
rect 2866 7896 2872 7908
rect 2924 7896 2930 7948
rect 4893 7939 4951 7945
rect 4893 7905 4905 7939
rect 4939 7936 4951 7939
rect 5074 7936 5080 7948
rect 4939 7908 5080 7936
rect 4939 7905 4951 7908
rect 4893 7899 4951 7905
rect 5074 7896 5080 7908
rect 5132 7896 5138 7948
rect 5552 7945 5580 7976
rect 5828 7976 11897 8004
rect 5537 7939 5595 7945
rect 5537 7905 5549 7939
rect 5583 7905 5595 7939
rect 5537 7899 5595 7905
rect 3050 7868 3056 7880
rect 3011 7840 3056 7868
rect 3050 7828 3056 7840
rect 3108 7828 3114 7880
rect 3970 7828 3976 7880
rect 4028 7868 4034 7880
rect 5828 7877 5856 7976
rect 11885 7973 11897 7976
rect 11931 7973 11943 8007
rect 11885 7967 11943 7973
rect 14550 7964 14556 8016
rect 14608 8004 14614 8016
rect 17865 8007 17923 8013
rect 17865 8004 17877 8007
rect 14608 7976 17877 8004
rect 14608 7964 14614 7976
rect 17865 7973 17877 7976
rect 17911 7973 17923 8007
rect 19518 8004 19524 8016
rect 17865 7967 17923 7973
rect 18340 7976 19524 8004
rect 7098 7896 7104 7948
rect 7156 7936 7162 7948
rect 7156 7908 7201 7936
rect 7156 7896 7162 7908
rect 8110 7896 8116 7948
rect 8168 7936 8174 7948
rect 8389 7939 8447 7945
rect 8389 7936 8401 7939
rect 8168 7908 8401 7936
rect 8168 7896 8174 7908
rect 8389 7905 8401 7908
rect 8435 7905 8447 7939
rect 8389 7899 8447 7905
rect 9309 7939 9367 7945
rect 9309 7905 9321 7939
rect 9355 7936 9367 7939
rect 10870 7936 10876 7948
rect 9355 7908 10876 7936
rect 9355 7905 9367 7908
rect 9309 7899 9367 7905
rect 10870 7896 10876 7908
rect 10928 7896 10934 7948
rect 11241 7939 11299 7945
rect 11241 7905 11253 7939
rect 11287 7936 11299 7939
rect 11330 7936 11336 7948
rect 11287 7908 11336 7936
rect 11287 7905 11299 7908
rect 11241 7899 11299 7905
rect 11330 7896 11336 7908
rect 11388 7896 11394 7948
rect 12526 7936 12532 7948
rect 12487 7908 12532 7936
rect 12526 7896 12532 7908
rect 12584 7896 12590 7948
rect 12986 7896 12992 7948
rect 13044 7936 13050 7948
rect 15194 7936 15200 7948
rect 13044 7908 15200 7936
rect 13044 7896 13050 7908
rect 15194 7896 15200 7908
rect 15252 7896 15258 7948
rect 16669 7939 16727 7945
rect 16669 7905 16681 7939
rect 16715 7936 16727 7939
rect 18340 7936 18368 7976
rect 19518 7964 19524 7976
rect 19576 7964 19582 8016
rect 16715 7908 18368 7936
rect 18509 7939 18567 7945
rect 16715 7905 16727 7908
rect 16669 7899 16727 7905
rect 18509 7905 18521 7939
rect 18555 7936 18567 7939
rect 19996 7936 20024 8044
rect 21542 8032 21548 8044
rect 21600 8032 21606 8084
rect 18555 7908 20024 7936
rect 18555 7905 18567 7908
rect 18509 7899 18567 7905
rect 21266 7896 21272 7948
rect 21324 7936 21330 7948
rect 21361 7939 21419 7945
rect 21361 7936 21373 7939
rect 21324 7908 21373 7936
rect 21324 7896 21330 7908
rect 21361 7905 21373 7908
rect 21407 7905 21419 7939
rect 21361 7899 21419 7905
rect 5813 7871 5871 7877
rect 4028 7840 5580 7868
rect 4028 7828 4034 7840
rect 3329 7803 3387 7809
rect 3329 7800 3341 7803
rect 1964 7772 3341 7800
rect 3329 7769 3341 7772
rect 3375 7800 3387 7803
rect 4614 7800 4620 7812
rect 3375 7772 4620 7800
rect 3375 7769 3387 7772
rect 3329 7763 3387 7769
rect 4614 7760 4620 7772
rect 4672 7760 4678 7812
rect 4706 7760 4712 7812
rect 4764 7800 4770 7812
rect 5169 7803 5227 7809
rect 5169 7800 5181 7803
rect 4764 7772 5181 7800
rect 4764 7760 4770 7772
rect 5169 7769 5181 7772
rect 5215 7800 5227 7803
rect 5258 7800 5264 7812
rect 5215 7772 5264 7800
rect 5215 7769 5227 7772
rect 5169 7763 5227 7769
rect 5258 7760 5264 7772
rect 5316 7760 5322 7812
rect 5552 7800 5580 7840
rect 5813 7837 5825 7871
rect 5859 7837 5871 7871
rect 6362 7868 6368 7880
rect 6323 7840 6368 7868
rect 5813 7831 5871 7837
rect 6362 7828 6368 7840
rect 6420 7828 6426 7880
rect 6914 7868 6920 7880
rect 6875 7840 6920 7868
rect 6914 7828 6920 7840
rect 6972 7828 6978 7880
rect 9401 7871 9459 7877
rect 9401 7837 9413 7871
rect 9447 7868 9459 7871
rect 15102 7868 15108 7880
rect 9447 7840 15108 7868
rect 9447 7837 9459 7840
rect 9401 7831 9459 7837
rect 15102 7828 15108 7840
rect 15160 7828 15166 7880
rect 15746 7828 15752 7880
rect 15804 7868 15810 7880
rect 16393 7871 16451 7877
rect 16393 7868 16405 7871
rect 15804 7840 16405 7868
rect 15804 7828 15810 7840
rect 16393 7837 16405 7840
rect 16439 7837 16451 7871
rect 18325 7871 18383 7877
rect 18325 7868 18337 7871
rect 16393 7831 16451 7837
rect 17512 7840 18337 7868
rect 6089 7803 6147 7809
rect 6089 7800 6101 7803
rect 5552 7772 6101 7800
rect 6089 7769 6101 7772
rect 6135 7769 6147 7803
rect 7834 7800 7840 7812
rect 6089 7763 6147 7769
rect 6748 7772 7840 7800
rect 1762 7692 1768 7744
rect 1820 7732 1826 7744
rect 2133 7735 2191 7741
rect 2133 7732 2145 7735
rect 1820 7704 2145 7732
rect 1820 7692 1826 7704
rect 2133 7701 2145 7704
rect 2179 7701 2191 7735
rect 2498 7732 2504 7744
rect 2459 7704 2504 7732
rect 2133 7695 2191 7701
rect 2498 7692 2504 7704
rect 2556 7692 2562 7744
rect 4982 7732 4988 7744
rect 4943 7704 4988 7732
rect 4982 7692 4988 7704
rect 5040 7692 5046 7744
rect 5074 7692 5080 7744
rect 5132 7732 5138 7744
rect 6748 7732 6776 7772
rect 7834 7760 7840 7772
rect 7892 7760 7898 7812
rect 8205 7803 8263 7809
rect 8205 7769 8217 7803
rect 8251 7800 8263 7803
rect 9306 7800 9312 7812
rect 8251 7772 9312 7800
rect 8251 7769 8263 7772
rect 8205 7763 8263 7769
rect 9306 7760 9312 7772
rect 9364 7760 9370 7812
rect 9493 7803 9551 7809
rect 9493 7800 9505 7803
rect 9416 7772 9505 7800
rect 9416 7744 9444 7772
rect 9493 7769 9505 7772
rect 9539 7800 9551 7803
rect 9953 7803 10011 7809
rect 9953 7800 9965 7803
rect 9539 7772 9965 7800
rect 9539 7769 9551 7772
rect 9493 7763 9551 7769
rect 9953 7769 9965 7772
rect 9999 7769 10011 7803
rect 10410 7800 10416 7812
rect 10371 7772 10416 7800
rect 9953 7763 10011 7769
rect 10410 7760 10416 7772
rect 10468 7760 10474 7812
rect 10502 7760 10508 7812
rect 10560 7800 10566 7812
rect 10689 7803 10747 7809
rect 10689 7800 10701 7803
rect 10560 7772 10701 7800
rect 10560 7760 10566 7772
rect 10689 7769 10701 7772
rect 10735 7769 10747 7803
rect 10962 7800 10968 7812
rect 10923 7772 10968 7800
rect 10689 7763 10747 7769
rect 5132 7704 6776 7732
rect 5132 7692 5138 7704
rect 6822 7692 6828 7744
rect 6880 7732 6886 7744
rect 6880 7704 6925 7732
rect 6880 7692 6886 7704
rect 7098 7692 7104 7744
rect 7156 7732 7162 7744
rect 7285 7735 7343 7741
rect 7285 7732 7297 7735
rect 7156 7704 7297 7732
rect 7156 7692 7162 7704
rect 7285 7701 7297 7704
rect 7331 7701 7343 7735
rect 7558 7732 7564 7744
rect 7519 7704 7564 7732
rect 7285 7695 7343 7701
rect 7558 7692 7564 7704
rect 7616 7692 7622 7744
rect 8297 7735 8355 7741
rect 8297 7701 8309 7735
rect 8343 7732 8355 7735
rect 8386 7732 8392 7744
rect 8343 7704 8392 7732
rect 8343 7701 8355 7704
rect 8297 7695 8355 7701
rect 8386 7692 8392 7704
rect 8444 7692 8450 7744
rect 8570 7692 8576 7744
rect 8628 7732 8634 7744
rect 8665 7735 8723 7741
rect 8665 7732 8677 7735
rect 8628 7704 8677 7732
rect 8628 7692 8634 7704
rect 8665 7701 8677 7704
rect 8711 7701 8723 7735
rect 8665 7695 8723 7701
rect 9398 7692 9404 7744
rect 9456 7692 9462 7744
rect 9582 7692 9588 7744
rect 9640 7732 9646 7744
rect 9861 7735 9919 7741
rect 9861 7732 9873 7735
rect 9640 7704 9873 7732
rect 9640 7692 9646 7704
rect 9861 7701 9873 7704
rect 9907 7701 9919 7735
rect 10704 7732 10732 7763
rect 10962 7760 10968 7772
rect 11020 7800 11026 7812
rect 11425 7803 11483 7809
rect 11425 7800 11437 7803
rect 11020 7772 11437 7800
rect 11020 7760 11026 7772
rect 11425 7769 11437 7772
rect 11471 7769 11483 7803
rect 14182 7800 14188 7812
rect 11425 7763 11483 7769
rect 11808 7772 14188 7800
rect 11808 7741 11836 7772
rect 14182 7760 14188 7772
rect 14240 7760 14246 7812
rect 14366 7760 14372 7812
rect 14424 7800 14430 7812
rect 14424 7772 16068 7800
rect 14424 7760 14430 7772
rect 11333 7735 11391 7741
rect 11333 7732 11345 7735
rect 10704 7704 11345 7732
rect 9861 7695 9919 7701
rect 11333 7701 11345 7704
rect 11379 7701 11391 7735
rect 11333 7695 11391 7701
rect 11793 7735 11851 7741
rect 11793 7701 11805 7735
rect 11839 7701 11851 7735
rect 11793 7695 11851 7701
rect 12066 7692 12072 7744
rect 12124 7732 12130 7744
rect 12253 7735 12311 7741
rect 12253 7732 12265 7735
rect 12124 7704 12265 7732
rect 12124 7692 12130 7704
rect 12253 7701 12265 7704
rect 12299 7701 12311 7735
rect 12253 7695 12311 7701
rect 12345 7735 12403 7741
rect 12345 7701 12357 7735
rect 12391 7732 12403 7735
rect 12434 7732 12440 7744
rect 12391 7704 12440 7732
rect 12391 7701 12403 7704
rect 12345 7695 12403 7701
rect 12434 7692 12440 7704
rect 12492 7692 12498 7744
rect 14274 7732 14280 7744
rect 14235 7704 14280 7732
rect 14274 7692 14280 7704
rect 14332 7692 14338 7744
rect 15746 7692 15752 7744
rect 15804 7732 15810 7744
rect 16040 7741 16068 7772
rect 15841 7735 15899 7741
rect 15841 7732 15853 7735
rect 15804 7704 15853 7732
rect 15804 7692 15810 7704
rect 15841 7701 15853 7704
rect 15887 7701 15899 7735
rect 15841 7695 15899 7701
rect 16025 7735 16083 7741
rect 16025 7701 16037 7735
rect 16071 7701 16083 7735
rect 16025 7695 16083 7701
rect 16390 7692 16396 7744
rect 16448 7732 16454 7744
rect 16485 7735 16543 7741
rect 16485 7732 16497 7735
rect 16448 7704 16497 7732
rect 16448 7692 16454 7704
rect 16485 7701 16497 7704
rect 16531 7701 16543 7735
rect 16485 7695 16543 7701
rect 17218 7692 17224 7744
rect 17276 7732 17282 7744
rect 17512 7741 17540 7840
rect 18325 7837 18337 7840
rect 18371 7837 18383 7871
rect 18325 7831 18383 7837
rect 19521 7871 19579 7877
rect 19521 7837 19533 7871
rect 19567 7868 19579 7871
rect 21284 7868 21312 7896
rect 19567 7840 21312 7868
rect 19567 7837 19579 7840
rect 19521 7831 19579 7837
rect 17586 7760 17592 7812
rect 17644 7800 17650 7812
rect 21002 7803 21060 7809
rect 21002 7800 21014 7803
rect 17644 7772 21014 7800
rect 17644 7760 17650 7772
rect 21002 7769 21014 7772
rect 21048 7769 21060 7803
rect 21002 7763 21060 7769
rect 17497 7735 17555 7741
rect 17497 7732 17509 7735
rect 17276 7704 17509 7732
rect 17276 7692 17282 7704
rect 17497 7701 17509 7704
rect 17543 7701 17555 7735
rect 17678 7732 17684 7744
rect 17639 7704 17684 7732
rect 17497 7695 17555 7701
rect 17678 7692 17684 7704
rect 17736 7732 17742 7744
rect 18233 7735 18291 7741
rect 18233 7732 18245 7735
rect 17736 7704 18245 7732
rect 17736 7692 17742 7704
rect 18233 7701 18245 7704
rect 18279 7701 18291 7735
rect 18233 7695 18291 7701
rect 1104 7642 22056 7664
rect 1104 7590 6148 7642
rect 6200 7590 6212 7642
rect 6264 7590 6276 7642
rect 6328 7590 6340 7642
rect 6392 7590 6404 7642
rect 6456 7590 11346 7642
rect 11398 7590 11410 7642
rect 11462 7590 11474 7642
rect 11526 7590 11538 7642
rect 11590 7590 11602 7642
rect 11654 7590 16544 7642
rect 16596 7590 16608 7642
rect 16660 7590 16672 7642
rect 16724 7590 16736 7642
rect 16788 7590 16800 7642
rect 16852 7590 21742 7642
rect 21794 7590 21806 7642
rect 21858 7590 21870 7642
rect 21922 7590 21934 7642
rect 21986 7590 21998 7642
rect 22050 7590 22056 7642
rect 1104 7568 22056 7590
rect 1673 7531 1731 7537
rect 1673 7497 1685 7531
rect 1719 7528 1731 7531
rect 2038 7528 2044 7540
rect 1719 7500 2044 7528
rect 1719 7497 1731 7500
rect 1673 7491 1731 7497
rect 2038 7488 2044 7500
rect 2096 7488 2102 7540
rect 4246 7528 4252 7540
rect 4207 7500 4252 7528
rect 4246 7488 4252 7500
rect 4304 7528 4310 7540
rect 4893 7531 4951 7537
rect 4893 7528 4905 7531
rect 4304 7500 4905 7528
rect 4304 7488 4310 7500
rect 4893 7497 4905 7500
rect 4939 7528 4951 7531
rect 4982 7528 4988 7540
rect 4939 7500 4988 7528
rect 4939 7497 4951 7500
rect 4893 7491 4951 7497
rect 4982 7488 4988 7500
rect 5040 7488 5046 7540
rect 6181 7531 6239 7537
rect 6181 7497 6193 7531
rect 6227 7528 6239 7531
rect 6638 7528 6644 7540
rect 6227 7500 6644 7528
rect 6227 7497 6239 7500
rect 6181 7491 6239 7497
rect 6638 7488 6644 7500
rect 6696 7488 6702 7540
rect 7282 7488 7288 7540
rect 7340 7528 7346 7540
rect 7561 7531 7619 7537
rect 7561 7528 7573 7531
rect 7340 7500 7573 7528
rect 7340 7488 7346 7500
rect 7561 7497 7573 7500
rect 7607 7497 7619 7531
rect 7561 7491 7619 7497
rect 9125 7531 9183 7537
rect 9125 7497 9137 7531
rect 9171 7497 9183 7531
rect 9582 7528 9588 7540
rect 9543 7500 9588 7528
rect 9125 7491 9183 7497
rect 1489 7463 1547 7469
rect 1489 7429 1501 7463
rect 1535 7460 1547 7463
rect 1762 7460 1768 7472
rect 1535 7432 1768 7460
rect 1535 7429 1547 7432
rect 1489 7423 1547 7429
rect 1762 7420 1768 7432
rect 1820 7420 1826 7472
rect 3050 7420 3056 7472
rect 3108 7460 3114 7472
rect 9140 7460 9168 7491
rect 9582 7488 9588 7500
rect 9640 7488 9646 7540
rect 10505 7531 10563 7537
rect 10505 7497 10517 7531
rect 10551 7497 10563 7531
rect 12066 7528 12072 7540
rect 12027 7500 12072 7528
rect 10505 7491 10563 7497
rect 3108 7432 9168 7460
rect 9493 7463 9551 7469
rect 3108 7420 3114 7432
rect 9493 7429 9505 7463
rect 9539 7460 9551 7463
rect 10520 7460 10548 7491
rect 12066 7488 12072 7500
rect 12124 7488 12130 7540
rect 13449 7531 13507 7537
rect 13449 7528 13461 7531
rect 12406 7500 13461 7528
rect 9539 7432 10548 7460
rect 9539 7429 9551 7432
rect 9493 7423 9551 7429
rect 10594 7420 10600 7472
rect 10652 7460 10658 7472
rect 12406 7460 12434 7500
rect 13449 7497 13461 7500
rect 13495 7497 13507 7531
rect 13449 7491 13507 7497
rect 14274 7488 14280 7540
rect 14332 7528 14338 7540
rect 14645 7531 14703 7537
rect 14645 7528 14657 7531
rect 14332 7500 14657 7528
rect 14332 7488 14338 7500
rect 14645 7497 14657 7500
rect 14691 7497 14703 7531
rect 15102 7528 15108 7540
rect 15063 7500 15108 7528
rect 14645 7491 14703 7497
rect 15102 7488 15108 7500
rect 15160 7488 15166 7540
rect 15470 7488 15476 7540
rect 15528 7528 15534 7540
rect 15565 7531 15623 7537
rect 15565 7528 15577 7531
rect 15528 7500 15577 7528
rect 15528 7488 15534 7500
rect 15565 7497 15577 7500
rect 15611 7497 15623 7531
rect 15565 7491 15623 7497
rect 10652 7432 12434 7460
rect 10652 7420 10658 7432
rect 13722 7420 13728 7472
rect 13780 7460 13786 7472
rect 14737 7463 14795 7469
rect 14737 7460 14749 7463
rect 13780 7432 14749 7460
rect 13780 7420 13786 7432
rect 14737 7429 14749 7432
rect 14783 7429 14795 7463
rect 15580 7460 15608 7491
rect 17770 7488 17776 7540
rect 17828 7528 17834 7540
rect 19337 7531 19395 7537
rect 19337 7528 19349 7531
rect 17828 7500 19349 7528
rect 17828 7488 17834 7500
rect 19337 7497 19349 7500
rect 19383 7497 19395 7531
rect 19337 7491 19395 7497
rect 20901 7531 20959 7537
rect 20901 7497 20913 7531
rect 20947 7528 20959 7531
rect 21266 7528 21272 7540
rect 20947 7500 21272 7528
rect 20947 7497 20959 7500
rect 20901 7491 20959 7497
rect 17862 7460 17868 7472
rect 15580 7432 17868 7460
rect 14737 7423 14795 7429
rect 17862 7420 17868 7432
rect 17920 7420 17926 7472
rect 20806 7460 20812 7472
rect 20640 7432 20812 7460
rect 4522 7392 4528 7404
rect 4483 7364 4528 7392
rect 4522 7352 4528 7364
rect 4580 7392 4586 7404
rect 4985 7395 5043 7401
rect 4985 7392 4997 7395
rect 4580 7364 4997 7392
rect 4580 7352 4586 7364
rect 4985 7361 4997 7364
rect 5031 7361 5043 7395
rect 5810 7392 5816 7404
rect 5771 7364 5816 7392
rect 4985 7355 5043 7361
rect 5810 7352 5816 7364
rect 5868 7352 5874 7404
rect 6825 7395 6883 7401
rect 6825 7361 6837 7395
rect 6871 7392 6883 7395
rect 7285 7395 7343 7401
rect 7285 7392 7297 7395
rect 6871 7364 7297 7392
rect 6871 7361 6883 7364
rect 6825 7355 6883 7361
rect 7285 7361 7297 7364
rect 7331 7361 7343 7395
rect 7926 7392 7932 7404
rect 7887 7364 7932 7392
rect 7285 7355 7343 7361
rect 7926 7352 7932 7364
rect 7984 7352 7990 7404
rect 8021 7395 8079 7401
rect 8021 7361 8033 7395
rect 8067 7392 8079 7395
rect 8662 7392 8668 7404
rect 8067 7364 8668 7392
rect 8067 7361 8079 7364
rect 8021 7355 8079 7361
rect 8662 7352 8668 7364
rect 8720 7352 8726 7404
rect 10873 7395 10931 7401
rect 10873 7361 10885 7395
rect 10919 7392 10931 7395
rect 11517 7395 11575 7401
rect 11517 7392 11529 7395
rect 10919 7364 11529 7392
rect 10919 7361 10931 7364
rect 10873 7355 10931 7361
rect 11517 7361 11529 7364
rect 11563 7361 11575 7395
rect 11517 7355 11575 7361
rect 12437 7395 12495 7401
rect 12437 7361 12449 7395
rect 12483 7392 12495 7395
rect 12897 7395 12955 7401
rect 12897 7392 12909 7395
rect 12483 7364 12909 7392
rect 12483 7361 12495 7364
rect 12437 7355 12495 7361
rect 12897 7361 12909 7364
rect 12943 7361 12955 7395
rect 12897 7355 12955 7361
rect 13817 7395 13875 7401
rect 13817 7361 13829 7395
rect 13863 7392 13875 7395
rect 15470 7392 15476 7404
rect 13863 7364 14320 7392
rect 15431 7364 15476 7392
rect 13863 7361 13875 7364
rect 13817 7355 13875 7361
rect 4801 7327 4859 7333
rect 4801 7293 4813 7327
rect 4847 7324 4859 7327
rect 5166 7324 5172 7336
rect 4847 7296 5172 7324
rect 4847 7293 4859 7296
rect 4801 7287 4859 7293
rect 5166 7284 5172 7296
rect 5224 7284 5230 7336
rect 5442 7284 5448 7336
rect 5500 7324 5506 7336
rect 5537 7327 5595 7333
rect 5537 7324 5549 7327
rect 5500 7296 5549 7324
rect 5500 7284 5506 7296
rect 5537 7293 5549 7296
rect 5583 7293 5595 7327
rect 5537 7287 5595 7293
rect 5721 7327 5779 7333
rect 5721 7293 5733 7327
rect 5767 7324 5779 7327
rect 5902 7324 5908 7336
rect 5767 7296 5908 7324
rect 5767 7293 5779 7296
rect 5721 7287 5779 7293
rect 5902 7284 5908 7296
rect 5960 7284 5966 7336
rect 6086 7284 6092 7336
rect 6144 7324 6150 7336
rect 6917 7327 6975 7333
rect 6917 7324 6929 7327
rect 6144 7296 6929 7324
rect 6144 7284 6150 7296
rect 6917 7293 6929 7296
rect 6963 7293 6975 7327
rect 7098 7324 7104 7336
rect 7059 7296 7104 7324
rect 6917 7287 6975 7293
rect 3970 7216 3976 7268
rect 4028 7256 4034 7268
rect 4028 7228 5948 7256
rect 4028 7216 4034 7228
rect 5353 7191 5411 7197
rect 5353 7157 5365 7191
rect 5399 7188 5411 7191
rect 5442 7188 5448 7200
rect 5399 7160 5448 7188
rect 5399 7157 5411 7160
rect 5353 7151 5411 7157
rect 5442 7148 5448 7160
rect 5500 7148 5506 7200
rect 5920 7188 5948 7228
rect 5994 7216 6000 7268
rect 6052 7256 6058 7268
rect 6457 7259 6515 7265
rect 6457 7256 6469 7259
rect 6052 7228 6469 7256
rect 6052 7216 6058 7228
rect 6457 7225 6469 7228
rect 6503 7225 6515 7259
rect 6932 7256 6960 7287
rect 7098 7284 7104 7296
rect 7156 7284 7162 7336
rect 8202 7324 8208 7336
rect 8163 7296 8208 7324
rect 8202 7284 8208 7296
rect 8260 7284 8266 7336
rect 9582 7284 9588 7336
rect 9640 7324 9646 7336
rect 9677 7327 9735 7333
rect 9677 7324 9689 7327
rect 9640 7296 9689 7324
rect 9640 7284 9646 7296
rect 9677 7293 9689 7296
rect 9723 7293 9735 7327
rect 10965 7327 11023 7333
rect 10965 7324 10977 7327
rect 9677 7287 9735 7293
rect 10336 7296 10977 7324
rect 7558 7256 7564 7268
rect 6932 7228 7564 7256
rect 6457 7219 6515 7225
rect 7558 7216 7564 7228
rect 7616 7216 7622 7268
rect 10336 7200 10364 7296
rect 10965 7293 10977 7296
rect 11011 7293 11023 7327
rect 10965 7287 11023 7293
rect 11057 7327 11115 7333
rect 11057 7293 11069 7327
rect 11103 7293 11115 7327
rect 12529 7327 12587 7333
rect 12529 7324 12541 7327
rect 11057 7287 11115 7293
rect 11900 7296 12541 7324
rect 10870 7216 10876 7268
rect 10928 7256 10934 7268
rect 11072 7256 11100 7287
rect 10928 7228 11100 7256
rect 10928 7216 10934 7228
rect 7190 7188 7196 7200
rect 5920 7160 7196 7188
rect 7190 7148 7196 7160
rect 7248 7148 7254 7200
rect 9858 7148 9864 7200
rect 9916 7188 9922 7200
rect 9953 7191 10011 7197
rect 9953 7188 9965 7191
rect 9916 7160 9965 7188
rect 9916 7148 9922 7160
rect 9953 7157 9965 7160
rect 9999 7157 10011 7191
rect 10318 7188 10324 7200
rect 10279 7160 10324 7188
rect 9953 7151 10011 7157
rect 10318 7148 10324 7160
rect 10376 7148 10382 7200
rect 11054 7148 11060 7200
rect 11112 7188 11118 7200
rect 11900 7197 11928 7296
rect 12529 7293 12541 7296
rect 12575 7293 12587 7327
rect 12529 7287 12587 7293
rect 12713 7327 12771 7333
rect 12713 7293 12725 7327
rect 12759 7324 12771 7327
rect 12986 7324 12992 7336
rect 12759 7296 12992 7324
rect 12759 7293 12771 7296
rect 12713 7287 12771 7293
rect 12986 7284 12992 7296
rect 13044 7284 13050 7336
rect 13909 7327 13967 7333
rect 13909 7324 13921 7327
rect 13832 7296 13921 7324
rect 13832 7268 13860 7296
rect 13909 7293 13921 7296
rect 13955 7293 13967 7327
rect 13909 7287 13967 7293
rect 14093 7327 14151 7333
rect 14093 7293 14105 7327
rect 14139 7293 14151 7327
rect 14093 7287 14151 7293
rect 12250 7216 12256 7268
rect 12308 7256 12314 7268
rect 12894 7256 12900 7268
rect 12308 7228 12900 7256
rect 12308 7216 12314 7228
rect 12894 7216 12900 7228
rect 12952 7216 12958 7268
rect 13814 7216 13820 7268
rect 13872 7216 13878 7268
rect 11885 7191 11943 7197
rect 11885 7188 11897 7191
rect 11112 7160 11897 7188
rect 11112 7148 11118 7160
rect 11885 7157 11897 7160
rect 11931 7157 11943 7191
rect 14108 7188 14136 7287
rect 14292 7265 14320 7364
rect 15470 7352 15476 7364
rect 15528 7352 15534 7404
rect 20450 7395 20508 7401
rect 20450 7392 20462 7395
rect 15764 7364 20462 7392
rect 14921 7327 14979 7333
rect 14921 7293 14933 7327
rect 14967 7324 14979 7327
rect 15010 7324 15016 7336
rect 14967 7296 15016 7324
rect 14967 7293 14979 7296
rect 14921 7287 14979 7293
rect 15010 7284 15016 7296
rect 15068 7284 15074 7336
rect 15764 7333 15792 7364
rect 20450 7361 20462 7364
rect 20496 7392 20508 7395
rect 20640 7392 20668 7432
rect 20806 7420 20812 7432
rect 20864 7420 20870 7472
rect 20496 7364 20668 7392
rect 20717 7395 20775 7401
rect 20496 7361 20508 7364
rect 20450 7355 20508 7361
rect 20717 7361 20729 7395
rect 20763 7392 20775 7395
rect 20916 7392 20944 7491
rect 21266 7488 21272 7500
rect 21324 7488 21330 7540
rect 20763 7364 20944 7392
rect 20763 7361 20775 7364
rect 20717 7355 20775 7361
rect 15749 7327 15807 7333
rect 15749 7293 15761 7327
rect 15795 7293 15807 7327
rect 15749 7287 15807 7293
rect 14277 7259 14335 7265
rect 14277 7225 14289 7259
rect 14323 7225 14335 7259
rect 14277 7219 14335 7225
rect 14918 7188 14924 7200
rect 14108 7160 14924 7188
rect 11885 7151 11943 7157
rect 14918 7148 14924 7160
rect 14976 7148 14982 7200
rect 1104 7098 21896 7120
rect 1104 7046 3549 7098
rect 3601 7046 3613 7098
rect 3665 7046 3677 7098
rect 3729 7046 3741 7098
rect 3793 7046 3805 7098
rect 3857 7046 8747 7098
rect 8799 7046 8811 7098
rect 8863 7046 8875 7098
rect 8927 7046 8939 7098
rect 8991 7046 9003 7098
rect 9055 7046 13945 7098
rect 13997 7046 14009 7098
rect 14061 7046 14073 7098
rect 14125 7046 14137 7098
rect 14189 7046 14201 7098
rect 14253 7046 19143 7098
rect 19195 7046 19207 7098
rect 19259 7046 19271 7098
rect 19323 7046 19335 7098
rect 19387 7046 19399 7098
rect 19451 7046 21896 7098
rect 1104 7024 21896 7046
rect 5810 6944 5816 6996
rect 5868 6984 5874 6996
rect 6457 6987 6515 6993
rect 6457 6984 6469 6987
rect 5868 6956 6469 6984
rect 5868 6944 5874 6956
rect 6457 6953 6469 6956
rect 6503 6953 6515 6987
rect 7098 6984 7104 6996
rect 6457 6947 6515 6953
rect 7024 6956 7104 6984
rect 5626 6876 5632 6928
rect 5684 6916 5690 6928
rect 6822 6916 6828 6928
rect 5684 6888 6828 6916
rect 5684 6876 5690 6888
rect 6822 6876 6828 6888
rect 6880 6876 6886 6928
rect 3970 6848 3976 6860
rect 3931 6820 3976 6848
rect 3970 6808 3976 6820
rect 4028 6808 4034 6860
rect 4154 6848 4160 6860
rect 4115 6820 4160 6848
rect 4154 6808 4160 6820
rect 4212 6808 4218 6860
rect 7024 6857 7052 6956
rect 7098 6944 7104 6956
rect 7156 6984 7162 6996
rect 7377 6987 7435 6993
rect 7377 6984 7389 6987
rect 7156 6956 7389 6984
rect 7156 6944 7162 6956
rect 7377 6953 7389 6956
rect 7423 6984 7435 6987
rect 8386 6984 8392 6996
rect 7423 6956 7972 6984
rect 8347 6956 8392 6984
rect 7423 6953 7435 6956
rect 7377 6947 7435 6953
rect 7944 6916 7972 6956
rect 8386 6944 8392 6956
rect 8444 6944 8450 6996
rect 9306 6984 9312 6996
rect 9267 6956 9312 6984
rect 9306 6944 9312 6956
rect 9364 6944 9370 6996
rect 10502 6944 10508 6996
rect 10560 6984 10566 6996
rect 11698 6984 11704 6996
rect 10560 6956 11704 6984
rect 10560 6944 10566 6956
rect 11698 6944 11704 6956
rect 11756 6944 11762 6996
rect 13814 6944 13820 6996
rect 13872 6984 13878 6996
rect 14093 6987 14151 6993
rect 14093 6984 14105 6987
rect 13872 6956 14105 6984
rect 13872 6944 13878 6956
rect 14093 6953 14105 6956
rect 14139 6953 14151 6987
rect 14093 6947 14151 6953
rect 12250 6916 12256 6928
rect 7944 6888 12256 6916
rect 12250 6876 12256 6888
rect 12308 6876 12314 6928
rect 12986 6876 12992 6928
rect 13044 6876 13050 6928
rect 15010 6916 15016 6928
rect 14660 6888 15016 6916
rect 7009 6851 7067 6857
rect 7009 6817 7021 6851
rect 7055 6817 7067 6851
rect 7742 6848 7748 6860
rect 7703 6820 7748 6848
rect 7009 6811 7067 6817
rect 7742 6808 7748 6820
rect 7800 6808 7806 6860
rect 8570 6848 8576 6860
rect 8531 6820 8576 6848
rect 8570 6808 8576 6820
rect 8628 6848 8634 6860
rect 9030 6848 9036 6860
rect 8628 6820 9036 6848
rect 8628 6808 8634 6820
rect 9030 6808 9036 6820
rect 9088 6808 9094 6860
rect 9766 6808 9772 6860
rect 9824 6848 9830 6860
rect 9861 6851 9919 6857
rect 9861 6848 9873 6851
rect 9824 6820 9873 6848
rect 9824 6808 9830 6820
rect 9861 6817 9873 6820
rect 9907 6817 9919 6851
rect 9861 6811 9919 6817
rect 10229 6851 10287 6857
rect 10229 6817 10241 6851
rect 10275 6848 10287 6851
rect 10686 6848 10692 6860
rect 10275 6820 10692 6848
rect 10275 6817 10287 6820
rect 10229 6811 10287 6817
rect 10686 6808 10692 6820
rect 10744 6808 10750 6860
rect 11977 6851 12035 6857
rect 11977 6817 11989 6851
rect 12023 6848 12035 6851
rect 13004 6848 13032 6876
rect 14550 6848 14556 6860
rect 12023 6820 13032 6848
rect 14511 6820 14556 6848
rect 12023 6817 12035 6820
rect 11977 6811 12035 6817
rect 14550 6808 14556 6820
rect 14608 6808 14614 6860
rect 14660 6857 14688 6888
rect 15010 6876 15016 6888
rect 15068 6876 15074 6928
rect 14645 6851 14703 6857
rect 14645 6817 14657 6851
rect 14691 6817 14703 6851
rect 14645 6811 14703 6817
rect 14734 6808 14740 6860
rect 14792 6848 14798 6860
rect 14921 6851 14979 6857
rect 14921 6848 14933 6851
rect 14792 6820 14933 6848
rect 14792 6808 14798 6820
rect 14921 6817 14933 6820
rect 14967 6848 14979 6851
rect 15470 6848 15476 6860
rect 14967 6820 15476 6848
rect 14967 6817 14979 6820
rect 14921 6811 14979 6817
rect 15470 6808 15476 6820
rect 15528 6808 15534 6860
rect 3418 6780 3424 6792
rect 3331 6752 3424 6780
rect 3418 6740 3424 6752
rect 3476 6780 3482 6792
rect 4172 6780 4200 6808
rect 3476 6752 4200 6780
rect 4249 6783 4307 6789
rect 3476 6740 3482 6752
rect 4249 6749 4261 6783
rect 4295 6780 4307 6783
rect 4430 6780 4436 6792
rect 4295 6752 4436 6780
rect 4295 6749 4307 6752
rect 4249 6743 4307 6749
rect 3605 6715 3663 6721
rect 3605 6681 3617 6715
rect 3651 6712 3663 6715
rect 4264 6712 4292 6743
rect 4430 6740 4436 6752
rect 4488 6740 4494 6792
rect 5718 6740 5724 6792
rect 5776 6780 5782 6792
rect 6825 6783 6883 6789
rect 6825 6780 6837 6783
rect 5776 6752 6837 6780
rect 5776 6740 5782 6752
rect 6825 6749 6837 6752
rect 6871 6780 6883 6783
rect 8941 6783 8999 6789
rect 8941 6780 8953 6783
rect 6871 6752 8953 6780
rect 6871 6749 6883 6752
rect 6825 6743 6883 6749
rect 8941 6749 8953 6752
rect 8987 6780 8999 6783
rect 9677 6783 9735 6789
rect 9677 6780 9689 6783
rect 8987 6752 9689 6780
rect 8987 6749 8999 6752
rect 8941 6743 8999 6749
rect 9677 6749 9689 6752
rect 9723 6780 9735 6783
rect 10318 6780 10324 6792
rect 9723 6752 10324 6780
rect 9723 6749 9735 6752
rect 9677 6743 9735 6749
rect 10318 6740 10324 6752
rect 10376 6740 10382 6792
rect 12069 6783 12127 6789
rect 10704 6752 12020 6780
rect 10704 6724 10732 6752
rect 9950 6712 9956 6724
rect 3651 6684 4292 6712
rect 4632 6684 9956 6712
rect 3651 6681 3663 6684
rect 3605 6675 3663 6681
rect 4632 6653 4660 6684
rect 9950 6672 9956 6684
rect 10008 6672 10014 6724
rect 10505 6715 10563 6721
rect 10505 6712 10517 6715
rect 10060 6684 10517 6712
rect 4617 6647 4675 6653
rect 4617 6613 4629 6647
rect 4663 6613 4675 6647
rect 4617 6607 4675 6613
rect 4801 6647 4859 6653
rect 4801 6613 4813 6647
rect 4847 6644 4859 6647
rect 4982 6644 4988 6656
rect 4847 6616 4988 6644
rect 4847 6613 4859 6616
rect 4801 6607 4859 6613
rect 4982 6604 4988 6616
rect 5040 6604 5046 6656
rect 5166 6604 5172 6656
rect 5224 6644 5230 6656
rect 5537 6647 5595 6653
rect 5537 6644 5549 6647
rect 5224 6616 5549 6644
rect 5224 6604 5230 6616
rect 5537 6613 5549 6616
rect 5583 6613 5595 6647
rect 5718 6644 5724 6656
rect 5679 6616 5724 6644
rect 5537 6607 5595 6613
rect 5718 6604 5724 6616
rect 5776 6604 5782 6656
rect 5810 6604 5816 6656
rect 5868 6644 5874 6656
rect 5905 6647 5963 6653
rect 5905 6644 5917 6647
rect 5868 6616 5917 6644
rect 5868 6604 5874 6616
rect 5905 6613 5917 6616
rect 5951 6613 5963 6647
rect 5905 6607 5963 6613
rect 5994 6604 6000 6656
rect 6052 6644 6058 6656
rect 6089 6647 6147 6653
rect 6089 6644 6101 6647
rect 6052 6616 6101 6644
rect 6052 6604 6058 6616
rect 6089 6613 6101 6616
rect 6135 6613 6147 6647
rect 6362 6644 6368 6656
rect 6323 6616 6368 6644
rect 6089 6607 6147 6613
rect 6362 6604 6368 6616
rect 6420 6604 6426 6656
rect 6822 6604 6828 6656
rect 6880 6644 6886 6656
rect 6917 6647 6975 6653
rect 6917 6644 6929 6647
rect 6880 6616 6929 6644
rect 6880 6604 6886 6616
rect 6917 6613 6929 6616
rect 6963 6613 6975 6647
rect 6917 6607 6975 6613
rect 7190 6604 7196 6656
rect 7248 6644 7254 6656
rect 7469 6647 7527 6653
rect 7469 6644 7481 6647
rect 7248 6616 7481 6644
rect 7248 6604 7254 6616
rect 7469 6613 7481 6616
rect 7515 6613 7527 6647
rect 7469 6607 7527 6613
rect 7650 6604 7656 6656
rect 7708 6644 7714 6656
rect 7929 6647 7987 6653
rect 7929 6644 7941 6647
rect 7708 6616 7941 6644
rect 7708 6604 7714 6616
rect 7929 6613 7941 6616
rect 7975 6613 7987 6647
rect 7929 6607 7987 6613
rect 8021 6647 8079 6653
rect 8021 6613 8033 6647
rect 8067 6644 8079 6647
rect 8110 6644 8116 6656
rect 8067 6616 8116 6644
rect 8067 6613 8079 6616
rect 8021 6607 8079 6613
rect 8110 6604 8116 6616
rect 8168 6604 8174 6656
rect 9122 6644 9128 6656
rect 9083 6616 9128 6644
rect 9122 6604 9128 6616
rect 9180 6644 9186 6656
rect 9769 6647 9827 6653
rect 9769 6644 9781 6647
rect 9180 6616 9781 6644
rect 9180 6604 9186 6616
rect 9769 6613 9781 6616
rect 9815 6613 9827 6647
rect 9769 6607 9827 6613
rect 9858 6604 9864 6656
rect 9916 6644 9922 6656
rect 10060 6644 10088 6684
rect 10505 6681 10517 6684
rect 10551 6681 10563 6715
rect 10505 6675 10563 6681
rect 10686 6672 10692 6724
rect 10744 6672 10750 6724
rect 11790 6712 11796 6724
rect 10888 6684 11796 6712
rect 10410 6644 10416 6656
rect 9916 6616 10088 6644
rect 10371 6616 10416 6644
rect 9916 6604 9922 6616
rect 10410 6604 10416 6616
rect 10468 6604 10474 6656
rect 10888 6653 10916 6684
rect 11790 6672 11796 6684
rect 11848 6672 11854 6724
rect 11992 6712 12020 6752
rect 12069 6749 12081 6783
rect 12115 6780 12127 6783
rect 14366 6780 14372 6792
rect 12115 6752 14372 6780
rect 12115 6749 12127 6752
rect 12069 6743 12127 6749
rect 14366 6740 14372 6752
rect 14424 6740 14430 6792
rect 14642 6712 14648 6724
rect 11992 6684 14648 6712
rect 14642 6672 14648 6684
rect 14700 6672 14706 6724
rect 10873 6647 10931 6653
rect 10873 6613 10885 6647
rect 10919 6613 10931 6647
rect 10873 6607 10931 6613
rect 10962 6604 10968 6656
rect 11020 6644 11026 6656
rect 11609 6647 11667 6653
rect 11609 6644 11621 6647
rect 11020 6616 11621 6644
rect 11020 6604 11026 6616
rect 11609 6613 11621 6616
rect 11655 6644 11667 6647
rect 12161 6647 12219 6653
rect 12161 6644 12173 6647
rect 11655 6616 12173 6644
rect 11655 6613 11667 6616
rect 11609 6607 11667 6613
rect 12161 6613 12173 6616
rect 12207 6613 12219 6647
rect 12161 6607 12219 6613
rect 12434 6604 12440 6656
rect 12492 6644 12498 6656
rect 12529 6647 12587 6653
rect 12529 6644 12541 6647
rect 12492 6616 12541 6644
rect 12492 6604 12498 6616
rect 12529 6613 12541 6616
rect 12575 6613 12587 6647
rect 13814 6644 13820 6656
rect 13775 6616 13820 6644
rect 12529 6607 12587 6613
rect 13814 6604 13820 6616
rect 13872 6644 13878 6656
rect 14461 6647 14519 6653
rect 14461 6644 14473 6647
rect 13872 6616 14473 6644
rect 13872 6604 13878 6616
rect 14461 6613 14473 6616
rect 14507 6613 14519 6647
rect 14461 6607 14519 6613
rect 1104 6554 22056 6576
rect 1104 6502 6148 6554
rect 6200 6502 6212 6554
rect 6264 6502 6276 6554
rect 6328 6502 6340 6554
rect 6392 6502 6404 6554
rect 6456 6502 11346 6554
rect 11398 6502 11410 6554
rect 11462 6502 11474 6554
rect 11526 6502 11538 6554
rect 11590 6502 11602 6554
rect 11654 6502 16544 6554
rect 16596 6502 16608 6554
rect 16660 6502 16672 6554
rect 16724 6502 16736 6554
rect 16788 6502 16800 6554
rect 16852 6502 21742 6554
rect 21794 6502 21806 6554
rect 21858 6502 21870 6554
rect 21922 6502 21934 6554
rect 21986 6502 21998 6554
rect 22050 6502 22056 6554
rect 1104 6480 22056 6502
rect 2409 6443 2467 6449
rect 2409 6409 2421 6443
rect 2455 6440 2467 6443
rect 5169 6443 5227 6449
rect 5169 6440 5181 6443
rect 2455 6412 5181 6440
rect 2455 6409 2467 6412
rect 2409 6403 2467 6409
rect 5169 6409 5181 6412
rect 5215 6409 5227 6443
rect 5169 6403 5227 6409
rect 5629 6443 5687 6449
rect 5629 6409 5641 6443
rect 5675 6440 5687 6443
rect 7101 6443 7159 6449
rect 5675 6412 7052 6440
rect 5675 6409 5687 6412
rect 5629 6403 5687 6409
rect 3973 6375 4031 6381
rect 3973 6341 3985 6375
rect 4019 6372 4031 6375
rect 4338 6372 4344 6384
rect 4019 6344 4344 6372
rect 4019 6341 4031 6344
rect 3973 6335 4031 6341
rect 4338 6332 4344 6344
rect 4396 6332 4402 6384
rect 4433 6375 4491 6381
rect 4433 6341 4445 6375
rect 4479 6372 4491 6375
rect 5721 6375 5779 6381
rect 5721 6372 5733 6375
rect 4479 6344 5733 6372
rect 4479 6341 4491 6344
rect 4433 6335 4491 6341
rect 5721 6341 5733 6344
rect 5767 6341 5779 6375
rect 7024 6372 7052 6412
rect 7101 6409 7113 6443
rect 7147 6440 7159 6443
rect 7374 6440 7380 6452
rect 7147 6412 7380 6440
rect 7147 6409 7159 6412
rect 7101 6403 7159 6409
rect 7374 6400 7380 6412
rect 7432 6400 7438 6452
rect 7469 6443 7527 6449
rect 7469 6409 7481 6443
rect 7515 6440 7527 6443
rect 7929 6443 7987 6449
rect 7929 6440 7941 6443
rect 7515 6412 7941 6440
rect 7515 6409 7527 6412
rect 7469 6403 7527 6409
rect 7929 6409 7941 6412
rect 7975 6409 7987 6443
rect 7929 6403 7987 6409
rect 8110 6400 8116 6452
rect 8168 6440 8174 6452
rect 8389 6443 8447 6449
rect 8389 6440 8401 6443
rect 8168 6412 8401 6440
rect 8168 6400 8174 6412
rect 8389 6409 8401 6412
rect 8435 6409 8447 6443
rect 8389 6403 8447 6409
rect 8662 6400 8668 6452
rect 8720 6440 8726 6452
rect 8757 6443 8815 6449
rect 8757 6440 8769 6443
rect 8720 6412 8769 6440
rect 8720 6400 8726 6412
rect 8757 6409 8769 6412
rect 8803 6409 8815 6443
rect 8757 6403 8815 6409
rect 9030 6400 9036 6452
rect 9088 6440 9094 6452
rect 9217 6443 9275 6449
rect 9217 6440 9229 6443
rect 9088 6412 9229 6440
rect 9088 6400 9094 6412
rect 9217 6409 9229 6412
rect 9263 6409 9275 6443
rect 9950 6440 9956 6452
rect 9911 6412 9956 6440
rect 9217 6403 9275 6409
rect 9950 6400 9956 6412
rect 10008 6400 10014 6452
rect 10410 6400 10416 6452
rect 10468 6440 10474 6452
rect 12253 6443 12311 6449
rect 12253 6440 12265 6443
rect 10468 6412 12265 6440
rect 10468 6400 10474 6412
rect 12253 6409 12265 6412
rect 12299 6409 12311 6443
rect 12253 6403 12311 6409
rect 12618 6400 12624 6452
rect 12676 6440 12682 6452
rect 12713 6443 12771 6449
rect 12713 6440 12725 6443
rect 12676 6412 12725 6440
rect 12676 6400 12682 6412
rect 12713 6409 12725 6412
rect 12759 6409 12771 6443
rect 12713 6403 12771 6409
rect 13262 6400 13268 6452
rect 13320 6440 13326 6452
rect 14185 6443 14243 6449
rect 14185 6440 14197 6443
rect 13320 6412 14197 6440
rect 13320 6400 13326 6412
rect 14185 6409 14197 6412
rect 14231 6409 14243 6443
rect 14185 6403 14243 6409
rect 14277 6443 14335 6449
rect 14277 6409 14289 6443
rect 14323 6440 14335 6443
rect 14458 6440 14464 6452
rect 14323 6412 14464 6440
rect 14323 6409 14335 6412
rect 14277 6403 14335 6409
rect 14458 6400 14464 6412
rect 14516 6400 14522 6452
rect 10594 6372 10600 6384
rect 7024 6344 10600 6372
rect 5721 6335 5779 6341
rect 10594 6332 10600 6344
rect 10652 6332 10658 6384
rect 11330 6372 11336 6384
rect 11072 6344 11336 6372
rect 1486 6264 1492 6316
rect 1544 6304 1550 6316
rect 2041 6307 2099 6313
rect 2041 6304 2053 6307
rect 1544 6276 2053 6304
rect 1544 6264 1550 6276
rect 2041 6273 2053 6276
rect 2087 6273 2099 6307
rect 2041 6267 2099 6273
rect 4246 6264 4252 6316
rect 4304 6304 4310 6316
rect 5261 6307 5319 6313
rect 5261 6304 5273 6307
rect 4304 6276 5273 6304
rect 4304 6264 4310 6276
rect 5261 6273 5273 6276
rect 5307 6273 5319 6307
rect 5261 6267 5319 6273
rect 5626 6264 5632 6316
rect 5684 6304 5690 6316
rect 5994 6304 6000 6316
rect 5684 6276 6000 6304
rect 5684 6264 5690 6276
rect 5994 6264 6000 6276
rect 6052 6264 6058 6316
rect 6181 6307 6239 6313
rect 6181 6273 6193 6307
rect 6227 6304 6239 6307
rect 6914 6304 6920 6316
rect 6227 6276 6920 6304
rect 6227 6273 6239 6276
rect 6181 6267 6239 6273
rect 6914 6264 6920 6276
rect 6972 6264 6978 6316
rect 7009 6307 7067 6313
rect 7009 6273 7021 6307
rect 7055 6304 7067 6307
rect 7098 6304 7104 6316
rect 7055 6276 7104 6304
rect 7055 6273 7067 6276
rect 7009 6267 7067 6273
rect 7098 6264 7104 6276
rect 7156 6264 7162 6316
rect 7374 6304 7380 6316
rect 7208 6276 7380 6304
rect 1854 6236 1860 6248
rect 1815 6208 1860 6236
rect 1854 6196 1860 6208
rect 1912 6196 1918 6248
rect 1949 6239 2007 6245
rect 1949 6205 1961 6239
rect 1995 6205 2007 6239
rect 1949 6199 2007 6205
rect 1394 6060 1400 6112
rect 1452 6100 1458 6112
rect 1489 6103 1547 6109
rect 1489 6100 1501 6103
rect 1452 6072 1501 6100
rect 1452 6060 1458 6072
rect 1489 6069 1501 6072
rect 1535 6100 1547 6103
rect 1964 6100 1992 6199
rect 3970 6196 3976 6248
rect 4028 6236 4034 6248
rect 4157 6239 4215 6245
rect 4157 6236 4169 6239
rect 4028 6208 4169 6236
rect 4028 6196 4034 6208
rect 4157 6205 4169 6208
rect 4203 6236 4215 6239
rect 4982 6236 4988 6248
rect 4203 6208 4988 6236
rect 4203 6205 4215 6208
rect 4157 6199 4215 6205
rect 4982 6196 4988 6208
rect 5040 6196 5046 6248
rect 5077 6239 5135 6245
rect 5077 6205 5089 6239
rect 5123 6236 5135 6239
rect 7208 6236 7236 6276
rect 7374 6264 7380 6276
rect 7432 6264 7438 6316
rect 8018 6264 8024 6316
rect 8076 6304 8082 6316
rect 8297 6307 8355 6313
rect 8297 6304 8309 6307
rect 8076 6276 8309 6304
rect 8076 6264 8082 6276
rect 8297 6273 8309 6276
rect 8343 6273 8355 6307
rect 8297 6267 8355 6273
rect 8386 6264 8392 6316
rect 8444 6304 8450 6316
rect 9125 6307 9183 6313
rect 9125 6304 9137 6307
rect 8444 6276 9137 6304
rect 8444 6264 8450 6276
rect 9125 6273 9137 6276
rect 9171 6273 9183 6307
rect 9125 6267 9183 6273
rect 10045 6307 10103 6313
rect 10045 6273 10057 6307
rect 10091 6273 10103 6307
rect 10045 6267 10103 6273
rect 10965 6307 11023 6313
rect 10965 6273 10977 6307
rect 11011 6304 11023 6307
rect 11072 6304 11100 6344
rect 11330 6332 11336 6344
rect 11388 6332 11394 6384
rect 14734 6372 14740 6384
rect 12544 6344 14740 6372
rect 12544 6304 12572 6344
rect 14734 6332 14740 6344
rect 14792 6332 14798 6384
rect 11011 6276 11100 6304
rect 11256 6276 12572 6304
rect 12621 6307 12679 6313
rect 11011 6273 11023 6276
rect 10965 6267 11023 6273
rect 7558 6236 7564 6248
rect 5123 6208 7236 6236
rect 7519 6208 7564 6236
rect 5123 6205 5135 6208
rect 5077 6199 5135 6205
rect 7558 6196 7564 6208
rect 7616 6196 7622 6248
rect 7745 6239 7803 6245
rect 7745 6205 7757 6239
rect 7791 6236 7803 6239
rect 8202 6236 8208 6248
rect 7791 6208 8208 6236
rect 7791 6205 7803 6208
rect 7745 6199 7803 6205
rect 8202 6196 8208 6208
rect 8260 6196 8266 6248
rect 8478 6196 8484 6248
rect 8536 6236 8542 6248
rect 8573 6239 8631 6245
rect 8573 6236 8585 6239
rect 8536 6208 8585 6236
rect 8536 6196 8542 6208
rect 8573 6205 8585 6208
rect 8619 6236 8631 6239
rect 9401 6239 9459 6245
rect 9401 6236 9413 6239
rect 8619 6208 9413 6236
rect 8619 6205 8631 6208
rect 8573 6199 8631 6205
rect 9401 6205 9413 6208
rect 9447 6236 9459 6239
rect 9582 6236 9588 6248
rect 9447 6208 9588 6236
rect 9447 6205 9459 6208
rect 9401 6199 9459 6205
rect 9582 6196 9588 6208
rect 9640 6196 9646 6248
rect 9858 6236 9864 6248
rect 9819 6208 9864 6236
rect 9858 6196 9864 6208
rect 9916 6196 9922 6248
rect 4801 6171 4859 6177
rect 4801 6137 4813 6171
rect 4847 6168 4859 6171
rect 10060 6168 10088 6267
rect 10686 6236 10692 6248
rect 10647 6208 10692 6236
rect 10686 6196 10692 6208
rect 10744 6196 10750 6248
rect 10870 6196 10876 6248
rect 10928 6236 10934 6248
rect 10928 6208 10973 6236
rect 10928 6196 10934 6208
rect 4847 6140 10088 6168
rect 10413 6171 10471 6177
rect 4847 6137 4859 6140
rect 4801 6131 4859 6137
rect 10413 6137 10425 6171
rect 10459 6168 10471 6171
rect 11256 6168 11284 6276
rect 12621 6273 12633 6307
rect 12667 6273 12679 6307
rect 15562 6304 15568 6316
rect 12621 6267 12679 6273
rect 12820 6276 15568 6304
rect 11514 6236 11520 6248
rect 11475 6208 11520 6236
rect 11514 6196 11520 6208
rect 11572 6196 11578 6248
rect 11701 6239 11759 6245
rect 11701 6205 11713 6239
rect 11747 6236 11759 6239
rect 11790 6236 11796 6248
rect 11747 6208 11796 6236
rect 11747 6205 11759 6208
rect 11701 6199 11759 6205
rect 11790 6196 11796 6208
rect 11848 6196 11854 6248
rect 12434 6236 12440 6248
rect 11992 6208 12440 6236
rect 10459 6140 11284 6168
rect 11333 6171 11391 6177
rect 10459 6137 10471 6140
rect 10413 6131 10471 6137
rect 11333 6137 11345 6171
rect 11379 6168 11391 6171
rect 11992 6168 12020 6208
rect 12434 6196 12440 6208
rect 12492 6196 12498 6248
rect 12526 6196 12532 6248
rect 12584 6236 12590 6248
rect 12636 6236 12664 6267
rect 12820 6245 12848 6276
rect 15562 6264 15568 6276
rect 15620 6264 15626 6316
rect 12584 6208 12664 6236
rect 12805 6239 12863 6245
rect 12584 6196 12590 6208
rect 12805 6205 12817 6239
rect 12851 6205 12863 6239
rect 12805 6199 12863 6205
rect 14093 6239 14151 6245
rect 14093 6205 14105 6239
rect 14139 6236 14151 6239
rect 19702 6236 19708 6248
rect 14139 6208 19708 6236
rect 14139 6205 14151 6208
rect 14093 6199 14151 6205
rect 19702 6196 19708 6208
rect 19760 6196 19766 6248
rect 11379 6140 12020 6168
rect 11379 6137 11391 6140
rect 11333 6131 11391 6137
rect 12158 6128 12164 6180
rect 12216 6168 12222 6180
rect 16298 6168 16304 6180
rect 12216 6140 16304 6168
rect 12216 6128 12222 6140
rect 16298 6128 16304 6140
rect 16356 6128 16362 6180
rect 1535 6072 1992 6100
rect 1535 6069 1547 6072
rect 1489 6063 1547 6069
rect 6270 6060 6276 6112
rect 6328 6100 6334 6112
rect 6365 6103 6423 6109
rect 6365 6100 6377 6103
rect 6328 6072 6377 6100
rect 6328 6060 6334 6072
rect 6365 6069 6377 6072
rect 6411 6069 6423 6103
rect 6365 6063 6423 6069
rect 7282 6060 7288 6112
rect 7340 6100 7346 6112
rect 12069 6103 12127 6109
rect 12069 6100 12081 6103
rect 7340 6072 12081 6100
rect 7340 6060 7346 6072
rect 12069 6069 12081 6072
rect 12115 6100 12127 6103
rect 12526 6100 12532 6112
rect 12115 6072 12532 6100
rect 12115 6069 12127 6072
rect 12069 6063 12127 6069
rect 12526 6060 12532 6072
rect 12584 6060 12590 6112
rect 14645 6103 14703 6109
rect 14645 6069 14657 6103
rect 14691 6100 14703 6103
rect 15838 6100 15844 6112
rect 14691 6072 15844 6100
rect 14691 6069 14703 6072
rect 14645 6063 14703 6069
rect 15838 6060 15844 6072
rect 15896 6060 15902 6112
rect 1104 6010 21896 6032
rect 1104 5958 3549 6010
rect 3601 5958 3613 6010
rect 3665 5958 3677 6010
rect 3729 5958 3741 6010
rect 3793 5958 3805 6010
rect 3857 5958 8747 6010
rect 8799 5958 8811 6010
rect 8863 5958 8875 6010
rect 8927 5958 8939 6010
rect 8991 5958 9003 6010
rect 9055 5958 13945 6010
rect 13997 5958 14009 6010
rect 14061 5958 14073 6010
rect 14125 5958 14137 6010
rect 14189 5958 14201 6010
rect 14253 5958 19143 6010
rect 19195 5958 19207 6010
rect 19259 5958 19271 6010
rect 19323 5958 19335 6010
rect 19387 5958 19399 6010
rect 19451 5958 21896 6010
rect 1104 5936 21896 5958
rect 1486 5896 1492 5908
rect 1447 5868 1492 5896
rect 1486 5856 1492 5868
rect 1544 5856 1550 5908
rect 5353 5899 5411 5905
rect 5353 5865 5365 5899
rect 5399 5896 5411 5899
rect 5534 5896 5540 5908
rect 5399 5868 5540 5896
rect 5399 5865 5411 5868
rect 5353 5859 5411 5865
rect 5534 5856 5540 5868
rect 5592 5896 5598 5908
rect 5810 5896 5816 5908
rect 5592 5868 5816 5896
rect 5592 5856 5598 5868
rect 5810 5856 5816 5868
rect 5868 5856 5874 5908
rect 7006 5896 7012 5908
rect 5920 5868 7012 5896
rect 5258 5720 5264 5772
rect 5316 5760 5322 5772
rect 5721 5763 5779 5769
rect 5721 5760 5733 5763
rect 5316 5732 5733 5760
rect 5316 5720 5322 5732
rect 5721 5729 5733 5732
rect 5767 5729 5779 5763
rect 5721 5723 5779 5729
rect 5442 5652 5448 5704
rect 5500 5692 5506 5704
rect 5920 5701 5948 5868
rect 7006 5856 7012 5868
rect 7064 5856 7070 5908
rect 7193 5899 7251 5905
rect 7193 5865 7205 5899
rect 7239 5896 7251 5899
rect 7558 5896 7564 5908
rect 7239 5868 7564 5896
rect 7239 5865 7251 5868
rect 7193 5859 7251 5865
rect 7558 5856 7564 5868
rect 7616 5856 7622 5908
rect 7742 5896 7748 5908
rect 7703 5868 7748 5896
rect 7742 5856 7748 5868
rect 7800 5896 7806 5908
rect 8110 5896 8116 5908
rect 7800 5868 8116 5896
rect 7800 5856 7806 5868
rect 8110 5856 8116 5868
rect 8168 5856 8174 5908
rect 8757 5899 8815 5905
rect 8757 5865 8769 5899
rect 8803 5896 8815 5899
rect 10870 5896 10876 5908
rect 8803 5868 10876 5896
rect 8803 5865 8815 5868
rect 8757 5859 8815 5865
rect 10870 5856 10876 5868
rect 10928 5856 10934 5908
rect 11149 5899 11207 5905
rect 11149 5865 11161 5899
rect 11195 5896 11207 5899
rect 13262 5896 13268 5908
rect 11195 5868 13032 5896
rect 13223 5868 13268 5896
rect 11195 5865 11207 5868
rect 11149 5859 11207 5865
rect 7466 5788 7472 5840
rect 7524 5828 7530 5840
rect 7653 5831 7711 5837
rect 7653 5828 7665 5831
rect 7524 5800 7665 5828
rect 7524 5788 7530 5800
rect 7653 5797 7665 5800
rect 7699 5828 7711 5831
rect 8018 5828 8024 5840
rect 7699 5800 8024 5828
rect 7699 5797 7711 5800
rect 7653 5791 7711 5797
rect 8018 5788 8024 5800
rect 8076 5788 8082 5840
rect 8386 5788 8392 5840
rect 8444 5828 8450 5840
rect 8941 5831 8999 5837
rect 8941 5828 8953 5831
rect 8444 5800 8953 5828
rect 8444 5788 8450 5800
rect 8941 5797 8953 5800
rect 8987 5797 8999 5831
rect 8941 5791 8999 5797
rect 9030 5788 9036 5840
rect 9088 5828 9094 5840
rect 9125 5831 9183 5837
rect 9125 5828 9137 5831
rect 9088 5800 9137 5828
rect 9088 5788 9094 5800
rect 9125 5797 9137 5800
rect 9171 5797 9183 5831
rect 9125 5791 9183 5797
rect 9858 5788 9864 5840
rect 9916 5828 9922 5840
rect 9916 5800 11744 5828
rect 9916 5788 9922 5800
rect 6546 5760 6552 5772
rect 6507 5732 6552 5760
rect 6546 5720 6552 5732
rect 6604 5720 6610 5772
rect 7374 5720 7380 5772
rect 7432 5760 7438 5772
rect 8205 5763 8263 5769
rect 8205 5760 8217 5763
rect 7432 5732 8217 5760
rect 7432 5720 7438 5732
rect 8205 5729 8217 5732
rect 8251 5760 8263 5763
rect 8251 5732 8524 5760
rect 8251 5729 8263 5732
rect 8205 5723 8263 5729
rect 5905 5695 5963 5701
rect 5905 5692 5917 5695
rect 5500 5664 5917 5692
rect 5500 5652 5506 5664
rect 5905 5661 5917 5664
rect 5951 5661 5963 5695
rect 8496 5692 8524 5732
rect 8570 5720 8576 5772
rect 8628 5760 8634 5772
rect 9490 5760 9496 5772
rect 8628 5732 9496 5760
rect 8628 5720 8634 5732
rect 9490 5720 9496 5732
rect 9548 5760 9554 5772
rect 9677 5763 9735 5769
rect 9677 5760 9689 5763
rect 9548 5732 9689 5760
rect 9548 5720 9554 5732
rect 9677 5729 9689 5732
rect 9723 5729 9735 5763
rect 9677 5723 9735 5729
rect 10597 5763 10655 5769
rect 10597 5729 10609 5763
rect 10643 5760 10655 5763
rect 11609 5763 11667 5769
rect 11609 5760 11621 5763
rect 10643 5732 11621 5760
rect 10643 5729 10655 5732
rect 10597 5723 10655 5729
rect 11609 5729 11621 5732
rect 11655 5729 11667 5763
rect 11716 5760 11744 5800
rect 12526 5760 12532 5772
rect 11716 5732 12532 5760
rect 11609 5723 11667 5729
rect 10778 5692 10784 5704
rect 8496 5664 10784 5692
rect 5905 5655 5963 5661
rect 10778 5652 10784 5664
rect 10836 5652 10842 5704
rect 4522 5584 4528 5636
rect 4580 5624 4586 5636
rect 6270 5624 6276 5636
rect 4580 5596 6276 5624
rect 4580 5584 4586 5596
rect 6270 5584 6276 5596
rect 6328 5624 6334 5636
rect 6825 5627 6883 5633
rect 6825 5624 6837 5627
rect 6328 5596 6837 5624
rect 6328 5584 6334 5596
rect 6825 5593 6837 5596
rect 6871 5593 6883 5627
rect 6825 5587 6883 5593
rect 8297 5627 8355 5633
rect 8297 5593 8309 5627
rect 8343 5624 8355 5627
rect 8938 5624 8944 5636
rect 8343 5596 8944 5624
rect 8343 5593 8355 5596
rect 8297 5587 8355 5593
rect 8938 5584 8944 5596
rect 8996 5584 9002 5636
rect 9048 5596 9260 5624
rect 4982 5556 4988 5568
rect 4943 5528 4988 5556
rect 4982 5516 4988 5528
rect 5040 5516 5046 5568
rect 5166 5556 5172 5568
rect 5127 5528 5172 5556
rect 5166 5516 5172 5528
rect 5224 5516 5230 5568
rect 5442 5556 5448 5568
rect 5403 5528 5448 5556
rect 5442 5516 5448 5528
rect 5500 5516 5506 5568
rect 5810 5516 5816 5568
rect 5868 5556 5874 5568
rect 5997 5559 6055 5565
rect 5997 5556 6009 5559
rect 5868 5528 6009 5556
rect 5868 5516 5874 5528
rect 5997 5525 6009 5528
rect 6043 5525 6055 5559
rect 5997 5519 6055 5525
rect 6365 5559 6423 5565
rect 6365 5525 6377 5559
rect 6411 5556 6423 5559
rect 6638 5556 6644 5568
rect 6411 5528 6644 5556
rect 6411 5525 6423 5528
rect 6365 5519 6423 5525
rect 6638 5516 6644 5528
rect 6696 5516 6702 5568
rect 6733 5559 6791 5565
rect 6733 5525 6745 5559
rect 6779 5556 6791 5559
rect 6914 5556 6920 5568
rect 6779 5528 6920 5556
rect 6779 5525 6791 5528
rect 6733 5519 6791 5525
rect 6914 5516 6920 5528
rect 6972 5516 6978 5568
rect 7374 5516 7380 5568
rect 7432 5556 7438 5568
rect 8389 5559 8447 5565
rect 8389 5556 8401 5559
rect 7432 5528 8401 5556
rect 7432 5516 7438 5528
rect 8389 5525 8401 5528
rect 8435 5525 8447 5559
rect 8389 5519 8447 5525
rect 8846 5516 8852 5568
rect 8904 5556 8910 5568
rect 9048 5556 9076 5596
rect 8904 5528 9076 5556
rect 9232 5556 9260 5596
rect 9306 5584 9312 5636
rect 9364 5624 9370 5636
rect 9585 5627 9643 5633
rect 9585 5624 9597 5627
rect 9364 5596 9597 5624
rect 9364 5584 9370 5596
rect 9585 5593 9597 5596
rect 9631 5593 9643 5627
rect 9585 5587 9643 5593
rect 10134 5584 10140 5636
rect 10192 5624 10198 5636
rect 10594 5624 10600 5636
rect 10192 5596 10600 5624
rect 10192 5584 10198 5596
rect 10594 5584 10600 5596
rect 10652 5584 10658 5636
rect 11624 5624 11652 5723
rect 12526 5720 12532 5732
rect 12584 5720 12590 5772
rect 12713 5763 12771 5769
rect 12713 5729 12725 5763
rect 12759 5760 12771 5763
rect 12802 5760 12808 5772
rect 12759 5732 12808 5760
rect 12759 5729 12771 5732
rect 12713 5723 12771 5729
rect 12802 5720 12808 5732
rect 12860 5720 12866 5772
rect 13004 5760 13032 5868
rect 13262 5856 13268 5868
rect 13320 5856 13326 5908
rect 19610 5896 19616 5908
rect 16684 5868 19616 5896
rect 16684 5769 16712 5868
rect 19610 5856 19616 5868
rect 19668 5856 19674 5908
rect 17313 5831 17371 5837
rect 17313 5797 17325 5831
rect 17359 5828 17371 5831
rect 19058 5828 19064 5840
rect 17359 5800 19064 5828
rect 17359 5797 17371 5800
rect 17313 5791 17371 5797
rect 19058 5788 19064 5800
rect 19116 5788 19122 5840
rect 20622 5828 20628 5840
rect 19168 5800 20628 5828
rect 16669 5763 16727 5769
rect 13004 5732 14044 5760
rect 11790 5692 11796 5704
rect 11751 5664 11796 5692
rect 11790 5652 11796 5664
rect 11848 5652 11854 5704
rect 12434 5652 12440 5704
rect 12492 5692 12498 5704
rect 13357 5695 13415 5701
rect 13357 5692 13369 5695
rect 12492 5664 13369 5692
rect 12492 5652 12498 5664
rect 13357 5661 13369 5664
rect 13403 5661 13415 5695
rect 14016 5692 14044 5732
rect 16669 5729 16681 5763
rect 16715 5729 16727 5763
rect 16669 5723 16727 5729
rect 17494 5720 17500 5772
rect 17552 5760 17558 5772
rect 17589 5763 17647 5769
rect 17589 5760 17601 5763
rect 17552 5732 17601 5760
rect 17552 5720 17558 5732
rect 17589 5729 17601 5732
rect 17635 5760 17647 5763
rect 19168 5760 19196 5800
rect 20622 5788 20628 5800
rect 20680 5788 20686 5840
rect 17635 5732 19196 5760
rect 20165 5763 20223 5769
rect 17635 5729 17647 5732
rect 17589 5723 17647 5729
rect 20165 5729 20177 5763
rect 20211 5760 20223 5763
rect 21174 5760 21180 5772
rect 20211 5732 21180 5760
rect 20211 5729 20223 5732
rect 20165 5723 20223 5729
rect 21174 5720 21180 5732
rect 21232 5720 21238 5772
rect 16853 5695 16911 5701
rect 16853 5692 16865 5695
rect 14016 5664 16865 5692
rect 13357 5655 13415 5661
rect 16853 5661 16865 5664
rect 16899 5661 16911 5695
rect 16853 5655 16911 5661
rect 13633 5627 13691 5633
rect 11624 5596 13584 5624
rect 9493 5559 9551 5565
rect 9493 5556 9505 5559
rect 9232 5528 9505 5556
rect 8904 5516 8910 5528
rect 9493 5525 9505 5528
rect 9539 5525 9551 5559
rect 10686 5556 10692 5568
rect 10647 5528 10692 5556
rect 9493 5519 9551 5525
rect 10686 5516 10692 5528
rect 10744 5516 10750 5568
rect 10778 5516 10784 5568
rect 10836 5556 10842 5568
rect 11698 5556 11704 5568
rect 10836 5528 10881 5556
rect 11659 5528 11704 5556
rect 10836 5516 10842 5528
rect 11698 5516 11704 5528
rect 11756 5516 11762 5568
rect 12161 5559 12219 5565
rect 12161 5525 12173 5559
rect 12207 5556 12219 5559
rect 12434 5556 12440 5568
rect 12207 5528 12440 5556
rect 12207 5525 12219 5528
rect 12161 5519 12219 5525
rect 12434 5516 12440 5528
rect 12492 5516 12498 5568
rect 12802 5556 12808 5568
rect 12763 5528 12808 5556
rect 12802 5516 12808 5528
rect 12860 5516 12866 5568
rect 12894 5516 12900 5568
rect 12952 5556 12958 5568
rect 13556 5556 13584 5596
rect 13633 5593 13645 5627
rect 13679 5624 13691 5627
rect 14274 5624 14280 5636
rect 13679 5596 14280 5624
rect 13679 5593 13691 5596
rect 13633 5587 13691 5593
rect 14274 5584 14280 5596
rect 14332 5584 14338 5636
rect 14366 5584 14372 5636
rect 14424 5624 14430 5636
rect 17681 5627 17739 5633
rect 17681 5624 17693 5627
rect 14424 5596 17693 5624
rect 14424 5584 14430 5596
rect 17681 5593 17693 5596
rect 17727 5593 17739 5627
rect 20349 5627 20407 5633
rect 20349 5624 20361 5627
rect 17681 5587 17739 5593
rect 18156 5596 20361 5624
rect 15654 5556 15660 5568
rect 12952 5528 12997 5556
rect 13556 5528 15660 5556
rect 12952 5516 12958 5528
rect 15654 5516 15660 5528
rect 15712 5516 15718 5568
rect 16390 5516 16396 5568
rect 16448 5556 16454 5568
rect 16945 5559 17003 5565
rect 16945 5556 16957 5559
rect 16448 5528 16957 5556
rect 16448 5516 16454 5528
rect 16945 5525 16957 5528
rect 16991 5525 17003 5559
rect 16945 5519 17003 5525
rect 17770 5516 17776 5568
rect 17828 5556 17834 5568
rect 18156 5565 18184 5596
rect 20349 5593 20361 5596
rect 20395 5593 20407 5627
rect 20349 5587 20407 5593
rect 18141 5559 18199 5565
rect 17828 5528 17873 5556
rect 17828 5516 17834 5528
rect 18141 5525 18153 5559
rect 18187 5525 18199 5559
rect 20254 5556 20260 5568
rect 20215 5528 20260 5556
rect 18141 5519 18199 5525
rect 20254 5516 20260 5528
rect 20312 5516 20318 5568
rect 20622 5516 20628 5568
rect 20680 5556 20686 5568
rect 20717 5559 20775 5565
rect 20717 5556 20729 5559
rect 20680 5528 20729 5556
rect 20680 5516 20686 5528
rect 20717 5525 20729 5528
rect 20763 5525 20775 5559
rect 20717 5519 20775 5525
rect 1104 5466 22056 5488
rect 1104 5414 6148 5466
rect 6200 5414 6212 5466
rect 6264 5414 6276 5466
rect 6328 5414 6340 5466
rect 6392 5414 6404 5466
rect 6456 5414 11346 5466
rect 11398 5414 11410 5466
rect 11462 5414 11474 5466
rect 11526 5414 11538 5466
rect 11590 5414 11602 5466
rect 11654 5414 16544 5466
rect 16596 5414 16608 5466
rect 16660 5414 16672 5466
rect 16724 5414 16736 5466
rect 16788 5414 16800 5466
rect 16852 5414 21742 5466
rect 21794 5414 21806 5466
rect 21858 5414 21870 5466
rect 21922 5414 21934 5466
rect 21986 5414 21998 5466
rect 22050 5414 22056 5466
rect 1104 5392 22056 5414
rect 1765 5355 1823 5361
rect 1765 5321 1777 5355
rect 1811 5352 1823 5355
rect 2133 5355 2191 5361
rect 2133 5352 2145 5355
rect 1811 5324 2145 5352
rect 1811 5321 1823 5324
rect 1765 5315 1823 5321
rect 2133 5321 2145 5324
rect 2179 5352 2191 5355
rect 2958 5352 2964 5364
rect 2179 5324 2964 5352
rect 2179 5321 2191 5324
rect 2133 5315 2191 5321
rect 2958 5312 2964 5324
rect 3016 5312 3022 5364
rect 3786 5312 3792 5364
rect 3844 5352 3850 5364
rect 4706 5352 4712 5364
rect 3844 5324 4712 5352
rect 3844 5312 3850 5324
rect 4706 5312 4712 5324
rect 4764 5312 4770 5364
rect 5074 5352 5080 5364
rect 5035 5324 5080 5352
rect 5074 5312 5080 5324
rect 5132 5312 5138 5364
rect 6638 5352 6644 5364
rect 6599 5324 6644 5352
rect 6638 5312 6644 5324
rect 6696 5312 6702 5364
rect 7101 5355 7159 5361
rect 7101 5321 7113 5355
rect 7147 5321 7159 5355
rect 7926 5352 7932 5364
rect 7887 5324 7932 5352
rect 7101 5315 7159 5321
rect 5537 5287 5595 5293
rect 5537 5284 5549 5287
rect 4632 5256 5549 5284
rect 2225 5219 2283 5225
rect 2225 5185 2237 5219
rect 2271 5216 2283 5219
rect 2685 5219 2743 5225
rect 2685 5216 2697 5219
rect 2271 5188 2697 5216
rect 2271 5185 2283 5188
rect 2225 5179 2283 5185
rect 2685 5185 2697 5188
rect 2731 5185 2743 5219
rect 2685 5179 2743 5185
rect 4062 5176 4068 5228
rect 4120 5216 4126 5228
rect 4632 5225 4660 5256
rect 5537 5253 5549 5256
rect 5583 5253 5595 5287
rect 5537 5247 5595 5253
rect 4617 5219 4675 5225
rect 4617 5216 4629 5219
rect 4120 5188 4629 5216
rect 4120 5176 4126 5188
rect 4617 5185 4629 5188
rect 4663 5185 4675 5219
rect 5166 5216 5172 5228
rect 4617 5179 4675 5185
rect 4724 5188 5172 5216
rect 4724 5160 4752 5188
rect 5166 5176 5172 5188
rect 5224 5176 5230 5228
rect 5810 5176 5816 5228
rect 5868 5216 5874 5228
rect 6733 5219 6791 5225
rect 6733 5216 6745 5219
rect 5868 5188 6745 5216
rect 5868 5176 5874 5188
rect 6733 5185 6745 5188
rect 6779 5185 6791 5219
rect 7116 5216 7144 5315
rect 7926 5312 7932 5324
rect 7984 5312 7990 5364
rect 8389 5355 8447 5361
rect 8389 5352 8401 5355
rect 8036 5324 8401 5352
rect 7742 5244 7748 5296
rect 7800 5284 7806 5296
rect 8036 5284 8064 5324
rect 8389 5321 8401 5324
rect 8435 5321 8447 5355
rect 8389 5315 8447 5321
rect 8938 5312 8944 5364
rect 8996 5352 9002 5364
rect 9033 5355 9091 5361
rect 9033 5352 9045 5355
rect 8996 5324 9045 5352
rect 8996 5312 9002 5324
rect 9033 5321 9045 5324
rect 9079 5321 9091 5355
rect 9033 5315 9091 5321
rect 9398 5312 9404 5364
rect 9456 5352 9462 5364
rect 9677 5355 9735 5361
rect 9677 5352 9689 5355
rect 9456 5324 9689 5352
rect 9456 5312 9462 5324
rect 9677 5321 9689 5324
rect 9723 5321 9735 5355
rect 9677 5315 9735 5321
rect 10137 5355 10195 5361
rect 10137 5321 10149 5355
rect 10183 5352 10195 5355
rect 10686 5352 10692 5364
rect 10183 5324 10692 5352
rect 10183 5321 10195 5324
rect 10137 5315 10195 5321
rect 10686 5312 10692 5324
rect 10744 5312 10750 5364
rect 10965 5355 11023 5361
rect 10965 5321 10977 5355
rect 11011 5352 11023 5355
rect 11885 5355 11943 5361
rect 11885 5352 11897 5355
rect 11011 5324 11897 5352
rect 11011 5321 11023 5324
rect 10965 5315 11023 5321
rect 11885 5321 11897 5324
rect 11931 5321 11943 5355
rect 11885 5315 11943 5321
rect 12802 5312 12808 5364
rect 12860 5352 12866 5364
rect 13173 5355 13231 5361
rect 13173 5352 13185 5355
rect 12860 5324 13185 5352
rect 12860 5312 12866 5324
rect 13173 5321 13185 5324
rect 13219 5321 13231 5355
rect 13173 5315 13231 5321
rect 13446 5312 13452 5364
rect 13504 5352 13510 5364
rect 13817 5355 13875 5361
rect 13817 5352 13829 5355
rect 13504 5324 13829 5352
rect 13504 5312 13510 5324
rect 13817 5321 13829 5324
rect 13863 5321 13875 5355
rect 13817 5315 13875 5321
rect 17221 5355 17279 5361
rect 17221 5321 17233 5355
rect 17267 5352 17279 5355
rect 17770 5352 17776 5364
rect 17267 5324 17776 5352
rect 17267 5321 17279 5324
rect 17221 5315 17279 5321
rect 17770 5312 17776 5324
rect 17828 5312 17834 5364
rect 11977 5287 12035 5293
rect 11977 5284 11989 5287
rect 7800 5256 8064 5284
rect 8220 5256 11989 5284
rect 7800 5244 7806 5256
rect 8220 5216 8248 5256
rect 11977 5253 11989 5256
rect 12023 5253 12035 5287
rect 11977 5247 12035 5253
rect 12526 5244 12532 5296
rect 12584 5284 12590 5296
rect 17034 5284 17040 5296
rect 12584 5256 17040 5284
rect 12584 5244 12590 5256
rect 7116 5188 8248 5216
rect 8297 5219 8355 5225
rect 6733 5179 6791 5185
rect 8297 5185 8309 5219
rect 8343 5216 8355 5219
rect 8757 5219 8815 5225
rect 8757 5216 8769 5219
rect 8343 5188 8769 5216
rect 8343 5185 8355 5188
rect 8297 5179 8355 5185
rect 8757 5185 8769 5188
rect 8803 5185 8815 5219
rect 9769 5219 9827 5225
rect 9769 5216 9781 5219
rect 8757 5179 8815 5185
rect 9324 5188 9781 5216
rect 9324 5160 9352 5188
rect 9769 5185 9781 5188
rect 9815 5185 9827 5219
rect 9769 5179 9827 5185
rect 9950 5176 9956 5228
rect 10008 5216 10014 5228
rect 10597 5219 10655 5225
rect 10597 5216 10609 5219
rect 10008 5188 10609 5216
rect 10008 5176 10014 5188
rect 10597 5185 10609 5188
rect 10643 5185 10655 5219
rect 10597 5179 10655 5185
rect 12066 5176 12072 5228
rect 12124 5216 12130 5228
rect 12250 5216 12256 5228
rect 12124 5188 12256 5216
rect 12124 5176 12130 5188
rect 12250 5176 12256 5188
rect 12308 5216 12314 5228
rect 12805 5219 12863 5225
rect 12805 5216 12817 5219
rect 12308 5188 12817 5216
rect 12308 5176 12314 5188
rect 12805 5185 12817 5188
rect 12851 5185 12863 5219
rect 12805 5179 12863 5185
rect 13265 5219 13323 5225
rect 13265 5185 13277 5219
rect 13311 5185 13323 5219
rect 13265 5179 13323 5185
rect 2038 5148 2044 5160
rect 1999 5120 2044 5148
rect 2038 5108 2044 5120
rect 2096 5108 2102 5160
rect 3786 5148 3792 5160
rect 3747 5120 3792 5148
rect 3786 5108 3792 5120
rect 3844 5108 3850 5160
rect 4525 5151 4583 5157
rect 4525 5117 4537 5151
rect 4571 5148 4583 5151
rect 4706 5148 4712 5160
rect 4571 5120 4712 5148
rect 4571 5117 4583 5120
rect 4525 5111 4583 5117
rect 4706 5108 4712 5120
rect 4764 5108 4770 5160
rect 5261 5151 5319 5157
rect 5261 5117 5273 5151
rect 5307 5117 5319 5151
rect 5261 5111 5319 5117
rect 5445 5151 5503 5157
rect 5445 5117 5457 5151
rect 5491 5117 5503 5151
rect 5994 5148 6000 5160
rect 5955 5120 6000 5148
rect 5445 5111 5503 5117
rect 2593 5083 2651 5089
rect 2593 5049 2605 5083
rect 2639 5080 2651 5083
rect 4246 5080 4252 5092
rect 2639 5052 4252 5080
rect 2639 5049 2651 5052
rect 2593 5043 2651 5049
rect 4246 5040 4252 5052
rect 4304 5040 4310 5092
rect 5166 5040 5172 5092
rect 5224 5080 5230 5092
rect 5276 5080 5304 5111
rect 5224 5052 5304 5080
rect 5224 5040 5230 5052
rect 4062 5012 4068 5024
rect 4023 4984 4068 5012
rect 4062 4972 4068 4984
rect 4120 4972 4126 5024
rect 4154 4972 4160 5024
rect 4212 5012 4218 5024
rect 5460 5012 5488 5111
rect 5994 5108 6000 5120
rect 6052 5108 6058 5160
rect 6549 5151 6607 5157
rect 6549 5117 6561 5151
rect 6595 5148 6607 5151
rect 7558 5148 7564 5160
rect 6595 5120 7564 5148
rect 6595 5117 6607 5120
rect 6549 5111 6607 5117
rect 7558 5108 7564 5120
rect 7616 5108 7622 5160
rect 8478 5148 8484 5160
rect 8439 5120 8484 5148
rect 8478 5108 8484 5120
rect 8536 5108 8542 5160
rect 9306 5108 9312 5160
rect 9364 5108 9370 5160
rect 9493 5151 9551 5157
rect 9493 5117 9505 5151
rect 9539 5117 9551 5151
rect 10318 5148 10324 5160
rect 10279 5120 10324 5148
rect 9493 5111 9551 5117
rect 5905 5083 5963 5089
rect 5905 5049 5917 5083
rect 5951 5080 5963 5083
rect 7374 5080 7380 5092
rect 5951 5052 7380 5080
rect 5951 5049 5963 5052
rect 5905 5043 5963 5049
rect 7374 5040 7380 5052
rect 7432 5040 7438 5092
rect 7742 5080 7748 5092
rect 7703 5052 7748 5080
rect 7742 5040 7748 5052
rect 7800 5040 7806 5092
rect 8294 5040 8300 5092
rect 8352 5080 8358 5092
rect 8846 5080 8852 5092
rect 8352 5052 8852 5080
rect 8352 5040 8358 5052
rect 8846 5040 8852 5052
rect 8904 5040 8910 5092
rect 9508 5080 9536 5111
rect 10318 5108 10324 5120
rect 10376 5108 10382 5160
rect 10502 5148 10508 5160
rect 10463 5120 10508 5148
rect 10502 5108 10508 5120
rect 10560 5108 10566 5160
rect 11790 5148 11796 5160
rect 11751 5120 11796 5148
rect 11790 5108 11796 5120
rect 11848 5108 11854 5160
rect 12526 5148 12532 5160
rect 12487 5120 12532 5148
rect 12526 5108 12532 5120
rect 12584 5108 12590 5160
rect 12618 5108 12624 5160
rect 12676 5148 12682 5160
rect 12713 5151 12771 5157
rect 12713 5148 12725 5151
rect 12676 5120 12725 5148
rect 12676 5108 12682 5120
rect 12713 5117 12725 5120
rect 12759 5117 12771 5151
rect 12713 5111 12771 5117
rect 11149 5083 11207 5089
rect 11149 5080 11161 5083
rect 8956 5052 11161 5080
rect 5626 5012 5632 5024
rect 4212 4984 5632 5012
rect 4212 4972 4218 4984
rect 5626 4972 5632 4984
rect 5684 4972 5690 5024
rect 8478 4972 8484 5024
rect 8536 5012 8542 5024
rect 8956 5012 8984 5052
rect 11149 5049 11161 5052
rect 11195 5080 11207 5083
rect 12158 5080 12164 5092
rect 11195 5052 12164 5080
rect 11195 5049 11207 5052
rect 11149 5043 11207 5049
rect 12158 5040 12164 5052
rect 12216 5040 12222 5092
rect 12345 5083 12403 5089
rect 12345 5049 12357 5083
rect 12391 5080 12403 5083
rect 13280 5080 13308 5179
rect 15194 5176 15200 5228
rect 15252 5216 15258 5228
rect 15381 5219 15439 5225
rect 15381 5216 15393 5219
rect 15252 5188 15393 5216
rect 15252 5176 15258 5188
rect 15381 5185 15393 5188
rect 15427 5185 15439 5219
rect 15381 5179 15439 5185
rect 13446 5148 13452 5160
rect 13407 5120 13452 5148
rect 13446 5108 13452 5120
rect 13504 5108 13510 5160
rect 15470 5148 15476 5160
rect 15431 5120 15476 5148
rect 15470 5108 15476 5120
rect 15528 5108 15534 5160
rect 15580 5157 15608 5256
rect 17034 5244 17040 5256
rect 17092 5244 17098 5296
rect 15838 5216 15844 5228
rect 15799 5188 15844 5216
rect 15838 5176 15844 5188
rect 15896 5176 15902 5228
rect 20622 5216 20628 5228
rect 20583 5188 20628 5216
rect 20622 5176 20628 5188
rect 20680 5176 20686 5228
rect 15565 5151 15623 5157
rect 15565 5117 15577 5151
rect 15611 5117 15623 5151
rect 15565 5111 15623 5117
rect 16117 5151 16175 5157
rect 16117 5117 16129 5151
rect 16163 5148 16175 5151
rect 17034 5148 17040 5160
rect 16163 5120 17040 5148
rect 16163 5117 16175 5120
rect 16117 5111 16175 5117
rect 17034 5108 17040 5120
rect 17092 5108 17098 5160
rect 20898 5148 20904 5160
rect 20859 5120 20904 5148
rect 20898 5108 20904 5120
rect 20956 5108 20962 5160
rect 12391 5052 13308 5080
rect 12391 5049 12403 5052
rect 12345 5043 12403 5049
rect 8536 4984 8984 5012
rect 8536 4972 8542 4984
rect 9306 4972 9312 5024
rect 9364 5012 9370 5024
rect 9364 4984 9409 5012
rect 9364 4972 9370 4984
rect 12526 4972 12532 5024
rect 12584 5012 12590 5024
rect 13354 5012 13360 5024
rect 12584 4984 13360 5012
rect 12584 4972 12590 4984
rect 13354 4972 13360 4984
rect 13412 4972 13418 5024
rect 14826 4972 14832 5024
rect 14884 5012 14890 5024
rect 15013 5015 15071 5021
rect 15013 5012 15025 5015
rect 14884 4984 15025 5012
rect 14884 4972 14890 4984
rect 15013 4981 15025 4984
rect 15059 4981 15071 5015
rect 15013 4975 15071 4981
rect 1104 4922 21896 4944
rect 1104 4870 3549 4922
rect 3601 4870 3613 4922
rect 3665 4870 3677 4922
rect 3729 4870 3741 4922
rect 3793 4870 3805 4922
rect 3857 4870 8747 4922
rect 8799 4870 8811 4922
rect 8863 4870 8875 4922
rect 8927 4870 8939 4922
rect 8991 4870 9003 4922
rect 9055 4870 13945 4922
rect 13997 4870 14009 4922
rect 14061 4870 14073 4922
rect 14125 4870 14137 4922
rect 14189 4870 14201 4922
rect 14253 4870 19143 4922
rect 19195 4870 19207 4922
rect 19259 4870 19271 4922
rect 19323 4870 19335 4922
rect 19387 4870 19399 4922
rect 19451 4870 21896 4922
rect 1104 4848 21896 4870
rect 4709 4811 4767 4817
rect 4709 4777 4721 4811
rect 4755 4808 4767 4811
rect 4890 4808 4896 4820
rect 4755 4780 4896 4808
rect 4755 4777 4767 4780
rect 4709 4771 4767 4777
rect 4890 4768 4896 4780
rect 4948 4768 4954 4820
rect 5810 4808 5816 4820
rect 5771 4780 5816 4808
rect 5810 4768 5816 4780
rect 5868 4768 5874 4820
rect 5902 4768 5908 4820
rect 5960 4808 5966 4820
rect 6273 4811 6331 4817
rect 6273 4808 6285 4811
rect 5960 4780 6285 4808
rect 5960 4768 5966 4780
rect 6273 4777 6285 4780
rect 6319 4777 6331 4811
rect 7098 4808 7104 4820
rect 7059 4780 7104 4808
rect 6273 4771 6331 4777
rect 7098 4768 7104 4780
rect 7156 4768 7162 4820
rect 7926 4768 7932 4820
rect 7984 4808 7990 4820
rect 8665 4811 8723 4817
rect 8665 4808 8677 4811
rect 7984 4780 8677 4808
rect 7984 4768 7990 4780
rect 8665 4777 8677 4780
rect 8711 4808 8723 4811
rect 8754 4808 8760 4820
rect 8711 4780 8760 4808
rect 8711 4777 8723 4780
rect 8665 4771 8723 4777
rect 8754 4768 8760 4780
rect 8812 4768 8818 4820
rect 9030 4768 9036 4820
rect 9088 4808 9094 4820
rect 9769 4811 9827 4817
rect 9769 4808 9781 4811
rect 9088 4780 9781 4808
rect 9088 4768 9094 4780
rect 9769 4777 9781 4780
rect 9815 4777 9827 4811
rect 9769 4771 9827 4777
rect 10410 4768 10416 4820
rect 10468 4808 10474 4820
rect 10597 4811 10655 4817
rect 10597 4808 10609 4811
rect 10468 4780 10609 4808
rect 10468 4768 10474 4780
rect 10597 4777 10609 4780
rect 10643 4777 10655 4811
rect 10597 4771 10655 4777
rect 12250 4768 12256 4820
rect 12308 4808 12314 4820
rect 15470 4808 15476 4820
rect 12308 4780 12353 4808
rect 15431 4780 15476 4808
rect 12308 4768 12314 4780
rect 15470 4768 15476 4780
rect 15528 4768 15534 4820
rect 16942 4808 16948 4820
rect 16903 4780 16948 4808
rect 16942 4768 16948 4780
rect 17000 4768 17006 4820
rect 18049 4811 18107 4817
rect 18049 4777 18061 4811
rect 18095 4808 18107 4811
rect 20254 4808 20260 4820
rect 18095 4780 20260 4808
rect 18095 4777 18107 4780
rect 18049 4771 18107 4777
rect 20254 4768 20260 4780
rect 20312 4768 20318 4820
rect 3418 4700 3424 4752
rect 3476 4740 3482 4752
rect 7561 4743 7619 4749
rect 7561 4740 7573 4743
rect 3476 4712 7573 4740
rect 3476 4700 3482 4712
rect 7561 4709 7573 4712
rect 7607 4740 7619 4743
rect 8481 4743 8539 4749
rect 7607 4712 8064 4740
rect 7607 4709 7619 4712
rect 7561 4703 7619 4709
rect 5258 4672 5264 4684
rect 5219 4644 5264 4672
rect 5258 4632 5264 4644
rect 5316 4632 5322 4684
rect 5905 4675 5963 4681
rect 5905 4641 5917 4675
rect 5951 4672 5963 4675
rect 6546 4672 6552 4684
rect 5951 4644 6552 4672
rect 5951 4641 5963 4644
rect 5905 4635 5963 4641
rect 6546 4632 6552 4644
rect 6604 4672 6610 4684
rect 6730 4672 6736 4684
rect 6604 4644 6736 4672
rect 6604 4632 6610 4644
rect 6730 4632 6736 4644
rect 6788 4632 6794 4684
rect 6917 4675 6975 4681
rect 6917 4641 6929 4675
rect 6963 4672 6975 4675
rect 7098 4672 7104 4684
rect 6963 4644 7104 4672
rect 6963 4641 6975 4644
rect 6917 4635 6975 4641
rect 7098 4632 7104 4644
rect 7156 4632 7162 4684
rect 7926 4672 7932 4684
rect 7887 4644 7932 4672
rect 7926 4632 7932 4644
rect 7984 4632 7990 4684
rect 8036 4681 8064 4712
rect 8481 4709 8493 4743
rect 8527 4740 8539 4743
rect 11425 4743 11483 4749
rect 8527 4712 10548 4740
rect 8527 4709 8539 4712
rect 8481 4703 8539 4709
rect 8021 4675 8079 4681
rect 8021 4641 8033 4675
rect 8067 4672 8079 4675
rect 9677 4675 9735 4681
rect 9677 4672 9689 4675
rect 8067 4644 9689 4672
rect 8067 4641 8079 4644
rect 8021 4635 8079 4641
rect 9677 4641 9689 4644
rect 9723 4672 9735 4675
rect 10134 4672 10140 4684
rect 9723 4644 10140 4672
rect 9723 4641 9735 4644
rect 9677 4635 9735 4641
rect 10134 4632 10140 4644
rect 10192 4672 10198 4684
rect 10229 4675 10287 4681
rect 10229 4672 10241 4675
rect 10192 4644 10241 4672
rect 10192 4632 10198 4644
rect 10229 4641 10241 4644
rect 10275 4641 10287 4675
rect 10229 4635 10287 4641
rect 10413 4675 10471 4681
rect 10413 4641 10425 4675
rect 10459 4641 10471 4675
rect 10520 4672 10548 4712
rect 11425 4709 11437 4743
rect 11471 4740 11483 4743
rect 11882 4740 11888 4752
rect 11471 4712 11888 4740
rect 11471 4709 11483 4712
rect 11425 4703 11483 4709
rect 11882 4700 11888 4712
rect 11940 4740 11946 4752
rect 13078 4740 13084 4752
rect 11940 4712 13084 4740
rect 11940 4700 11946 4712
rect 13078 4700 13084 4712
rect 13136 4700 13142 4752
rect 17586 4740 17592 4752
rect 15028 4712 17592 4740
rect 12894 4672 12900 4684
rect 10520 4644 12900 4672
rect 10413 4635 10471 4641
rect 4890 4564 4896 4616
rect 4948 4604 4954 4616
rect 5353 4607 5411 4613
rect 5353 4604 5365 4607
rect 4948 4576 5365 4604
rect 4948 4564 4954 4576
rect 5353 4573 5365 4576
rect 5399 4573 5411 4607
rect 5353 4567 5411 4573
rect 5445 4607 5503 4613
rect 5445 4573 5457 4607
rect 5491 4604 5503 4607
rect 5994 4604 6000 4616
rect 5491 4576 6000 4604
rect 5491 4573 5503 4576
rect 5445 4567 5503 4573
rect 5994 4564 6000 4576
rect 6052 4564 6058 4616
rect 7650 4564 7656 4616
rect 7708 4604 7714 4616
rect 9306 4604 9312 4616
rect 7708 4576 9312 4604
rect 7708 4564 7714 4576
rect 9306 4564 9312 4576
rect 9364 4604 9370 4616
rect 9401 4607 9459 4613
rect 9401 4604 9413 4607
rect 9364 4576 9413 4604
rect 9364 4564 9370 4576
rect 9401 4573 9413 4576
rect 9447 4604 9459 4607
rect 9447 4576 9674 4604
rect 9447 4573 9459 4576
rect 9401 4567 9459 4573
rect 4062 4496 4068 4548
rect 4120 4536 4126 4548
rect 4801 4539 4859 4545
rect 4801 4536 4813 4539
rect 4120 4508 4813 4536
rect 4120 4496 4126 4508
rect 4801 4505 4813 4508
rect 4847 4505 4859 4539
rect 4801 4499 4859 4505
rect 5626 4496 5632 4548
rect 5684 4536 5690 4548
rect 7377 4539 7435 4545
rect 7377 4536 7389 4539
rect 5684 4508 7389 4536
rect 5684 4496 5690 4508
rect 7377 4505 7389 4508
rect 7423 4536 7435 4539
rect 8113 4539 8171 4545
rect 8113 4536 8125 4539
rect 7423 4508 8125 4536
rect 7423 4505 7435 4508
rect 7377 4499 7435 4505
rect 8113 4505 8125 4508
rect 8159 4505 8171 4539
rect 8113 4499 8171 4505
rect 8294 4496 8300 4548
rect 8352 4536 8358 4548
rect 9030 4536 9036 4548
rect 8352 4508 9036 4536
rect 8352 4496 8358 4508
rect 9030 4496 9036 4508
rect 9088 4496 9094 4548
rect 9646 4536 9674 4576
rect 10318 4564 10324 4616
rect 10376 4604 10382 4616
rect 10428 4604 10456 4635
rect 12894 4632 12900 4644
rect 12952 4632 12958 4684
rect 14826 4672 14832 4684
rect 14787 4644 14832 4672
rect 14826 4632 14832 4644
rect 14884 4632 14890 4684
rect 15028 4681 15056 4712
rect 17586 4700 17592 4712
rect 17644 4700 17650 4752
rect 15013 4675 15071 4681
rect 15013 4641 15025 4675
rect 15059 4641 15071 4675
rect 16022 4672 16028 4684
rect 15983 4644 16028 4672
rect 15013 4635 15071 4641
rect 16022 4632 16028 4644
rect 16080 4632 16086 4684
rect 16393 4675 16451 4681
rect 16393 4641 16405 4675
rect 16439 4672 16451 4675
rect 17494 4672 17500 4684
rect 16439 4644 17080 4672
rect 17455 4644 17500 4672
rect 16439 4641 16451 4644
rect 16393 4635 16451 4641
rect 12161 4607 12219 4613
rect 10376 4576 10732 4604
rect 10376 4564 10382 4576
rect 10137 4539 10195 4545
rect 10137 4536 10149 4539
rect 9646 4508 10149 4536
rect 10137 4505 10149 4508
rect 10183 4505 10195 4539
rect 10137 4499 10195 4505
rect 5994 4428 6000 4480
rect 6052 4468 6058 4480
rect 6089 4471 6147 4477
rect 6089 4468 6101 4471
rect 6052 4440 6101 4468
rect 6052 4428 6058 4440
rect 6089 4437 6101 4440
rect 6135 4468 6147 4471
rect 6641 4471 6699 4477
rect 6641 4468 6653 4471
rect 6135 4440 6653 4468
rect 6135 4437 6147 4440
rect 6089 4431 6147 4437
rect 6641 4437 6653 4440
rect 6687 4437 6699 4471
rect 6641 4431 6699 4437
rect 6730 4428 6736 4480
rect 6788 4468 6794 4480
rect 9490 4468 9496 4480
rect 6788 4440 9496 4468
rect 6788 4428 6794 4440
rect 9490 4428 9496 4440
rect 9548 4428 9554 4480
rect 10704 4468 10732 4576
rect 12161 4573 12173 4607
rect 12207 4604 12219 4607
rect 12618 4604 12624 4616
rect 12207 4576 12624 4604
rect 12207 4573 12219 4576
rect 12161 4567 12219 4573
rect 12618 4564 12624 4576
rect 12676 4604 12682 4616
rect 13630 4604 13636 4616
rect 12676 4576 13636 4604
rect 12676 4564 12682 4576
rect 13630 4564 13636 4576
rect 13688 4564 13694 4616
rect 14734 4604 14740 4616
rect 14695 4576 14740 4604
rect 14734 4564 14740 4576
rect 14792 4564 14798 4616
rect 15838 4604 15844 4616
rect 15751 4576 15844 4604
rect 15838 4564 15844 4576
rect 15896 4604 15902 4616
rect 16408 4604 16436 4635
rect 15896 4576 16436 4604
rect 16853 4607 16911 4613
rect 15896 4564 15902 4576
rect 16853 4573 16865 4607
rect 16899 4604 16911 4607
rect 16942 4604 16948 4616
rect 16899 4576 16948 4604
rect 16899 4573 16911 4576
rect 16853 4567 16911 4573
rect 16942 4564 16948 4576
rect 17000 4564 17006 4616
rect 17052 4604 17080 4644
rect 17494 4632 17500 4644
rect 17552 4632 17558 4684
rect 22462 4672 22468 4684
rect 17604 4644 22468 4672
rect 17604 4604 17632 4644
rect 22462 4632 22468 4644
rect 22520 4632 22526 4684
rect 17052 4576 17632 4604
rect 19058 4564 19064 4616
rect 19116 4604 19122 4616
rect 19245 4607 19303 4613
rect 19245 4604 19257 4607
rect 19116 4576 19257 4604
rect 19116 4564 19122 4576
rect 19245 4573 19257 4576
rect 19291 4573 19303 4607
rect 19245 4567 19303 4573
rect 12250 4496 12256 4548
rect 12308 4536 12314 4548
rect 17770 4536 17776 4548
rect 12308 4508 17776 4536
rect 12308 4496 12314 4508
rect 17770 4496 17776 4508
rect 17828 4496 17834 4548
rect 19521 4539 19579 4545
rect 19521 4505 19533 4539
rect 19567 4536 19579 4539
rect 19886 4536 19892 4548
rect 19567 4508 19892 4536
rect 19567 4505 19579 4508
rect 19521 4499 19579 4505
rect 19886 4496 19892 4508
rect 19944 4496 19950 4548
rect 13170 4468 13176 4480
rect 10704 4440 13176 4468
rect 13170 4428 13176 4440
rect 13228 4428 13234 4480
rect 14366 4468 14372 4480
rect 14327 4440 14372 4468
rect 14366 4428 14372 4440
rect 14424 4428 14430 4480
rect 15930 4428 15936 4480
rect 15988 4468 15994 4480
rect 15988 4440 16033 4468
rect 15988 4428 15994 4440
rect 16390 4428 16396 4480
rect 16448 4468 16454 4480
rect 16669 4471 16727 4477
rect 16669 4468 16681 4471
rect 16448 4440 16681 4468
rect 16448 4428 16454 4440
rect 16669 4437 16681 4440
rect 16715 4437 16727 4471
rect 17218 4468 17224 4480
rect 17179 4440 17224 4468
rect 16669 4431 16727 4437
rect 17218 4428 17224 4440
rect 17276 4468 17282 4480
rect 17402 4468 17408 4480
rect 17276 4440 17408 4468
rect 17276 4428 17282 4440
rect 17402 4428 17408 4440
rect 17460 4428 17466 4480
rect 17586 4468 17592 4480
rect 17547 4440 17592 4468
rect 17586 4428 17592 4440
rect 17644 4428 17650 4480
rect 17678 4428 17684 4480
rect 17736 4468 17742 4480
rect 17736 4440 17781 4468
rect 17736 4428 17742 4440
rect 1104 4378 22056 4400
rect 1104 4326 6148 4378
rect 6200 4326 6212 4378
rect 6264 4326 6276 4378
rect 6328 4326 6340 4378
rect 6392 4326 6404 4378
rect 6456 4326 11346 4378
rect 11398 4326 11410 4378
rect 11462 4326 11474 4378
rect 11526 4326 11538 4378
rect 11590 4326 11602 4378
rect 11654 4326 16544 4378
rect 16596 4326 16608 4378
rect 16660 4326 16672 4378
rect 16724 4326 16736 4378
rect 16788 4326 16800 4378
rect 16852 4326 21742 4378
rect 21794 4326 21806 4378
rect 21858 4326 21870 4378
rect 21922 4326 21934 4378
rect 21986 4326 21998 4378
rect 22050 4326 22056 4378
rect 1104 4304 22056 4326
rect 5258 4224 5264 4276
rect 5316 4264 5322 4276
rect 7834 4264 7840 4276
rect 5316 4236 7840 4264
rect 5316 4224 5322 4236
rect 7834 4224 7840 4236
rect 7892 4224 7898 4276
rect 8941 4267 8999 4273
rect 8941 4233 8953 4267
rect 8987 4264 8999 4267
rect 9122 4264 9128 4276
rect 8987 4236 9128 4264
rect 8987 4233 8999 4236
rect 8941 4227 8999 4233
rect 9122 4224 9128 4236
rect 9180 4224 9186 4276
rect 9490 4264 9496 4276
rect 9451 4236 9496 4264
rect 9490 4224 9496 4236
rect 9548 4224 9554 4276
rect 10502 4264 10508 4276
rect 10463 4236 10508 4264
rect 10502 4224 10508 4236
rect 10560 4224 10566 4276
rect 10870 4264 10876 4276
rect 10831 4236 10876 4264
rect 10870 4224 10876 4236
rect 10928 4224 10934 4276
rect 11882 4264 11888 4276
rect 11843 4236 11888 4264
rect 11882 4224 11888 4236
rect 11940 4224 11946 4276
rect 12066 4224 12072 4276
rect 12124 4264 12130 4276
rect 12437 4267 12495 4273
rect 12437 4264 12449 4267
rect 12124 4236 12449 4264
rect 12124 4224 12130 4236
rect 12437 4233 12449 4236
rect 12483 4264 12495 4267
rect 13262 4264 13268 4276
rect 12483 4236 13268 4264
rect 12483 4233 12495 4236
rect 12437 4227 12495 4233
rect 13262 4224 13268 4236
rect 13320 4224 13326 4276
rect 17586 4264 17592 4276
rect 17547 4236 17592 4264
rect 17586 4224 17592 4236
rect 17644 4224 17650 4276
rect 5813 4199 5871 4205
rect 5813 4165 5825 4199
rect 5859 4196 5871 4199
rect 6365 4199 6423 4205
rect 6365 4196 6377 4199
rect 5859 4168 6377 4196
rect 5859 4165 5871 4168
rect 5813 4159 5871 4165
rect 6365 4165 6377 4168
rect 6411 4165 6423 4199
rect 6365 4159 6423 4165
rect 6546 4156 6552 4208
rect 6604 4196 6610 4208
rect 7193 4199 7251 4205
rect 7193 4196 7205 4199
rect 6604 4168 7205 4196
rect 6604 4156 6610 4168
rect 7193 4165 7205 4168
rect 7239 4196 7251 4199
rect 7653 4199 7711 4205
rect 7653 4196 7665 4199
rect 7239 4168 7665 4196
rect 7239 4165 7251 4168
rect 7193 4159 7251 4165
rect 7653 4165 7665 4168
rect 7699 4196 7711 4199
rect 7926 4196 7932 4208
rect 7699 4168 7932 4196
rect 7699 4165 7711 4168
rect 7653 4159 7711 4165
rect 7926 4156 7932 4168
rect 7984 4156 7990 4208
rect 8202 4156 8208 4208
rect 8260 4196 8266 4208
rect 8481 4199 8539 4205
rect 8481 4196 8493 4199
rect 8260 4168 8493 4196
rect 8260 4156 8266 4168
rect 8481 4165 8493 4168
rect 8527 4165 8539 4199
rect 8481 4159 8539 4165
rect 10045 4199 10103 4205
rect 10045 4165 10057 4199
rect 10091 4196 10103 4199
rect 10410 4196 10416 4208
rect 10091 4168 10416 4196
rect 10091 4165 10103 4168
rect 10045 4159 10103 4165
rect 10410 4156 10416 4168
rect 10468 4196 10474 4208
rect 15746 4196 15752 4208
rect 10468 4168 15752 4196
rect 10468 4156 10474 4168
rect 15746 4156 15752 4168
rect 15804 4156 15810 4208
rect 17129 4199 17187 4205
rect 17129 4196 17141 4199
rect 16960 4168 17141 4196
rect 16960 4140 16988 4168
rect 17129 4165 17141 4168
rect 17175 4165 17187 4199
rect 17129 4159 17187 4165
rect 17402 4156 17408 4208
rect 17460 4196 17466 4208
rect 17957 4199 18015 4205
rect 17957 4196 17969 4199
rect 17460 4168 17969 4196
rect 17460 4156 17466 4168
rect 17957 4165 17969 4168
rect 18003 4196 18015 4199
rect 19058 4196 19064 4208
rect 18003 4168 19064 4196
rect 18003 4165 18015 4168
rect 17957 4159 18015 4165
rect 19058 4156 19064 4168
rect 19116 4156 19122 4208
rect 3970 4088 3976 4140
rect 4028 4128 4034 4140
rect 5994 4128 6000 4140
rect 4028 4100 6000 4128
rect 4028 4088 4034 4100
rect 5994 4088 6000 4100
rect 6052 4088 6058 4140
rect 7745 4131 7803 4137
rect 7745 4097 7757 4131
rect 7791 4097 7803 4131
rect 7745 4091 7803 4097
rect 2222 4020 2228 4072
rect 2280 4060 2286 4072
rect 4154 4060 4160 4072
rect 2280 4032 4160 4060
rect 2280 4020 2286 4032
rect 4154 4020 4160 4032
rect 4212 4020 4218 4072
rect 5534 4060 5540 4072
rect 5495 4032 5540 4060
rect 5534 4020 5540 4032
rect 5592 4020 5598 4072
rect 5718 4060 5724 4072
rect 5679 4032 5724 4060
rect 5718 4020 5724 4032
rect 5776 4020 5782 4072
rect 7558 4060 7564 4072
rect 7519 4032 7564 4060
rect 7558 4020 7564 4032
rect 7616 4020 7622 4072
rect 3326 3952 3332 4004
rect 3384 3992 3390 4004
rect 5810 3992 5816 4004
rect 3384 3964 5816 3992
rect 3384 3952 3390 3964
rect 5810 3952 5816 3964
rect 5868 3952 5874 4004
rect 4614 3884 4620 3936
rect 4672 3924 4678 3936
rect 5442 3924 5448 3936
rect 4672 3896 5448 3924
rect 4672 3884 4678 3896
rect 5442 3884 5448 3896
rect 5500 3884 5506 3936
rect 6178 3924 6184 3936
rect 6139 3896 6184 3924
rect 6178 3884 6184 3896
rect 6236 3884 6242 3936
rect 6454 3884 6460 3936
rect 6512 3924 6518 3936
rect 7009 3927 7067 3933
rect 7009 3924 7021 3927
rect 6512 3896 7021 3924
rect 6512 3884 6518 3896
rect 7009 3893 7021 3896
rect 7055 3924 7067 3927
rect 7760 3924 7788 4091
rect 8570 4088 8576 4140
rect 8628 4128 8634 4140
rect 9674 4128 9680 4140
rect 8628 4100 8673 4128
rect 8772 4100 9680 4128
rect 8628 4088 8634 4100
rect 7834 4020 7840 4072
rect 7892 4060 7898 4072
rect 8389 4063 8447 4069
rect 8389 4060 8401 4063
rect 7892 4032 8401 4060
rect 7892 4020 7898 4032
rect 8389 4029 8401 4032
rect 8435 4029 8447 4063
rect 8389 4023 8447 4029
rect 8110 3992 8116 4004
rect 8071 3964 8116 3992
rect 8110 3952 8116 3964
rect 8168 3952 8174 4004
rect 8404 3992 8432 4023
rect 8772 3992 8800 4100
rect 9674 4088 9680 4100
rect 9732 4088 9738 4140
rect 10137 4131 10195 4137
rect 10137 4097 10149 4131
rect 10183 4097 10195 4131
rect 11977 4131 12035 4137
rect 11977 4128 11989 4131
rect 10137 4091 10195 4097
rect 11440 4100 11989 4128
rect 9490 4020 9496 4072
rect 9548 4060 9554 4072
rect 10152 4060 10180 4091
rect 11440 4072 11468 4100
rect 11977 4097 11989 4100
rect 12023 4128 12035 4131
rect 12023 4100 12296 4128
rect 12023 4097 12035 4100
rect 11977 4091 12035 4097
rect 10318 4060 10324 4072
rect 9548 4032 10180 4060
rect 10279 4032 10324 4060
rect 9548 4020 9554 4032
rect 8404 3964 8800 3992
rect 9214 3952 9220 4004
rect 9272 3992 9278 4004
rect 9677 3995 9735 4001
rect 9677 3992 9689 3995
rect 9272 3964 9689 3992
rect 9272 3952 9278 3964
rect 9677 3961 9689 3964
rect 9723 3961 9735 3995
rect 10152 3992 10180 4032
rect 10318 4020 10324 4032
rect 10376 4020 10382 4072
rect 10965 4063 11023 4069
rect 10965 4029 10977 4063
rect 11011 4029 11023 4063
rect 10965 4023 11023 4029
rect 10502 3992 10508 4004
rect 10152 3964 10508 3992
rect 9677 3955 9735 3961
rect 10502 3952 10508 3964
rect 10560 3952 10566 4004
rect 10980 3992 11008 4023
rect 11054 4020 11060 4072
rect 11112 4060 11118 4072
rect 11112 4032 11157 4060
rect 11112 4020 11118 4032
rect 11422 4020 11428 4072
rect 11480 4020 11486 4072
rect 12066 4060 12072 4072
rect 12027 4032 12072 4060
rect 12066 4020 12072 4032
rect 12124 4020 12130 4072
rect 11517 3995 11575 4001
rect 11517 3992 11529 3995
rect 10980 3964 11529 3992
rect 11517 3961 11529 3964
rect 11563 3961 11575 3995
rect 12268 3992 12296 4100
rect 12802 4088 12808 4140
rect 12860 4128 12866 4140
rect 13814 4128 13820 4140
rect 12860 4100 13820 4128
rect 12860 4088 12866 4100
rect 13814 4088 13820 4100
rect 13872 4088 13878 4140
rect 14366 4128 14372 4140
rect 14327 4100 14372 4128
rect 14366 4088 14372 4100
rect 14424 4088 14430 4140
rect 16393 4131 16451 4137
rect 16393 4097 16405 4131
rect 16439 4128 16451 4131
rect 16942 4128 16948 4140
rect 16439 4100 16948 4128
rect 16439 4097 16451 4100
rect 16393 4091 16451 4097
rect 16942 4088 16948 4100
rect 17000 4088 17006 4140
rect 17037 4131 17095 4137
rect 17037 4097 17049 4131
rect 17083 4128 17095 4131
rect 17083 4100 17117 4128
rect 17083 4097 17095 4100
rect 17037 4091 17095 4097
rect 14645 4063 14703 4069
rect 14645 4029 14657 4063
rect 14691 4060 14703 4063
rect 15378 4060 15384 4072
rect 14691 4032 15384 4060
rect 14691 4029 14703 4032
rect 14645 4023 14703 4029
rect 15378 4020 15384 4032
rect 15436 4020 15442 4072
rect 16209 4063 16267 4069
rect 16209 4029 16221 4063
rect 16255 4060 16267 4063
rect 17052 4060 17080 4091
rect 17862 4088 17868 4140
rect 17920 4128 17926 4140
rect 18049 4131 18107 4137
rect 18049 4128 18061 4131
rect 17920 4100 18061 4128
rect 17920 4088 17926 4100
rect 18049 4097 18061 4100
rect 18095 4097 18107 4131
rect 18049 4091 18107 4097
rect 17126 4060 17132 4072
rect 16255 4032 17132 4060
rect 16255 4029 16267 4032
rect 16209 4023 16267 4029
rect 17126 4020 17132 4032
rect 17184 4020 17190 4072
rect 17310 4060 17316 4072
rect 17271 4032 17316 4060
rect 17310 4020 17316 4032
rect 17368 4020 17374 4072
rect 18138 4020 18144 4072
rect 18196 4060 18202 4072
rect 18196 4032 18241 4060
rect 18196 4020 18202 4032
rect 14550 3992 14556 4004
rect 12268 3964 14556 3992
rect 11517 3955 11575 3961
rect 14550 3952 14556 3964
rect 14608 3952 14614 4004
rect 15930 3952 15936 4004
rect 15988 3992 15994 4004
rect 16669 3995 16727 4001
rect 16669 3992 16681 3995
rect 15988 3964 16681 3992
rect 15988 3952 15994 3964
rect 16669 3961 16681 3964
rect 16715 3961 16727 3995
rect 16669 3955 16727 3961
rect 8018 3924 8024 3936
rect 7055 3896 8024 3924
rect 7055 3893 7067 3896
rect 7009 3887 7067 3893
rect 8018 3884 8024 3896
rect 8076 3924 8082 3936
rect 8386 3924 8392 3936
rect 8076 3896 8392 3924
rect 8076 3884 8082 3896
rect 8386 3884 8392 3896
rect 8444 3884 8450 3936
rect 8570 3884 8576 3936
rect 8628 3924 8634 3936
rect 9125 3927 9183 3933
rect 9125 3924 9137 3927
rect 8628 3896 9137 3924
rect 8628 3884 8634 3896
rect 9125 3893 9137 3896
rect 9171 3924 9183 3927
rect 16022 3924 16028 3936
rect 9171 3896 16028 3924
rect 9171 3893 9183 3896
rect 9125 3887 9183 3893
rect 16022 3884 16028 3896
rect 16080 3924 16086 3936
rect 17218 3924 17224 3936
rect 16080 3896 17224 3924
rect 16080 3884 16086 3896
rect 17218 3884 17224 3896
rect 17276 3884 17282 3936
rect 1104 3834 21896 3856
rect 1104 3782 3549 3834
rect 3601 3782 3613 3834
rect 3665 3782 3677 3834
rect 3729 3782 3741 3834
rect 3793 3782 3805 3834
rect 3857 3782 8747 3834
rect 8799 3782 8811 3834
rect 8863 3782 8875 3834
rect 8927 3782 8939 3834
rect 8991 3782 9003 3834
rect 9055 3782 13945 3834
rect 13997 3782 14009 3834
rect 14061 3782 14073 3834
rect 14125 3782 14137 3834
rect 14189 3782 14201 3834
rect 14253 3782 19143 3834
rect 19195 3782 19207 3834
rect 19259 3782 19271 3834
rect 19323 3782 19335 3834
rect 19387 3782 19399 3834
rect 19451 3782 21896 3834
rect 1104 3760 21896 3782
rect 1762 3680 1768 3732
rect 1820 3720 1826 3732
rect 6089 3723 6147 3729
rect 6089 3720 6101 3723
rect 1820 3692 6101 3720
rect 1820 3680 1826 3692
rect 6089 3689 6101 3692
rect 6135 3720 6147 3723
rect 6546 3720 6552 3732
rect 6135 3692 6552 3720
rect 6135 3689 6147 3692
rect 6089 3683 6147 3689
rect 6546 3680 6552 3692
rect 6604 3680 6610 3732
rect 7742 3680 7748 3732
rect 7800 3720 7806 3732
rect 9766 3720 9772 3732
rect 7800 3692 9772 3720
rect 7800 3680 7806 3692
rect 9766 3680 9772 3692
rect 9824 3680 9830 3732
rect 10870 3720 10876 3732
rect 10831 3692 10876 3720
rect 10870 3680 10876 3692
rect 10928 3680 10934 3732
rect 11054 3680 11060 3732
rect 11112 3720 11118 3732
rect 12345 3723 12403 3729
rect 12345 3720 12357 3723
rect 11112 3692 12357 3720
rect 11112 3680 11118 3692
rect 12345 3689 12357 3692
rect 12391 3720 12403 3723
rect 15838 3720 15844 3732
rect 12391 3692 15844 3720
rect 12391 3689 12403 3692
rect 12345 3683 12403 3689
rect 15838 3680 15844 3692
rect 15896 3680 15902 3732
rect 16206 3680 16212 3732
rect 16264 3720 16270 3732
rect 17402 3720 17408 3732
rect 16264 3692 17408 3720
rect 16264 3680 16270 3692
rect 17402 3680 17408 3692
rect 17460 3680 17466 3732
rect 3142 3612 3148 3664
rect 3200 3652 3206 3664
rect 4525 3655 4583 3661
rect 4525 3652 4537 3655
rect 3200 3624 4537 3652
rect 3200 3612 3206 3624
rect 4525 3621 4537 3624
rect 4571 3621 4583 3655
rect 6454 3652 6460 3664
rect 4525 3615 4583 3621
rect 5368 3624 6460 3652
rect 4540 3516 4568 3615
rect 5261 3519 5319 3525
rect 5261 3516 5273 3519
rect 4540 3488 5273 3516
rect 5261 3485 5273 3488
rect 5307 3485 5319 3519
rect 5261 3479 5319 3485
rect 5368 3457 5396 3624
rect 6454 3612 6460 3624
rect 6512 3612 6518 3664
rect 6730 3612 6736 3664
rect 6788 3652 6794 3664
rect 7101 3655 7159 3661
rect 7101 3652 7113 3655
rect 6788 3624 7113 3652
rect 6788 3612 6794 3624
rect 7101 3621 7113 3624
rect 7147 3652 7159 3655
rect 7834 3652 7840 3664
rect 7147 3624 7840 3652
rect 7147 3621 7159 3624
rect 7101 3615 7159 3621
rect 7834 3612 7840 3624
rect 7892 3612 7898 3664
rect 8018 3652 8024 3664
rect 7979 3624 8024 3652
rect 8018 3612 8024 3624
rect 8076 3612 8082 3664
rect 10965 3655 11023 3661
rect 10965 3652 10977 3655
rect 10336 3624 10977 3652
rect 10336 3596 10364 3624
rect 10965 3621 10977 3624
rect 11011 3652 11023 3655
rect 12066 3652 12072 3664
rect 11011 3624 12072 3652
rect 11011 3621 11023 3624
rect 10965 3615 11023 3621
rect 12066 3612 12072 3624
rect 12124 3612 12130 3664
rect 17126 3612 17132 3664
rect 17184 3652 17190 3664
rect 18598 3652 18604 3664
rect 17184 3624 18604 3652
rect 17184 3612 17190 3624
rect 18598 3612 18604 3624
rect 18656 3612 18662 3664
rect 5442 3544 5448 3596
rect 5500 3584 5506 3596
rect 5500 3556 5545 3584
rect 5500 3544 5506 3556
rect 5626 3544 5632 3596
rect 5684 3584 5690 3596
rect 5902 3584 5908 3596
rect 5684 3556 5908 3584
rect 5684 3544 5690 3556
rect 5902 3544 5908 3556
rect 5960 3544 5966 3596
rect 6362 3584 6368 3596
rect 6104 3556 6368 3584
rect 5460 3516 5488 3544
rect 5721 3519 5779 3525
rect 5721 3516 5733 3519
rect 5460 3488 5733 3516
rect 5721 3485 5733 3488
rect 5767 3516 5779 3519
rect 5810 3516 5816 3528
rect 5767 3488 5816 3516
rect 5767 3485 5779 3488
rect 5721 3479 5779 3485
rect 5810 3476 5816 3488
rect 5868 3516 5874 3528
rect 6104 3516 6132 3556
rect 6362 3544 6368 3556
rect 6420 3544 6426 3596
rect 6546 3584 6552 3596
rect 6507 3556 6552 3584
rect 6546 3544 6552 3556
rect 6604 3544 6610 3596
rect 9125 3587 9183 3593
rect 9125 3553 9137 3587
rect 9171 3584 9183 3587
rect 9950 3584 9956 3596
rect 9171 3556 9956 3584
rect 9171 3553 9183 3556
rect 9125 3547 9183 3553
rect 9950 3544 9956 3556
rect 10008 3544 10014 3596
rect 10318 3584 10324 3596
rect 10231 3556 10324 3584
rect 10318 3544 10324 3556
rect 10376 3544 10382 3596
rect 10410 3544 10416 3596
rect 10468 3584 10474 3596
rect 11054 3584 11060 3596
rect 10468 3556 11060 3584
rect 10468 3544 10474 3556
rect 11054 3544 11060 3556
rect 11112 3544 11118 3596
rect 11238 3544 11244 3596
rect 11296 3584 11302 3596
rect 11517 3587 11575 3593
rect 11517 3584 11529 3587
rect 11296 3556 11529 3584
rect 11296 3544 11302 3556
rect 11517 3553 11529 3556
rect 11563 3553 11575 3587
rect 11517 3547 11575 3553
rect 13173 3587 13231 3593
rect 13173 3553 13185 3587
rect 13219 3584 13231 3587
rect 18506 3584 18512 3596
rect 13219 3556 18512 3584
rect 13219 3553 13231 3556
rect 13173 3547 13231 3553
rect 18506 3544 18512 3556
rect 18564 3544 18570 3596
rect 5868 3488 6132 3516
rect 5868 3476 5874 3488
rect 6178 3476 6184 3528
rect 6236 3516 6242 3528
rect 9309 3519 9367 3525
rect 9309 3516 9321 3519
rect 6236 3488 9321 3516
rect 6236 3476 6242 3488
rect 9309 3485 9321 3488
rect 9355 3485 9367 3519
rect 13357 3519 13415 3525
rect 13357 3516 13369 3519
rect 9309 3479 9367 3485
rect 9692 3488 13369 3516
rect 5353 3451 5411 3457
rect 5353 3448 5365 3451
rect 4724 3420 5365 3448
rect 3878 3340 3884 3392
rect 3936 3380 3942 3392
rect 4724 3389 4752 3420
rect 5353 3417 5365 3420
rect 5399 3417 5411 3451
rect 5353 3411 5411 3417
rect 5442 3408 5448 3460
rect 5500 3448 5506 3460
rect 9217 3451 9275 3457
rect 9217 3448 9229 3451
rect 5500 3420 9229 3448
rect 5500 3408 5506 3420
rect 9217 3417 9229 3420
rect 9263 3417 9275 3451
rect 9217 3411 9275 3417
rect 4709 3383 4767 3389
rect 4709 3380 4721 3383
rect 3936 3352 4721 3380
rect 3936 3340 3942 3352
rect 4709 3349 4721 3352
rect 4755 3349 4767 3383
rect 4709 3343 4767 3349
rect 4893 3383 4951 3389
rect 4893 3349 4905 3383
rect 4939 3380 4951 3383
rect 5074 3380 5080 3392
rect 4939 3352 5080 3380
rect 4939 3349 4951 3352
rect 4893 3343 4951 3349
rect 5074 3340 5080 3352
rect 5132 3340 5138 3392
rect 5902 3340 5908 3392
rect 5960 3380 5966 3392
rect 6641 3383 6699 3389
rect 6641 3380 6653 3383
rect 5960 3352 6653 3380
rect 5960 3340 5966 3352
rect 6641 3349 6653 3352
rect 6687 3349 6699 3383
rect 6641 3343 6699 3349
rect 6730 3340 6736 3392
rect 6788 3380 6794 3392
rect 9692 3389 9720 3488
rect 13357 3485 13369 3488
rect 13403 3485 13415 3519
rect 13357 3479 13415 3485
rect 13538 3476 13544 3528
rect 13596 3516 13602 3528
rect 14918 3516 14924 3528
rect 13596 3488 14924 3516
rect 13596 3476 13602 3488
rect 14918 3476 14924 3488
rect 14976 3476 14982 3528
rect 17313 3519 17371 3525
rect 17313 3485 17325 3519
rect 17359 3516 17371 3519
rect 17862 3516 17868 3528
rect 17359 3488 17868 3516
rect 17359 3485 17371 3488
rect 17313 3479 17371 3485
rect 17862 3476 17868 3488
rect 17920 3516 17926 3528
rect 18414 3516 18420 3528
rect 17920 3488 18420 3516
rect 17920 3476 17926 3488
rect 18414 3476 18420 3488
rect 18472 3476 18478 3528
rect 9766 3408 9772 3460
rect 9824 3448 9830 3460
rect 11793 3451 11851 3457
rect 11793 3448 11805 3451
rect 9824 3420 11805 3448
rect 9824 3408 9830 3420
rect 11793 3417 11805 3420
rect 11839 3417 11851 3451
rect 13265 3451 13323 3457
rect 13265 3448 13277 3451
rect 11793 3411 11851 3417
rect 12176 3420 13277 3448
rect 7009 3383 7067 3389
rect 7009 3380 7021 3383
rect 6788 3352 7021 3380
rect 6788 3340 6794 3352
rect 7009 3349 7021 3352
rect 7055 3349 7067 3383
rect 7009 3343 7067 3349
rect 9677 3383 9735 3389
rect 9677 3349 9689 3383
rect 9723 3349 9735 3383
rect 9950 3380 9956 3392
rect 9911 3352 9956 3380
rect 9677 3343 9735 3349
rect 9950 3340 9956 3352
rect 10008 3380 10014 3392
rect 10505 3383 10563 3389
rect 10505 3380 10517 3383
rect 10008 3352 10517 3380
rect 10008 3340 10014 3352
rect 10505 3349 10517 3352
rect 10551 3349 10563 3383
rect 10505 3343 10563 3349
rect 11054 3340 11060 3392
rect 11112 3380 11118 3392
rect 11149 3383 11207 3389
rect 11149 3380 11161 3383
rect 11112 3352 11161 3380
rect 11112 3340 11118 3352
rect 11149 3349 11161 3352
rect 11195 3380 11207 3383
rect 11422 3380 11428 3392
rect 11195 3352 11428 3380
rect 11195 3349 11207 3352
rect 11149 3343 11207 3349
rect 11422 3340 11428 3352
rect 11480 3340 11486 3392
rect 11698 3380 11704 3392
rect 11659 3352 11704 3380
rect 11698 3340 11704 3352
rect 11756 3340 11762 3392
rect 12176 3389 12204 3420
rect 13265 3417 13277 3420
rect 13311 3417 13323 3451
rect 13265 3411 13323 3417
rect 13630 3408 13636 3460
rect 13688 3448 13694 3460
rect 13688 3420 16252 3448
rect 13688 3408 13694 3420
rect 16224 3392 16252 3420
rect 16298 3408 16304 3460
rect 16356 3448 16362 3460
rect 20162 3448 20168 3460
rect 16356 3420 20168 3448
rect 16356 3408 16362 3420
rect 20162 3408 20168 3420
rect 20220 3408 20226 3460
rect 12161 3383 12219 3389
rect 12161 3349 12173 3383
rect 12207 3349 12219 3383
rect 13722 3380 13728 3392
rect 13683 3352 13728 3380
rect 12161 3343 12219 3349
rect 13722 3340 13728 3352
rect 13780 3340 13786 3392
rect 16206 3340 16212 3392
rect 16264 3380 16270 3392
rect 16577 3383 16635 3389
rect 16577 3380 16589 3383
rect 16264 3352 16589 3380
rect 16264 3340 16270 3352
rect 16577 3349 16589 3352
rect 16623 3349 16635 3383
rect 16577 3343 16635 3349
rect 18230 3340 18236 3392
rect 18288 3380 18294 3392
rect 21542 3380 21548 3392
rect 18288 3352 21548 3380
rect 18288 3340 18294 3352
rect 21542 3340 21548 3352
rect 21600 3340 21606 3392
rect 1104 3290 22056 3312
rect 1104 3238 6148 3290
rect 6200 3238 6212 3290
rect 6264 3238 6276 3290
rect 6328 3238 6340 3290
rect 6392 3238 6404 3290
rect 6456 3238 11346 3290
rect 11398 3238 11410 3290
rect 11462 3238 11474 3290
rect 11526 3238 11538 3290
rect 11590 3238 11602 3290
rect 11654 3238 16544 3290
rect 16596 3238 16608 3290
rect 16660 3238 16672 3290
rect 16724 3238 16736 3290
rect 16788 3238 16800 3290
rect 16852 3238 21742 3290
rect 21794 3238 21806 3290
rect 21858 3238 21870 3290
rect 21922 3238 21934 3290
rect 21986 3238 21998 3290
rect 22050 3238 22056 3290
rect 1104 3216 22056 3238
rect 5074 3176 5080 3188
rect 5035 3148 5080 3176
rect 5074 3136 5080 3148
rect 5132 3136 5138 3188
rect 5442 3176 5448 3188
rect 5403 3148 5448 3176
rect 5442 3136 5448 3148
rect 5500 3136 5506 3188
rect 6730 3176 6736 3188
rect 6691 3148 6736 3176
rect 6730 3136 6736 3148
rect 6788 3136 6794 3188
rect 7101 3179 7159 3185
rect 7101 3145 7113 3179
rect 7147 3176 7159 3179
rect 9766 3176 9772 3188
rect 7147 3148 9772 3176
rect 7147 3145 7159 3148
rect 7101 3139 7159 3145
rect 9766 3136 9772 3148
rect 9824 3136 9830 3188
rect 10045 3179 10103 3185
rect 10045 3145 10057 3179
rect 10091 3176 10103 3179
rect 10410 3176 10416 3188
rect 10091 3148 10416 3176
rect 10091 3145 10103 3148
rect 10045 3139 10103 3145
rect 10410 3136 10416 3148
rect 10468 3136 10474 3188
rect 10505 3179 10563 3185
rect 10505 3145 10517 3179
rect 10551 3176 10563 3179
rect 10965 3179 11023 3185
rect 10965 3176 10977 3179
rect 10551 3148 10977 3176
rect 10551 3145 10563 3148
rect 10505 3139 10563 3145
rect 10965 3145 10977 3148
rect 11011 3145 11023 3179
rect 10965 3139 11023 3145
rect 11333 3179 11391 3185
rect 11333 3145 11345 3179
rect 11379 3176 11391 3179
rect 11698 3176 11704 3188
rect 11379 3148 11704 3176
rect 11379 3145 11391 3148
rect 11333 3139 11391 3145
rect 11698 3136 11704 3148
rect 11756 3136 11762 3188
rect 11793 3179 11851 3185
rect 11793 3145 11805 3179
rect 11839 3176 11851 3179
rect 11974 3176 11980 3188
rect 11839 3148 11980 3176
rect 11839 3145 11851 3148
rect 11793 3139 11851 3145
rect 11974 3136 11980 3148
rect 12032 3136 12038 3188
rect 12069 3179 12127 3185
rect 12069 3145 12081 3179
rect 12115 3176 12127 3179
rect 15562 3176 15568 3188
rect 12115 3148 15568 3176
rect 12115 3145 12127 3148
rect 12069 3139 12127 3145
rect 15562 3136 15568 3148
rect 15620 3136 15626 3188
rect 15933 3179 15991 3185
rect 15933 3145 15945 3179
rect 15979 3145 15991 3179
rect 16298 3176 16304 3188
rect 16259 3148 16304 3176
rect 15933 3139 15991 3145
rect 6914 3068 6920 3120
rect 6972 3108 6978 3120
rect 7650 3108 7656 3120
rect 6972 3080 7656 3108
rect 6972 3068 6978 3080
rect 7650 3068 7656 3080
rect 7708 3068 7714 3120
rect 8570 3108 8576 3120
rect 8531 3080 8576 3108
rect 8570 3068 8576 3080
rect 8628 3068 8634 3120
rect 9217 3111 9275 3117
rect 9217 3108 9229 3111
rect 8772 3080 9229 3108
rect 5442 3000 5448 3052
rect 5500 3040 5506 3052
rect 7098 3040 7104 3052
rect 5500 3012 7104 3040
rect 5500 3000 5506 3012
rect 7098 3000 7104 3012
rect 7156 3000 7162 3052
rect 8772 3049 8800 3080
rect 9217 3077 9229 3080
rect 9263 3108 9275 3111
rect 10134 3108 10140 3120
rect 9263 3080 9674 3108
rect 10095 3080 10140 3108
rect 9263 3077 9275 3080
rect 9217 3071 9275 3077
rect 8757 3043 8815 3049
rect 8757 3040 8769 3043
rect 7760 3012 8769 3040
rect 4801 2975 4859 2981
rect 4801 2941 4813 2975
rect 4847 2941 4859 2975
rect 4982 2972 4988 2984
rect 4943 2944 4988 2972
rect 4801 2935 4859 2941
rect 382 2864 388 2916
rect 440 2904 446 2916
rect 3418 2904 3424 2916
rect 440 2876 3424 2904
rect 440 2864 446 2876
rect 3418 2864 3424 2876
rect 3476 2864 3482 2916
rect 4816 2904 4844 2935
rect 4982 2932 4988 2944
rect 5040 2932 5046 2984
rect 5534 2932 5540 2984
rect 5592 2972 5598 2984
rect 6546 2972 6552 2984
rect 5592 2944 6552 2972
rect 5592 2932 5598 2944
rect 6546 2932 6552 2944
rect 6604 2932 6610 2984
rect 6641 2975 6699 2981
rect 6641 2941 6653 2975
rect 6687 2972 6699 2975
rect 6687 2944 7328 2972
rect 6687 2941 6699 2944
rect 6641 2935 6699 2941
rect 5552 2904 5580 2932
rect 7300 2913 7328 2944
rect 7650 2932 7656 2984
rect 7708 2972 7714 2984
rect 7760 2981 7788 3012
rect 8757 3009 8769 3012
rect 8803 3009 8815 3043
rect 9306 3040 9312 3052
rect 9267 3012 9312 3040
rect 8757 3003 8815 3009
rect 9306 3000 9312 3012
rect 9364 3000 9370 3052
rect 7745 2975 7803 2981
rect 7745 2972 7757 2975
rect 7708 2944 7757 2972
rect 7708 2932 7714 2944
rect 7745 2941 7757 2944
rect 7791 2941 7803 2975
rect 7745 2935 7803 2941
rect 7834 2932 7840 2984
rect 7892 2972 7898 2984
rect 8113 2975 8171 2981
rect 8113 2972 8125 2975
rect 7892 2944 8125 2972
rect 7892 2932 7898 2944
rect 8113 2941 8125 2944
rect 8159 2972 8171 2975
rect 8159 2944 8708 2972
rect 8159 2941 8171 2944
rect 8113 2935 8171 2941
rect 4816 2876 5580 2904
rect 7285 2907 7343 2913
rect 7285 2873 7297 2907
rect 7331 2873 7343 2907
rect 8680 2904 8708 2944
rect 9122 2932 9128 2984
rect 9180 2972 9186 2984
rect 9646 2972 9674 3080
rect 10134 3068 10140 3080
rect 10192 3068 10198 3120
rect 11054 3068 11060 3120
rect 11112 3108 11118 3120
rect 11517 3111 11575 3117
rect 11517 3108 11529 3111
rect 11112 3080 11529 3108
rect 11112 3068 11118 3080
rect 11517 3077 11529 3080
rect 11563 3108 11575 3111
rect 12713 3111 12771 3117
rect 12713 3108 12725 3111
rect 11563 3080 12434 3108
rect 11563 3077 11575 3080
rect 11517 3071 11575 3077
rect 9950 3040 9956 3052
rect 9784 3012 9956 3040
rect 9784 2972 9812 3012
rect 9950 3000 9956 3012
rect 10008 3000 10014 3052
rect 10502 3000 10508 3052
rect 10560 3040 10566 3052
rect 11790 3040 11796 3052
rect 10560 3012 11796 3040
rect 10560 3000 10566 3012
rect 11790 3000 11796 3012
rect 11848 3040 11854 3052
rect 11885 3043 11943 3049
rect 11885 3040 11897 3043
rect 11848 3012 11897 3040
rect 11848 3000 11854 3012
rect 11885 3009 11897 3012
rect 11931 3009 11943 3043
rect 11885 3003 11943 3009
rect 11974 3000 11980 3052
rect 12032 3040 12038 3052
rect 12406 3040 12434 3080
rect 12544 3080 12725 3108
rect 12544 3040 12572 3080
rect 12713 3077 12725 3080
rect 12759 3108 12771 3111
rect 15948 3108 15976 3139
rect 16298 3136 16304 3148
rect 16356 3136 16362 3188
rect 17862 3136 17868 3188
rect 17920 3176 17926 3188
rect 18601 3179 18659 3185
rect 18601 3176 18613 3179
rect 17920 3148 18613 3176
rect 17920 3136 17926 3148
rect 18601 3145 18613 3148
rect 18647 3145 18659 3179
rect 18601 3139 18659 3145
rect 18782 3136 18788 3188
rect 18840 3176 18846 3188
rect 19242 3176 19248 3188
rect 18840 3148 19248 3176
rect 18840 3136 18846 3148
rect 19242 3136 19248 3148
rect 19300 3136 19306 3188
rect 19337 3179 19395 3185
rect 19337 3145 19349 3179
rect 19383 3145 19395 3179
rect 19337 3139 19395 3145
rect 19352 3108 19380 3139
rect 19426 3136 19432 3188
rect 19484 3176 19490 3188
rect 20717 3179 20775 3185
rect 20717 3176 20729 3179
rect 19484 3148 20729 3176
rect 19484 3136 19490 3148
rect 20717 3145 20729 3148
rect 20763 3145 20775 3179
rect 20717 3139 20775 3145
rect 22094 3108 22100 3120
rect 12759 3080 14964 3108
rect 15948 3080 19288 3108
rect 19352 3080 22100 3108
rect 12759 3077 12771 3080
rect 12713 3071 12771 3077
rect 14936 3052 14964 3080
rect 12032 3012 12296 3040
rect 12406 3012 12572 3040
rect 12621 3043 12679 3049
rect 12032 3000 12038 3012
rect 9180 2944 9225 2972
rect 9646 2944 9812 2972
rect 9861 2975 9919 2981
rect 9180 2932 9186 2944
rect 9861 2941 9873 2975
rect 9907 2941 9919 2975
rect 9861 2935 9919 2941
rect 9674 2904 9680 2916
rect 8680 2876 8800 2904
rect 9635 2876 9680 2904
rect 7285 2867 7343 2873
rect 8772 2836 8800 2876
rect 9674 2864 9680 2876
rect 9732 2864 9738 2916
rect 9876 2904 9904 2935
rect 10594 2932 10600 2984
rect 10652 2972 10658 2984
rect 10689 2975 10747 2981
rect 10689 2972 10701 2975
rect 10652 2944 10701 2972
rect 10652 2932 10658 2944
rect 10689 2941 10701 2944
rect 10735 2941 10747 2975
rect 10689 2935 10747 2941
rect 10873 2975 10931 2981
rect 10873 2941 10885 2975
rect 10919 2972 10931 2975
rect 12268 2972 12296 3012
rect 12621 3009 12633 3043
rect 12667 3040 12679 3043
rect 13446 3040 13452 3052
rect 12667 3012 13317 3040
rect 13407 3012 13452 3040
rect 12667 3009 12679 3012
rect 12621 3003 12679 3009
rect 12636 2972 12664 3003
rect 10919 2944 12204 2972
rect 12268 2944 12664 2972
rect 12897 2975 12955 2981
rect 10919 2941 10931 2944
rect 10873 2935 10931 2941
rect 9784 2876 9904 2904
rect 12176 2904 12204 2944
rect 12897 2941 12909 2975
rect 12943 2972 12955 2975
rect 13170 2972 13176 2984
rect 12943 2944 13176 2972
rect 12943 2941 12955 2944
rect 12897 2935 12955 2941
rect 12253 2907 12311 2913
rect 12253 2904 12265 2907
rect 12176 2876 12265 2904
rect 9784 2836 9812 2876
rect 12253 2873 12265 2876
rect 12299 2873 12311 2907
rect 12253 2867 12311 2873
rect 10870 2836 10876 2848
rect 8772 2808 10876 2836
rect 10870 2796 10876 2808
rect 10928 2836 10934 2848
rect 12912 2836 12940 2935
rect 13170 2932 13176 2944
rect 13228 2932 13234 2984
rect 13289 2904 13317 3012
rect 13446 3000 13452 3012
rect 13504 3000 13510 3052
rect 13538 3000 13544 3052
rect 13596 3040 13602 3052
rect 13722 3040 13728 3052
rect 13596 3012 13641 3040
rect 13683 3012 13728 3040
rect 13596 3000 13602 3012
rect 13722 3000 13728 3012
rect 13780 3000 13786 3052
rect 14274 3040 14280 3052
rect 14235 3012 14280 3040
rect 14274 3000 14280 3012
rect 14332 3000 14338 3052
rect 14550 3000 14556 3052
rect 14608 3040 14614 3052
rect 14645 3043 14703 3049
rect 14645 3040 14657 3043
rect 14608 3012 14657 3040
rect 14608 3000 14614 3012
rect 14645 3009 14657 3012
rect 14691 3009 14703 3043
rect 14645 3003 14703 3009
rect 14918 3000 14924 3052
rect 14976 3040 14982 3052
rect 15013 3043 15071 3049
rect 15013 3040 15025 3043
rect 14976 3012 15025 3040
rect 14976 3000 14982 3012
rect 15013 3009 15025 3012
rect 15059 3009 15071 3043
rect 15378 3040 15384 3052
rect 15339 3012 15384 3040
rect 15013 3003 15071 3009
rect 15378 3000 15384 3012
rect 15436 3000 15442 3052
rect 15746 3040 15752 3052
rect 15707 3012 15752 3040
rect 15746 3000 15752 3012
rect 15804 3000 15810 3052
rect 16117 3043 16175 3049
rect 16117 3009 16129 3043
rect 16163 3009 16175 3043
rect 16117 3003 16175 3009
rect 13814 2932 13820 2984
rect 13872 2972 13878 2984
rect 13909 2975 13967 2981
rect 13909 2972 13921 2975
rect 13872 2944 13921 2972
rect 13872 2932 13878 2944
rect 13909 2941 13921 2944
rect 13955 2941 13967 2975
rect 15930 2972 15936 2984
rect 13909 2935 13967 2941
rect 15028 2944 15936 2972
rect 15028 2904 15056 2944
rect 15930 2932 15936 2944
rect 15988 2972 15994 2984
rect 16132 2972 16160 3003
rect 16206 3000 16212 3052
rect 16264 3040 16270 3052
rect 16669 3043 16727 3049
rect 16669 3040 16681 3043
rect 16264 3012 16681 3040
rect 16264 3000 16270 3012
rect 16669 3009 16681 3012
rect 16715 3009 16727 3043
rect 17034 3040 17040 3052
rect 16995 3012 17040 3040
rect 16669 3003 16727 3009
rect 17034 3000 17040 3012
rect 17092 3000 17098 3052
rect 17770 3000 17776 3052
rect 17828 3040 17834 3052
rect 17957 3043 18015 3049
rect 17957 3040 17969 3043
rect 17828 3012 17969 3040
rect 17828 3000 17834 3012
rect 17957 3009 17969 3012
rect 18003 3040 18015 3043
rect 18049 3043 18107 3049
rect 18049 3040 18061 3043
rect 18003 3012 18061 3040
rect 18003 3009 18015 3012
rect 17957 3003 18015 3009
rect 18049 3009 18061 3012
rect 18095 3009 18107 3043
rect 18414 3040 18420 3052
rect 18375 3012 18420 3040
rect 18049 3003 18107 3009
rect 18414 3000 18420 3012
rect 18472 3000 18478 3052
rect 18598 3000 18604 3052
rect 18656 3040 18662 3052
rect 18785 3043 18843 3049
rect 18785 3040 18797 3043
rect 18656 3012 18797 3040
rect 18656 3000 18662 3012
rect 18785 3009 18797 3012
rect 18831 3009 18843 3043
rect 18785 3003 18843 3009
rect 19058 3000 19064 3052
rect 19116 3040 19122 3052
rect 19153 3043 19211 3049
rect 19153 3040 19165 3043
rect 19116 3012 19165 3040
rect 19116 3000 19122 3012
rect 19153 3009 19165 3012
rect 19199 3009 19211 3043
rect 19260 3040 19288 3080
rect 22094 3068 22100 3080
rect 22152 3068 22158 3120
rect 19518 3040 19524 3052
rect 19260 3012 19524 3040
rect 19153 3003 19211 3009
rect 19518 3000 19524 3012
rect 19576 3000 19582 3052
rect 19610 3000 19616 3052
rect 19668 3040 19674 3052
rect 19705 3043 19763 3049
rect 19705 3040 19717 3043
rect 19668 3012 19717 3040
rect 19668 3000 19674 3012
rect 19705 3009 19717 3012
rect 19751 3009 19763 3043
rect 19886 3040 19892 3052
rect 19847 3012 19892 3040
rect 19705 3003 19763 3009
rect 19886 3000 19892 3012
rect 19944 3000 19950 3052
rect 19978 3000 19984 3052
rect 20036 3040 20042 3052
rect 20257 3043 20315 3049
rect 20257 3040 20269 3043
rect 20036 3012 20269 3040
rect 20036 3000 20042 3012
rect 20257 3009 20269 3012
rect 20303 3009 20315 3043
rect 20898 3040 20904 3052
rect 20859 3012 20904 3040
rect 20257 3003 20315 3009
rect 20898 3000 20904 3012
rect 20956 3000 20962 3052
rect 21082 2972 21088 2984
rect 15988 2944 16160 2972
rect 18984 2944 21088 2972
rect 15988 2932 15994 2944
rect 13289 2876 15056 2904
rect 15102 2864 15108 2916
rect 15160 2904 15166 2916
rect 15565 2907 15623 2913
rect 15565 2904 15577 2907
rect 15160 2876 15577 2904
rect 15160 2864 15166 2876
rect 15565 2873 15577 2876
rect 15611 2873 15623 2907
rect 16022 2904 16028 2916
rect 15565 2867 15623 2873
rect 15856 2876 16028 2904
rect 13262 2836 13268 2848
rect 10928 2808 12940 2836
rect 13223 2808 13268 2836
rect 10928 2796 10934 2808
rect 13262 2796 13268 2808
rect 13320 2796 13326 2848
rect 13722 2796 13728 2848
rect 13780 2836 13786 2848
rect 14461 2839 14519 2845
rect 14461 2836 14473 2839
rect 13780 2808 14473 2836
rect 13780 2796 13786 2808
rect 14461 2805 14473 2808
rect 14507 2805 14519 2839
rect 14461 2799 14519 2805
rect 14642 2796 14648 2848
rect 14700 2836 14706 2848
rect 14829 2839 14887 2845
rect 14829 2836 14841 2839
rect 14700 2808 14841 2836
rect 14700 2796 14706 2808
rect 14829 2805 14841 2808
rect 14875 2805 14887 2839
rect 14829 2799 14887 2805
rect 15197 2839 15255 2845
rect 15197 2805 15209 2839
rect 15243 2836 15255 2839
rect 15856 2836 15884 2876
rect 16022 2864 16028 2876
rect 16080 2864 16086 2916
rect 16853 2907 16911 2913
rect 16853 2873 16865 2907
rect 16899 2904 16911 2907
rect 17402 2904 17408 2916
rect 16899 2876 17408 2904
rect 16899 2873 16911 2876
rect 16853 2867 16911 2873
rect 17402 2864 17408 2876
rect 17460 2864 17466 2916
rect 18230 2904 18236 2916
rect 18191 2876 18236 2904
rect 18230 2864 18236 2876
rect 18288 2864 18294 2916
rect 18984 2913 19012 2944
rect 21082 2932 21088 2944
rect 21140 2932 21146 2984
rect 18969 2907 19027 2913
rect 18969 2873 18981 2907
rect 19015 2873 19027 2907
rect 18969 2867 19027 2873
rect 19058 2864 19064 2916
rect 19116 2904 19122 2916
rect 20073 2907 20131 2913
rect 19116 2876 19840 2904
rect 19116 2864 19122 2876
rect 15243 2808 15884 2836
rect 15243 2805 15255 2808
rect 15197 2799 15255 2805
rect 16942 2796 16948 2848
rect 17000 2836 17006 2848
rect 17221 2839 17279 2845
rect 17221 2836 17233 2839
rect 17000 2808 17233 2836
rect 17000 2796 17006 2808
rect 17221 2805 17233 2808
rect 17267 2805 17279 2839
rect 17221 2799 17279 2805
rect 19150 2796 19156 2848
rect 19208 2836 19214 2848
rect 19521 2839 19579 2845
rect 19521 2836 19533 2839
rect 19208 2808 19533 2836
rect 19208 2796 19214 2808
rect 19521 2805 19533 2808
rect 19567 2805 19579 2839
rect 19812 2836 19840 2876
rect 20073 2873 20085 2907
rect 20119 2904 20131 2907
rect 20622 2904 20628 2916
rect 20119 2876 20628 2904
rect 20119 2873 20131 2876
rect 20073 2867 20131 2873
rect 20622 2864 20628 2876
rect 20680 2864 20686 2916
rect 20441 2839 20499 2845
rect 20441 2836 20453 2839
rect 19812 2808 20453 2836
rect 19521 2799 19579 2805
rect 20441 2805 20453 2808
rect 20487 2805 20499 2839
rect 20441 2799 20499 2805
rect 1104 2746 21896 2768
rect 1104 2694 3549 2746
rect 3601 2694 3613 2746
rect 3665 2694 3677 2746
rect 3729 2694 3741 2746
rect 3793 2694 3805 2746
rect 3857 2694 8747 2746
rect 8799 2694 8811 2746
rect 8863 2694 8875 2746
rect 8927 2694 8939 2746
rect 8991 2694 9003 2746
rect 9055 2694 13945 2746
rect 13997 2694 14009 2746
rect 14061 2694 14073 2746
rect 14125 2694 14137 2746
rect 14189 2694 14201 2746
rect 14253 2694 19143 2746
rect 19195 2694 19207 2746
rect 19259 2694 19271 2746
rect 19323 2694 19335 2746
rect 19387 2694 19399 2746
rect 19451 2694 21896 2746
rect 1104 2672 21896 2694
rect 4982 2632 4988 2644
rect 4943 2604 4988 2632
rect 4982 2592 4988 2604
rect 5040 2592 5046 2644
rect 5810 2632 5816 2644
rect 5771 2604 5816 2632
rect 5810 2592 5816 2604
rect 5868 2592 5874 2644
rect 8110 2592 8116 2644
rect 8168 2632 8174 2644
rect 8941 2635 8999 2641
rect 8941 2632 8953 2635
rect 8168 2604 8953 2632
rect 8168 2592 8174 2604
rect 8941 2601 8953 2604
rect 8987 2601 8999 2635
rect 8941 2595 8999 2601
rect 9861 2635 9919 2641
rect 9861 2601 9873 2635
rect 9907 2632 9919 2635
rect 10134 2632 10140 2644
rect 9907 2604 10140 2632
rect 9907 2601 9919 2604
rect 9861 2595 9919 2601
rect 10134 2592 10140 2604
rect 10192 2592 10198 2644
rect 10410 2592 10416 2644
rect 10468 2632 10474 2644
rect 10597 2635 10655 2641
rect 10597 2632 10609 2635
rect 10468 2604 10609 2632
rect 10468 2592 10474 2604
rect 10597 2601 10609 2604
rect 10643 2601 10655 2635
rect 10870 2632 10876 2644
rect 10831 2604 10876 2632
rect 10597 2595 10655 2601
rect 10870 2592 10876 2604
rect 10928 2592 10934 2644
rect 11790 2632 11796 2644
rect 11751 2604 11796 2632
rect 11790 2592 11796 2604
rect 11848 2592 11854 2644
rect 14550 2632 14556 2644
rect 14511 2604 14556 2632
rect 14550 2592 14556 2604
rect 14608 2592 14614 2644
rect 14918 2632 14924 2644
rect 14879 2604 14924 2632
rect 14918 2592 14924 2604
rect 14976 2592 14982 2644
rect 15657 2635 15715 2641
rect 15657 2601 15669 2635
rect 15703 2632 15715 2635
rect 15746 2632 15752 2644
rect 15703 2604 15752 2632
rect 15703 2601 15715 2604
rect 15657 2595 15715 2601
rect 15746 2592 15752 2604
rect 15804 2592 15810 2644
rect 15930 2632 15936 2644
rect 15891 2604 15936 2632
rect 15930 2592 15936 2604
rect 15988 2592 15994 2644
rect 17954 2592 17960 2644
rect 18012 2632 18018 2644
rect 18417 2635 18475 2641
rect 18417 2632 18429 2635
rect 18012 2604 18429 2632
rect 18012 2592 18018 2604
rect 3418 2524 3424 2576
rect 3476 2564 3482 2576
rect 8662 2564 8668 2576
rect 3476 2536 8668 2564
rect 3476 2524 3482 2536
rect 8662 2524 8668 2536
rect 8720 2524 8726 2576
rect 10045 2567 10103 2573
rect 10045 2564 10057 2567
rect 9600 2536 10057 2564
rect 5629 2499 5687 2505
rect 5629 2465 5641 2499
rect 5675 2496 5687 2499
rect 5810 2496 5816 2508
rect 5675 2468 5816 2496
rect 5675 2465 5687 2468
rect 5629 2459 5687 2465
rect 5810 2456 5816 2468
rect 5868 2456 5874 2508
rect 9600 2505 9628 2536
rect 10045 2533 10057 2536
rect 10091 2564 10103 2567
rect 10318 2564 10324 2576
rect 10091 2536 10324 2564
rect 10091 2533 10103 2536
rect 10045 2527 10103 2533
rect 10318 2524 10324 2536
rect 10376 2524 10382 2576
rect 9401 2499 9459 2505
rect 9401 2465 9413 2499
rect 9447 2465 9459 2499
rect 9401 2459 9459 2465
rect 9585 2499 9643 2505
rect 9585 2465 9597 2499
rect 9631 2465 9643 2499
rect 9585 2459 9643 2465
rect 842 2388 848 2440
rect 900 2428 906 2440
rect 7101 2431 7159 2437
rect 7101 2428 7113 2431
rect 900 2400 7113 2428
rect 900 2388 906 2400
rect 7101 2397 7113 2400
rect 7147 2428 7159 2431
rect 7650 2428 7656 2440
rect 7147 2400 7656 2428
rect 7147 2397 7159 2400
rect 7101 2391 7159 2397
rect 7650 2388 7656 2400
rect 7708 2388 7714 2440
rect 7926 2388 7932 2440
rect 7984 2428 7990 2440
rect 8665 2431 8723 2437
rect 8665 2428 8677 2431
rect 7984 2400 8677 2428
rect 7984 2388 7990 2400
rect 8665 2397 8677 2400
rect 8711 2428 8723 2431
rect 9416 2428 9444 2459
rect 8711 2400 9444 2428
rect 8711 2397 8723 2400
rect 8665 2391 8723 2397
rect 13814 2388 13820 2440
rect 13872 2428 13878 2440
rect 14093 2431 14151 2437
rect 14093 2428 14105 2431
rect 13872 2400 14105 2428
rect 13872 2388 13878 2400
rect 14093 2397 14105 2400
rect 14139 2397 14151 2431
rect 18248 2428 18276 2604
rect 18417 2601 18429 2604
rect 18463 2601 18475 2635
rect 18417 2595 18475 2601
rect 18322 2524 18328 2576
rect 18380 2564 18386 2576
rect 18785 2567 18843 2573
rect 18785 2564 18797 2567
rect 18380 2536 18797 2564
rect 18380 2524 18386 2536
rect 18785 2533 18797 2536
rect 18831 2533 18843 2567
rect 18785 2527 18843 2533
rect 18601 2431 18659 2437
rect 18601 2428 18613 2431
rect 18248 2400 18613 2428
rect 14093 2391 14151 2397
rect 18601 2397 18613 2400
rect 18647 2397 18659 2431
rect 18601 2391 18659 2397
rect 2682 2320 2688 2372
rect 2740 2360 2746 2372
rect 4801 2363 4859 2369
rect 4801 2360 4813 2363
rect 2740 2332 4813 2360
rect 2740 2320 2746 2332
rect 4801 2329 4813 2332
rect 4847 2360 4859 2363
rect 5445 2363 5503 2369
rect 5445 2360 5457 2363
rect 4847 2332 5457 2360
rect 4847 2329 4859 2332
rect 4801 2323 4859 2329
rect 5445 2329 5457 2332
rect 5491 2360 5503 2363
rect 8481 2363 8539 2369
rect 8481 2360 8493 2363
rect 5491 2332 8493 2360
rect 5491 2329 5503 2332
rect 5445 2323 5503 2329
rect 8481 2329 8493 2332
rect 8527 2360 8539 2363
rect 8570 2360 8576 2372
rect 8527 2332 8576 2360
rect 8527 2329 8539 2332
rect 8481 2323 8539 2329
rect 8570 2320 8576 2332
rect 8628 2360 8634 2372
rect 9306 2360 9312 2372
rect 8628 2332 9312 2360
rect 8628 2320 8634 2332
rect 9306 2320 9312 2332
rect 9364 2320 9370 2372
rect 18325 2363 18383 2369
rect 18325 2329 18337 2363
rect 18371 2360 18383 2363
rect 18414 2360 18420 2372
rect 18371 2332 18420 2360
rect 18371 2329 18383 2332
rect 18325 2323 18383 2329
rect 18414 2320 18420 2332
rect 18472 2320 18478 2372
rect 3142 2252 3148 2304
rect 3200 2292 3206 2304
rect 4062 2292 4068 2304
rect 3200 2264 4068 2292
rect 3200 2252 3206 2264
rect 4062 2252 4068 2264
rect 4120 2292 4126 2304
rect 4617 2295 4675 2301
rect 4617 2292 4629 2295
rect 4120 2264 4629 2292
rect 4120 2252 4126 2264
rect 4617 2261 4629 2264
rect 4663 2292 4675 2295
rect 5353 2295 5411 2301
rect 5353 2292 5365 2295
rect 4663 2264 5365 2292
rect 4663 2261 4675 2264
rect 4617 2255 4675 2261
rect 5353 2261 5365 2264
rect 5399 2261 5411 2295
rect 6914 2292 6920 2304
rect 6875 2264 6920 2292
rect 5353 2255 5411 2261
rect 6914 2252 6920 2264
rect 6972 2252 6978 2304
rect 14182 2252 14188 2304
rect 14240 2292 14246 2304
rect 14277 2295 14335 2301
rect 14277 2292 14289 2295
rect 14240 2264 14289 2292
rect 14240 2252 14246 2264
rect 14277 2261 14289 2264
rect 14323 2261 14335 2295
rect 14277 2255 14335 2261
rect 1104 2202 22056 2224
rect 1104 2150 6148 2202
rect 6200 2150 6212 2202
rect 6264 2150 6276 2202
rect 6328 2150 6340 2202
rect 6392 2150 6404 2202
rect 6456 2150 11346 2202
rect 11398 2150 11410 2202
rect 11462 2150 11474 2202
rect 11526 2150 11538 2202
rect 11590 2150 11602 2202
rect 11654 2150 16544 2202
rect 16596 2150 16608 2202
rect 16660 2150 16672 2202
rect 16724 2150 16736 2202
rect 16788 2150 16800 2202
rect 16852 2150 21742 2202
rect 21794 2150 21806 2202
rect 21858 2150 21870 2202
rect 21922 2150 21934 2202
rect 21986 2150 21998 2202
rect 22050 2150 22056 2202
rect 1104 2128 22056 2150
rect 3418 2048 3424 2100
rect 3476 2088 3482 2100
rect 7558 2088 7564 2100
rect 3476 2060 7564 2088
rect 3476 2048 3482 2060
rect 7558 2048 7564 2060
rect 7616 2048 7622 2100
rect 1302 1980 1308 2032
rect 1360 2020 1366 2032
rect 6914 2020 6920 2032
rect 1360 1992 6920 2020
rect 1360 1980 1366 1992
rect 6914 1980 6920 1992
rect 6972 1980 6978 2032
<< via1 >>
rect 11244 20952 11296 21004
rect 11704 20952 11756 21004
rect 6148 20646 6200 20698
rect 6212 20646 6264 20698
rect 6276 20646 6328 20698
rect 6340 20646 6392 20698
rect 6404 20646 6456 20698
rect 11346 20646 11398 20698
rect 11410 20646 11462 20698
rect 11474 20646 11526 20698
rect 11538 20646 11590 20698
rect 11602 20646 11654 20698
rect 16544 20646 16596 20698
rect 16608 20646 16660 20698
rect 16672 20646 16724 20698
rect 16736 20646 16788 20698
rect 16800 20646 16852 20698
rect 21742 20646 21794 20698
rect 21806 20646 21858 20698
rect 21870 20646 21922 20698
rect 21934 20646 21986 20698
rect 21998 20646 22050 20698
rect 7748 20544 7800 20596
rect 15844 20544 15896 20596
rect 11060 20476 11112 20528
rect 14004 20476 14056 20528
rect 9220 20315 9272 20324
rect 9220 20281 9229 20315
rect 9229 20281 9263 20315
rect 9263 20281 9272 20315
rect 9220 20272 9272 20281
rect 10692 20408 10744 20460
rect 22284 20408 22336 20460
rect 9680 20340 9732 20392
rect 14464 20340 14516 20392
rect 21548 20340 21600 20392
rect 11152 20272 11204 20324
rect 12532 20272 12584 20324
rect 17224 20272 17276 20324
rect 8116 20204 8168 20256
rect 20444 20204 20496 20256
rect 3549 20102 3601 20154
rect 3613 20102 3665 20154
rect 3677 20102 3729 20154
rect 3741 20102 3793 20154
rect 3805 20102 3857 20154
rect 8747 20102 8799 20154
rect 8811 20102 8863 20154
rect 8875 20102 8927 20154
rect 8939 20102 8991 20154
rect 9003 20102 9055 20154
rect 13945 20102 13997 20154
rect 14009 20102 14061 20154
rect 14073 20102 14125 20154
rect 14137 20102 14189 20154
rect 14201 20102 14253 20154
rect 19143 20102 19195 20154
rect 19207 20102 19259 20154
rect 19271 20102 19323 20154
rect 19335 20102 19387 20154
rect 19399 20102 19451 20154
rect 2780 20043 2832 20052
rect 2780 20009 2789 20043
rect 2789 20009 2823 20043
rect 2823 20009 2832 20043
rect 7748 20043 7800 20052
rect 2780 20000 2832 20009
rect 7748 20009 7757 20043
rect 7757 20009 7791 20043
rect 7791 20009 7800 20043
rect 7748 20000 7800 20009
rect 9680 20000 9732 20052
rect 13544 20000 13596 20052
rect 19064 20000 19116 20052
rect 11060 19864 11112 19916
rect 6736 19660 6788 19712
rect 7656 19796 7708 19848
rect 8392 19839 8444 19848
rect 8392 19805 8401 19839
rect 8401 19805 8435 19839
rect 8435 19805 8444 19839
rect 8392 19796 8444 19805
rect 9404 19839 9456 19848
rect 8116 19728 8168 19780
rect 9404 19805 9413 19839
rect 9413 19805 9447 19839
rect 9447 19805 9456 19839
rect 9404 19796 9456 19805
rect 9772 19839 9824 19848
rect 9772 19805 9781 19839
rect 9781 19805 9815 19839
rect 9815 19805 9824 19839
rect 9772 19796 9824 19805
rect 9956 19796 10008 19848
rect 10048 19796 10100 19848
rect 10600 19839 10652 19848
rect 10600 19805 10609 19839
rect 10609 19805 10643 19839
rect 10643 19805 10652 19839
rect 10600 19796 10652 19805
rect 21364 20000 21416 20052
rect 21548 19907 21600 19916
rect 21548 19873 21557 19907
rect 21557 19873 21591 19907
rect 21591 19873 21600 19907
rect 21548 19864 21600 19873
rect 12900 19796 12952 19848
rect 13084 19796 13136 19848
rect 13636 19796 13688 19848
rect 14832 19796 14884 19848
rect 12440 19728 12492 19780
rect 7380 19703 7432 19712
rect 7380 19669 7389 19703
rect 7389 19669 7423 19703
rect 7423 19669 7432 19703
rect 7380 19660 7432 19669
rect 10140 19660 10192 19712
rect 10416 19703 10468 19712
rect 10416 19669 10425 19703
rect 10425 19669 10459 19703
rect 10459 19669 10468 19703
rect 10416 19660 10468 19669
rect 11060 19660 11112 19712
rect 11888 19660 11940 19712
rect 14372 19728 14424 19780
rect 14464 19728 14516 19780
rect 21088 19728 21140 19780
rect 13084 19703 13136 19712
rect 13084 19669 13093 19703
rect 13093 19669 13127 19703
rect 13127 19669 13136 19703
rect 13084 19660 13136 19669
rect 16948 19660 17000 19712
rect 20168 19703 20220 19712
rect 20168 19669 20177 19703
rect 20177 19669 20211 19703
rect 20211 19669 20220 19703
rect 20168 19660 20220 19669
rect 6148 19558 6200 19610
rect 6212 19558 6264 19610
rect 6276 19558 6328 19610
rect 6340 19558 6392 19610
rect 6404 19558 6456 19610
rect 11346 19558 11398 19610
rect 11410 19558 11462 19610
rect 11474 19558 11526 19610
rect 11538 19558 11590 19610
rect 11602 19558 11654 19610
rect 16544 19558 16596 19610
rect 16608 19558 16660 19610
rect 16672 19558 16724 19610
rect 16736 19558 16788 19610
rect 16800 19558 16852 19610
rect 21742 19558 21794 19610
rect 21806 19558 21858 19610
rect 21870 19558 21922 19610
rect 21934 19558 21986 19610
rect 21998 19558 22050 19610
rect 8300 19499 8352 19508
rect 8300 19465 8309 19499
rect 8309 19465 8343 19499
rect 8343 19465 8352 19499
rect 8300 19456 8352 19465
rect 11888 19456 11940 19508
rect 12440 19456 12492 19508
rect 19616 19456 19668 19508
rect 21548 19499 21600 19508
rect 8668 19320 8720 19372
rect 9128 19252 9180 19304
rect 8576 19159 8628 19168
rect 8576 19125 8585 19159
rect 8585 19125 8619 19159
rect 8619 19125 8628 19159
rect 8576 19116 8628 19125
rect 12532 19388 12584 19440
rect 12808 19388 12860 19440
rect 10048 19363 10100 19372
rect 10048 19329 10057 19363
rect 10057 19329 10091 19363
rect 10091 19329 10100 19363
rect 10048 19320 10100 19329
rect 13084 19320 13136 19372
rect 13820 19320 13872 19372
rect 9496 19116 9548 19168
rect 10140 19184 10192 19236
rect 10876 19116 10928 19168
rect 12900 19116 12952 19168
rect 14648 19252 14700 19304
rect 17040 19252 17092 19304
rect 21548 19465 21557 19499
rect 21557 19465 21591 19499
rect 21591 19465 21600 19499
rect 21548 19456 21600 19465
rect 20996 19320 21048 19372
rect 20904 19252 20956 19304
rect 16304 19184 16356 19236
rect 16948 19184 17000 19236
rect 14740 19116 14792 19168
rect 18144 19116 18196 19168
rect 21640 19116 21692 19168
rect 3549 19014 3601 19066
rect 3613 19014 3665 19066
rect 3677 19014 3729 19066
rect 3741 19014 3793 19066
rect 3805 19014 3857 19066
rect 8747 19014 8799 19066
rect 8811 19014 8863 19066
rect 8875 19014 8927 19066
rect 8939 19014 8991 19066
rect 9003 19014 9055 19066
rect 13945 19014 13997 19066
rect 14009 19014 14061 19066
rect 14073 19014 14125 19066
rect 14137 19014 14189 19066
rect 14201 19014 14253 19066
rect 19143 19014 19195 19066
rect 19207 19014 19259 19066
rect 19271 19014 19323 19066
rect 19335 19014 19387 19066
rect 19399 19014 19451 19066
rect 8944 18912 8996 18964
rect 9956 18912 10008 18964
rect 10416 18912 10468 18964
rect 9864 18844 9916 18896
rect 10048 18844 10100 18896
rect 12900 18912 12952 18964
rect 17500 18912 17552 18964
rect 20996 18955 21048 18964
rect 20996 18921 21005 18955
rect 21005 18921 21039 18955
rect 21039 18921 21048 18955
rect 20996 18912 21048 18921
rect 14740 18844 14792 18896
rect 9404 18819 9456 18828
rect 9404 18785 9413 18819
rect 9413 18785 9447 18819
rect 9447 18785 9456 18819
rect 9404 18776 9456 18785
rect 9772 18776 9824 18828
rect 10508 18776 10560 18828
rect 13360 18776 13412 18828
rect 14188 18776 14240 18828
rect 14556 18776 14608 18828
rect 8576 18708 8628 18760
rect 9128 18708 9180 18760
rect 9220 18751 9272 18760
rect 9220 18717 9229 18751
rect 9229 18717 9263 18751
rect 9263 18717 9272 18751
rect 9220 18708 9272 18717
rect 10968 18708 11020 18760
rect 11060 18708 11112 18760
rect 13176 18708 13228 18760
rect 13728 18708 13780 18760
rect 14648 18708 14700 18760
rect 16396 18708 16448 18760
rect 204 18572 256 18624
rect 4620 18572 4672 18624
rect 8300 18615 8352 18624
rect 8300 18581 8309 18615
rect 8309 18581 8343 18615
rect 8343 18581 8352 18615
rect 8300 18572 8352 18581
rect 10140 18640 10192 18692
rect 10416 18615 10468 18624
rect 10416 18581 10425 18615
rect 10425 18581 10459 18615
rect 10459 18581 10468 18615
rect 10416 18572 10468 18581
rect 11980 18640 12032 18692
rect 14280 18640 14332 18692
rect 14372 18640 14424 18692
rect 17868 18683 17920 18692
rect 17868 18649 17886 18683
rect 17886 18649 17920 18683
rect 17868 18640 17920 18649
rect 19708 18708 19760 18760
rect 22744 18708 22796 18760
rect 20352 18640 20404 18692
rect 12532 18572 12584 18624
rect 13544 18572 13596 18624
rect 16120 18615 16172 18624
rect 16120 18581 16129 18615
rect 16129 18581 16163 18615
rect 16163 18581 16172 18615
rect 16120 18572 16172 18581
rect 16948 18572 17000 18624
rect 18236 18615 18288 18624
rect 18236 18581 18245 18615
rect 18245 18581 18279 18615
rect 18279 18581 18288 18615
rect 18236 18572 18288 18581
rect 19892 18572 19944 18624
rect 6148 18470 6200 18522
rect 6212 18470 6264 18522
rect 6276 18470 6328 18522
rect 6340 18470 6392 18522
rect 6404 18470 6456 18522
rect 11346 18470 11398 18522
rect 11410 18470 11462 18522
rect 11474 18470 11526 18522
rect 11538 18470 11590 18522
rect 11602 18470 11654 18522
rect 16544 18470 16596 18522
rect 16608 18470 16660 18522
rect 16672 18470 16724 18522
rect 16736 18470 16788 18522
rect 16800 18470 16852 18522
rect 21742 18470 21794 18522
rect 21806 18470 21858 18522
rect 21870 18470 21922 18522
rect 21934 18470 21986 18522
rect 21998 18470 22050 18522
rect 2872 18368 2924 18420
rect 4344 18368 4396 18420
rect 9036 18368 9088 18420
rect 2504 18300 2556 18352
rect 4436 18300 4488 18352
rect 3148 18232 3200 18284
rect 3884 18232 3936 18284
rect 5080 18232 5132 18284
rect 8024 18232 8076 18284
rect 2044 18164 2096 18216
rect 4344 18164 4396 18216
rect 6092 18164 6144 18216
rect 9036 18232 9088 18284
rect 9634 18275 9686 18284
rect 9634 18241 9658 18275
rect 9658 18241 9686 18275
rect 9634 18232 9686 18241
rect 10140 18368 10192 18420
rect 14188 18368 14240 18420
rect 14648 18411 14700 18420
rect 10232 18300 10284 18352
rect 10416 18300 10468 18352
rect 13360 18300 13412 18352
rect 14372 18300 14424 18352
rect 8852 18207 8904 18216
rect 8852 18173 8861 18207
rect 8861 18173 8895 18207
rect 8895 18173 8904 18207
rect 8852 18164 8904 18173
rect 9404 18207 9456 18216
rect 9404 18173 9413 18207
rect 9413 18173 9447 18207
rect 9447 18173 9456 18207
rect 9404 18164 9456 18173
rect 13728 18232 13780 18284
rect 14188 18275 14240 18284
rect 14648 18377 14657 18411
rect 14657 18377 14691 18411
rect 14691 18377 14700 18411
rect 14648 18368 14700 18377
rect 14188 18241 14206 18275
rect 14206 18241 14240 18275
rect 14188 18232 14240 18241
rect 1584 18096 1636 18148
rect 4160 18096 4212 18148
rect 4804 18096 4856 18148
rect 6828 18096 6880 18148
rect 7012 18096 7064 18148
rect 8944 18096 8996 18148
rect 1124 18028 1176 18080
rect 3884 18028 3936 18080
rect 5356 18028 5408 18080
rect 6092 18071 6144 18080
rect 6092 18037 6101 18071
rect 6101 18037 6135 18071
rect 6135 18037 6144 18071
rect 6092 18028 6144 18037
rect 8024 18028 8076 18080
rect 8208 18071 8260 18080
rect 8208 18037 8217 18071
rect 8217 18037 8251 18071
rect 8251 18037 8260 18071
rect 8208 18028 8260 18037
rect 8484 18028 8536 18080
rect 10508 18164 10560 18216
rect 9956 18096 10008 18148
rect 11336 18071 11388 18080
rect 11336 18037 11345 18071
rect 11345 18037 11379 18071
rect 11379 18037 11388 18071
rect 11336 18028 11388 18037
rect 11980 18028 12032 18080
rect 13084 18071 13136 18080
rect 13084 18037 13093 18071
rect 13093 18037 13127 18071
rect 13127 18037 13136 18071
rect 13084 18028 13136 18037
rect 13176 18028 13228 18080
rect 17868 18368 17920 18420
rect 20996 18368 21048 18420
rect 16396 18232 16448 18284
rect 17776 18275 17828 18284
rect 18236 18300 18288 18352
rect 17776 18241 17794 18275
rect 17794 18241 17828 18275
rect 17776 18232 17828 18241
rect 18972 18232 19024 18284
rect 16120 18028 16172 18080
rect 20904 18096 20956 18148
rect 3549 17926 3601 17978
rect 3613 17926 3665 17978
rect 3677 17926 3729 17978
rect 3741 17926 3793 17978
rect 3805 17926 3857 17978
rect 8747 17926 8799 17978
rect 8811 17926 8863 17978
rect 8875 17926 8927 17978
rect 8939 17926 8991 17978
rect 9003 17926 9055 17978
rect 13945 17926 13997 17978
rect 14009 17926 14061 17978
rect 14073 17926 14125 17978
rect 14137 17926 14189 17978
rect 14201 17926 14253 17978
rect 19143 17926 19195 17978
rect 19207 17926 19259 17978
rect 19271 17926 19323 17978
rect 19335 17926 19387 17978
rect 19399 17926 19451 17978
rect 3056 17824 3108 17876
rect 3424 17824 3476 17876
rect 4528 17824 4580 17876
rect 7012 17824 7064 17876
rect 9220 17824 9272 17876
rect 9956 17824 10008 17876
rect 10968 17824 11020 17876
rect 11336 17824 11388 17876
rect 6920 17756 6972 17808
rect 11612 17756 11664 17808
rect 5172 17731 5224 17740
rect 5172 17697 5181 17731
rect 5181 17697 5215 17731
rect 5215 17697 5224 17731
rect 5172 17688 5224 17697
rect 5356 17731 5408 17740
rect 5356 17697 5365 17731
rect 5365 17697 5399 17731
rect 5399 17697 5408 17731
rect 5356 17688 5408 17697
rect 3424 17620 3476 17672
rect 4988 17620 5040 17672
rect 6092 17688 6144 17740
rect 13452 17867 13504 17876
rect 13452 17833 13461 17867
rect 13461 17833 13495 17867
rect 13495 17833 13504 17867
rect 13452 17824 13504 17833
rect 16856 17824 16908 17876
rect 5724 17620 5776 17672
rect 6644 17620 6696 17672
rect 7472 17620 7524 17672
rect 9128 17620 9180 17672
rect 9864 17620 9916 17672
rect 12808 17688 12860 17740
rect 13268 17688 13320 17740
rect 13544 17756 13596 17808
rect 13728 17688 13780 17740
rect 3516 17552 3568 17604
rect 7380 17552 7432 17604
rect 9220 17552 9272 17604
rect 4988 17484 5040 17536
rect 5724 17484 5776 17536
rect 5908 17527 5960 17536
rect 5908 17493 5917 17527
rect 5917 17493 5951 17527
rect 5951 17493 5960 17527
rect 5908 17484 5960 17493
rect 6552 17484 6604 17536
rect 7932 17484 7984 17536
rect 9128 17484 9180 17536
rect 12348 17552 12400 17604
rect 12532 17620 12584 17672
rect 14372 17688 14424 17740
rect 15108 17688 15160 17740
rect 16396 17688 16448 17740
rect 20996 17824 21048 17876
rect 19892 17620 19944 17672
rect 12532 17484 12584 17536
rect 12992 17484 13044 17536
rect 19708 17552 19760 17604
rect 18972 17484 19024 17536
rect 21088 17484 21140 17536
rect 6148 17382 6200 17434
rect 6212 17382 6264 17434
rect 6276 17382 6328 17434
rect 6340 17382 6392 17434
rect 6404 17382 6456 17434
rect 11346 17382 11398 17434
rect 11410 17382 11462 17434
rect 11474 17382 11526 17434
rect 11538 17382 11590 17434
rect 11602 17382 11654 17434
rect 16544 17382 16596 17434
rect 16608 17382 16660 17434
rect 16672 17382 16724 17434
rect 16736 17382 16788 17434
rect 16800 17382 16852 17434
rect 21742 17382 21794 17434
rect 21806 17382 21858 17434
rect 21870 17382 21922 17434
rect 21934 17382 21986 17434
rect 21998 17382 22050 17434
rect 2964 17280 3016 17332
rect 3332 17280 3384 17332
rect 4068 17280 4120 17332
rect 4528 17323 4580 17332
rect 4528 17289 4537 17323
rect 4537 17289 4571 17323
rect 4571 17289 4580 17323
rect 4528 17280 4580 17289
rect 4988 17280 5040 17332
rect 5816 17280 5868 17332
rect 7380 17323 7432 17332
rect 7380 17289 7389 17323
rect 7389 17289 7423 17323
rect 7423 17289 7432 17323
rect 7380 17280 7432 17289
rect 7932 17323 7984 17332
rect 7932 17289 7941 17323
rect 7941 17289 7975 17323
rect 7975 17289 7984 17323
rect 7932 17280 7984 17289
rect 8392 17280 8444 17332
rect 9128 17323 9180 17332
rect 9128 17289 9137 17323
rect 9137 17289 9171 17323
rect 9171 17289 9180 17323
rect 9128 17280 9180 17289
rect 3424 17255 3476 17264
rect 3424 17221 3433 17255
rect 3433 17221 3467 17255
rect 3467 17221 3476 17255
rect 3424 17212 3476 17221
rect 4160 17212 4212 17264
rect 5724 17212 5776 17264
rect 8208 17212 8260 17264
rect 9312 17212 9364 17264
rect 2964 17144 3016 17196
rect 3148 17187 3200 17196
rect 3148 17153 3157 17187
rect 3157 17153 3191 17187
rect 3191 17153 3200 17187
rect 3148 17144 3200 17153
rect 5540 17187 5592 17196
rect 2780 17008 2832 17060
rect 3240 17008 3292 17060
rect 5540 17153 5549 17187
rect 5549 17153 5583 17187
rect 5583 17153 5592 17187
rect 5540 17144 5592 17153
rect 8392 17144 8444 17196
rect 4896 17076 4948 17128
rect 5172 17076 5224 17128
rect 5448 17076 5500 17128
rect 6920 17076 6972 17128
rect 7196 17076 7248 17128
rect 7748 17119 7800 17128
rect 7748 17085 7757 17119
rect 7757 17085 7791 17119
rect 7791 17085 7800 17119
rect 7748 17076 7800 17085
rect 13176 17280 13228 17332
rect 13360 17280 13412 17332
rect 10692 17255 10744 17264
rect 10692 17221 10701 17255
rect 10701 17221 10735 17255
rect 10735 17221 10744 17255
rect 10692 17212 10744 17221
rect 10968 17212 11020 17264
rect 12808 17212 12860 17264
rect 10416 17187 10468 17196
rect 10416 17153 10425 17187
rect 10425 17153 10459 17187
rect 10459 17153 10468 17187
rect 10416 17144 10468 17153
rect 15844 17212 15896 17264
rect 16396 17212 16448 17264
rect 14372 17144 14424 17196
rect 16212 17187 16264 17196
rect 16212 17153 16230 17187
rect 16230 17153 16264 17187
rect 16212 17144 16264 17153
rect 20168 17280 20220 17332
rect 20996 17280 21048 17332
rect 2872 16940 2924 16992
rect 4620 16940 4672 16992
rect 6552 16940 6604 16992
rect 8392 16983 8444 16992
rect 8392 16949 8401 16983
rect 8401 16949 8435 16983
rect 8435 16949 8444 16983
rect 8392 16940 8444 16949
rect 9128 16940 9180 16992
rect 9772 16940 9824 16992
rect 10692 16940 10744 16992
rect 10968 16983 11020 16992
rect 10968 16949 10977 16983
rect 10977 16949 11011 16983
rect 11011 16949 11020 16983
rect 10968 16940 11020 16949
rect 11520 16983 11572 16992
rect 11520 16949 11529 16983
rect 11529 16949 11563 16983
rect 11563 16949 11572 16983
rect 11520 16940 11572 16949
rect 18052 17119 18104 17128
rect 15108 17051 15160 17060
rect 15108 17017 15117 17051
rect 15117 17017 15151 17051
rect 15151 17017 15160 17051
rect 15108 17008 15160 17017
rect 18052 17085 18061 17119
rect 18061 17085 18095 17119
rect 18095 17085 18104 17119
rect 19064 17144 19116 17196
rect 18052 17076 18104 17085
rect 15476 16940 15528 16992
rect 17776 16940 17828 16992
rect 20352 16983 20404 16992
rect 20352 16949 20361 16983
rect 20361 16949 20395 16983
rect 20395 16949 20404 16983
rect 20352 16940 20404 16949
rect 3549 16838 3601 16890
rect 3613 16838 3665 16890
rect 3677 16838 3729 16890
rect 3741 16838 3793 16890
rect 3805 16838 3857 16890
rect 8747 16838 8799 16890
rect 8811 16838 8863 16890
rect 8875 16838 8927 16890
rect 8939 16838 8991 16890
rect 9003 16838 9055 16890
rect 13945 16838 13997 16890
rect 14009 16838 14061 16890
rect 14073 16838 14125 16890
rect 14137 16838 14189 16890
rect 14201 16838 14253 16890
rect 19143 16838 19195 16890
rect 19207 16838 19259 16890
rect 19271 16838 19323 16890
rect 19335 16838 19387 16890
rect 19399 16838 19451 16890
rect 3884 16779 3936 16788
rect 3884 16745 3893 16779
rect 3893 16745 3927 16779
rect 3927 16745 3936 16779
rect 3884 16736 3936 16745
rect 4344 16736 4396 16788
rect 6552 16779 6604 16788
rect 6552 16745 6561 16779
rect 6561 16745 6595 16779
rect 6595 16745 6604 16779
rect 6552 16736 6604 16745
rect 664 16668 716 16720
rect 3424 16668 3476 16720
rect 2964 16600 3016 16652
rect 4896 16600 4948 16652
rect 6184 16643 6236 16652
rect 2780 16575 2832 16584
rect 2780 16541 2789 16575
rect 2789 16541 2823 16575
rect 2823 16541 2832 16575
rect 2780 16532 2832 16541
rect 3608 16575 3660 16584
rect 3608 16541 3617 16575
rect 3617 16541 3651 16575
rect 3651 16541 3660 16575
rect 3608 16532 3660 16541
rect 5540 16532 5592 16584
rect 4160 16464 4212 16516
rect 6184 16609 6193 16643
rect 6193 16609 6227 16643
rect 6227 16609 6236 16643
rect 6184 16600 6236 16609
rect 7564 16643 7616 16652
rect 7564 16609 7573 16643
rect 7573 16609 7607 16643
rect 7607 16609 7616 16643
rect 7564 16600 7616 16609
rect 9128 16668 9180 16720
rect 8116 16643 8168 16652
rect 8116 16609 8125 16643
rect 8125 16609 8159 16643
rect 8159 16609 8168 16643
rect 8116 16600 8168 16609
rect 10692 16668 10744 16720
rect 12532 16736 12584 16788
rect 13820 16736 13872 16788
rect 15844 16779 15896 16788
rect 15844 16745 15853 16779
rect 15853 16745 15887 16779
rect 15887 16745 15896 16779
rect 15844 16736 15896 16745
rect 18052 16736 18104 16788
rect 5724 16532 5776 16584
rect 8668 16532 8720 16584
rect 9496 16575 9548 16584
rect 9496 16541 9505 16575
rect 9505 16541 9539 16575
rect 9539 16541 9548 16575
rect 9496 16532 9548 16541
rect 3884 16396 3936 16448
rect 4896 16439 4948 16448
rect 4896 16405 4905 16439
rect 4905 16405 4939 16439
rect 4939 16405 4948 16439
rect 4896 16396 4948 16405
rect 5356 16396 5408 16448
rect 5540 16439 5592 16448
rect 5540 16405 5549 16439
rect 5549 16405 5583 16439
rect 5583 16405 5592 16439
rect 5540 16396 5592 16405
rect 5908 16439 5960 16448
rect 5908 16405 5917 16439
rect 5917 16405 5951 16439
rect 5951 16405 5960 16439
rect 5908 16396 5960 16405
rect 6000 16439 6052 16448
rect 6000 16405 6009 16439
rect 6009 16405 6043 16439
rect 6043 16405 6052 16439
rect 8300 16507 8352 16516
rect 8300 16473 8309 16507
rect 8309 16473 8343 16507
rect 8343 16473 8352 16507
rect 8300 16464 8352 16473
rect 6000 16396 6052 16405
rect 9128 16464 9180 16516
rect 9312 16464 9364 16516
rect 11152 16532 11204 16584
rect 12256 16600 12308 16652
rect 9772 16464 9824 16516
rect 9404 16396 9456 16448
rect 10324 16439 10376 16448
rect 10324 16405 10333 16439
rect 10333 16405 10367 16439
rect 10367 16405 10376 16439
rect 10324 16396 10376 16405
rect 12992 16507 13044 16516
rect 12992 16473 13010 16507
rect 13010 16473 13044 16507
rect 14740 16600 14792 16652
rect 20996 16736 21048 16788
rect 21456 16736 21508 16788
rect 13360 16532 13412 16584
rect 12992 16464 13044 16473
rect 13728 16464 13780 16516
rect 15200 16464 15252 16516
rect 15384 16464 15436 16516
rect 16396 16464 16448 16516
rect 17960 16507 18012 16516
rect 17960 16473 17978 16507
rect 17978 16473 18012 16507
rect 17960 16464 18012 16473
rect 11060 16396 11112 16448
rect 11980 16396 12032 16448
rect 12072 16396 12124 16448
rect 13820 16396 13872 16448
rect 14740 16396 14792 16448
rect 18972 16396 19024 16448
rect 21364 16396 21416 16448
rect 6148 16294 6200 16346
rect 6212 16294 6264 16346
rect 6276 16294 6328 16346
rect 6340 16294 6392 16346
rect 6404 16294 6456 16346
rect 11346 16294 11398 16346
rect 11410 16294 11462 16346
rect 11474 16294 11526 16346
rect 11538 16294 11590 16346
rect 11602 16294 11654 16346
rect 16544 16294 16596 16346
rect 16608 16294 16660 16346
rect 16672 16294 16724 16346
rect 16736 16294 16788 16346
rect 16800 16294 16852 16346
rect 21742 16294 21794 16346
rect 21806 16294 21858 16346
rect 21870 16294 21922 16346
rect 21934 16294 21986 16346
rect 21998 16294 22050 16346
rect 4068 16235 4120 16244
rect 4068 16201 4077 16235
rect 4077 16201 4111 16235
rect 4111 16201 4120 16235
rect 4068 16192 4120 16201
rect 4344 16235 4396 16244
rect 4344 16201 4353 16235
rect 4353 16201 4387 16235
rect 4387 16201 4396 16235
rect 4344 16192 4396 16201
rect 5908 16192 5960 16244
rect 9312 16192 9364 16244
rect 3056 16167 3108 16176
rect 3056 16133 3065 16167
rect 3065 16133 3099 16167
rect 3099 16133 3108 16167
rect 3056 16124 3108 16133
rect 3148 16124 3200 16176
rect 5540 16124 5592 16176
rect 6552 16124 6604 16176
rect 9956 16124 10008 16176
rect 10784 16192 10836 16244
rect 11060 16235 11112 16244
rect 11060 16201 11069 16235
rect 11069 16201 11103 16235
rect 11103 16201 11112 16235
rect 11060 16192 11112 16201
rect 11152 16192 11204 16244
rect 14832 16192 14884 16244
rect 3884 16099 3936 16108
rect 3884 16065 3893 16099
rect 3893 16065 3927 16099
rect 3927 16065 3936 16099
rect 3884 16056 3936 16065
rect 5172 16056 5224 16108
rect 6368 16056 6420 16108
rect 7840 16099 7892 16108
rect 7840 16065 7849 16099
rect 7849 16065 7883 16099
rect 7883 16065 7892 16099
rect 7840 16056 7892 16065
rect 10048 16099 10100 16108
rect 10048 16065 10057 16099
rect 10057 16065 10091 16099
rect 10091 16065 10100 16099
rect 10048 16056 10100 16065
rect 11612 16124 11664 16176
rect 15384 16124 15436 16176
rect 3976 15988 4028 16040
rect 5264 15988 5316 16040
rect 6000 15988 6052 16040
rect 10508 16031 10560 16040
rect 5816 15920 5868 15972
rect 6920 15920 6972 15972
rect 8668 15920 8720 15972
rect 9128 15920 9180 15972
rect 10508 15997 10517 16031
rect 10517 15997 10551 16031
rect 10551 15997 10560 16031
rect 10508 15988 10560 15997
rect 12072 16056 12124 16108
rect 12532 16056 12584 16108
rect 15108 16056 15160 16108
rect 18972 16099 19024 16108
rect 18972 16065 18990 16099
rect 18990 16065 19024 16099
rect 18972 16056 19024 16065
rect 21180 16099 21232 16108
rect 21180 16065 21198 16099
rect 21198 16065 21232 16099
rect 21456 16099 21508 16108
rect 21180 16056 21232 16065
rect 21456 16065 21465 16099
rect 21465 16065 21499 16099
rect 21499 16065 21508 16099
rect 21456 16056 21508 16065
rect 11152 16031 11204 16040
rect 9772 15920 9824 15972
rect 11152 15997 11161 16031
rect 11161 15997 11195 16031
rect 11195 15997 11204 16031
rect 11152 15988 11204 15997
rect 15200 16031 15252 16040
rect 10784 15920 10836 15972
rect 12348 15920 12400 15972
rect 15200 15997 15209 16031
rect 15209 15997 15243 16031
rect 15243 15997 15252 16031
rect 15200 15988 15252 15997
rect 3884 15852 3936 15904
rect 4988 15852 5040 15904
rect 6368 15895 6420 15904
rect 6368 15861 6377 15895
rect 6377 15861 6411 15895
rect 6411 15861 6420 15895
rect 6368 15852 6420 15861
rect 7932 15852 7984 15904
rect 8300 15895 8352 15904
rect 8300 15861 8309 15895
rect 8309 15861 8343 15895
rect 8343 15861 8352 15895
rect 9220 15895 9272 15904
rect 8300 15852 8352 15861
rect 9220 15861 9229 15895
rect 9229 15861 9263 15895
rect 9263 15861 9272 15895
rect 9220 15852 9272 15861
rect 9312 15852 9364 15904
rect 9956 15852 10008 15904
rect 11612 15852 11664 15904
rect 13728 15895 13780 15904
rect 13728 15861 13737 15895
rect 13737 15861 13771 15895
rect 13771 15861 13780 15895
rect 13728 15852 13780 15861
rect 14832 15852 14884 15904
rect 15844 15852 15896 15904
rect 20076 15895 20128 15904
rect 20076 15861 20085 15895
rect 20085 15861 20119 15895
rect 20119 15861 20128 15895
rect 20076 15852 20128 15861
rect 3549 15750 3601 15802
rect 3613 15750 3665 15802
rect 3677 15750 3729 15802
rect 3741 15750 3793 15802
rect 3805 15750 3857 15802
rect 8747 15750 8799 15802
rect 8811 15750 8863 15802
rect 8875 15750 8927 15802
rect 8939 15750 8991 15802
rect 9003 15750 9055 15802
rect 13945 15750 13997 15802
rect 14009 15750 14061 15802
rect 14073 15750 14125 15802
rect 14137 15750 14189 15802
rect 14201 15750 14253 15802
rect 19143 15750 19195 15802
rect 19207 15750 19259 15802
rect 19271 15750 19323 15802
rect 19335 15750 19387 15802
rect 19399 15750 19451 15802
rect 1952 15691 2004 15700
rect 1952 15657 1961 15691
rect 1961 15657 1995 15691
rect 1995 15657 2004 15691
rect 1952 15648 2004 15657
rect 2320 15691 2372 15700
rect 2320 15657 2329 15691
rect 2329 15657 2363 15691
rect 2363 15657 2372 15691
rect 2320 15648 2372 15657
rect 2688 15691 2740 15700
rect 2688 15657 2697 15691
rect 2697 15657 2731 15691
rect 2731 15657 2740 15691
rect 2688 15648 2740 15657
rect 3332 15648 3384 15700
rect 4068 15648 4120 15700
rect 4804 15648 4856 15700
rect 5172 15691 5224 15700
rect 5172 15657 5181 15691
rect 5181 15657 5215 15691
rect 5215 15657 5224 15691
rect 5172 15648 5224 15657
rect 6000 15691 6052 15700
rect 6000 15657 6009 15691
rect 6009 15657 6043 15691
rect 6043 15657 6052 15691
rect 6000 15648 6052 15657
rect 6092 15691 6144 15700
rect 6092 15657 6101 15691
rect 6101 15657 6135 15691
rect 6135 15657 6144 15691
rect 6092 15648 6144 15657
rect 7840 15648 7892 15700
rect 9128 15648 9180 15700
rect 10232 15691 10284 15700
rect 10232 15657 10241 15691
rect 10241 15657 10275 15691
rect 10275 15657 10284 15691
rect 10232 15648 10284 15657
rect 3884 15580 3936 15632
rect 4252 15512 4304 15564
rect 8116 15580 8168 15632
rect 8484 15580 8536 15632
rect 19892 15648 19944 15700
rect 15844 15623 15896 15632
rect 5632 15512 5684 15564
rect 6920 15512 6972 15564
rect 7748 15555 7800 15564
rect 7748 15521 7757 15555
rect 7757 15521 7791 15555
rect 7791 15521 7800 15555
rect 7748 15512 7800 15521
rect 7932 15555 7984 15564
rect 7932 15521 7941 15555
rect 7941 15521 7975 15555
rect 7975 15521 7984 15555
rect 7932 15512 7984 15521
rect 9404 15555 9456 15564
rect 9404 15521 9413 15555
rect 9413 15521 9447 15555
rect 9447 15521 9456 15555
rect 9404 15512 9456 15521
rect 3240 15376 3292 15428
rect 4712 15444 4764 15496
rect 4804 15487 4856 15496
rect 4804 15453 4813 15487
rect 4813 15453 4847 15487
rect 4847 15453 4856 15487
rect 4804 15444 4856 15453
rect 5540 15444 5592 15496
rect 9956 15512 10008 15564
rect 4620 15376 4672 15428
rect 3424 15351 3476 15360
rect 3424 15317 3433 15351
rect 3433 15317 3467 15351
rect 3467 15317 3476 15351
rect 3424 15308 3476 15317
rect 4068 15308 4120 15360
rect 4344 15308 4396 15360
rect 5264 15376 5316 15428
rect 5816 15376 5868 15428
rect 8208 15376 8260 15428
rect 8760 15376 8812 15428
rect 10692 15512 10744 15564
rect 15844 15589 15853 15623
rect 15853 15589 15887 15623
rect 15887 15589 15896 15623
rect 15844 15580 15896 15589
rect 11152 15444 11204 15496
rect 13728 15444 13780 15496
rect 14924 15444 14976 15496
rect 14648 15376 14700 15428
rect 15384 15376 15436 15428
rect 20720 15444 20772 15496
rect 21456 15444 21508 15496
rect 15568 15376 15620 15428
rect 21272 15419 21324 15428
rect 21272 15385 21290 15419
rect 21290 15385 21324 15419
rect 21272 15376 21324 15385
rect 6368 15308 6420 15360
rect 7012 15308 7064 15360
rect 9404 15308 9456 15360
rect 10692 15351 10744 15360
rect 10692 15317 10701 15351
rect 10701 15317 10735 15351
rect 10735 15317 10744 15351
rect 11060 15351 11112 15360
rect 10692 15308 10744 15317
rect 11060 15317 11069 15351
rect 11069 15317 11103 15351
rect 11103 15317 11112 15351
rect 11060 15308 11112 15317
rect 12532 15308 12584 15360
rect 13728 15308 13780 15360
rect 13820 15308 13872 15360
rect 14740 15308 14792 15360
rect 17500 15351 17552 15360
rect 17500 15317 17509 15351
rect 17509 15317 17543 15351
rect 17543 15317 17552 15351
rect 17500 15308 17552 15317
rect 20536 15308 20588 15360
rect 6148 15206 6200 15258
rect 6212 15206 6264 15258
rect 6276 15206 6328 15258
rect 6340 15206 6392 15258
rect 6404 15206 6456 15258
rect 11346 15206 11398 15258
rect 11410 15206 11462 15258
rect 11474 15206 11526 15258
rect 11538 15206 11590 15258
rect 11602 15206 11654 15258
rect 16544 15206 16596 15258
rect 16608 15206 16660 15258
rect 16672 15206 16724 15258
rect 16736 15206 16788 15258
rect 16800 15206 16852 15258
rect 21742 15206 21794 15258
rect 21806 15206 21858 15258
rect 21870 15206 21922 15258
rect 21934 15206 21986 15258
rect 21998 15206 22050 15258
rect 1860 15104 1912 15156
rect 2596 15104 2648 15156
rect 3332 15147 3384 15156
rect 3332 15113 3341 15147
rect 3341 15113 3375 15147
rect 3375 15113 3384 15147
rect 3332 15104 3384 15113
rect 3424 15104 3476 15156
rect 4436 15104 4488 15156
rect 2136 15011 2188 15020
rect 2136 14977 2145 15011
rect 2145 14977 2179 15011
rect 2179 14977 2188 15011
rect 2136 14968 2188 14977
rect 4344 15036 4396 15088
rect 3976 14968 4028 15020
rect 4068 14968 4120 15020
rect 5632 15104 5684 15156
rect 7104 15104 7156 15156
rect 7472 15147 7524 15156
rect 7472 15113 7481 15147
rect 7481 15113 7515 15147
rect 7515 15113 7524 15147
rect 7472 15104 7524 15113
rect 7564 15104 7616 15156
rect 8208 15147 8260 15156
rect 8208 15113 8217 15147
rect 8217 15113 8251 15147
rect 8251 15113 8260 15147
rect 8208 15104 8260 15113
rect 8668 15104 8720 15156
rect 3884 14943 3936 14952
rect 3884 14909 3893 14943
rect 3893 14909 3927 14943
rect 3927 14909 3936 14943
rect 4804 14968 4856 15020
rect 8392 15036 8444 15088
rect 9128 15104 9180 15156
rect 9680 15104 9732 15156
rect 10692 15104 10744 15156
rect 10968 15104 11020 15156
rect 12624 15104 12676 15156
rect 14556 15104 14608 15156
rect 16396 15104 16448 15156
rect 3884 14900 3936 14909
rect 4620 14832 4672 14884
rect 4804 14832 4856 14884
rect 3240 14764 3292 14816
rect 4068 14764 4120 14816
rect 4436 14764 4488 14816
rect 5356 14900 5408 14952
rect 5724 14968 5776 15020
rect 9864 15011 9916 15020
rect 5540 14832 5592 14884
rect 5632 14764 5684 14816
rect 7288 14900 7340 14952
rect 7748 14900 7800 14952
rect 9864 14977 9873 15011
rect 9873 14977 9907 15011
rect 9907 14977 9916 15011
rect 9864 14968 9916 14977
rect 7196 14832 7248 14884
rect 8208 14832 8260 14884
rect 8668 14900 8720 14952
rect 9128 14900 9180 14952
rect 12900 15036 12952 15088
rect 13544 15036 13596 15088
rect 10508 14832 10560 14884
rect 9404 14807 9456 14816
rect 9404 14773 9413 14807
rect 9413 14773 9447 14807
rect 9447 14773 9456 14807
rect 9404 14764 9456 14773
rect 10232 14764 10284 14816
rect 13360 14968 13412 15020
rect 15016 15011 15068 15020
rect 15016 14977 15034 15011
rect 15034 14977 15068 15011
rect 15016 14968 15068 14977
rect 15200 14968 15252 15020
rect 13728 14900 13780 14952
rect 13452 14832 13504 14884
rect 12072 14807 12124 14816
rect 12072 14773 12081 14807
rect 12081 14773 12115 14807
rect 12115 14773 12124 14807
rect 12072 14764 12124 14773
rect 12532 14764 12584 14816
rect 13636 14764 13688 14816
rect 20076 15104 20128 15156
rect 18052 14943 18104 14952
rect 18052 14909 18061 14943
rect 18061 14909 18095 14943
rect 18095 14909 18104 14943
rect 19800 15011 19852 15020
rect 20168 15036 20220 15088
rect 19800 14977 19818 15011
rect 19818 14977 19852 15011
rect 19800 14968 19852 14977
rect 20720 14968 20772 15020
rect 18052 14900 18104 14909
rect 16212 14875 16264 14884
rect 16212 14841 16221 14875
rect 16221 14841 16255 14875
rect 16255 14841 16264 14875
rect 16212 14832 16264 14841
rect 18696 14807 18748 14816
rect 18696 14773 18705 14807
rect 18705 14773 18739 14807
rect 18739 14773 18748 14807
rect 18696 14764 18748 14773
rect 3549 14662 3601 14714
rect 3613 14662 3665 14714
rect 3677 14662 3729 14714
rect 3741 14662 3793 14714
rect 3805 14662 3857 14714
rect 8747 14662 8799 14714
rect 8811 14662 8863 14714
rect 8875 14662 8927 14714
rect 8939 14662 8991 14714
rect 9003 14662 9055 14714
rect 13945 14662 13997 14714
rect 14009 14662 14061 14714
rect 14073 14662 14125 14714
rect 14137 14662 14189 14714
rect 14201 14662 14253 14714
rect 19143 14662 19195 14714
rect 19207 14662 19259 14714
rect 19271 14662 19323 14714
rect 19335 14662 19387 14714
rect 19399 14662 19451 14714
rect 4160 14560 4212 14612
rect 4896 14560 4948 14612
rect 4436 14492 4488 14544
rect 3424 14424 3476 14476
rect 5632 14492 5684 14544
rect 9128 14560 9180 14612
rect 10048 14560 10100 14612
rect 10508 14560 10560 14612
rect 5264 14424 5316 14476
rect 7748 14492 7800 14544
rect 8392 14535 8444 14544
rect 4160 14356 4212 14408
rect 7380 14424 7432 14476
rect 7656 14424 7708 14476
rect 7840 14424 7892 14476
rect 8392 14501 8401 14535
rect 8401 14501 8435 14535
rect 8435 14501 8444 14535
rect 8392 14492 8444 14501
rect 11060 14560 11112 14612
rect 12532 14560 12584 14612
rect 8208 14467 8260 14476
rect 8208 14433 8217 14467
rect 8217 14433 8251 14467
rect 8251 14433 8260 14467
rect 8208 14424 8260 14433
rect 8300 14424 8352 14476
rect 9128 14424 9180 14476
rect 9404 14424 9456 14476
rect 7104 14356 7156 14408
rect 4528 14288 4580 14340
rect 7472 14288 7524 14340
rect 11244 14492 11296 14544
rect 14924 14560 14976 14612
rect 15200 14560 15252 14612
rect 13636 14492 13688 14544
rect 10324 14399 10376 14408
rect 10324 14365 10333 14399
rect 10333 14365 10367 14399
rect 10367 14365 10376 14399
rect 10324 14356 10376 14365
rect 10508 14356 10560 14408
rect 11796 14356 11848 14408
rect 6552 14220 6604 14272
rect 7748 14220 7800 14272
rect 7840 14220 7892 14272
rect 8024 14220 8076 14272
rect 8208 14220 8260 14272
rect 9128 14220 9180 14272
rect 9588 14220 9640 14272
rect 13728 14424 13780 14476
rect 12532 14356 12584 14408
rect 13820 14356 13872 14408
rect 13452 14288 13504 14340
rect 13544 14288 13596 14340
rect 16396 14424 16448 14476
rect 18052 14560 18104 14612
rect 20720 14560 20772 14612
rect 21456 14603 21508 14612
rect 21456 14569 21465 14603
rect 21465 14569 21499 14603
rect 21499 14569 21508 14603
rect 21456 14560 21508 14569
rect 15568 14399 15620 14408
rect 15568 14365 15597 14399
rect 15597 14365 15620 14399
rect 15568 14356 15620 14365
rect 16212 14356 16264 14408
rect 20352 14356 20404 14408
rect 10048 14220 10100 14272
rect 10324 14220 10376 14272
rect 11888 14220 11940 14272
rect 12348 14220 12400 14272
rect 12716 14220 12768 14272
rect 13176 14220 13228 14272
rect 13636 14263 13688 14272
rect 13636 14229 13645 14263
rect 13645 14229 13679 14263
rect 13679 14229 13688 14263
rect 13636 14220 13688 14229
rect 17224 14288 17276 14340
rect 20812 14331 20864 14340
rect 20812 14297 20830 14331
rect 20830 14297 20864 14331
rect 20812 14288 20864 14297
rect 16212 14263 16264 14272
rect 16212 14229 16221 14263
rect 16221 14229 16255 14263
rect 16255 14229 16264 14263
rect 16212 14220 16264 14229
rect 19064 14220 19116 14272
rect 19800 14220 19852 14272
rect 6148 14118 6200 14170
rect 6212 14118 6264 14170
rect 6276 14118 6328 14170
rect 6340 14118 6392 14170
rect 6404 14118 6456 14170
rect 11346 14118 11398 14170
rect 11410 14118 11462 14170
rect 11474 14118 11526 14170
rect 11538 14118 11590 14170
rect 11602 14118 11654 14170
rect 16544 14118 16596 14170
rect 16608 14118 16660 14170
rect 16672 14118 16724 14170
rect 16736 14118 16788 14170
rect 16800 14118 16852 14170
rect 21742 14118 21794 14170
rect 21806 14118 21858 14170
rect 21870 14118 21922 14170
rect 21934 14118 21986 14170
rect 21998 14118 22050 14170
rect 2136 14016 2188 14068
rect 4160 14016 4212 14068
rect 4528 14059 4580 14068
rect 4528 14025 4537 14059
rect 4537 14025 4571 14059
rect 4571 14025 4580 14059
rect 4528 14016 4580 14025
rect 5356 14059 5408 14068
rect 5356 14025 5365 14059
rect 5365 14025 5399 14059
rect 5399 14025 5408 14059
rect 5356 14016 5408 14025
rect 5724 14059 5776 14068
rect 5724 14025 5733 14059
rect 5733 14025 5767 14059
rect 5767 14025 5776 14059
rect 5724 14016 5776 14025
rect 6552 14016 6604 14068
rect 7288 14059 7340 14068
rect 7288 14025 7297 14059
rect 7297 14025 7331 14059
rect 7331 14025 7340 14059
rect 7288 14016 7340 14025
rect 7748 14059 7800 14068
rect 7748 14025 7757 14059
rect 7757 14025 7791 14059
rect 7791 14025 7800 14059
rect 7748 14016 7800 14025
rect 7196 13948 7248 14000
rect 8668 13948 8720 14000
rect 6736 13923 6788 13932
rect 6736 13889 6745 13923
rect 6745 13889 6779 13923
rect 6779 13889 6788 13923
rect 6736 13880 6788 13889
rect 7656 13923 7708 13932
rect 5172 13812 5224 13864
rect 6092 13855 6144 13864
rect 6092 13821 6101 13855
rect 6101 13821 6135 13855
rect 6135 13821 6144 13855
rect 6092 13812 6144 13821
rect 5448 13744 5500 13796
rect 4804 13676 4856 13728
rect 7656 13889 7665 13923
rect 7665 13889 7699 13923
rect 7699 13889 7708 13923
rect 7656 13880 7708 13889
rect 9772 14016 9824 14068
rect 10416 14016 10468 14068
rect 11060 14059 11112 14068
rect 11060 14025 11069 14059
rect 11069 14025 11103 14059
rect 11103 14025 11112 14059
rect 11060 14016 11112 14025
rect 11244 14059 11296 14068
rect 11244 14025 11253 14059
rect 11253 14025 11287 14059
rect 11287 14025 11296 14059
rect 11244 14016 11296 14025
rect 10324 13948 10376 14000
rect 7380 13812 7432 13864
rect 9772 13880 9824 13932
rect 12532 14016 12584 14068
rect 13636 14016 13688 14068
rect 15108 14059 15160 14068
rect 15108 14025 15117 14059
rect 15117 14025 15151 14059
rect 15151 14025 15160 14059
rect 15108 14016 15160 14025
rect 17224 14016 17276 14068
rect 12348 13948 12400 14000
rect 10232 13855 10284 13864
rect 7288 13676 7340 13728
rect 7564 13676 7616 13728
rect 10232 13821 10241 13855
rect 10241 13821 10275 13855
rect 10275 13821 10284 13855
rect 10232 13812 10284 13821
rect 10508 13812 10560 13864
rect 10876 13812 10928 13864
rect 11796 13812 11848 13864
rect 11980 13812 12032 13864
rect 13544 13880 13596 13932
rect 18696 13948 18748 14000
rect 18972 13948 19024 14000
rect 16396 13880 16448 13932
rect 20720 14016 20772 14068
rect 21272 14016 21324 14068
rect 21548 14059 21600 14068
rect 21548 14025 21557 14059
rect 21557 14025 21591 14059
rect 21591 14025 21600 14059
rect 21548 14016 21600 14025
rect 20260 13880 20312 13932
rect 13360 13812 13412 13864
rect 9680 13744 9732 13796
rect 10048 13787 10100 13796
rect 10048 13753 10057 13787
rect 10057 13753 10091 13787
rect 10091 13753 10100 13787
rect 10048 13744 10100 13753
rect 17960 13812 18012 13864
rect 10600 13676 10652 13728
rect 10876 13719 10928 13728
rect 10876 13685 10885 13719
rect 10885 13685 10919 13719
rect 10919 13685 10928 13719
rect 10876 13676 10928 13685
rect 12256 13676 12308 13728
rect 13544 13676 13596 13728
rect 14280 13676 14332 13728
rect 3549 13574 3601 13626
rect 3613 13574 3665 13626
rect 3677 13574 3729 13626
rect 3741 13574 3793 13626
rect 3805 13574 3857 13626
rect 8747 13574 8799 13626
rect 8811 13574 8863 13626
rect 8875 13574 8927 13626
rect 8939 13574 8991 13626
rect 9003 13574 9055 13626
rect 13945 13574 13997 13626
rect 14009 13574 14061 13626
rect 14073 13574 14125 13626
rect 14137 13574 14189 13626
rect 14201 13574 14253 13626
rect 19143 13574 19195 13626
rect 19207 13574 19259 13626
rect 19271 13574 19323 13626
rect 19335 13574 19387 13626
rect 19399 13574 19451 13626
rect 4804 13472 4856 13524
rect 5540 13472 5592 13524
rect 6828 13472 6880 13524
rect 7104 13515 7156 13524
rect 7104 13481 7113 13515
rect 7113 13481 7147 13515
rect 7147 13481 7156 13515
rect 7104 13472 7156 13481
rect 9680 13472 9732 13524
rect 5080 13404 5132 13456
rect 5448 13404 5500 13456
rect 4712 13379 4764 13388
rect 4712 13345 4721 13379
rect 4721 13345 4755 13379
rect 4755 13345 4764 13379
rect 4712 13336 4764 13345
rect 6552 13379 6604 13388
rect 6552 13345 6561 13379
rect 6561 13345 6595 13379
rect 6595 13345 6604 13379
rect 6552 13336 6604 13345
rect 7748 13404 7800 13456
rect 7472 13379 7524 13388
rect 7472 13345 7481 13379
rect 7481 13345 7515 13379
rect 7515 13345 7524 13379
rect 7472 13336 7524 13345
rect 3332 13268 3384 13320
rect 9496 13404 9548 13456
rect 8668 13379 8720 13388
rect 8668 13345 8677 13379
rect 8677 13345 8711 13379
rect 8711 13345 8720 13379
rect 8668 13336 8720 13345
rect 8208 13268 8260 13320
rect 5356 13200 5408 13252
rect 6920 13200 6972 13252
rect 10968 13336 11020 13388
rect 12440 13404 12492 13456
rect 13820 13472 13872 13524
rect 14372 13472 14424 13524
rect 15016 13472 15068 13524
rect 21456 13515 21508 13524
rect 21456 13481 21465 13515
rect 21465 13481 21499 13515
rect 21499 13481 21508 13515
rect 21456 13472 21508 13481
rect 15568 13404 15620 13456
rect 11980 13336 12032 13388
rect 11520 13311 11572 13320
rect 11520 13277 11529 13311
rect 11529 13277 11563 13311
rect 11563 13277 11572 13311
rect 11520 13268 11572 13277
rect 12532 13311 12584 13320
rect 12532 13277 12541 13311
rect 12541 13277 12575 13311
rect 12575 13277 12584 13311
rect 12532 13268 12584 13277
rect 12808 13243 12860 13252
rect 12808 13209 12842 13243
rect 12842 13209 12860 13243
rect 17408 13268 17460 13320
rect 12808 13200 12860 13209
rect 18052 13200 18104 13252
rect 19708 13268 19760 13320
rect 20720 13268 20772 13320
rect 20628 13200 20680 13252
rect 1952 13175 2004 13184
rect 1952 13141 1961 13175
rect 1961 13141 1995 13175
rect 1995 13141 2004 13175
rect 1952 13132 2004 13141
rect 6736 13175 6788 13184
rect 6736 13141 6745 13175
rect 6745 13141 6779 13175
rect 6779 13141 6788 13175
rect 6736 13132 6788 13141
rect 7564 13175 7616 13184
rect 7564 13141 7573 13175
rect 7573 13141 7607 13175
rect 7607 13141 7616 13175
rect 8392 13175 8444 13184
rect 7564 13132 7616 13141
rect 8392 13141 8401 13175
rect 8401 13141 8435 13175
rect 8435 13141 8444 13175
rect 8392 13132 8444 13141
rect 9312 13132 9364 13184
rect 9404 13132 9456 13184
rect 9588 13132 9640 13184
rect 9680 13132 9732 13184
rect 10416 13132 10468 13184
rect 10876 13132 10928 13184
rect 11244 13132 11296 13184
rect 11980 13132 12032 13184
rect 14096 13132 14148 13184
rect 14280 13132 14332 13184
rect 15936 13175 15988 13184
rect 15936 13141 15945 13175
rect 15945 13141 15979 13175
rect 15979 13141 15988 13175
rect 15936 13132 15988 13141
rect 17408 13132 17460 13184
rect 18144 13175 18196 13184
rect 18144 13141 18153 13175
rect 18153 13141 18187 13175
rect 18187 13141 18196 13175
rect 18144 13132 18196 13141
rect 20904 13132 20956 13184
rect 21180 13132 21232 13184
rect 6148 13030 6200 13082
rect 6212 13030 6264 13082
rect 6276 13030 6328 13082
rect 6340 13030 6392 13082
rect 6404 13030 6456 13082
rect 11346 13030 11398 13082
rect 11410 13030 11462 13082
rect 11474 13030 11526 13082
rect 11538 13030 11590 13082
rect 11602 13030 11654 13082
rect 16544 13030 16596 13082
rect 16608 13030 16660 13082
rect 16672 13030 16724 13082
rect 16736 13030 16788 13082
rect 16800 13030 16852 13082
rect 21742 13030 21794 13082
rect 21806 13030 21858 13082
rect 21870 13030 21922 13082
rect 21934 13030 21986 13082
rect 21998 13030 22050 13082
rect 6828 12928 6880 12980
rect 3332 12903 3384 12912
rect 3332 12869 3341 12903
rect 3341 12869 3375 12903
rect 3375 12869 3384 12903
rect 3332 12860 3384 12869
rect 4252 12903 4304 12912
rect 4252 12869 4261 12903
rect 4261 12869 4295 12903
rect 4295 12869 4304 12903
rect 4252 12860 4304 12869
rect 4528 12835 4580 12844
rect 4528 12801 4537 12835
rect 4537 12801 4571 12835
rect 4571 12801 4580 12835
rect 4528 12792 4580 12801
rect 5632 12792 5684 12844
rect 5816 12835 5868 12844
rect 5816 12801 5825 12835
rect 5825 12801 5859 12835
rect 5859 12801 5868 12835
rect 5816 12792 5868 12801
rect 5264 12767 5316 12776
rect 5264 12733 5273 12767
rect 5273 12733 5307 12767
rect 5307 12733 5316 12767
rect 5264 12724 5316 12733
rect 5448 12724 5500 12776
rect 6552 12724 6604 12776
rect 7104 12724 7156 12776
rect 8208 12928 8260 12980
rect 8392 12928 8444 12980
rect 9956 12971 10008 12980
rect 9956 12937 9965 12971
rect 9965 12937 9999 12971
rect 9999 12937 10008 12971
rect 9956 12928 10008 12937
rect 10416 12971 10468 12980
rect 10416 12937 10425 12971
rect 10425 12937 10459 12971
rect 10459 12937 10468 12971
rect 10416 12928 10468 12937
rect 14096 12928 14148 12980
rect 14832 12928 14884 12980
rect 18052 12971 18104 12980
rect 14280 12860 14332 12912
rect 18052 12937 18061 12971
rect 18061 12937 18095 12971
rect 18095 12937 18104 12971
rect 18052 12928 18104 12937
rect 19524 12971 19576 12980
rect 19524 12937 19533 12971
rect 19533 12937 19567 12971
rect 19567 12937 19576 12971
rect 19524 12928 19576 12937
rect 20720 12928 20772 12980
rect 8392 12792 8444 12844
rect 9588 12792 9640 12844
rect 12072 12792 12124 12844
rect 14372 12792 14424 12844
rect 15936 12792 15988 12844
rect 16672 12835 16724 12844
rect 16672 12801 16681 12835
rect 16681 12801 16715 12835
rect 16715 12801 16724 12835
rect 16672 12792 16724 12801
rect 17500 12792 17552 12844
rect 7748 12767 7800 12776
rect 7748 12733 7757 12767
rect 7757 12733 7791 12767
rect 7791 12733 7800 12767
rect 7748 12724 7800 12733
rect 7840 12724 7892 12776
rect 8300 12724 8352 12776
rect 5540 12656 5592 12708
rect 6736 12656 6788 12708
rect 9772 12656 9824 12708
rect 11888 12724 11940 12776
rect 14280 12724 14332 12776
rect 10876 12656 10928 12708
rect 3332 12588 3384 12640
rect 4252 12588 4304 12640
rect 6552 12588 6604 12640
rect 12256 12588 12308 12640
rect 12532 12631 12584 12640
rect 12532 12597 12541 12631
rect 12541 12597 12575 12631
rect 12575 12597 12584 12631
rect 12532 12588 12584 12597
rect 12716 12631 12768 12640
rect 12716 12597 12725 12631
rect 12725 12597 12759 12631
rect 12759 12597 12768 12631
rect 12716 12588 12768 12597
rect 14556 12588 14608 12640
rect 20904 12792 20956 12844
rect 21272 12928 21324 12980
rect 18144 12767 18196 12776
rect 18144 12733 18153 12767
rect 18153 12733 18187 12767
rect 18187 12733 18196 12767
rect 18144 12724 18196 12733
rect 19616 12631 19668 12640
rect 19616 12597 19625 12631
rect 19625 12597 19659 12631
rect 19659 12597 19668 12631
rect 19616 12588 19668 12597
rect 3549 12486 3601 12538
rect 3613 12486 3665 12538
rect 3677 12486 3729 12538
rect 3741 12486 3793 12538
rect 3805 12486 3857 12538
rect 8747 12486 8799 12538
rect 8811 12486 8863 12538
rect 8875 12486 8927 12538
rect 8939 12486 8991 12538
rect 9003 12486 9055 12538
rect 13945 12486 13997 12538
rect 14009 12486 14061 12538
rect 14073 12486 14125 12538
rect 14137 12486 14189 12538
rect 14201 12486 14253 12538
rect 19143 12486 19195 12538
rect 19207 12486 19259 12538
rect 19271 12486 19323 12538
rect 19335 12486 19387 12538
rect 19399 12486 19451 12538
rect 2872 12384 2924 12436
rect 5632 12427 5684 12436
rect 5632 12393 5641 12427
rect 5641 12393 5675 12427
rect 5675 12393 5684 12427
rect 5632 12384 5684 12393
rect 6828 12384 6880 12436
rect 7288 12384 7340 12436
rect 7656 12384 7708 12436
rect 7748 12384 7800 12436
rect 8300 12384 8352 12436
rect 9312 12384 9364 12436
rect 10600 12384 10652 12436
rect 4528 12316 4580 12368
rect 10968 12316 11020 12368
rect 11152 12316 11204 12368
rect 14648 12316 14700 12368
rect 4988 12248 5040 12300
rect 6552 12248 6604 12300
rect 6644 12248 6696 12300
rect 8024 12291 8076 12300
rect 8024 12257 8033 12291
rect 8033 12257 8067 12291
rect 8067 12257 8076 12291
rect 8024 12248 8076 12257
rect 9496 12291 9548 12300
rect 9496 12257 9505 12291
rect 9505 12257 9539 12291
rect 9539 12257 9548 12291
rect 9496 12248 9548 12257
rect 9588 12248 9640 12300
rect 10876 12291 10928 12300
rect 10876 12257 10885 12291
rect 10885 12257 10919 12291
rect 10919 12257 10928 12291
rect 10876 12248 10928 12257
rect 12532 12291 12584 12300
rect 12532 12257 12541 12291
rect 12541 12257 12575 12291
rect 12575 12257 12584 12291
rect 12532 12248 12584 12257
rect 16672 12291 16724 12300
rect 16672 12257 16681 12291
rect 16681 12257 16715 12291
rect 16715 12257 16724 12291
rect 16672 12248 16724 12257
rect 18236 12427 18288 12436
rect 18236 12393 18245 12427
rect 18245 12393 18279 12427
rect 18279 12393 18288 12427
rect 18236 12384 18288 12393
rect 19708 12427 19760 12436
rect 19708 12393 19717 12427
rect 19717 12393 19751 12427
rect 19751 12393 19760 12427
rect 19708 12384 19760 12393
rect 21272 12427 21324 12436
rect 21272 12393 21281 12427
rect 21281 12393 21315 12427
rect 21315 12393 21324 12427
rect 21272 12384 21324 12393
rect 4068 12180 4120 12232
rect 9312 12180 9364 12232
rect 11152 12180 11204 12232
rect 11796 12180 11848 12232
rect 11888 12180 11940 12232
rect 13912 12180 13964 12232
rect 14372 12180 14424 12232
rect 14924 12180 14976 12232
rect 5448 12112 5500 12164
rect 7196 12112 7248 12164
rect 7656 12112 7708 12164
rect 6000 12087 6052 12096
rect 6000 12053 6009 12087
rect 6009 12053 6043 12087
rect 6043 12053 6052 12087
rect 6000 12044 6052 12053
rect 6552 12044 6604 12096
rect 7288 12087 7340 12096
rect 7288 12053 7297 12087
rect 7297 12053 7331 12087
rect 7331 12053 7340 12087
rect 7288 12044 7340 12053
rect 8300 12044 8352 12096
rect 9128 12044 9180 12096
rect 10048 12044 10100 12096
rect 11704 12112 11756 12164
rect 11980 12112 12032 12164
rect 12256 12112 12308 12164
rect 12624 12112 12676 12164
rect 14648 12112 14700 12164
rect 16580 12112 16632 12164
rect 12532 12044 12584 12096
rect 12992 12044 13044 12096
rect 13912 12087 13964 12096
rect 13912 12053 13921 12087
rect 13921 12053 13955 12087
rect 13955 12053 13964 12087
rect 13912 12044 13964 12053
rect 14188 12087 14240 12096
rect 14188 12053 14197 12087
rect 14197 12053 14231 12087
rect 14231 12053 14240 12087
rect 14188 12044 14240 12053
rect 14740 12044 14792 12096
rect 6148 11942 6200 11994
rect 6212 11942 6264 11994
rect 6276 11942 6328 11994
rect 6340 11942 6392 11994
rect 6404 11942 6456 11994
rect 11346 11942 11398 11994
rect 11410 11942 11462 11994
rect 11474 11942 11526 11994
rect 11538 11942 11590 11994
rect 11602 11942 11654 11994
rect 16544 11942 16596 11994
rect 16608 11942 16660 11994
rect 16672 11942 16724 11994
rect 16736 11942 16788 11994
rect 16800 11942 16852 11994
rect 21742 11942 21794 11994
rect 21806 11942 21858 11994
rect 21870 11942 21922 11994
rect 21934 11942 21986 11994
rect 21998 11942 22050 11994
rect 5448 11883 5500 11892
rect 5448 11849 5457 11883
rect 5457 11849 5491 11883
rect 5491 11849 5500 11883
rect 5448 11840 5500 11849
rect 6552 11840 6604 11892
rect 4160 11815 4212 11824
rect 4160 11781 4169 11815
rect 4169 11781 4203 11815
rect 4203 11781 4212 11815
rect 4160 11772 4212 11781
rect 4436 11747 4488 11756
rect 4436 11713 4445 11747
rect 4445 11713 4479 11747
rect 4479 11713 4488 11747
rect 4436 11704 4488 11713
rect 6920 11840 6972 11892
rect 7104 11840 7156 11892
rect 9312 11883 9364 11892
rect 9312 11849 9321 11883
rect 9321 11849 9355 11883
rect 9355 11849 9364 11883
rect 9312 11840 9364 11849
rect 10968 11840 11020 11892
rect 11244 11840 11296 11892
rect 7932 11772 7984 11824
rect 8208 11772 8260 11824
rect 11060 11772 11112 11824
rect 11704 11772 11756 11824
rect 8024 11747 8076 11756
rect 4988 11636 5040 11688
rect 6644 11636 6696 11688
rect 8024 11713 8033 11747
rect 8033 11713 8067 11747
rect 8067 11713 8076 11747
rect 8024 11704 8076 11713
rect 9680 11747 9732 11756
rect 9680 11713 9689 11747
rect 9689 11713 9723 11747
rect 9723 11713 9732 11747
rect 9680 11704 9732 11713
rect 10692 11704 10744 11756
rect 13820 11840 13872 11892
rect 18236 11840 18288 11892
rect 11980 11772 12032 11824
rect 14556 11772 14608 11824
rect 11888 11747 11940 11756
rect 11888 11713 11897 11747
rect 11897 11713 11931 11747
rect 11931 11713 11940 11747
rect 11888 11704 11940 11713
rect 12716 11704 12768 11756
rect 5632 11568 5684 11620
rect 7104 11636 7156 11688
rect 7472 11636 7524 11688
rect 7932 11679 7984 11688
rect 7932 11645 7941 11679
rect 7941 11645 7975 11679
rect 7975 11645 7984 11679
rect 7932 11636 7984 11645
rect 9956 11679 10008 11688
rect 9956 11645 9965 11679
rect 9965 11645 9999 11679
rect 9999 11645 10008 11679
rect 9956 11636 10008 11645
rect 10784 11679 10836 11688
rect 10784 11645 10793 11679
rect 10793 11645 10827 11679
rect 10827 11645 10836 11679
rect 10784 11636 10836 11645
rect 11336 11636 11388 11688
rect 12256 11636 12308 11688
rect 15108 11704 15160 11756
rect 16396 11704 16448 11756
rect 19892 11704 19944 11756
rect 21272 11840 21324 11892
rect 9864 11568 9916 11620
rect 10968 11568 11020 11620
rect 6368 11500 6420 11552
rect 7748 11500 7800 11552
rect 8300 11500 8352 11552
rect 9036 11500 9088 11552
rect 10232 11500 10284 11552
rect 11152 11543 11204 11552
rect 11152 11509 11161 11543
rect 11161 11509 11195 11543
rect 11195 11509 11204 11543
rect 11152 11500 11204 11509
rect 11796 11568 11848 11620
rect 12072 11500 12124 11552
rect 13728 11500 13780 11552
rect 14188 11636 14240 11688
rect 16304 11500 16356 11552
rect 18880 11543 18932 11552
rect 18880 11509 18889 11543
rect 18889 11509 18923 11543
rect 18923 11509 18932 11543
rect 18880 11500 18932 11509
rect 18972 11500 19024 11552
rect 3549 11398 3601 11450
rect 3613 11398 3665 11450
rect 3677 11398 3729 11450
rect 3741 11398 3793 11450
rect 3805 11398 3857 11450
rect 8747 11398 8799 11450
rect 8811 11398 8863 11450
rect 8875 11398 8927 11450
rect 8939 11398 8991 11450
rect 9003 11398 9055 11450
rect 13945 11398 13997 11450
rect 14009 11398 14061 11450
rect 14073 11398 14125 11450
rect 14137 11398 14189 11450
rect 14201 11398 14253 11450
rect 19143 11398 19195 11450
rect 19207 11398 19259 11450
rect 19271 11398 19323 11450
rect 19335 11398 19387 11450
rect 19399 11398 19451 11450
rect 2780 11296 2832 11348
rect 5540 11296 5592 11348
rect 6000 11296 6052 11348
rect 7012 11339 7064 11348
rect 7012 11305 7021 11339
rect 7021 11305 7055 11339
rect 7055 11305 7064 11339
rect 7012 11296 7064 11305
rect 7104 11296 7156 11348
rect 10048 11339 10100 11348
rect 10048 11305 10057 11339
rect 10057 11305 10091 11339
rect 10091 11305 10100 11339
rect 10048 11296 10100 11305
rect 10968 11296 11020 11348
rect 11336 11339 11388 11348
rect 11336 11305 11345 11339
rect 11345 11305 11379 11339
rect 11379 11305 11388 11339
rect 11336 11296 11388 11305
rect 3056 11228 3108 11280
rect 4436 11228 4488 11280
rect 9312 11228 9364 11280
rect 4344 11160 4396 11212
rect 5448 11160 5500 11212
rect 5632 11203 5684 11212
rect 5632 11169 5641 11203
rect 5641 11169 5675 11203
rect 5675 11169 5684 11203
rect 5632 11160 5684 11169
rect 6000 11160 6052 11212
rect 9404 11160 9456 11212
rect 10508 11203 10560 11212
rect 3056 11092 3108 11144
rect 4436 11092 4488 11144
rect 6552 11092 6604 11144
rect 6644 11092 6696 11144
rect 8300 11092 8352 11144
rect 8576 11092 8628 11144
rect 10508 11169 10517 11203
rect 10517 11169 10551 11203
rect 10551 11169 10560 11203
rect 10508 11160 10560 11169
rect 10692 11228 10744 11280
rect 12440 11296 12492 11348
rect 14280 11296 14332 11348
rect 20260 11296 20312 11348
rect 13176 11228 13228 11280
rect 13544 11228 13596 11280
rect 14740 11228 14792 11280
rect 16764 11228 16816 11280
rect 12532 11160 12584 11212
rect 14372 11160 14424 11212
rect 12808 11092 12860 11144
rect 15108 11092 15160 11144
rect 16304 11135 16356 11144
rect 16304 11101 16313 11135
rect 16313 11101 16347 11135
rect 16347 11101 16356 11135
rect 16304 11092 16356 11101
rect 3240 11024 3292 11076
rect 4252 11067 4304 11076
rect 4252 11033 4261 11067
rect 4261 11033 4295 11067
rect 4295 11033 4304 11067
rect 4252 11024 4304 11033
rect 4988 11067 5040 11076
rect 4988 11033 4997 11067
rect 4997 11033 5031 11067
rect 5031 11033 5040 11067
rect 4988 11024 5040 11033
rect 9772 11024 9824 11076
rect 9956 11024 10008 11076
rect 11060 11067 11112 11076
rect 4804 10956 4856 11008
rect 6368 10956 6420 11008
rect 6552 10999 6604 11008
rect 6552 10965 6561 10999
rect 6561 10965 6595 10999
rect 6595 10965 6604 10999
rect 6552 10956 6604 10965
rect 6644 10999 6696 11008
rect 6644 10965 6653 10999
rect 6653 10965 6687 10999
rect 6687 10965 6696 10999
rect 8576 10999 8628 11008
rect 6644 10956 6696 10965
rect 8576 10965 8585 10999
rect 8585 10965 8619 10999
rect 8619 10965 8628 10999
rect 8576 10956 8628 10965
rect 9404 10999 9456 11008
rect 9404 10965 9413 10999
rect 9413 10965 9447 10999
rect 9447 10965 9456 10999
rect 9404 10956 9456 10965
rect 10232 10956 10284 11008
rect 11060 11033 11069 11067
rect 11069 11033 11103 11067
rect 11103 11033 11112 11067
rect 11060 11024 11112 11033
rect 11244 11024 11296 11076
rect 12256 11024 12308 11076
rect 12716 11024 12768 11076
rect 14464 11024 14516 11076
rect 11980 10956 12032 11008
rect 12440 10956 12492 11008
rect 15200 10956 15252 11008
rect 17684 11024 17736 11076
rect 18144 11067 18196 11076
rect 18144 11033 18153 11067
rect 18153 11033 18187 11067
rect 18187 11033 18196 11067
rect 18144 11024 18196 11033
rect 20996 11203 21048 11212
rect 20996 11169 21005 11203
rect 21005 11169 21039 11203
rect 21039 11169 21048 11203
rect 21272 11296 21324 11348
rect 20996 11160 21048 11169
rect 19524 11024 19576 11076
rect 6148 10854 6200 10906
rect 6212 10854 6264 10906
rect 6276 10854 6328 10906
rect 6340 10854 6392 10906
rect 6404 10854 6456 10906
rect 11346 10854 11398 10906
rect 11410 10854 11462 10906
rect 11474 10854 11526 10906
rect 11538 10854 11590 10906
rect 11602 10854 11654 10906
rect 16544 10854 16596 10906
rect 16608 10854 16660 10906
rect 16672 10854 16724 10906
rect 16736 10854 16788 10906
rect 16800 10854 16852 10906
rect 21742 10854 21794 10906
rect 21806 10854 21858 10906
rect 21870 10854 21922 10906
rect 21934 10854 21986 10906
rect 21998 10854 22050 10906
rect 3424 10752 3476 10804
rect 5172 10752 5224 10804
rect 6644 10752 6696 10804
rect 3332 10684 3384 10736
rect 7932 10752 7984 10804
rect 8484 10752 8536 10804
rect 8576 10752 8628 10804
rect 9036 10795 9088 10804
rect 9036 10761 9045 10795
rect 9045 10761 9079 10795
rect 9079 10761 9088 10795
rect 9036 10752 9088 10761
rect 9404 10752 9456 10804
rect 9680 10752 9732 10804
rect 10692 10752 10744 10804
rect 16396 10752 16448 10804
rect 10140 10684 10192 10736
rect 10508 10684 10560 10736
rect 5540 10659 5592 10668
rect 5540 10625 5549 10659
rect 5549 10625 5583 10659
rect 5583 10625 5592 10659
rect 5540 10616 5592 10625
rect 5724 10616 5776 10668
rect 2780 10548 2832 10600
rect 4436 10591 4488 10600
rect 4436 10557 4445 10591
rect 4445 10557 4479 10591
rect 4479 10557 4488 10591
rect 4436 10548 4488 10557
rect 5448 10591 5500 10600
rect 5448 10557 5457 10591
rect 5457 10557 5491 10591
rect 5491 10557 5500 10591
rect 5448 10548 5500 10557
rect 6920 10616 6972 10668
rect 7196 10616 7248 10668
rect 5908 10480 5960 10532
rect 6828 10548 6880 10600
rect 8392 10548 8444 10600
rect 9312 10616 9364 10668
rect 10048 10616 10100 10668
rect 8576 10591 8628 10600
rect 8576 10557 8585 10591
rect 8585 10557 8619 10591
rect 8619 10557 8628 10591
rect 8576 10548 8628 10557
rect 9588 10548 9640 10600
rect 10784 10591 10836 10600
rect 9128 10480 9180 10532
rect 10784 10557 10793 10591
rect 10793 10557 10827 10591
rect 10827 10557 10836 10591
rect 10784 10548 10836 10557
rect 10876 10591 10928 10600
rect 10876 10557 10885 10591
rect 10885 10557 10919 10591
rect 10919 10557 10928 10591
rect 12440 10684 12492 10736
rect 12808 10684 12860 10736
rect 13728 10684 13780 10736
rect 14464 10727 14516 10736
rect 14464 10693 14473 10727
rect 14473 10693 14507 10727
rect 14507 10693 14516 10727
rect 14464 10684 14516 10693
rect 15568 10684 15620 10736
rect 13636 10616 13688 10668
rect 15108 10659 15160 10668
rect 15108 10625 15117 10659
rect 15117 10625 15151 10659
rect 15151 10625 15160 10659
rect 15108 10616 15160 10625
rect 16304 10616 16356 10668
rect 16948 10752 17000 10804
rect 20996 10795 21048 10804
rect 20996 10761 21005 10795
rect 21005 10761 21039 10795
rect 21039 10761 21048 10795
rect 20996 10752 21048 10761
rect 10876 10548 10928 10557
rect 11704 10548 11756 10600
rect 20076 10616 20128 10668
rect 3976 10455 4028 10464
rect 3976 10421 3985 10455
rect 3985 10421 4019 10455
rect 4019 10421 4028 10455
rect 3976 10412 4028 10421
rect 7196 10412 7248 10464
rect 9312 10412 9364 10464
rect 9864 10412 9916 10464
rect 11612 10412 11664 10464
rect 12992 10412 13044 10464
rect 13728 10412 13780 10464
rect 14648 10412 14700 10464
rect 17960 10548 18012 10600
rect 19708 10480 19760 10532
rect 19524 10412 19576 10464
rect 3549 10310 3601 10362
rect 3613 10310 3665 10362
rect 3677 10310 3729 10362
rect 3741 10310 3793 10362
rect 3805 10310 3857 10362
rect 8747 10310 8799 10362
rect 8811 10310 8863 10362
rect 8875 10310 8927 10362
rect 8939 10310 8991 10362
rect 9003 10310 9055 10362
rect 13945 10310 13997 10362
rect 14009 10310 14061 10362
rect 14073 10310 14125 10362
rect 14137 10310 14189 10362
rect 14201 10310 14253 10362
rect 19143 10310 19195 10362
rect 19207 10310 19259 10362
rect 19271 10310 19323 10362
rect 19335 10310 19387 10362
rect 19399 10310 19451 10362
rect 1768 10208 1820 10260
rect 2964 10208 3016 10260
rect 3332 10208 3384 10260
rect 4068 10208 4120 10260
rect 4436 10208 4488 10260
rect 5448 10208 5500 10260
rect 5816 10208 5868 10260
rect 6552 10208 6604 10260
rect 7104 10208 7156 10260
rect 7564 10208 7616 10260
rect 8024 10208 8076 10260
rect 10140 10251 10192 10260
rect 10140 10217 10149 10251
rect 10149 10217 10183 10251
rect 10183 10217 10192 10251
rect 10140 10208 10192 10217
rect 11612 10208 11664 10260
rect 12532 10208 12584 10260
rect 13728 10208 13780 10260
rect 3792 10072 3844 10124
rect 2780 10047 2832 10056
rect 2780 10013 2789 10047
rect 2789 10013 2823 10047
rect 2823 10013 2832 10047
rect 2780 10004 2832 10013
rect 3700 10004 3752 10056
rect 4620 10072 4672 10124
rect 5540 10115 5592 10124
rect 5540 10081 5549 10115
rect 5549 10081 5583 10115
rect 5583 10081 5592 10115
rect 5540 10072 5592 10081
rect 6000 10072 6052 10124
rect 5080 10004 5132 10056
rect 5264 10047 5316 10056
rect 5264 10013 5273 10047
rect 5273 10013 5307 10047
rect 5307 10013 5316 10047
rect 5264 10004 5316 10013
rect 9312 10140 9364 10192
rect 12164 10140 12216 10192
rect 12348 10140 12400 10192
rect 13452 10140 13504 10192
rect 6644 10115 6696 10124
rect 6644 10081 6653 10115
rect 6653 10081 6687 10115
rect 6687 10081 6696 10115
rect 6644 10072 6696 10081
rect 6736 10072 6788 10124
rect 8116 10115 8168 10124
rect 8116 10081 8125 10115
rect 8125 10081 8159 10115
rect 8159 10081 8168 10115
rect 8116 10072 8168 10081
rect 8576 10072 8628 10124
rect 9404 10115 9456 10124
rect 9404 10081 9413 10115
rect 9413 10081 9447 10115
rect 9447 10081 9456 10115
rect 9404 10072 9456 10081
rect 9588 10115 9640 10124
rect 9588 10081 9597 10115
rect 9597 10081 9631 10115
rect 9631 10081 9640 10115
rect 9588 10072 9640 10081
rect 13728 10072 13780 10124
rect 8392 10047 8444 10056
rect 8392 10013 8401 10047
rect 8401 10013 8435 10047
rect 8435 10013 8444 10047
rect 8392 10004 8444 10013
rect 10048 10004 10100 10056
rect 12072 10004 12124 10056
rect 12440 10004 12492 10056
rect 14464 10208 14516 10260
rect 14924 10208 14976 10260
rect 20996 10251 21048 10260
rect 20996 10217 21005 10251
rect 21005 10217 21039 10251
rect 21039 10217 21048 10251
rect 20996 10208 21048 10217
rect 14464 10047 14516 10056
rect 14464 10013 14498 10047
rect 14498 10013 14516 10047
rect 14464 10004 14516 10013
rect 15292 10004 15344 10056
rect 3424 9936 3476 9988
rect 4988 9936 5040 9988
rect 1768 9868 1820 9920
rect 2964 9868 3016 9920
rect 5540 9868 5592 9920
rect 6092 9911 6144 9920
rect 6092 9877 6101 9911
rect 6101 9877 6135 9911
rect 6135 9877 6144 9911
rect 6092 9868 6144 9877
rect 6276 9936 6328 9988
rect 8024 9936 8076 9988
rect 7012 9868 7064 9920
rect 7748 9911 7800 9920
rect 7748 9877 7757 9911
rect 7757 9877 7791 9911
rect 7791 9877 7800 9911
rect 7748 9868 7800 9877
rect 8208 9868 8260 9920
rect 10784 9936 10836 9988
rect 9772 9911 9824 9920
rect 9772 9877 9781 9911
rect 9781 9877 9815 9911
rect 9815 9877 9824 9911
rect 9772 9868 9824 9877
rect 10600 9911 10652 9920
rect 10600 9877 10609 9911
rect 10609 9877 10643 9911
rect 10643 9877 10652 9911
rect 10600 9868 10652 9877
rect 12716 9868 12768 9920
rect 13360 9936 13412 9988
rect 16304 9936 16356 9988
rect 16948 10004 17000 10056
rect 17960 10004 18012 10056
rect 19616 10072 19668 10124
rect 13912 9868 13964 9920
rect 15568 9911 15620 9920
rect 15568 9877 15577 9911
rect 15577 9877 15611 9911
rect 15611 9877 15620 9911
rect 15568 9868 15620 9877
rect 15660 9911 15712 9920
rect 15660 9877 15669 9911
rect 15669 9877 15703 9911
rect 15703 9877 15712 9911
rect 19892 10004 19944 10056
rect 19340 9936 19392 9988
rect 20536 9936 20588 9988
rect 18512 9911 18564 9920
rect 15660 9868 15712 9877
rect 18512 9877 18521 9911
rect 18521 9877 18555 9911
rect 18555 9877 18564 9911
rect 18512 9868 18564 9877
rect 19156 9868 19208 9920
rect 6148 9766 6200 9818
rect 6212 9766 6264 9818
rect 6276 9766 6328 9818
rect 6340 9766 6392 9818
rect 6404 9766 6456 9818
rect 11346 9766 11398 9818
rect 11410 9766 11462 9818
rect 11474 9766 11526 9818
rect 11538 9766 11590 9818
rect 11602 9766 11654 9818
rect 16544 9766 16596 9818
rect 16608 9766 16660 9818
rect 16672 9766 16724 9818
rect 16736 9766 16788 9818
rect 16800 9766 16852 9818
rect 21742 9766 21794 9818
rect 21806 9766 21858 9818
rect 21870 9766 21922 9818
rect 21934 9766 21986 9818
rect 21998 9766 22050 9818
rect 2780 9664 2832 9716
rect 3792 9664 3844 9716
rect 3884 9664 3936 9716
rect 9404 9664 9456 9716
rect 2136 9571 2188 9580
rect 2136 9537 2145 9571
rect 2145 9537 2179 9571
rect 2179 9537 2188 9571
rect 2136 9528 2188 9537
rect 6184 9596 6236 9648
rect 6368 9596 6420 9648
rect 9772 9596 9824 9648
rect 10784 9664 10836 9716
rect 12072 9707 12124 9716
rect 10968 9596 11020 9648
rect 12072 9673 12081 9707
rect 12081 9673 12115 9707
rect 12115 9673 12124 9707
rect 12072 9664 12124 9673
rect 13636 9707 13688 9716
rect 13636 9673 13645 9707
rect 13645 9673 13679 9707
rect 13679 9673 13688 9707
rect 13636 9664 13688 9673
rect 15016 9664 15068 9716
rect 19340 9664 19392 9716
rect 14648 9596 14700 9648
rect 2872 9571 2924 9580
rect 2872 9537 2881 9571
rect 2881 9537 2915 9571
rect 2915 9537 2924 9571
rect 2872 9528 2924 9537
rect 4160 9528 4212 9580
rect 3792 9503 3844 9512
rect 3792 9469 3801 9503
rect 3801 9469 3835 9503
rect 3835 9469 3844 9503
rect 3792 9460 3844 9469
rect 4344 9460 4396 9512
rect 1584 9435 1636 9444
rect 1584 9401 1593 9435
rect 1593 9401 1627 9435
rect 1627 9401 1636 9435
rect 1584 9392 1636 9401
rect 1860 9392 1912 9444
rect 3148 9392 3200 9444
rect 4436 9392 4488 9444
rect 5264 9528 5316 9580
rect 5540 9528 5592 9580
rect 6092 9571 6144 9580
rect 6092 9537 6101 9571
rect 6101 9537 6135 9571
rect 6135 9537 6144 9571
rect 6092 9528 6144 9537
rect 6276 9528 6328 9580
rect 5632 9460 5684 9512
rect 9128 9503 9180 9512
rect 5356 9392 5408 9444
rect 5816 9392 5868 9444
rect 6368 9392 6420 9444
rect 9128 9469 9137 9503
rect 9137 9469 9171 9503
rect 9171 9469 9180 9503
rect 9128 9460 9180 9469
rect 12440 9528 12492 9580
rect 12716 9528 12768 9580
rect 13636 9528 13688 9580
rect 15108 9528 15160 9580
rect 15660 9528 15712 9580
rect 16488 9571 16540 9580
rect 16488 9537 16497 9571
rect 16497 9537 16531 9571
rect 16531 9537 16540 9571
rect 16488 9528 16540 9537
rect 17776 9571 17828 9580
rect 19616 9596 19668 9648
rect 20168 9596 20220 9648
rect 17776 9537 17794 9571
rect 17794 9537 17828 9571
rect 17776 9528 17828 9537
rect 18880 9528 18932 9580
rect 6736 9392 6788 9444
rect 7840 9392 7892 9444
rect 3700 9324 3752 9376
rect 3884 9324 3936 9376
rect 4988 9324 5040 9376
rect 5632 9324 5684 9376
rect 7012 9324 7064 9376
rect 7748 9324 7800 9376
rect 8392 9324 8444 9376
rect 8484 9324 8536 9376
rect 9680 9435 9732 9444
rect 9680 9401 9689 9435
rect 9689 9401 9723 9435
rect 9723 9401 9732 9435
rect 9680 9392 9732 9401
rect 10048 9392 10100 9444
rect 10140 9324 10192 9376
rect 10876 9460 10928 9512
rect 11060 9392 11112 9444
rect 11888 9392 11940 9444
rect 12256 9392 12308 9444
rect 11612 9324 11664 9376
rect 12164 9367 12216 9376
rect 12164 9333 12173 9367
rect 12173 9333 12207 9367
rect 12207 9333 12216 9367
rect 12164 9324 12216 9333
rect 13820 9460 13872 9512
rect 18052 9503 18104 9512
rect 18052 9469 18061 9503
rect 18061 9469 18095 9503
rect 18095 9469 18104 9503
rect 18052 9460 18104 9469
rect 19156 9460 19208 9512
rect 14004 9392 14056 9444
rect 13912 9324 13964 9376
rect 14832 9324 14884 9376
rect 16948 9324 17000 9376
rect 20812 9324 20864 9376
rect 21272 9367 21324 9376
rect 21272 9333 21281 9367
rect 21281 9333 21315 9367
rect 21315 9333 21324 9367
rect 21272 9324 21324 9333
rect 3549 9222 3601 9274
rect 3613 9222 3665 9274
rect 3677 9222 3729 9274
rect 3741 9222 3793 9274
rect 3805 9222 3857 9274
rect 8747 9222 8799 9274
rect 8811 9222 8863 9274
rect 8875 9222 8927 9274
rect 8939 9222 8991 9274
rect 9003 9222 9055 9274
rect 13945 9222 13997 9274
rect 14009 9222 14061 9274
rect 14073 9222 14125 9274
rect 14137 9222 14189 9274
rect 14201 9222 14253 9274
rect 19143 9222 19195 9274
rect 19207 9222 19259 9274
rect 19271 9222 19323 9274
rect 19335 9222 19387 9274
rect 19399 9222 19451 9274
rect 1676 9163 1728 9172
rect 1676 9129 1685 9163
rect 1685 9129 1719 9163
rect 1719 9129 1728 9163
rect 1676 9120 1728 9129
rect 2044 9120 2096 9172
rect 2228 9052 2280 9104
rect 2504 8984 2556 9036
rect 1676 8916 1728 8968
rect 5908 9120 5960 9172
rect 6552 9120 6604 9172
rect 8024 9120 8076 9172
rect 9588 9120 9640 9172
rect 9864 9120 9916 9172
rect 3240 9027 3292 9036
rect 3240 8993 3249 9027
rect 3249 8993 3283 9027
rect 3283 8993 3292 9027
rect 3240 8984 3292 8993
rect 3976 8984 4028 9036
rect 4620 9027 4672 9036
rect 4344 8959 4396 8968
rect 4344 8925 4353 8959
rect 4353 8925 4387 8959
rect 4387 8925 4396 8959
rect 4344 8916 4396 8925
rect 4620 8993 4629 9027
rect 4629 8993 4663 9027
rect 4663 8993 4672 9027
rect 4620 8984 4672 8993
rect 5080 9052 5132 9104
rect 7840 9052 7892 9104
rect 8208 9052 8260 9104
rect 11796 9120 11848 9172
rect 3148 8848 3200 8900
rect 3424 8848 3476 8900
rect 5080 8848 5132 8900
rect 6092 8984 6144 9036
rect 6828 9027 6880 9036
rect 6828 8993 6837 9027
rect 6837 8993 6871 9027
rect 6871 8993 6880 9027
rect 6828 8984 6880 8993
rect 7656 9027 7708 9036
rect 7656 8993 7665 9027
rect 7665 8993 7699 9027
rect 7699 8993 7708 9027
rect 7656 8984 7708 8993
rect 8116 8984 8168 9036
rect 9588 8984 9640 9036
rect 7472 8916 7524 8968
rect 9956 8916 10008 8968
rect 10140 9027 10192 9036
rect 10140 8993 10149 9027
rect 10149 8993 10183 9027
rect 10183 8993 10192 9027
rect 10324 9027 10376 9036
rect 10140 8984 10192 8993
rect 10324 8993 10333 9027
rect 10333 8993 10367 9027
rect 10367 8993 10376 9027
rect 10324 8984 10376 8993
rect 10692 9027 10744 9036
rect 10692 8993 10701 9027
rect 10701 8993 10735 9027
rect 10735 8993 10744 9027
rect 10692 8984 10744 8993
rect 13636 9120 13688 9172
rect 10600 8916 10652 8968
rect 5724 8891 5776 8900
rect 5724 8857 5733 8891
rect 5733 8857 5767 8891
rect 5767 8857 5776 8891
rect 5724 8848 5776 8857
rect 3700 8780 3752 8832
rect 7288 8848 7340 8900
rect 6184 8823 6236 8832
rect 6184 8789 6193 8823
rect 6193 8789 6227 8823
rect 6227 8789 6236 8823
rect 6184 8780 6236 8789
rect 6552 8823 6604 8832
rect 6552 8789 6561 8823
rect 6561 8789 6595 8823
rect 6595 8789 6604 8823
rect 6552 8780 6604 8789
rect 6644 8823 6696 8832
rect 6644 8789 6653 8823
rect 6653 8789 6687 8823
rect 6687 8789 6696 8823
rect 7472 8823 7524 8832
rect 6644 8780 6696 8789
rect 7472 8789 7481 8823
rect 7481 8789 7515 8823
rect 7515 8789 7524 8823
rect 7472 8780 7524 8789
rect 9128 8848 9180 8900
rect 9496 8848 9548 8900
rect 9588 8848 9640 8900
rect 13820 9027 13872 9036
rect 13820 8993 13829 9027
rect 13829 8993 13863 9027
rect 13863 8993 13872 9027
rect 15752 9120 15804 9172
rect 16488 9120 16540 9172
rect 18052 9120 18104 9172
rect 19064 9120 19116 9172
rect 13820 8984 13872 8993
rect 18880 8916 18932 8968
rect 8208 8823 8260 8832
rect 8208 8789 8217 8823
rect 8217 8789 8251 8823
rect 8251 8789 8260 8823
rect 8208 8780 8260 8789
rect 8576 8780 8628 8832
rect 8668 8823 8720 8832
rect 8668 8789 8677 8823
rect 8677 8789 8711 8823
rect 8711 8789 8720 8823
rect 8668 8780 8720 8789
rect 10508 8780 10560 8832
rect 10876 8823 10928 8832
rect 10876 8789 10885 8823
rect 10885 8789 10919 8823
rect 10919 8789 10928 8823
rect 10876 8780 10928 8789
rect 13268 8848 13320 8900
rect 13544 8848 13596 8900
rect 11336 8823 11388 8832
rect 11336 8789 11345 8823
rect 11345 8789 11379 8823
rect 11379 8789 11388 8823
rect 11796 8823 11848 8832
rect 11336 8780 11388 8789
rect 11796 8789 11805 8823
rect 11805 8789 11839 8823
rect 11839 8789 11848 8823
rect 11796 8780 11848 8789
rect 12440 8780 12492 8832
rect 16212 8848 16264 8900
rect 15292 8780 15344 8832
rect 16948 8848 17000 8900
rect 20076 8916 20128 8968
rect 19708 8848 19760 8900
rect 17040 8780 17092 8832
rect 17592 8780 17644 8832
rect 18880 8780 18932 8832
rect 21272 8780 21324 8832
rect 6148 8678 6200 8730
rect 6212 8678 6264 8730
rect 6276 8678 6328 8730
rect 6340 8678 6392 8730
rect 6404 8678 6456 8730
rect 11346 8678 11398 8730
rect 11410 8678 11462 8730
rect 11474 8678 11526 8730
rect 11538 8678 11590 8730
rect 11602 8678 11654 8730
rect 16544 8678 16596 8730
rect 16608 8678 16660 8730
rect 16672 8678 16724 8730
rect 16736 8678 16788 8730
rect 16800 8678 16852 8730
rect 21742 8678 21794 8730
rect 21806 8678 21858 8730
rect 21870 8678 21922 8730
rect 21934 8678 21986 8730
rect 21998 8678 22050 8730
rect 1492 8576 1544 8628
rect 2136 8508 2188 8560
rect 1400 8304 1452 8356
rect 2780 8440 2832 8492
rect 5172 8508 5224 8560
rect 6552 8576 6604 8628
rect 6828 8576 6880 8628
rect 7932 8576 7984 8628
rect 8668 8576 8720 8628
rect 9956 8619 10008 8628
rect 9956 8585 9965 8619
rect 9965 8585 9999 8619
rect 9999 8585 10008 8619
rect 9956 8576 10008 8585
rect 10508 8619 10560 8628
rect 10508 8585 10517 8619
rect 10517 8585 10551 8619
rect 10551 8585 10560 8619
rect 10508 8576 10560 8585
rect 10600 8576 10652 8628
rect 13820 8619 13872 8628
rect 13820 8585 13829 8619
rect 13829 8585 13863 8619
rect 13863 8585 13872 8619
rect 13820 8576 13872 8585
rect 14556 8576 14608 8628
rect 15108 8576 15160 8628
rect 15752 8619 15804 8628
rect 15752 8585 15761 8619
rect 15761 8585 15795 8619
rect 15795 8585 15804 8619
rect 15752 8576 15804 8585
rect 18880 8576 18932 8628
rect 1676 8347 1728 8356
rect 1676 8313 1685 8347
rect 1685 8313 1719 8347
rect 1719 8313 1728 8347
rect 1676 8304 1728 8313
rect 2780 8304 2832 8356
rect 3332 8440 3384 8492
rect 3976 8483 4028 8492
rect 3424 8372 3476 8424
rect 3700 8415 3752 8424
rect 3700 8381 3709 8415
rect 3709 8381 3743 8415
rect 3743 8381 3752 8415
rect 3700 8372 3752 8381
rect 3976 8449 3985 8483
rect 3985 8449 4019 8483
rect 4019 8449 4028 8483
rect 3976 8440 4028 8449
rect 6000 8440 6052 8492
rect 6920 8440 6972 8492
rect 7288 8483 7340 8492
rect 7288 8449 7297 8483
rect 7297 8449 7331 8483
rect 7331 8449 7340 8483
rect 7288 8440 7340 8449
rect 7656 8508 7708 8560
rect 7840 8508 7892 8560
rect 15384 8483 15436 8492
rect 15384 8449 15402 8483
rect 15402 8449 15436 8483
rect 15384 8440 15436 8449
rect 18972 8508 19024 8560
rect 20628 8576 20680 8628
rect 17316 8440 17368 8492
rect 4620 8372 4672 8424
rect 5080 8372 5132 8424
rect 5448 8372 5500 8424
rect 5724 8415 5776 8424
rect 5724 8381 5733 8415
rect 5733 8381 5767 8415
rect 5767 8381 5776 8415
rect 5724 8372 5776 8381
rect 7380 8415 7432 8424
rect 7380 8381 7389 8415
rect 7389 8381 7423 8415
rect 7423 8381 7432 8415
rect 7380 8372 7432 8381
rect 7564 8415 7616 8424
rect 7564 8381 7573 8415
rect 7573 8381 7607 8415
rect 7607 8381 7616 8415
rect 7564 8372 7616 8381
rect 5080 8236 5132 8288
rect 5816 8236 5868 8288
rect 6828 8279 6880 8288
rect 6828 8245 6837 8279
rect 6837 8245 6871 8279
rect 6871 8245 6880 8279
rect 6828 8236 6880 8245
rect 7748 8236 7800 8288
rect 8208 8304 8260 8356
rect 8668 8372 8720 8424
rect 9128 8372 9180 8424
rect 9772 8372 9824 8424
rect 9864 8415 9916 8424
rect 9864 8381 9873 8415
rect 9873 8381 9907 8415
rect 9907 8381 9916 8415
rect 11060 8415 11112 8424
rect 9864 8372 9916 8381
rect 11060 8381 11069 8415
rect 11069 8381 11103 8415
rect 11103 8381 11112 8415
rect 11060 8372 11112 8381
rect 8576 8279 8628 8288
rect 8576 8245 8585 8279
rect 8585 8245 8619 8279
rect 8619 8245 8628 8279
rect 8576 8236 8628 8245
rect 9864 8236 9916 8288
rect 10324 8236 10376 8288
rect 14464 8372 14516 8424
rect 13268 8304 13320 8356
rect 18144 8304 18196 8356
rect 12532 8236 12584 8288
rect 12808 8236 12860 8288
rect 13452 8236 13504 8288
rect 13728 8236 13780 8288
rect 16488 8236 16540 8288
rect 17408 8236 17460 8288
rect 21272 8236 21324 8288
rect 3549 8134 3601 8186
rect 3613 8134 3665 8186
rect 3677 8134 3729 8186
rect 3741 8134 3793 8186
rect 3805 8134 3857 8186
rect 8747 8134 8799 8186
rect 8811 8134 8863 8186
rect 8875 8134 8927 8186
rect 8939 8134 8991 8186
rect 9003 8134 9055 8186
rect 13945 8134 13997 8186
rect 14009 8134 14061 8186
rect 14073 8134 14125 8186
rect 14137 8134 14189 8186
rect 14201 8134 14253 8186
rect 19143 8134 19195 8186
rect 19207 8134 19259 8186
rect 19271 8134 19323 8186
rect 19335 8134 19387 8186
rect 19399 8134 19451 8186
rect 1492 8075 1544 8084
rect 1492 8041 1501 8075
rect 1501 8041 1535 8075
rect 1535 8041 1544 8075
rect 1492 8032 1544 8041
rect 2780 8032 2832 8084
rect 3884 8032 3936 8084
rect 4988 8032 5040 8084
rect 5632 8032 5684 8084
rect 5724 8032 5776 8084
rect 7472 8032 7524 8084
rect 8208 8032 8260 8084
rect 12624 8032 12676 8084
rect 13728 8032 13780 8084
rect 15108 8032 15160 8084
rect 15476 8032 15528 8084
rect 16396 8032 16448 8084
rect 16488 8032 16540 8084
rect 3056 7964 3108 8016
rect 2044 7939 2096 7948
rect 2044 7905 2053 7939
rect 2053 7905 2087 7939
rect 2087 7905 2096 7939
rect 2872 7939 2924 7948
rect 2044 7896 2096 7905
rect 2872 7905 2881 7939
rect 2881 7905 2915 7939
rect 2915 7905 2924 7939
rect 2872 7896 2924 7905
rect 5080 7896 5132 7948
rect 3056 7871 3108 7880
rect 3056 7837 3065 7871
rect 3065 7837 3099 7871
rect 3099 7837 3108 7871
rect 3056 7828 3108 7837
rect 3976 7828 4028 7880
rect 14556 7964 14608 8016
rect 7104 7939 7156 7948
rect 7104 7905 7113 7939
rect 7113 7905 7147 7939
rect 7147 7905 7156 7939
rect 7104 7896 7156 7905
rect 8116 7896 8168 7948
rect 10876 7896 10928 7948
rect 11336 7896 11388 7948
rect 12532 7939 12584 7948
rect 12532 7905 12541 7939
rect 12541 7905 12575 7939
rect 12575 7905 12584 7939
rect 12532 7896 12584 7905
rect 12992 7896 13044 7948
rect 15200 7896 15252 7948
rect 19524 7964 19576 8016
rect 21548 8032 21600 8084
rect 21272 7939 21324 7948
rect 21272 7905 21281 7939
rect 21281 7905 21315 7939
rect 21315 7905 21324 7939
rect 21272 7896 21324 7905
rect 4620 7760 4672 7812
rect 4712 7760 4764 7812
rect 5264 7760 5316 7812
rect 6368 7871 6420 7880
rect 6368 7837 6377 7871
rect 6377 7837 6411 7871
rect 6411 7837 6420 7871
rect 6368 7828 6420 7837
rect 6920 7871 6972 7880
rect 6920 7837 6929 7871
rect 6929 7837 6963 7871
rect 6963 7837 6972 7871
rect 6920 7828 6972 7837
rect 15108 7828 15160 7880
rect 15752 7828 15804 7880
rect 1768 7692 1820 7744
rect 2504 7735 2556 7744
rect 2504 7701 2513 7735
rect 2513 7701 2547 7735
rect 2547 7701 2556 7735
rect 2504 7692 2556 7701
rect 4988 7735 5040 7744
rect 4988 7701 4997 7735
rect 4997 7701 5031 7735
rect 5031 7701 5040 7735
rect 4988 7692 5040 7701
rect 5080 7692 5132 7744
rect 7840 7760 7892 7812
rect 9312 7760 9364 7812
rect 10416 7803 10468 7812
rect 10416 7769 10425 7803
rect 10425 7769 10459 7803
rect 10459 7769 10468 7803
rect 10416 7760 10468 7769
rect 10508 7760 10560 7812
rect 10968 7803 11020 7812
rect 6828 7735 6880 7744
rect 6828 7701 6837 7735
rect 6837 7701 6871 7735
rect 6871 7701 6880 7735
rect 6828 7692 6880 7701
rect 7104 7692 7156 7744
rect 7564 7735 7616 7744
rect 7564 7701 7573 7735
rect 7573 7701 7607 7735
rect 7607 7701 7616 7735
rect 7564 7692 7616 7701
rect 8392 7692 8444 7744
rect 8576 7692 8628 7744
rect 9404 7692 9456 7744
rect 9588 7692 9640 7744
rect 10968 7769 10977 7803
rect 10977 7769 11011 7803
rect 11011 7769 11020 7803
rect 10968 7760 11020 7769
rect 14188 7760 14240 7812
rect 14372 7760 14424 7812
rect 12072 7692 12124 7744
rect 12440 7692 12492 7744
rect 14280 7735 14332 7744
rect 14280 7701 14289 7735
rect 14289 7701 14323 7735
rect 14323 7701 14332 7735
rect 14280 7692 14332 7701
rect 15752 7692 15804 7744
rect 16396 7692 16448 7744
rect 17224 7692 17276 7744
rect 17592 7760 17644 7812
rect 17684 7735 17736 7744
rect 17684 7701 17693 7735
rect 17693 7701 17727 7735
rect 17727 7701 17736 7735
rect 17684 7692 17736 7701
rect 6148 7590 6200 7642
rect 6212 7590 6264 7642
rect 6276 7590 6328 7642
rect 6340 7590 6392 7642
rect 6404 7590 6456 7642
rect 11346 7590 11398 7642
rect 11410 7590 11462 7642
rect 11474 7590 11526 7642
rect 11538 7590 11590 7642
rect 11602 7590 11654 7642
rect 16544 7590 16596 7642
rect 16608 7590 16660 7642
rect 16672 7590 16724 7642
rect 16736 7590 16788 7642
rect 16800 7590 16852 7642
rect 21742 7590 21794 7642
rect 21806 7590 21858 7642
rect 21870 7590 21922 7642
rect 21934 7590 21986 7642
rect 21998 7590 22050 7642
rect 2044 7488 2096 7540
rect 4252 7531 4304 7540
rect 4252 7497 4261 7531
rect 4261 7497 4295 7531
rect 4295 7497 4304 7531
rect 4252 7488 4304 7497
rect 4988 7488 5040 7540
rect 6644 7488 6696 7540
rect 7288 7488 7340 7540
rect 9588 7531 9640 7540
rect 1768 7420 1820 7472
rect 3056 7420 3108 7472
rect 9588 7497 9597 7531
rect 9597 7497 9631 7531
rect 9631 7497 9640 7531
rect 9588 7488 9640 7497
rect 12072 7531 12124 7540
rect 12072 7497 12081 7531
rect 12081 7497 12115 7531
rect 12115 7497 12124 7531
rect 12072 7488 12124 7497
rect 10600 7420 10652 7472
rect 14280 7488 14332 7540
rect 15108 7531 15160 7540
rect 15108 7497 15117 7531
rect 15117 7497 15151 7531
rect 15151 7497 15160 7531
rect 15108 7488 15160 7497
rect 15476 7488 15528 7540
rect 13728 7420 13780 7472
rect 17776 7488 17828 7540
rect 17868 7420 17920 7472
rect 4528 7395 4580 7404
rect 4528 7361 4537 7395
rect 4537 7361 4571 7395
rect 4571 7361 4580 7395
rect 4528 7352 4580 7361
rect 5816 7395 5868 7404
rect 5816 7361 5825 7395
rect 5825 7361 5859 7395
rect 5859 7361 5868 7395
rect 5816 7352 5868 7361
rect 7932 7395 7984 7404
rect 7932 7361 7941 7395
rect 7941 7361 7975 7395
rect 7975 7361 7984 7395
rect 7932 7352 7984 7361
rect 8668 7352 8720 7404
rect 15476 7395 15528 7404
rect 5172 7284 5224 7336
rect 5448 7284 5500 7336
rect 5908 7284 5960 7336
rect 6092 7284 6144 7336
rect 7104 7327 7156 7336
rect 3976 7216 4028 7268
rect 5448 7148 5500 7200
rect 6000 7216 6052 7268
rect 7104 7293 7113 7327
rect 7113 7293 7147 7327
rect 7147 7293 7156 7327
rect 7104 7284 7156 7293
rect 8208 7327 8260 7336
rect 8208 7293 8217 7327
rect 8217 7293 8251 7327
rect 8251 7293 8260 7327
rect 8208 7284 8260 7293
rect 9588 7284 9640 7336
rect 7564 7216 7616 7268
rect 10876 7216 10928 7268
rect 7196 7148 7248 7200
rect 9864 7148 9916 7200
rect 10324 7191 10376 7200
rect 10324 7157 10333 7191
rect 10333 7157 10367 7191
rect 10367 7157 10376 7191
rect 10324 7148 10376 7157
rect 11060 7148 11112 7200
rect 12992 7284 13044 7336
rect 12256 7216 12308 7268
rect 12900 7216 12952 7268
rect 13820 7216 13872 7268
rect 15476 7361 15485 7395
rect 15485 7361 15519 7395
rect 15519 7361 15528 7395
rect 15476 7352 15528 7361
rect 15016 7284 15068 7336
rect 20812 7420 20864 7472
rect 21272 7488 21324 7540
rect 14924 7148 14976 7200
rect 3549 7046 3601 7098
rect 3613 7046 3665 7098
rect 3677 7046 3729 7098
rect 3741 7046 3793 7098
rect 3805 7046 3857 7098
rect 8747 7046 8799 7098
rect 8811 7046 8863 7098
rect 8875 7046 8927 7098
rect 8939 7046 8991 7098
rect 9003 7046 9055 7098
rect 13945 7046 13997 7098
rect 14009 7046 14061 7098
rect 14073 7046 14125 7098
rect 14137 7046 14189 7098
rect 14201 7046 14253 7098
rect 19143 7046 19195 7098
rect 19207 7046 19259 7098
rect 19271 7046 19323 7098
rect 19335 7046 19387 7098
rect 19399 7046 19451 7098
rect 5816 6944 5868 6996
rect 5632 6876 5684 6928
rect 6828 6876 6880 6928
rect 3976 6851 4028 6860
rect 3976 6817 3985 6851
rect 3985 6817 4019 6851
rect 4019 6817 4028 6851
rect 3976 6808 4028 6817
rect 4160 6851 4212 6860
rect 4160 6817 4169 6851
rect 4169 6817 4203 6851
rect 4203 6817 4212 6851
rect 4160 6808 4212 6817
rect 7104 6944 7156 6996
rect 8392 6987 8444 6996
rect 8392 6953 8401 6987
rect 8401 6953 8435 6987
rect 8435 6953 8444 6987
rect 8392 6944 8444 6953
rect 9312 6987 9364 6996
rect 9312 6953 9321 6987
rect 9321 6953 9355 6987
rect 9355 6953 9364 6987
rect 9312 6944 9364 6953
rect 10508 6944 10560 6996
rect 11704 6944 11756 6996
rect 13820 6944 13872 6996
rect 12256 6876 12308 6928
rect 12992 6876 13044 6928
rect 7748 6851 7800 6860
rect 7748 6817 7757 6851
rect 7757 6817 7791 6851
rect 7791 6817 7800 6851
rect 7748 6808 7800 6817
rect 8576 6851 8628 6860
rect 8576 6817 8585 6851
rect 8585 6817 8619 6851
rect 8619 6817 8628 6851
rect 8576 6808 8628 6817
rect 9036 6808 9088 6860
rect 9772 6808 9824 6860
rect 10692 6808 10744 6860
rect 14556 6851 14608 6860
rect 14556 6817 14565 6851
rect 14565 6817 14599 6851
rect 14599 6817 14608 6851
rect 14556 6808 14608 6817
rect 15016 6876 15068 6928
rect 14740 6808 14792 6860
rect 15476 6808 15528 6860
rect 3424 6783 3476 6792
rect 3424 6749 3433 6783
rect 3433 6749 3467 6783
rect 3467 6749 3476 6783
rect 3424 6740 3476 6749
rect 4436 6740 4488 6792
rect 5724 6740 5776 6792
rect 10324 6740 10376 6792
rect 9956 6672 10008 6724
rect 4988 6604 5040 6656
rect 5172 6604 5224 6656
rect 5724 6647 5776 6656
rect 5724 6613 5733 6647
rect 5733 6613 5767 6647
rect 5767 6613 5776 6647
rect 5724 6604 5776 6613
rect 5816 6604 5868 6656
rect 6000 6604 6052 6656
rect 6368 6647 6420 6656
rect 6368 6613 6377 6647
rect 6377 6613 6411 6647
rect 6411 6613 6420 6647
rect 6368 6604 6420 6613
rect 6828 6604 6880 6656
rect 7196 6604 7248 6656
rect 7656 6604 7708 6656
rect 8116 6604 8168 6656
rect 9128 6647 9180 6656
rect 9128 6613 9137 6647
rect 9137 6613 9171 6647
rect 9171 6613 9180 6647
rect 9128 6604 9180 6613
rect 9864 6604 9916 6656
rect 10692 6672 10744 6724
rect 10416 6647 10468 6656
rect 10416 6613 10425 6647
rect 10425 6613 10459 6647
rect 10459 6613 10468 6647
rect 10416 6604 10468 6613
rect 11796 6672 11848 6724
rect 14372 6740 14424 6792
rect 14648 6672 14700 6724
rect 10968 6604 11020 6656
rect 12440 6604 12492 6656
rect 13820 6647 13872 6656
rect 13820 6613 13829 6647
rect 13829 6613 13863 6647
rect 13863 6613 13872 6647
rect 13820 6604 13872 6613
rect 6148 6502 6200 6554
rect 6212 6502 6264 6554
rect 6276 6502 6328 6554
rect 6340 6502 6392 6554
rect 6404 6502 6456 6554
rect 11346 6502 11398 6554
rect 11410 6502 11462 6554
rect 11474 6502 11526 6554
rect 11538 6502 11590 6554
rect 11602 6502 11654 6554
rect 16544 6502 16596 6554
rect 16608 6502 16660 6554
rect 16672 6502 16724 6554
rect 16736 6502 16788 6554
rect 16800 6502 16852 6554
rect 21742 6502 21794 6554
rect 21806 6502 21858 6554
rect 21870 6502 21922 6554
rect 21934 6502 21986 6554
rect 21998 6502 22050 6554
rect 4344 6375 4396 6384
rect 4344 6341 4353 6375
rect 4353 6341 4387 6375
rect 4387 6341 4396 6375
rect 4344 6332 4396 6341
rect 7380 6400 7432 6452
rect 8116 6400 8168 6452
rect 8668 6400 8720 6452
rect 9036 6400 9088 6452
rect 9956 6443 10008 6452
rect 9956 6409 9965 6443
rect 9965 6409 9999 6443
rect 9999 6409 10008 6443
rect 9956 6400 10008 6409
rect 10416 6400 10468 6452
rect 12624 6400 12676 6452
rect 13268 6400 13320 6452
rect 14464 6400 14516 6452
rect 10600 6332 10652 6384
rect 1492 6264 1544 6316
rect 4252 6264 4304 6316
rect 5632 6264 5684 6316
rect 6000 6264 6052 6316
rect 6920 6264 6972 6316
rect 7104 6264 7156 6316
rect 1860 6239 1912 6248
rect 1860 6205 1869 6239
rect 1869 6205 1903 6239
rect 1903 6205 1912 6239
rect 1860 6196 1912 6205
rect 1400 6060 1452 6112
rect 3976 6196 4028 6248
rect 4988 6196 5040 6248
rect 7380 6264 7432 6316
rect 8024 6264 8076 6316
rect 8392 6264 8444 6316
rect 11336 6332 11388 6384
rect 14740 6332 14792 6384
rect 7564 6239 7616 6248
rect 7564 6205 7573 6239
rect 7573 6205 7607 6239
rect 7607 6205 7616 6239
rect 7564 6196 7616 6205
rect 8208 6196 8260 6248
rect 8484 6196 8536 6248
rect 9588 6196 9640 6248
rect 9864 6239 9916 6248
rect 9864 6205 9873 6239
rect 9873 6205 9907 6239
rect 9907 6205 9916 6239
rect 9864 6196 9916 6205
rect 10692 6239 10744 6248
rect 10692 6205 10701 6239
rect 10701 6205 10735 6239
rect 10735 6205 10744 6239
rect 10692 6196 10744 6205
rect 10876 6239 10928 6248
rect 10876 6205 10885 6239
rect 10885 6205 10919 6239
rect 10919 6205 10928 6239
rect 10876 6196 10928 6205
rect 11520 6239 11572 6248
rect 11520 6205 11529 6239
rect 11529 6205 11563 6239
rect 11563 6205 11572 6239
rect 11520 6196 11572 6205
rect 11796 6196 11848 6248
rect 12440 6196 12492 6248
rect 12532 6196 12584 6248
rect 15568 6264 15620 6316
rect 19708 6196 19760 6248
rect 12164 6128 12216 6180
rect 16304 6128 16356 6180
rect 6276 6060 6328 6112
rect 7288 6060 7340 6112
rect 12532 6060 12584 6112
rect 15844 6060 15896 6112
rect 3549 5958 3601 6010
rect 3613 5958 3665 6010
rect 3677 5958 3729 6010
rect 3741 5958 3793 6010
rect 3805 5958 3857 6010
rect 8747 5958 8799 6010
rect 8811 5958 8863 6010
rect 8875 5958 8927 6010
rect 8939 5958 8991 6010
rect 9003 5958 9055 6010
rect 13945 5958 13997 6010
rect 14009 5958 14061 6010
rect 14073 5958 14125 6010
rect 14137 5958 14189 6010
rect 14201 5958 14253 6010
rect 19143 5958 19195 6010
rect 19207 5958 19259 6010
rect 19271 5958 19323 6010
rect 19335 5958 19387 6010
rect 19399 5958 19451 6010
rect 1492 5899 1544 5908
rect 1492 5865 1501 5899
rect 1501 5865 1535 5899
rect 1535 5865 1544 5899
rect 1492 5856 1544 5865
rect 5540 5856 5592 5908
rect 5816 5856 5868 5908
rect 5264 5720 5316 5772
rect 5448 5652 5500 5704
rect 7012 5856 7064 5908
rect 7564 5856 7616 5908
rect 7748 5899 7800 5908
rect 7748 5865 7757 5899
rect 7757 5865 7791 5899
rect 7791 5865 7800 5899
rect 7748 5856 7800 5865
rect 8116 5856 8168 5908
rect 10876 5856 10928 5908
rect 13268 5899 13320 5908
rect 7472 5788 7524 5840
rect 8024 5788 8076 5840
rect 8392 5788 8444 5840
rect 9036 5788 9088 5840
rect 9864 5788 9916 5840
rect 6552 5763 6604 5772
rect 6552 5729 6561 5763
rect 6561 5729 6595 5763
rect 6595 5729 6604 5763
rect 6552 5720 6604 5729
rect 7380 5720 7432 5772
rect 8576 5720 8628 5772
rect 9496 5720 9548 5772
rect 10784 5652 10836 5704
rect 4528 5584 4580 5636
rect 6276 5584 6328 5636
rect 8944 5584 8996 5636
rect 4988 5559 5040 5568
rect 4988 5525 4997 5559
rect 4997 5525 5031 5559
rect 5031 5525 5040 5559
rect 4988 5516 5040 5525
rect 5172 5559 5224 5568
rect 5172 5525 5181 5559
rect 5181 5525 5215 5559
rect 5215 5525 5224 5559
rect 5172 5516 5224 5525
rect 5448 5559 5500 5568
rect 5448 5525 5457 5559
rect 5457 5525 5491 5559
rect 5491 5525 5500 5559
rect 5448 5516 5500 5525
rect 5816 5516 5868 5568
rect 6644 5516 6696 5568
rect 6920 5516 6972 5568
rect 7380 5516 7432 5568
rect 8852 5516 8904 5568
rect 9312 5584 9364 5636
rect 10140 5584 10192 5636
rect 10600 5584 10652 5636
rect 12532 5720 12584 5772
rect 12808 5720 12860 5772
rect 13268 5865 13277 5899
rect 13277 5865 13311 5899
rect 13311 5865 13320 5899
rect 13268 5856 13320 5865
rect 19616 5856 19668 5908
rect 19064 5788 19116 5840
rect 11796 5695 11848 5704
rect 11796 5661 11805 5695
rect 11805 5661 11839 5695
rect 11839 5661 11848 5695
rect 11796 5652 11848 5661
rect 12440 5652 12492 5704
rect 17500 5720 17552 5772
rect 20628 5788 20680 5840
rect 21180 5720 21232 5772
rect 10692 5559 10744 5568
rect 10692 5525 10701 5559
rect 10701 5525 10735 5559
rect 10735 5525 10744 5559
rect 10692 5516 10744 5525
rect 10784 5559 10836 5568
rect 10784 5525 10793 5559
rect 10793 5525 10827 5559
rect 10827 5525 10836 5559
rect 11704 5559 11756 5568
rect 10784 5516 10836 5525
rect 11704 5525 11713 5559
rect 11713 5525 11747 5559
rect 11747 5525 11756 5559
rect 11704 5516 11756 5525
rect 12440 5516 12492 5568
rect 12808 5559 12860 5568
rect 12808 5525 12817 5559
rect 12817 5525 12851 5559
rect 12851 5525 12860 5559
rect 12808 5516 12860 5525
rect 12900 5559 12952 5568
rect 12900 5525 12909 5559
rect 12909 5525 12943 5559
rect 12943 5525 12952 5559
rect 14280 5584 14332 5636
rect 14372 5584 14424 5636
rect 12900 5516 12952 5525
rect 15660 5516 15712 5568
rect 16396 5516 16448 5568
rect 17776 5559 17828 5568
rect 17776 5525 17785 5559
rect 17785 5525 17819 5559
rect 17819 5525 17828 5559
rect 17776 5516 17828 5525
rect 20260 5559 20312 5568
rect 20260 5525 20269 5559
rect 20269 5525 20303 5559
rect 20303 5525 20312 5559
rect 20260 5516 20312 5525
rect 20628 5516 20680 5568
rect 6148 5414 6200 5466
rect 6212 5414 6264 5466
rect 6276 5414 6328 5466
rect 6340 5414 6392 5466
rect 6404 5414 6456 5466
rect 11346 5414 11398 5466
rect 11410 5414 11462 5466
rect 11474 5414 11526 5466
rect 11538 5414 11590 5466
rect 11602 5414 11654 5466
rect 16544 5414 16596 5466
rect 16608 5414 16660 5466
rect 16672 5414 16724 5466
rect 16736 5414 16788 5466
rect 16800 5414 16852 5466
rect 21742 5414 21794 5466
rect 21806 5414 21858 5466
rect 21870 5414 21922 5466
rect 21934 5414 21986 5466
rect 21998 5414 22050 5466
rect 2964 5312 3016 5364
rect 3792 5312 3844 5364
rect 4712 5355 4764 5364
rect 4712 5321 4721 5355
rect 4721 5321 4755 5355
rect 4755 5321 4764 5355
rect 4712 5312 4764 5321
rect 5080 5355 5132 5364
rect 5080 5321 5089 5355
rect 5089 5321 5123 5355
rect 5123 5321 5132 5355
rect 5080 5312 5132 5321
rect 6644 5355 6696 5364
rect 6644 5321 6653 5355
rect 6653 5321 6687 5355
rect 6687 5321 6696 5355
rect 6644 5312 6696 5321
rect 7932 5355 7984 5364
rect 4068 5176 4120 5228
rect 5172 5176 5224 5228
rect 5816 5176 5868 5228
rect 7932 5321 7941 5355
rect 7941 5321 7975 5355
rect 7975 5321 7984 5355
rect 7932 5312 7984 5321
rect 7748 5244 7800 5296
rect 8944 5312 8996 5364
rect 9404 5312 9456 5364
rect 10692 5312 10744 5364
rect 12808 5312 12860 5364
rect 13452 5312 13504 5364
rect 17776 5312 17828 5364
rect 12532 5244 12584 5296
rect 9956 5176 10008 5228
rect 12072 5176 12124 5228
rect 12256 5176 12308 5228
rect 2044 5151 2096 5160
rect 2044 5117 2053 5151
rect 2053 5117 2087 5151
rect 2087 5117 2096 5151
rect 2044 5108 2096 5117
rect 3792 5151 3844 5160
rect 3792 5117 3801 5151
rect 3801 5117 3835 5151
rect 3835 5117 3844 5151
rect 3792 5108 3844 5117
rect 4712 5108 4764 5160
rect 6000 5151 6052 5160
rect 4252 5040 4304 5092
rect 5172 5040 5224 5092
rect 4068 5015 4120 5024
rect 4068 4981 4077 5015
rect 4077 4981 4111 5015
rect 4111 4981 4120 5015
rect 4068 4972 4120 4981
rect 4160 5015 4212 5024
rect 4160 4981 4169 5015
rect 4169 4981 4203 5015
rect 4203 4981 4212 5015
rect 6000 5117 6009 5151
rect 6009 5117 6043 5151
rect 6043 5117 6052 5151
rect 6000 5108 6052 5117
rect 7564 5108 7616 5160
rect 8484 5151 8536 5160
rect 8484 5117 8493 5151
rect 8493 5117 8527 5151
rect 8527 5117 8536 5151
rect 8484 5108 8536 5117
rect 9312 5108 9364 5160
rect 10324 5151 10376 5160
rect 7380 5040 7432 5092
rect 7748 5083 7800 5092
rect 7748 5049 7757 5083
rect 7757 5049 7791 5083
rect 7791 5049 7800 5083
rect 7748 5040 7800 5049
rect 8300 5040 8352 5092
rect 8852 5040 8904 5092
rect 10324 5117 10333 5151
rect 10333 5117 10367 5151
rect 10367 5117 10376 5151
rect 10324 5108 10376 5117
rect 10508 5151 10560 5160
rect 10508 5117 10517 5151
rect 10517 5117 10551 5151
rect 10551 5117 10560 5151
rect 10508 5108 10560 5117
rect 11796 5151 11848 5160
rect 11796 5117 11805 5151
rect 11805 5117 11839 5151
rect 11839 5117 11848 5151
rect 11796 5108 11848 5117
rect 12532 5151 12584 5160
rect 12532 5117 12541 5151
rect 12541 5117 12575 5151
rect 12575 5117 12584 5151
rect 12532 5108 12584 5117
rect 12624 5108 12676 5160
rect 4160 4972 4212 4981
rect 5632 4972 5684 5024
rect 8484 4972 8536 5024
rect 12164 5040 12216 5092
rect 15200 5176 15252 5228
rect 13452 5151 13504 5160
rect 13452 5117 13461 5151
rect 13461 5117 13495 5151
rect 13495 5117 13504 5151
rect 13452 5108 13504 5117
rect 15476 5151 15528 5160
rect 15476 5117 15485 5151
rect 15485 5117 15519 5151
rect 15519 5117 15528 5151
rect 15476 5108 15528 5117
rect 17040 5244 17092 5296
rect 15844 5219 15896 5228
rect 15844 5185 15853 5219
rect 15853 5185 15887 5219
rect 15887 5185 15896 5219
rect 15844 5176 15896 5185
rect 20628 5219 20680 5228
rect 20628 5185 20637 5219
rect 20637 5185 20671 5219
rect 20671 5185 20680 5219
rect 20628 5176 20680 5185
rect 17040 5108 17092 5160
rect 20904 5151 20956 5160
rect 20904 5117 20913 5151
rect 20913 5117 20947 5151
rect 20947 5117 20956 5151
rect 20904 5108 20956 5117
rect 9312 5015 9364 5024
rect 9312 4981 9321 5015
rect 9321 4981 9355 5015
rect 9355 4981 9364 5015
rect 9312 4972 9364 4981
rect 12532 4972 12584 5024
rect 13360 4972 13412 5024
rect 14832 4972 14884 5024
rect 3549 4870 3601 4922
rect 3613 4870 3665 4922
rect 3677 4870 3729 4922
rect 3741 4870 3793 4922
rect 3805 4870 3857 4922
rect 8747 4870 8799 4922
rect 8811 4870 8863 4922
rect 8875 4870 8927 4922
rect 8939 4870 8991 4922
rect 9003 4870 9055 4922
rect 13945 4870 13997 4922
rect 14009 4870 14061 4922
rect 14073 4870 14125 4922
rect 14137 4870 14189 4922
rect 14201 4870 14253 4922
rect 19143 4870 19195 4922
rect 19207 4870 19259 4922
rect 19271 4870 19323 4922
rect 19335 4870 19387 4922
rect 19399 4870 19451 4922
rect 4896 4768 4948 4820
rect 5816 4811 5868 4820
rect 5816 4777 5825 4811
rect 5825 4777 5859 4811
rect 5859 4777 5868 4811
rect 5816 4768 5868 4777
rect 5908 4768 5960 4820
rect 7104 4811 7156 4820
rect 7104 4777 7113 4811
rect 7113 4777 7147 4811
rect 7147 4777 7156 4811
rect 7104 4768 7156 4777
rect 7932 4768 7984 4820
rect 8760 4768 8812 4820
rect 9036 4768 9088 4820
rect 10416 4768 10468 4820
rect 12256 4811 12308 4820
rect 12256 4777 12265 4811
rect 12265 4777 12299 4811
rect 12299 4777 12308 4811
rect 15476 4811 15528 4820
rect 12256 4768 12308 4777
rect 15476 4777 15485 4811
rect 15485 4777 15519 4811
rect 15519 4777 15528 4811
rect 15476 4768 15528 4777
rect 16948 4811 17000 4820
rect 16948 4777 16957 4811
rect 16957 4777 16991 4811
rect 16991 4777 17000 4811
rect 16948 4768 17000 4777
rect 20260 4768 20312 4820
rect 3424 4700 3476 4752
rect 5264 4675 5316 4684
rect 5264 4641 5273 4675
rect 5273 4641 5307 4675
rect 5307 4641 5316 4675
rect 5264 4632 5316 4641
rect 6552 4632 6604 4684
rect 6736 4675 6788 4684
rect 6736 4641 6745 4675
rect 6745 4641 6779 4675
rect 6779 4641 6788 4675
rect 6736 4632 6788 4641
rect 7104 4632 7156 4684
rect 7932 4675 7984 4684
rect 7932 4641 7941 4675
rect 7941 4641 7975 4675
rect 7975 4641 7984 4675
rect 7932 4632 7984 4641
rect 10140 4632 10192 4684
rect 11888 4700 11940 4752
rect 13084 4700 13136 4752
rect 4896 4564 4948 4616
rect 6000 4564 6052 4616
rect 7656 4564 7708 4616
rect 9312 4564 9364 4616
rect 4068 4496 4120 4548
rect 5632 4496 5684 4548
rect 8300 4496 8352 4548
rect 9036 4496 9088 4548
rect 10324 4564 10376 4616
rect 12900 4632 12952 4684
rect 14832 4675 14884 4684
rect 14832 4641 14841 4675
rect 14841 4641 14875 4675
rect 14875 4641 14884 4675
rect 14832 4632 14884 4641
rect 17592 4700 17644 4752
rect 16028 4675 16080 4684
rect 16028 4641 16037 4675
rect 16037 4641 16071 4675
rect 16071 4641 16080 4675
rect 16028 4632 16080 4641
rect 17500 4675 17552 4684
rect 6000 4428 6052 4480
rect 6736 4428 6788 4480
rect 9496 4428 9548 4480
rect 12624 4564 12676 4616
rect 13636 4564 13688 4616
rect 14740 4607 14792 4616
rect 14740 4573 14749 4607
rect 14749 4573 14783 4607
rect 14783 4573 14792 4607
rect 14740 4564 14792 4573
rect 15844 4607 15896 4616
rect 15844 4573 15853 4607
rect 15853 4573 15887 4607
rect 15887 4573 15896 4607
rect 15844 4564 15896 4573
rect 16948 4564 17000 4616
rect 17500 4641 17509 4675
rect 17509 4641 17543 4675
rect 17543 4641 17552 4675
rect 17500 4632 17552 4641
rect 22468 4632 22520 4684
rect 19064 4564 19116 4616
rect 12256 4496 12308 4548
rect 17776 4496 17828 4548
rect 19892 4496 19944 4548
rect 13176 4428 13228 4480
rect 14372 4471 14424 4480
rect 14372 4437 14381 4471
rect 14381 4437 14415 4471
rect 14415 4437 14424 4471
rect 14372 4428 14424 4437
rect 15936 4471 15988 4480
rect 15936 4437 15945 4471
rect 15945 4437 15979 4471
rect 15979 4437 15988 4471
rect 15936 4428 15988 4437
rect 16396 4428 16448 4480
rect 17224 4471 17276 4480
rect 17224 4437 17233 4471
rect 17233 4437 17267 4471
rect 17267 4437 17276 4471
rect 17224 4428 17276 4437
rect 17408 4428 17460 4480
rect 17592 4471 17644 4480
rect 17592 4437 17601 4471
rect 17601 4437 17635 4471
rect 17635 4437 17644 4471
rect 17592 4428 17644 4437
rect 17684 4471 17736 4480
rect 17684 4437 17693 4471
rect 17693 4437 17727 4471
rect 17727 4437 17736 4471
rect 17684 4428 17736 4437
rect 6148 4326 6200 4378
rect 6212 4326 6264 4378
rect 6276 4326 6328 4378
rect 6340 4326 6392 4378
rect 6404 4326 6456 4378
rect 11346 4326 11398 4378
rect 11410 4326 11462 4378
rect 11474 4326 11526 4378
rect 11538 4326 11590 4378
rect 11602 4326 11654 4378
rect 16544 4326 16596 4378
rect 16608 4326 16660 4378
rect 16672 4326 16724 4378
rect 16736 4326 16788 4378
rect 16800 4326 16852 4378
rect 21742 4326 21794 4378
rect 21806 4326 21858 4378
rect 21870 4326 21922 4378
rect 21934 4326 21986 4378
rect 21998 4326 22050 4378
rect 5264 4224 5316 4276
rect 7840 4224 7892 4276
rect 9128 4224 9180 4276
rect 9496 4267 9548 4276
rect 9496 4233 9505 4267
rect 9505 4233 9539 4267
rect 9539 4233 9548 4267
rect 9496 4224 9548 4233
rect 10508 4267 10560 4276
rect 10508 4233 10517 4267
rect 10517 4233 10551 4267
rect 10551 4233 10560 4267
rect 10508 4224 10560 4233
rect 10876 4267 10928 4276
rect 10876 4233 10885 4267
rect 10885 4233 10919 4267
rect 10919 4233 10928 4267
rect 10876 4224 10928 4233
rect 11888 4267 11940 4276
rect 11888 4233 11897 4267
rect 11897 4233 11931 4267
rect 11931 4233 11940 4267
rect 11888 4224 11940 4233
rect 12072 4224 12124 4276
rect 13268 4224 13320 4276
rect 17592 4267 17644 4276
rect 17592 4233 17601 4267
rect 17601 4233 17635 4267
rect 17635 4233 17644 4267
rect 17592 4224 17644 4233
rect 6552 4156 6604 4208
rect 7932 4156 7984 4208
rect 8208 4156 8260 4208
rect 10416 4156 10468 4208
rect 15752 4156 15804 4208
rect 17408 4156 17460 4208
rect 19064 4156 19116 4208
rect 3976 4088 4028 4140
rect 6000 4088 6052 4140
rect 2228 4020 2280 4072
rect 4160 4020 4212 4072
rect 5540 4063 5592 4072
rect 5540 4029 5549 4063
rect 5549 4029 5583 4063
rect 5583 4029 5592 4063
rect 5540 4020 5592 4029
rect 5724 4063 5776 4072
rect 5724 4029 5733 4063
rect 5733 4029 5767 4063
rect 5767 4029 5776 4063
rect 5724 4020 5776 4029
rect 7564 4063 7616 4072
rect 7564 4029 7573 4063
rect 7573 4029 7607 4063
rect 7607 4029 7616 4063
rect 7564 4020 7616 4029
rect 3332 3952 3384 4004
rect 5816 3952 5868 4004
rect 4620 3884 4672 3936
rect 5448 3884 5500 3936
rect 6184 3927 6236 3936
rect 6184 3893 6193 3927
rect 6193 3893 6227 3927
rect 6227 3893 6236 3927
rect 6184 3884 6236 3893
rect 6460 3884 6512 3936
rect 8576 4131 8628 4140
rect 8576 4097 8585 4131
rect 8585 4097 8619 4131
rect 8619 4097 8628 4131
rect 8576 4088 8628 4097
rect 7840 4020 7892 4072
rect 8116 3995 8168 4004
rect 8116 3961 8125 3995
rect 8125 3961 8159 3995
rect 8159 3961 8168 3995
rect 8116 3952 8168 3961
rect 9680 4088 9732 4140
rect 9496 4020 9548 4072
rect 10324 4063 10376 4072
rect 9220 3952 9272 4004
rect 10324 4029 10333 4063
rect 10333 4029 10367 4063
rect 10367 4029 10376 4063
rect 10324 4020 10376 4029
rect 10508 3952 10560 4004
rect 11060 4063 11112 4072
rect 11060 4029 11069 4063
rect 11069 4029 11103 4063
rect 11103 4029 11112 4063
rect 11060 4020 11112 4029
rect 11428 4020 11480 4072
rect 12072 4063 12124 4072
rect 12072 4029 12081 4063
rect 12081 4029 12115 4063
rect 12115 4029 12124 4063
rect 12072 4020 12124 4029
rect 12808 4088 12860 4140
rect 13820 4088 13872 4140
rect 14372 4131 14424 4140
rect 14372 4097 14381 4131
rect 14381 4097 14415 4131
rect 14415 4097 14424 4131
rect 14372 4088 14424 4097
rect 16948 4088 17000 4140
rect 15384 4020 15436 4072
rect 17868 4088 17920 4140
rect 17132 4020 17184 4072
rect 17316 4063 17368 4072
rect 17316 4029 17325 4063
rect 17325 4029 17359 4063
rect 17359 4029 17368 4063
rect 17316 4020 17368 4029
rect 18144 4063 18196 4072
rect 18144 4029 18153 4063
rect 18153 4029 18187 4063
rect 18187 4029 18196 4063
rect 18144 4020 18196 4029
rect 14556 3952 14608 4004
rect 15936 3952 15988 4004
rect 8024 3884 8076 3936
rect 8392 3884 8444 3936
rect 8576 3884 8628 3936
rect 16028 3884 16080 3936
rect 17224 3884 17276 3936
rect 3549 3782 3601 3834
rect 3613 3782 3665 3834
rect 3677 3782 3729 3834
rect 3741 3782 3793 3834
rect 3805 3782 3857 3834
rect 8747 3782 8799 3834
rect 8811 3782 8863 3834
rect 8875 3782 8927 3834
rect 8939 3782 8991 3834
rect 9003 3782 9055 3834
rect 13945 3782 13997 3834
rect 14009 3782 14061 3834
rect 14073 3782 14125 3834
rect 14137 3782 14189 3834
rect 14201 3782 14253 3834
rect 19143 3782 19195 3834
rect 19207 3782 19259 3834
rect 19271 3782 19323 3834
rect 19335 3782 19387 3834
rect 19399 3782 19451 3834
rect 1768 3680 1820 3732
rect 6552 3680 6604 3732
rect 7748 3680 7800 3732
rect 9772 3680 9824 3732
rect 10876 3723 10928 3732
rect 10876 3689 10885 3723
rect 10885 3689 10919 3723
rect 10919 3689 10928 3723
rect 10876 3680 10928 3689
rect 11060 3680 11112 3732
rect 15844 3680 15896 3732
rect 16212 3680 16264 3732
rect 17408 3723 17460 3732
rect 17408 3689 17417 3723
rect 17417 3689 17451 3723
rect 17451 3689 17460 3723
rect 17408 3680 17460 3689
rect 3148 3612 3200 3664
rect 6460 3612 6512 3664
rect 6736 3612 6788 3664
rect 7840 3612 7892 3664
rect 8024 3655 8076 3664
rect 8024 3621 8033 3655
rect 8033 3621 8067 3655
rect 8067 3621 8076 3655
rect 8024 3612 8076 3621
rect 12072 3612 12124 3664
rect 17132 3612 17184 3664
rect 18604 3655 18656 3664
rect 18604 3621 18613 3655
rect 18613 3621 18647 3655
rect 18647 3621 18656 3655
rect 18604 3612 18656 3621
rect 5448 3587 5500 3596
rect 5448 3553 5457 3587
rect 5457 3553 5491 3587
rect 5491 3553 5500 3587
rect 5448 3544 5500 3553
rect 5632 3544 5684 3596
rect 5908 3587 5960 3596
rect 5908 3553 5917 3587
rect 5917 3553 5951 3587
rect 5951 3553 5960 3587
rect 5908 3544 5960 3553
rect 6368 3587 6420 3596
rect 5816 3476 5868 3528
rect 6368 3553 6377 3587
rect 6377 3553 6411 3587
rect 6411 3553 6420 3587
rect 6368 3544 6420 3553
rect 6552 3587 6604 3596
rect 6552 3553 6561 3587
rect 6561 3553 6595 3587
rect 6595 3553 6604 3587
rect 6552 3544 6604 3553
rect 9956 3544 10008 3596
rect 10324 3587 10376 3596
rect 10324 3553 10333 3587
rect 10333 3553 10367 3587
rect 10367 3553 10376 3587
rect 10324 3544 10376 3553
rect 10416 3587 10468 3596
rect 10416 3553 10425 3587
rect 10425 3553 10459 3587
rect 10459 3553 10468 3587
rect 10416 3544 10468 3553
rect 11060 3544 11112 3596
rect 11244 3544 11296 3596
rect 18512 3544 18564 3596
rect 6184 3476 6236 3528
rect 3884 3340 3936 3392
rect 5448 3408 5500 3460
rect 5080 3340 5132 3392
rect 5908 3340 5960 3392
rect 6736 3340 6788 3392
rect 13544 3476 13596 3528
rect 14924 3476 14976 3528
rect 17868 3476 17920 3528
rect 18420 3476 18472 3528
rect 9772 3408 9824 3460
rect 9956 3383 10008 3392
rect 9956 3349 9965 3383
rect 9965 3349 9999 3383
rect 9999 3349 10008 3383
rect 9956 3340 10008 3349
rect 11060 3340 11112 3392
rect 11428 3340 11480 3392
rect 11704 3383 11756 3392
rect 11704 3349 11713 3383
rect 11713 3349 11747 3383
rect 11747 3349 11756 3383
rect 11704 3340 11756 3349
rect 13636 3408 13688 3460
rect 16304 3408 16356 3460
rect 20168 3408 20220 3460
rect 13728 3383 13780 3392
rect 13728 3349 13737 3383
rect 13737 3349 13771 3383
rect 13771 3349 13780 3383
rect 13728 3340 13780 3349
rect 16212 3340 16264 3392
rect 18236 3340 18288 3392
rect 21548 3340 21600 3392
rect 6148 3238 6200 3290
rect 6212 3238 6264 3290
rect 6276 3238 6328 3290
rect 6340 3238 6392 3290
rect 6404 3238 6456 3290
rect 11346 3238 11398 3290
rect 11410 3238 11462 3290
rect 11474 3238 11526 3290
rect 11538 3238 11590 3290
rect 11602 3238 11654 3290
rect 16544 3238 16596 3290
rect 16608 3238 16660 3290
rect 16672 3238 16724 3290
rect 16736 3238 16788 3290
rect 16800 3238 16852 3290
rect 21742 3238 21794 3290
rect 21806 3238 21858 3290
rect 21870 3238 21922 3290
rect 21934 3238 21986 3290
rect 21998 3238 22050 3290
rect 5080 3179 5132 3188
rect 5080 3145 5089 3179
rect 5089 3145 5123 3179
rect 5123 3145 5132 3179
rect 5080 3136 5132 3145
rect 5448 3179 5500 3188
rect 5448 3145 5457 3179
rect 5457 3145 5491 3179
rect 5491 3145 5500 3179
rect 5448 3136 5500 3145
rect 6736 3179 6788 3188
rect 6736 3145 6745 3179
rect 6745 3145 6779 3179
rect 6779 3145 6788 3179
rect 6736 3136 6788 3145
rect 9772 3136 9824 3188
rect 10416 3136 10468 3188
rect 11704 3136 11756 3188
rect 11980 3136 12032 3188
rect 15568 3136 15620 3188
rect 16304 3179 16356 3188
rect 6920 3068 6972 3120
rect 7656 3111 7708 3120
rect 7656 3077 7665 3111
rect 7665 3077 7699 3111
rect 7699 3077 7708 3111
rect 7656 3068 7708 3077
rect 8576 3111 8628 3120
rect 8576 3077 8585 3111
rect 8585 3077 8619 3111
rect 8619 3077 8628 3111
rect 8576 3068 8628 3077
rect 5448 3000 5500 3052
rect 7104 3000 7156 3052
rect 10140 3111 10192 3120
rect 4988 2975 5040 2984
rect 388 2864 440 2916
rect 3424 2864 3476 2916
rect 4988 2941 4997 2975
rect 4997 2941 5031 2975
rect 5031 2941 5040 2975
rect 4988 2932 5040 2941
rect 5540 2932 5592 2984
rect 6552 2975 6604 2984
rect 6552 2941 6561 2975
rect 6561 2941 6595 2975
rect 6595 2941 6604 2975
rect 6552 2932 6604 2941
rect 7656 2932 7708 2984
rect 9312 3043 9364 3052
rect 9312 3009 9321 3043
rect 9321 3009 9355 3043
rect 9355 3009 9364 3043
rect 9312 3000 9364 3009
rect 7840 2975 7892 2984
rect 7840 2941 7849 2975
rect 7849 2941 7883 2975
rect 7883 2941 7892 2975
rect 7840 2932 7892 2941
rect 9128 2975 9180 2984
rect 9128 2941 9137 2975
rect 9137 2941 9171 2975
rect 9171 2941 9180 2975
rect 10140 3077 10149 3111
rect 10149 3077 10183 3111
rect 10183 3077 10192 3111
rect 10140 3068 10192 3077
rect 11060 3068 11112 3120
rect 9956 3000 10008 3052
rect 10508 3000 10560 3052
rect 11796 3000 11848 3052
rect 11980 3000 12032 3052
rect 16304 3145 16313 3179
rect 16313 3145 16347 3179
rect 16347 3145 16356 3179
rect 16304 3136 16356 3145
rect 17868 3136 17920 3188
rect 18788 3136 18840 3188
rect 19248 3136 19300 3188
rect 19432 3136 19484 3188
rect 9128 2932 9180 2941
rect 9680 2907 9732 2916
rect 9680 2873 9689 2907
rect 9689 2873 9723 2907
rect 9723 2873 9732 2907
rect 9680 2864 9732 2873
rect 10600 2932 10652 2984
rect 13452 3043 13504 3052
rect 10876 2796 10928 2848
rect 13176 2932 13228 2984
rect 13452 3009 13461 3043
rect 13461 3009 13495 3043
rect 13495 3009 13504 3043
rect 13452 3000 13504 3009
rect 13544 3043 13596 3052
rect 13544 3009 13553 3043
rect 13553 3009 13587 3043
rect 13587 3009 13596 3043
rect 13728 3043 13780 3052
rect 13544 3000 13596 3009
rect 13728 3009 13737 3043
rect 13737 3009 13771 3043
rect 13771 3009 13780 3043
rect 13728 3000 13780 3009
rect 14280 3043 14332 3052
rect 14280 3009 14289 3043
rect 14289 3009 14323 3043
rect 14323 3009 14332 3043
rect 14280 3000 14332 3009
rect 14556 3000 14608 3052
rect 14924 3000 14976 3052
rect 15384 3043 15436 3052
rect 15384 3009 15393 3043
rect 15393 3009 15427 3043
rect 15427 3009 15436 3043
rect 15384 3000 15436 3009
rect 15752 3043 15804 3052
rect 15752 3009 15761 3043
rect 15761 3009 15795 3043
rect 15795 3009 15804 3043
rect 15752 3000 15804 3009
rect 13820 2932 13872 2984
rect 15936 2932 15988 2984
rect 16212 3000 16264 3052
rect 17040 3043 17092 3052
rect 17040 3009 17049 3043
rect 17049 3009 17083 3043
rect 17083 3009 17092 3043
rect 17040 3000 17092 3009
rect 17776 3000 17828 3052
rect 18420 3043 18472 3052
rect 18420 3009 18429 3043
rect 18429 3009 18463 3043
rect 18463 3009 18472 3043
rect 18420 3000 18472 3009
rect 18604 3000 18656 3052
rect 19064 3000 19116 3052
rect 22100 3068 22152 3120
rect 19524 3000 19576 3052
rect 19616 3000 19668 3052
rect 19892 3043 19944 3052
rect 19892 3009 19901 3043
rect 19901 3009 19935 3043
rect 19935 3009 19944 3043
rect 19892 3000 19944 3009
rect 19984 3000 20036 3052
rect 20904 3043 20956 3052
rect 20904 3009 20913 3043
rect 20913 3009 20947 3043
rect 20947 3009 20956 3043
rect 20904 3000 20956 3009
rect 15108 2864 15160 2916
rect 13268 2839 13320 2848
rect 13268 2805 13277 2839
rect 13277 2805 13311 2839
rect 13311 2805 13320 2839
rect 13268 2796 13320 2805
rect 13728 2796 13780 2848
rect 14648 2796 14700 2848
rect 16028 2864 16080 2916
rect 17408 2864 17460 2916
rect 18236 2907 18288 2916
rect 18236 2873 18245 2907
rect 18245 2873 18279 2907
rect 18279 2873 18288 2907
rect 18236 2864 18288 2873
rect 21088 2932 21140 2984
rect 19064 2864 19116 2916
rect 16948 2796 17000 2848
rect 19156 2796 19208 2848
rect 20628 2864 20680 2916
rect 3549 2694 3601 2746
rect 3613 2694 3665 2746
rect 3677 2694 3729 2746
rect 3741 2694 3793 2746
rect 3805 2694 3857 2746
rect 8747 2694 8799 2746
rect 8811 2694 8863 2746
rect 8875 2694 8927 2746
rect 8939 2694 8991 2746
rect 9003 2694 9055 2746
rect 13945 2694 13997 2746
rect 14009 2694 14061 2746
rect 14073 2694 14125 2746
rect 14137 2694 14189 2746
rect 14201 2694 14253 2746
rect 19143 2694 19195 2746
rect 19207 2694 19259 2746
rect 19271 2694 19323 2746
rect 19335 2694 19387 2746
rect 19399 2694 19451 2746
rect 4988 2635 5040 2644
rect 4988 2601 4997 2635
rect 4997 2601 5031 2635
rect 5031 2601 5040 2635
rect 4988 2592 5040 2601
rect 5816 2635 5868 2644
rect 5816 2601 5825 2635
rect 5825 2601 5859 2635
rect 5859 2601 5868 2635
rect 5816 2592 5868 2601
rect 8116 2592 8168 2644
rect 10140 2592 10192 2644
rect 10416 2592 10468 2644
rect 10876 2635 10928 2644
rect 10876 2601 10885 2635
rect 10885 2601 10919 2635
rect 10919 2601 10928 2635
rect 10876 2592 10928 2601
rect 11796 2635 11848 2644
rect 11796 2601 11805 2635
rect 11805 2601 11839 2635
rect 11839 2601 11848 2635
rect 11796 2592 11848 2601
rect 14556 2635 14608 2644
rect 14556 2601 14565 2635
rect 14565 2601 14599 2635
rect 14599 2601 14608 2635
rect 14556 2592 14608 2601
rect 14924 2635 14976 2644
rect 14924 2601 14933 2635
rect 14933 2601 14967 2635
rect 14967 2601 14976 2635
rect 14924 2592 14976 2601
rect 15752 2592 15804 2644
rect 15936 2635 15988 2644
rect 15936 2601 15945 2635
rect 15945 2601 15979 2635
rect 15979 2601 15988 2635
rect 15936 2592 15988 2601
rect 17960 2592 18012 2644
rect 3424 2524 3476 2576
rect 8668 2524 8720 2576
rect 5816 2456 5868 2508
rect 10324 2524 10376 2576
rect 848 2388 900 2440
rect 7656 2388 7708 2440
rect 7932 2388 7984 2440
rect 13820 2388 13872 2440
rect 18328 2524 18380 2576
rect 2688 2320 2740 2372
rect 8576 2320 8628 2372
rect 9312 2363 9364 2372
rect 9312 2329 9321 2363
rect 9321 2329 9355 2363
rect 9355 2329 9364 2363
rect 9312 2320 9364 2329
rect 18420 2320 18472 2372
rect 3148 2252 3200 2304
rect 4068 2252 4120 2304
rect 6920 2295 6972 2304
rect 6920 2261 6929 2295
rect 6929 2261 6963 2295
rect 6963 2261 6972 2295
rect 6920 2252 6972 2261
rect 14188 2252 14240 2304
rect 6148 2150 6200 2202
rect 6212 2150 6264 2202
rect 6276 2150 6328 2202
rect 6340 2150 6392 2202
rect 6404 2150 6456 2202
rect 11346 2150 11398 2202
rect 11410 2150 11462 2202
rect 11474 2150 11526 2202
rect 11538 2150 11590 2202
rect 11602 2150 11654 2202
rect 16544 2150 16596 2202
rect 16608 2150 16660 2202
rect 16672 2150 16724 2202
rect 16736 2150 16788 2202
rect 16800 2150 16852 2202
rect 21742 2150 21794 2202
rect 21806 2150 21858 2202
rect 21870 2150 21922 2202
rect 21934 2150 21986 2202
rect 21998 2150 22050 2202
rect 3424 2048 3476 2100
rect 7564 2048 7616 2100
rect 1308 1980 1360 2032
rect 6920 1980 6972 2032
<< metal2 >>
rect 202 22200 258 23000
rect 662 22200 718 23000
rect 1122 22200 1178 23000
rect 1582 22200 1638 23000
rect 2042 22200 2098 23000
rect 2502 22200 2558 23000
rect 2962 22200 3018 23000
rect 3068 22222 3372 22250
rect 216 18630 244 22200
rect 204 18624 256 18630
rect 204 18566 256 18572
rect 676 16726 704 22200
rect 1136 18086 1164 22200
rect 1596 18154 1624 22200
rect 2056 18222 2084 22200
rect 2516 18358 2544 22200
rect 2976 22114 3004 22200
rect 3068 22114 3096 22222
rect 2976 22086 3096 22114
rect 2778 21040 2834 21049
rect 2778 20975 2834 20984
rect 2792 20058 2820 20975
rect 2870 20632 2926 20641
rect 2870 20567 2926 20576
rect 2780 20052 2832 20058
rect 2780 19994 2832 20000
rect 2778 19408 2834 19417
rect 2778 19343 2834 19352
rect 2504 18352 2556 18358
rect 2504 18294 2556 18300
rect 2044 18216 2096 18222
rect 2044 18158 2096 18164
rect 2594 18184 2650 18193
rect 1584 18148 1636 18154
rect 2594 18119 2650 18128
rect 1584 18090 1636 18096
rect 1124 18080 1176 18086
rect 1124 18022 1176 18028
rect 2318 17776 2374 17785
rect 2318 17711 2374 17720
rect 1950 16960 2006 16969
rect 1950 16895 2006 16904
rect 664 16720 716 16726
rect 664 16662 716 16668
rect 1858 16552 1914 16561
rect 1858 16487 1914 16496
rect 1872 15162 1900 16487
rect 1964 15706 1992 16895
rect 2332 15706 2360 17711
rect 1952 15700 2004 15706
rect 1952 15642 2004 15648
rect 2320 15700 2372 15706
rect 2320 15642 2372 15648
rect 2608 15162 2636 18119
rect 2686 17368 2742 17377
rect 2686 17303 2742 17312
rect 2700 15706 2728 17303
rect 2792 17218 2820 19343
rect 2884 18426 2912 20567
rect 2962 20224 3018 20233
rect 2962 20159 3018 20168
rect 2872 18420 2924 18426
rect 2872 18362 2924 18368
rect 2976 17338 3004 20159
rect 3054 19816 3110 19825
rect 3054 19751 3110 19760
rect 3068 17882 3096 19751
rect 3238 19000 3294 19009
rect 3238 18935 3294 18944
rect 3148 18284 3200 18290
rect 3148 18226 3200 18232
rect 3056 17876 3108 17882
rect 3056 17818 3108 17824
rect 3160 17354 3188 18226
rect 2964 17332 3016 17338
rect 2964 17274 3016 17280
rect 3068 17326 3188 17354
rect 2792 17190 2912 17218
rect 2780 17060 2832 17066
rect 2780 17002 2832 17008
rect 2792 16590 2820 17002
rect 2884 16998 2912 17190
rect 2964 17196 3016 17202
rect 2964 17138 3016 17144
rect 2872 16992 2924 16998
rect 2872 16934 2924 16940
rect 2976 16658 3004 17138
rect 2964 16652 3016 16658
rect 2964 16594 3016 16600
rect 2780 16584 2832 16590
rect 2780 16526 2832 16532
rect 3068 16182 3096 17326
rect 3148 17196 3200 17202
rect 3148 17138 3200 17144
rect 3160 16182 3188 17138
rect 3252 17066 3280 18935
rect 3344 17338 3372 22222
rect 3422 22200 3478 23000
rect 3882 22200 3938 23000
rect 4342 22200 4398 23000
rect 4802 22200 4858 23000
rect 5262 22200 5318 23000
rect 5722 22200 5778 23000
rect 6182 22200 6238 23000
rect 6642 22200 6698 23000
rect 7102 22200 7158 23000
rect 7562 22200 7618 23000
rect 8022 22200 8078 23000
rect 8482 22200 8538 23000
rect 8942 22200 8998 23000
rect 9048 22222 9352 22250
rect 3436 17882 3464 22200
rect 3549 20156 3857 20165
rect 3549 20154 3555 20156
rect 3611 20154 3635 20156
rect 3691 20154 3715 20156
rect 3771 20154 3795 20156
rect 3851 20154 3857 20156
rect 3611 20102 3613 20154
rect 3793 20102 3795 20154
rect 3549 20100 3555 20102
rect 3611 20100 3635 20102
rect 3691 20100 3715 20102
rect 3771 20100 3795 20102
rect 3851 20100 3857 20102
rect 3549 20091 3857 20100
rect 3549 19068 3857 19077
rect 3549 19066 3555 19068
rect 3611 19066 3635 19068
rect 3691 19066 3715 19068
rect 3771 19066 3795 19068
rect 3851 19066 3857 19068
rect 3611 19014 3613 19066
rect 3793 19014 3795 19066
rect 3549 19012 3555 19014
rect 3611 19012 3635 19014
rect 3691 19012 3715 19014
rect 3771 19012 3795 19014
rect 3851 19012 3857 19014
rect 3549 19003 3857 19012
rect 3896 18290 3924 22200
rect 4356 18426 4384 22200
rect 4620 18624 4672 18630
rect 4620 18566 4672 18572
rect 4344 18420 4396 18426
rect 4344 18362 4396 18368
rect 4436 18352 4488 18358
rect 4436 18294 4488 18300
rect 3884 18284 3936 18290
rect 3884 18226 3936 18232
rect 4344 18216 4396 18222
rect 4344 18158 4396 18164
rect 4160 18148 4212 18154
rect 4160 18090 4212 18096
rect 3884 18080 3936 18086
rect 3884 18022 3936 18028
rect 3549 17980 3857 17989
rect 3549 17978 3555 17980
rect 3611 17978 3635 17980
rect 3691 17978 3715 17980
rect 3771 17978 3795 17980
rect 3851 17978 3857 17980
rect 3611 17926 3613 17978
rect 3793 17926 3795 17978
rect 3549 17924 3555 17926
rect 3611 17924 3635 17926
rect 3691 17924 3715 17926
rect 3771 17924 3795 17926
rect 3851 17924 3857 17926
rect 3549 17915 3857 17924
rect 3424 17876 3476 17882
rect 3424 17818 3476 17824
rect 3424 17672 3476 17678
rect 3424 17614 3476 17620
rect 3332 17332 3384 17338
rect 3332 17274 3384 17280
rect 3436 17270 3464 17614
rect 3516 17604 3568 17610
rect 3516 17546 3568 17552
rect 3424 17264 3476 17270
rect 3424 17206 3476 17212
rect 3528 17082 3556 17546
rect 3240 17060 3292 17066
rect 3240 17002 3292 17008
rect 3436 17054 3556 17082
rect 3436 16726 3464 17054
rect 3549 16892 3857 16901
rect 3549 16890 3555 16892
rect 3611 16890 3635 16892
rect 3691 16890 3715 16892
rect 3771 16890 3795 16892
rect 3851 16890 3857 16892
rect 3611 16838 3613 16890
rect 3793 16838 3795 16890
rect 3549 16836 3555 16838
rect 3611 16836 3635 16838
rect 3691 16836 3715 16838
rect 3771 16836 3795 16838
rect 3851 16836 3857 16838
rect 3549 16827 3857 16836
rect 3896 16794 3924 18022
rect 4068 17332 4120 17338
rect 4068 17274 4120 17280
rect 3884 16788 3936 16794
rect 3884 16730 3936 16736
rect 3424 16720 3476 16726
rect 3424 16662 3476 16668
rect 3056 16176 3108 16182
rect 2870 16144 2926 16153
rect 3056 16118 3108 16124
rect 3148 16176 3200 16182
rect 3148 16118 3200 16124
rect 2870 16079 2926 16088
rect 2688 15700 2740 15706
rect 2688 15642 2740 15648
rect 1860 15156 1912 15162
rect 1860 15098 1912 15104
rect 2596 15156 2648 15162
rect 2596 15098 2648 15104
rect 2136 15020 2188 15026
rect 2136 14962 2188 14968
rect 1858 14104 1914 14113
rect 2148 14074 2176 14962
rect 2778 14512 2834 14521
rect 2778 14447 2834 14456
rect 1858 14039 1914 14048
rect 2136 14068 2188 14074
rect 1582 13696 1638 13705
rect 1582 13631 1638 13640
rect 1596 9450 1624 13631
rect 1766 12064 1822 12073
rect 1766 11999 1822 12008
rect 1780 10266 1808 11999
rect 1768 10260 1820 10266
rect 1768 10202 1820 10208
rect 1780 9926 1808 10202
rect 1768 9920 1820 9926
rect 1768 9862 1820 9868
rect 1584 9444 1636 9450
rect 1584 9386 1636 9392
rect 1674 9208 1730 9217
rect 1674 9143 1676 9152
rect 1728 9143 1730 9152
rect 1676 9114 1728 9120
rect 1676 8968 1728 8974
rect 1676 8910 1728 8916
rect 1490 8800 1546 8809
rect 1490 8735 1546 8744
rect 1504 8634 1532 8735
rect 1492 8628 1544 8634
rect 1492 8570 1544 8576
rect 1400 8356 1452 8362
rect 1400 8298 1452 8304
rect 1412 6118 1440 8298
rect 1504 8090 1532 8570
rect 1688 8362 1716 8910
rect 1676 8356 1728 8362
rect 1676 8298 1728 8304
rect 1492 8084 1544 8090
rect 1492 8026 1544 8032
rect 1504 6914 1532 8026
rect 1504 6886 1624 6914
rect 1596 6338 1624 6886
rect 1688 6633 1716 8298
rect 1780 7750 1808 9862
rect 1872 9450 1900 14039
rect 2136 14010 2188 14016
rect 2226 13832 2282 13841
rect 2226 13767 2282 13776
rect 1950 13288 2006 13297
rect 1950 13223 2006 13232
rect 1964 13190 1992 13223
rect 1952 13184 2004 13190
rect 1952 13126 2004 13132
rect 2136 9580 2188 9586
rect 2136 9522 2188 9528
rect 1860 9444 1912 9450
rect 1860 9386 1912 9392
rect 2044 9172 2096 9178
rect 2044 9114 2096 9120
rect 2056 7954 2084 9114
rect 2148 8566 2176 9522
rect 2240 9110 2268 13767
rect 2792 11354 2820 14447
rect 2884 12442 2912 16079
rect 3054 15736 3110 15745
rect 3054 15671 3110 15680
rect 3332 15700 3384 15706
rect 2962 14920 3018 14929
rect 2962 14855 3018 14864
rect 2872 12436 2924 12442
rect 2872 12378 2924 12384
rect 2870 11656 2926 11665
rect 2870 11591 2926 11600
rect 2780 11348 2832 11354
rect 2780 11290 2832 11296
rect 2780 10600 2832 10606
rect 2780 10542 2832 10548
rect 2792 10062 2820 10542
rect 2780 10056 2832 10062
rect 2780 9998 2832 10004
rect 2884 9908 2912 11591
rect 2976 10266 3004 14855
rect 3068 11286 3096 15671
rect 3332 15642 3384 15648
rect 3240 15428 3292 15434
rect 3240 15370 3292 15376
rect 3146 15328 3202 15337
rect 3146 15263 3202 15272
rect 3056 11280 3108 11286
rect 3056 11222 3108 11228
rect 3056 11144 3108 11150
rect 3056 11086 3108 11092
rect 2964 10260 3016 10266
rect 2964 10202 3016 10208
rect 2964 9920 3016 9926
rect 2884 9880 2964 9908
rect 2964 9862 3016 9868
rect 2780 9716 2832 9722
rect 2780 9658 2832 9664
rect 2228 9104 2280 9110
rect 2792 9058 2820 9658
rect 2872 9580 2924 9586
rect 2872 9522 2924 9528
rect 2228 9046 2280 9052
rect 2516 9042 2820 9058
rect 2504 9036 2820 9042
rect 2556 9030 2820 9036
rect 2504 8978 2556 8984
rect 2136 8560 2188 8566
rect 2136 8502 2188 8508
rect 2792 8498 2820 9030
rect 2780 8492 2832 8498
rect 2780 8434 2832 8440
rect 2780 8356 2832 8362
rect 2780 8298 2832 8304
rect 2792 8090 2820 8298
rect 2780 8084 2832 8090
rect 2780 8026 2832 8032
rect 2884 7954 2912 9522
rect 2044 7948 2096 7954
rect 2044 7890 2096 7896
rect 2872 7948 2924 7954
rect 2872 7890 2924 7896
rect 1768 7744 1820 7750
rect 1768 7686 1820 7692
rect 1780 7478 1808 7686
rect 2056 7546 2084 7890
rect 2504 7744 2556 7750
rect 2504 7686 2556 7692
rect 2044 7540 2096 7546
rect 2044 7482 2096 7488
rect 1768 7472 1820 7478
rect 1768 7414 1820 7420
rect 1674 6624 1730 6633
rect 1674 6559 1730 6568
rect 1504 6322 1624 6338
rect 1492 6316 1624 6322
rect 1544 6310 1624 6316
rect 1492 6258 1544 6264
rect 1400 6112 1452 6118
rect 1400 6054 1452 6060
rect 1412 5953 1440 6054
rect 1398 5944 1454 5953
rect 1504 5914 1532 6258
rect 1398 5879 1454 5888
rect 1492 5908 1544 5914
rect 1492 5850 1544 5856
rect 388 2916 440 2922
rect 388 2858 440 2864
rect 400 800 428 2858
rect 848 2440 900 2446
rect 848 2382 900 2388
rect 860 800 888 2382
rect 1688 2281 1716 6559
rect 1860 6248 1912 6254
rect 1912 6208 2084 6236
rect 1860 6190 1912 6196
rect 2056 5273 2084 6208
rect 2042 5264 2098 5273
rect 2042 5199 2098 5208
rect 2056 5166 2084 5199
rect 2044 5160 2096 5166
rect 2044 5102 2096 5108
rect 2228 4072 2280 4078
rect 2516 4049 2544 7686
rect 2870 7440 2926 7449
rect 2870 7375 2926 7384
rect 2228 4014 2280 4020
rect 2502 4040 2558 4049
rect 1768 3732 1820 3738
rect 1768 3674 1820 3680
rect 1674 2272 1730 2281
rect 1674 2207 1730 2216
rect 1308 2032 1360 2038
rect 1308 1974 1360 1980
rect 1320 800 1348 1974
rect 1780 800 1808 3674
rect 2240 800 2268 4014
rect 2502 3975 2558 3984
rect 2884 3097 2912 7375
rect 2976 5370 3004 9862
rect 3068 8022 3096 11086
rect 3160 9450 3188 15263
rect 3252 14822 3280 15370
rect 3344 15162 3372 15642
rect 3436 15366 3464 16662
rect 3608 16584 3660 16590
rect 3606 16552 3608 16561
rect 3660 16552 3662 16561
rect 3606 16487 3662 16496
rect 3896 16454 3924 16730
rect 3884 16448 3936 16454
rect 3884 16390 3936 16396
rect 3896 16266 3924 16390
rect 3896 16238 4016 16266
rect 4080 16250 4108 17274
rect 4172 17270 4200 18090
rect 4160 17264 4212 17270
rect 4160 17206 4212 17212
rect 4172 16522 4200 17206
rect 4356 16794 4384 18158
rect 4344 16788 4396 16794
rect 4344 16730 4396 16736
rect 4160 16516 4212 16522
rect 4160 16458 4212 16464
rect 3884 16108 3936 16114
rect 3884 16050 3936 16056
rect 3896 16017 3924 16050
rect 3988 16046 4016 16238
rect 4068 16244 4120 16250
rect 4068 16186 4120 16192
rect 3976 16040 4028 16046
rect 3882 16008 3938 16017
rect 3976 15982 4028 15988
rect 3882 15943 3938 15952
rect 3884 15904 3936 15910
rect 3884 15846 3936 15852
rect 3549 15804 3857 15813
rect 3549 15802 3555 15804
rect 3611 15802 3635 15804
rect 3691 15802 3715 15804
rect 3771 15802 3795 15804
rect 3851 15802 3857 15804
rect 3611 15750 3613 15802
rect 3793 15750 3795 15802
rect 3549 15748 3555 15750
rect 3611 15748 3635 15750
rect 3691 15748 3715 15750
rect 3771 15748 3795 15750
rect 3851 15748 3857 15750
rect 3549 15739 3857 15748
rect 3896 15638 3924 15846
rect 3884 15632 3936 15638
rect 3884 15574 3936 15580
rect 3424 15360 3476 15366
rect 3424 15302 3476 15308
rect 3436 15162 3464 15302
rect 3332 15156 3384 15162
rect 3332 15098 3384 15104
rect 3424 15156 3476 15162
rect 3424 15098 3476 15104
rect 3240 14816 3292 14822
rect 3240 14758 3292 14764
rect 3252 11665 3280 14758
rect 3436 14482 3464 15098
rect 3988 15026 4016 15982
rect 4080 15706 4108 16186
rect 4068 15700 4120 15706
rect 4068 15642 4120 15648
rect 4068 15360 4120 15366
rect 4068 15302 4120 15308
rect 4080 15026 4108 15302
rect 3976 15020 4028 15026
rect 3976 14962 4028 14968
rect 4068 15020 4120 15026
rect 4068 14962 4120 14968
rect 3884 14952 3936 14958
rect 3884 14894 3936 14900
rect 3549 14716 3857 14725
rect 3549 14714 3555 14716
rect 3611 14714 3635 14716
rect 3691 14714 3715 14716
rect 3771 14714 3795 14716
rect 3851 14714 3857 14716
rect 3611 14662 3613 14714
rect 3793 14662 3795 14714
rect 3549 14660 3555 14662
rect 3611 14660 3635 14662
rect 3691 14660 3715 14662
rect 3771 14660 3795 14662
rect 3851 14660 3857 14662
rect 3549 14651 3857 14660
rect 3424 14476 3476 14482
rect 3424 14418 3476 14424
rect 3549 13628 3857 13637
rect 3549 13626 3555 13628
rect 3611 13626 3635 13628
rect 3691 13626 3715 13628
rect 3771 13626 3795 13628
rect 3851 13626 3857 13628
rect 3611 13574 3613 13626
rect 3793 13574 3795 13626
rect 3549 13572 3555 13574
rect 3611 13572 3635 13574
rect 3691 13572 3715 13574
rect 3771 13572 3795 13574
rect 3851 13572 3857 13574
rect 3549 13563 3857 13572
rect 3332 13320 3384 13326
rect 3332 13262 3384 13268
rect 3344 12918 3372 13262
rect 3332 12912 3384 12918
rect 3332 12854 3384 12860
rect 3422 12880 3478 12889
rect 3422 12815 3478 12824
rect 3332 12640 3384 12646
rect 3332 12582 3384 12588
rect 3344 12481 3372 12582
rect 3330 12472 3386 12481
rect 3330 12407 3386 12416
rect 3238 11656 3294 11665
rect 3238 11591 3294 11600
rect 3240 11076 3292 11082
rect 3240 11018 3292 11024
rect 3148 9444 3200 9450
rect 3148 9386 3200 9392
rect 3252 9042 3280 11018
rect 3436 10810 3464 12815
rect 3549 12540 3857 12549
rect 3549 12538 3555 12540
rect 3611 12538 3635 12540
rect 3691 12538 3715 12540
rect 3771 12538 3795 12540
rect 3851 12538 3857 12540
rect 3611 12486 3613 12538
rect 3793 12486 3795 12538
rect 3549 12484 3555 12486
rect 3611 12484 3635 12486
rect 3691 12484 3715 12486
rect 3771 12484 3795 12486
rect 3851 12484 3857 12486
rect 3549 12475 3857 12484
rect 3549 11452 3857 11461
rect 3549 11450 3555 11452
rect 3611 11450 3635 11452
rect 3691 11450 3715 11452
rect 3771 11450 3795 11452
rect 3851 11450 3857 11452
rect 3611 11398 3613 11450
rect 3793 11398 3795 11450
rect 3549 11396 3555 11398
rect 3611 11396 3635 11398
rect 3691 11396 3715 11398
rect 3771 11396 3795 11398
rect 3851 11396 3857 11398
rect 3549 11387 3857 11396
rect 3424 10804 3476 10810
rect 3424 10746 3476 10752
rect 3332 10736 3384 10742
rect 3332 10678 3384 10684
rect 3344 10266 3372 10678
rect 3332 10260 3384 10266
rect 3332 10202 3384 10208
rect 3436 10146 3464 10746
rect 3549 10364 3857 10373
rect 3549 10362 3555 10364
rect 3611 10362 3635 10364
rect 3691 10362 3715 10364
rect 3771 10362 3795 10364
rect 3851 10362 3857 10364
rect 3611 10310 3613 10362
rect 3793 10310 3795 10362
rect 3549 10308 3555 10310
rect 3611 10308 3635 10310
rect 3691 10308 3715 10310
rect 3771 10308 3795 10310
rect 3851 10308 3857 10310
rect 3549 10299 3857 10308
rect 3896 10146 3924 14894
rect 4068 14816 4120 14822
rect 4068 14758 4120 14764
rect 4080 13297 4108 14758
rect 4172 14618 4200 16458
rect 4356 16250 4384 16730
rect 4344 16244 4396 16250
rect 4344 16186 4396 16192
rect 4252 15564 4304 15570
rect 4252 15506 4304 15512
rect 4160 14612 4212 14618
rect 4160 14554 4212 14560
rect 4172 14414 4200 14554
rect 4160 14408 4212 14414
rect 4160 14350 4212 14356
rect 4160 14068 4212 14074
rect 4160 14010 4212 14016
rect 4066 13288 4122 13297
rect 4066 13223 4122 13232
rect 4068 12232 4120 12238
rect 4068 12174 4120 12180
rect 4080 10962 4108 12174
rect 4172 11830 4200 14010
rect 4264 12918 4292 15506
rect 4356 15366 4384 16186
rect 4344 15360 4396 15366
rect 4344 15302 4396 15308
rect 4448 15162 4476 18294
rect 4528 17876 4580 17882
rect 4528 17818 4580 17824
rect 4540 17338 4568 17818
rect 4528 17332 4580 17338
rect 4528 17274 4580 17280
rect 4436 15156 4488 15162
rect 4436 15098 4488 15104
rect 4344 15088 4396 15094
rect 4344 15030 4396 15036
rect 4356 13682 4384 15030
rect 4448 14822 4476 15098
rect 4436 14816 4488 14822
rect 4436 14758 4488 14764
rect 4448 14550 4476 14758
rect 4436 14544 4488 14550
rect 4436 14486 4488 14492
rect 4540 14346 4568 17274
rect 4632 16998 4660 18566
rect 4816 18154 4844 22200
rect 5080 18284 5132 18290
rect 5080 18226 5132 18232
rect 4804 18148 4856 18154
rect 4804 18090 4856 18096
rect 4988 17672 5040 17678
rect 4908 17632 4988 17660
rect 4908 17134 4936 17632
rect 4988 17614 5040 17620
rect 4988 17536 5040 17542
rect 4988 17478 5040 17484
rect 5000 17338 5028 17478
rect 4988 17332 5040 17338
rect 4988 17274 5040 17280
rect 4896 17128 4948 17134
rect 4896 17070 4948 17076
rect 4620 16992 4672 16998
rect 4620 16934 4672 16940
rect 4632 15586 4660 16934
rect 4908 16658 4936 17070
rect 4896 16652 4948 16658
rect 4896 16594 4948 16600
rect 4908 16454 4936 16594
rect 4896 16448 4948 16454
rect 4896 16390 4948 16396
rect 4988 15904 5040 15910
rect 4988 15846 5040 15852
rect 4804 15700 4856 15706
rect 4804 15642 4856 15648
rect 4632 15558 4752 15586
rect 4724 15502 4752 15558
rect 4816 15502 4844 15642
rect 4712 15496 4764 15502
rect 4712 15438 4764 15444
rect 4804 15496 4856 15502
rect 4804 15438 4856 15444
rect 4620 15428 4672 15434
rect 4620 15370 4672 15376
rect 4632 15178 4660 15370
rect 4632 15150 4752 15178
rect 4620 14884 4672 14890
rect 4620 14826 4672 14832
rect 4632 14793 4660 14826
rect 4618 14784 4674 14793
rect 4618 14719 4674 14728
rect 4528 14340 4580 14346
rect 4528 14282 4580 14288
rect 4540 14074 4568 14282
rect 4528 14068 4580 14074
rect 4528 14010 4580 14016
rect 4356 13654 4660 13682
rect 4252 12912 4304 12918
rect 4252 12854 4304 12860
rect 4528 12844 4580 12850
rect 4528 12786 4580 12792
rect 4252 12640 4304 12646
rect 4252 12582 4304 12588
rect 4160 11824 4212 11830
rect 4160 11766 4212 11772
rect 4264 11082 4292 12582
rect 4540 12374 4568 12786
rect 4528 12368 4580 12374
rect 4528 12310 4580 12316
rect 4436 11756 4488 11762
rect 4436 11698 4488 11704
rect 4448 11286 4476 11698
rect 4436 11280 4488 11286
rect 4436 11222 4488 11228
rect 4344 11212 4396 11218
rect 4344 11154 4396 11160
rect 4252 11076 4304 11082
rect 4252 11018 4304 11024
rect 4080 10934 4200 10962
rect 4066 10840 4122 10849
rect 4066 10775 4122 10784
rect 3976 10464 4028 10470
rect 3976 10406 4028 10412
rect 3344 10118 3464 10146
rect 3804 10130 3924 10146
rect 3792 10124 3924 10130
rect 3240 9036 3292 9042
rect 3240 8978 3292 8984
rect 3148 8900 3200 8906
rect 3148 8842 3200 8848
rect 3056 8016 3108 8022
rect 3056 7958 3108 7964
rect 3056 7880 3108 7886
rect 3056 7822 3108 7828
rect 3068 7478 3096 7822
rect 3056 7472 3108 7478
rect 3056 7414 3108 7420
rect 3160 6361 3188 8842
rect 3344 8498 3372 10118
rect 3844 10118 3924 10124
rect 3792 10066 3844 10072
rect 3700 10056 3752 10062
rect 3700 9998 3752 10004
rect 3424 9988 3476 9994
rect 3424 9930 3476 9936
rect 3436 8906 3464 9930
rect 3712 9382 3740 9998
rect 3804 9722 3832 10066
rect 3988 10033 4016 10406
rect 4080 10266 4108 10775
rect 4068 10260 4120 10266
rect 4068 10202 4120 10208
rect 4172 10146 4200 10934
rect 4080 10118 4200 10146
rect 3974 10024 4030 10033
rect 3974 9959 4030 9968
rect 3882 9888 3938 9897
rect 3882 9823 3938 9832
rect 3896 9722 3924 9823
rect 3792 9716 3844 9722
rect 3792 9658 3844 9664
rect 3884 9716 3936 9722
rect 3884 9658 3936 9664
rect 3790 9616 3846 9625
rect 3790 9551 3846 9560
rect 3804 9518 3832 9551
rect 3792 9512 3844 9518
rect 3792 9454 3844 9460
rect 3700 9376 3752 9382
rect 3700 9318 3752 9324
rect 3884 9376 3936 9382
rect 3884 9318 3936 9324
rect 3549 9276 3857 9285
rect 3549 9274 3555 9276
rect 3611 9274 3635 9276
rect 3691 9274 3715 9276
rect 3771 9274 3795 9276
rect 3851 9274 3857 9276
rect 3611 9222 3613 9274
rect 3793 9222 3795 9274
rect 3549 9220 3555 9222
rect 3611 9220 3635 9222
rect 3691 9220 3715 9222
rect 3771 9220 3795 9222
rect 3851 9220 3857 9222
rect 3549 9211 3857 9220
rect 3424 8900 3476 8906
rect 3424 8842 3476 8848
rect 3700 8832 3752 8838
rect 3700 8774 3752 8780
rect 3332 8492 3384 8498
rect 3332 8434 3384 8440
rect 3712 8430 3740 8774
rect 3424 8424 3476 8430
rect 3424 8366 3476 8372
rect 3700 8424 3752 8430
rect 3700 8366 3752 8372
rect 3436 7177 3464 8366
rect 3549 8188 3857 8197
rect 3549 8186 3555 8188
rect 3611 8186 3635 8188
rect 3691 8186 3715 8188
rect 3771 8186 3795 8188
rect 3851 8186 3857 8188
rect 3611 8134 3613 8186
rect 3793 8134 3795 8186
rect 3549 8132 3555 8134
rect 3611 8132 3635 8134
rect 3691 8132 3715 8134
rect 3771 8132 3795 8134
rect 3851 8132 3857 8134
rect 3549 8123 3857 8132
rect 3896 8090 3924 9318
rect 3988 9042 4016 9959
rect 3976 9036 4028 9042
rect 3976 8978 4028 8984
rect 3988 8498 4016 8978
rect 3976 8492 4028 8498
rect 3976 8434 4028 8440
rect 3884 8084 3936 8090
rect 4080 8072 4108 10118
rect 4160 9580 4212 9586
rect 4160 9522 4212 9528
rect 3884 8026 3936 8032
rect 3988 8044 4108 8072
rect 3988 7886 4016 8044
rect 3976 7880 4028 7886
rect 3976 7822 4028 7828
rect 3974 7576 4030 7585
rect 3974 7511 4030 7520
rect 3988 7274 4016 7511
rect 3976 7268 4028 7274
rect 3976 7210 4028 7216
rect 3422 7168 3478 7177
rect 3422 7103 3478 7112
rect 3549 7100 3857 7109
rect 3549 7098 3555 7100
rect 3611 7098 3635 7100
rect 3691 7098 3715 7100
rect 3771 7098 3795 7100
rect 3851 7098 3857 7100
rect 3611 7046 3613 7098
rect 3793 7046 3795 7098
rect 3549 7044 3555 7046
rect 3611 7044 3635 7046
rect 3691 7044 3715 7046
rect 3771 7044 3795 7046
rect 3851 7044 3857 7046
rect 3549 7035 3857 7044
rect 4172 6866 4200 9522
rect 4264 8786 4292 11018
rect 4356 9518 4384 11154
rect 4436 11144 4488 11150
rect 4436 11086 4488 11092
rect 4448 10606 4476 11086
rect 4436 10600 4488 10606
rect 4436 10542 4488 10548
rect 4436 10260 4488 10266
rect 4488 10220 4568 10248
rect 4436 10202 4488 10208
rect 4344 9512 4396 9518
rect 4344 9454 4396 9460
rect 4436 9444 4488 9450
rect 4436 9386 4488 9392
rect 4344 8968 4396 8974
rect 4342 8936 4344 8945
rect 4396 8936 4398 8945
rect 4342 8871 4398 8880
rect 4264 8758 4384 8786
rect 4250 7984 4306 7993
rect 4250 7919 4306 7928
rect 4264 7546 4292 7919
rect 4252 7540 4304 7546
rect 4252 7482 4304 7488
rect 3976 6860 4028 6866
rect 3976 6802 4028 6808
rect 4160 6860 4212 6866
rect 4160 6802 4212 6808
rect 3424 6792 3476 6798
rect 3422 6760 3424 6769
rect 3476 6760 3478 6769
rect 3422 6695 3478 6704
rect 3146 6352 3202 6361
rect 3146 6287 3202 6296
rect 3330 6352 3386 6361
rect 3330 6287 3386 6296
rect 2964 5364 3016 5370
rect 2964 5306 3016 5312
rect 3160 3670 3188 6287
rect 3344 6202 3372 6287
rect 3988 6254 4016 6802
rect 4356 6390 4384 8758
rect 4448 6798 4476 9386
rect 4540 7410 4568 10220
rect 4632 10130 4660 13654
rect 4724 13394 4752 15150
rect 4816 15026 4936 15042
rect 4804 15020 4936 15026
rect 4856 15014 4936 15020
rect 4804 14962 4856 14968
rect 4804 14884 4856 14890
rect 4804 14826 4856 14832
rect 4816 13734 4844 14826
rect 4908 14618 4936 15014
rect 4896 14612 4948 14618
rect 4896 14554 4948 14560
rect 4804 13728 4856 13734
rect 4804 13670 4856 13676
rect 4804 13524 4856 13530
rect 4804 13466 4856 13472
rect 4712 13388 4764 13394
rect 4712 13330 4764 13336
rect 4816 11014 4844 13466
rect 5000 12306 5028 15846
rect 5092 13462 5120 18226
rect 5276 18170 5304 22200
rect 5276 18142 5672 18170
rect 5356 18080 5408 18086
rect 5356 18022 5408 18028
rect 5368 17746 5396 18022
rect 5172 17740 5224 17746
rect 5172 17682 5224 17688
rect 5356 17740 5408 17746
rect 5356 17682 5408 17688
rect 5184 17134 5212 17682
rect 5540 17196 5592 17202
rect 5540 17138 5592 17144
rect 5172 17128 5224 17134
rect 5172 17070 5224 17076
rect 5448 17128 5500 17134
rect 5448 17070 5500 17076
rect 5356 16448 5408 16454
rect 5356 16390 5408 16396
rect 5172 16108 5224 16114
rect 5172 16050 5224 16056
rect 5184 15706 5212 16050
rect 5264 16040 5316 16046
rect 5264 15982 5316 15988
rect 5172 15700 5224 15706
rect 5172 15642 5224 15648
rect 5276 15434 5304 15982
rect 5264 15428 5316 15434
rect 5264 15370 5316 15376
rect 5368 15065 5396 16390
rect 5354 15056 5410 15065
rect 5354 14991 5410 15000
rect 5356 14952 5408 14958
rect 5262 14920 5318 14929
rect 5356 14894 5408 14900
rect 5262 14855 5318 14864
rect 5276 14482 5304 14855
rect 5264 14476 5316 14482
rect 5264 14418 5316 14424
rect 5368 14074 5396 14894
rect 5356 14068 5408 14074
rect 5356 14010 5408 14016
rect 5172 13864 5224 13870
rect 5172 13806 5224 13812
rect 5080 13456 5132 13462
rect 5080 13398 5132 13404
rect 4988 12300 5040 12306
rect 4988 12242 5040 12248
rect 4988 11688 5040 11694
rect 4988 11630 5040 11636
rect 5078 11656 5134 11665
rect 4894 11248 4950 11257
rect 4894 11183 4950 11192
rect 4804 11008 4856 11014
rect 4804 10950 4856 10956
rect 4620 10124 4672 10130
rect 4620 10066 4672 10072
rect 4620 9036 4672 9042
rect 4620 8978 4672 8984
rect 4632 8430 4660 8978
rect 4620 8424 4672 8430
rect 4620 8366 4672 8372
rect 4620 7812 4672 7818
rect 4620 7754 4672 7760
rect 4712 7812 4764 7818
rect 4712 7754 4764 7760
rect 4528 7404 4580 7410
rect 4528 7346 4580 7352
rect 4436 6792 4488 6798
rect 4436 6734 4488 6740
rect 4344 6384 4396 6390
rect 4344 6326 4396 6332
rect 4252 6316 4304 6322
rect 4252 6258 4304 6264
rect 3252 6174 3372 6202
rect 3976 6248 4028 6254
rect 3976 6190 4028 6196
rect 3148 3664 3200 3670
rect 3148 3606 3200 3612
rect 3252 3505 3280 6174
rect 3549 6012 3857 6021
rect 3549 6010 3555 6012
rect 3611 6010 3635 6012
rect 3691 6010 3715 6012
rect 3771 6010 3795 6012
rect 3851 6010 3857 6012
rect 3611 5958 3613 6010
rect 3793 5958 3795 6010
rect 3549 5956 3555 5958
rect 3611 5956 3635 5958
rect 3691 5956 3715 5958
rect 3771 5956 3795 5958
rect 3851 5956 3857 5958
rect 3549 5947 3857 5956
rect 3974 5400 4030 5409
rect 3792 5364 3844 5370
rect 3974 5335 4030 5344
rect 3792 5306 3844 5312
rect 3804 5166 3832 5306
rect 3792 5160 3844 5166
rect 3790 5128 3792 5137
rect 3844 5128 3846 5137
rect 3790 5063 3846 5072
rect 3549 4924 3857 4933
rect 3549 4922 3555 4924
rect 3611 4922 3635 4924
rect 3691 4922 3715 4924
rect 3771 4922 3795 4924
rect 3851 4922 3857 4924
rect 3611 4870 3613 4922
rect 3793 4870 3795 4922
rect 3549 4868 3555 4870
rect 3611 4868 3635 4870
rect 3691 4868 3715 4870
rect 3771 4868 3795 4870
rect 3851 4868 3857 4870
rect 3549 4859 3857 4868
rect 3424 4752 3476 4758
rect 3988 4729 4016 5335
rect 4068 5228 4120 5234
rect 4068 5170 4120 5176
rect 4080 5030 4108 5170
rect 4264 5098 4292 6258
rect 4528 5636 4580 5642
rect 4528 5578 4580 5584
rect 4252 5092 4304 5098
rect 4252 5034 4304 5040
rect 4068 5024 4120 5030
rect 4068 4966 4120 4972
rect 4160 5024 4212 5030
rect 4160 4966 4212 4972
rect 3424 4694 3476 4700
rect 3974 4720 4030 4729
rect 3332 4004 3384 4010
rect 3332 3946 3384 3952
rect 3344 3913 3372 3946
rect 3330 3904 3386 3913
rect 3330 3839 3386 3848
rect 3238 3496 3294 3505
rect 3238 3431 3294 3440
rect 2870 3088 2926 3097
rect 2870 3023 2926 3032
rect 3436 2922 3464 4694
rect 3974 4655 4030 4664
rect 4080 4554 4108 4966
rect 4068 4548 4120 4554
rect 4068 4490 4120 4496
rect 3976 4140 4028 4146
rect 3976 4082 4028 4088
rect 3549 3836 3857 3845
rect 3549 3834 3555 3836
rect 3611 3834 3635 3836
rect 3691 3834 3715 3836
rect 3771 3834 3795 3836
rect 3851 3834 3857 3836
rect 3611 3782 3613 3834
rect 3793 3782 3795 3834
rect 3549 3780 3555 3782
rect 3611 3780 3635 3782
rect 3691 3780 3715 3782
rect 3771 3780 3795 3782
rect 3851 3780 3857 3782
rect 3549 3771 3857 3780
rect 3884 3392 3936 3398
rect 3884 3334 3936 3340
rect 3424 2916 3476 2922
rect 3424 2858 3476 2864
rect 3549 2748 3857 2757
rect 3549 2746 3555 2748
rect 3611 2746 3635 2748
rect 3691 2746 3715 2748
rect 3771 2746 3795 2748
rect 3851 2746 3857 2748
rect 3611 2694 3613 2746
rect 3793 2694 3795 2746
rect 3549 2692 3555 2694
rect 3611 2692 3635 2694
rect 3691 2692 3715 2694
rect 3771 2692 3795 2694
rect 3851 2692 3857 2694
rect 3422 2680 3478 2689
rect 3549 2683 3857 2692
rect 3422 2615 3478 2624
rect 3436 2582 3464 2615
rect 3424 2576 3476 2582
rect 3424 2518 3476 2524
rect 2688 2372 2740 2378
rect 2688 2314 2740 2320
rect 2700 800 2728 2314
rect 3148 2304 3200 2310
rect 3148 2246 3200 2252
rect 3160 800 3188 2246
rect 3424 2100 3476 2106
rect 3424 2042 3476 2048
rect 3436 1873 3464 2042
rect 3422 1864 3478 1873
rect 3422 1799 3478 1808
rect 3620 870 3740 898
rect 3620 800 3648 870
rect 386 0 442 800
rect 846 0 902 800
rect 1306 0 1362 800
rect 1766 0 1822 800
rect 2226 0 2282 800
rect 2686 0 2742 800
rect 3146 0 3202 800
rect 3606 0 3662 800
rect 3712 762 3740 870
rect 3896 762 3924 3334
rect 3988 2122 4016 4082
rect 4080 2310 4108 4490
rect 4172 4078 4200 4966
rect 4160 4072 4212 4078
rect 4160 4014 4212 4020
rect 4068 2304 4120 2310
rect 4068 2246 4120 2252
rect 3988 2094 4108 2122
rect 4080 800 4108 2094
rect 4540 800 4568 5578
rect 4632 3942 4660 7754
rect 4724 5370 4752 7754
rect 4712 5364 4764 5370
rect 4712 5306 4764 5312
rect 4712 5160 4764 5166
rect 4712 5102 4764 5108
rect 4724 4729 4752 5102
rect 4710 4720 4766 4729
rect 4710 4655 4766 4664
rect 4816 4321 4844 10950
rect 4908 9489 4936 11183
rect 5000 11082 5028 11630
rect 5078 11591 5134 11600
rect 5092 11257 5120 11591
rect 5078 11248 5134 11257
rect 5078 11183 5134 11192
rect 4988 11076 5040 11082
rect 4988 11018 5040 11024
rect 5092 10062 5120 11183
rect 5184 10810 5212 13806
rect 5460 13802 5488 17070
rect 5552 16590 5580 17138
rect 5540 16584 5592 16590
rect 5540 16526 5592 16532
rect 5540 16448 5592 16454
rect 5540 16390 5592 16396
rect 5552 16182 5580 16390
rect 5540 16176 5592 16182
rect 5540 16118 5592 16124
rect 5644 15570 5672 18142
rect 5736 17678 5764 22200
rect 6196 20890 6224 22200
rect 6012 20862 6224 20890
rect 5724 17672 5776 17678
rect 5724 17614 5776 17620
rect 5724 17536 5776 17542
rect 5724 17478 5776 17484
rect 5908 17536 5960 17542
rect 5908 17478 5960 17484
rect 5736 17270 5764 17478
rect 5920 17354 5948 17478
rect 5828 17338 5948 17354
rect 5816 17332 5948 17338
rect 5868 17326 5948 17332
rect 5816 17274 5868 17280
rect 5724 17264 5776 17270
rect 5724 17206 5776 17212
rect 6012 16697 6040 20862
rect 6148 20700 6456 20709
rect 6148 20698 6154 20700
rect 6210 20698 6234 20700
rect 6290 20698 6314 20700
rect 6370 20698 6394 20700
rect 6450 20698 6456 20700
rect 6210 20646 6212 20698
rect 6392 20646 6394 20698
rect 6148 20644 6154 20646
rect 6210 20644 6234 20646
rect 6290 20644 6314 20646
rect 6370 20644 6394 20646
rect 6450 20644 6456 20646
rect 6148 20635 6456 20644
rect 6148 19612 6456 19621
rect 6148 19610 6154 19612
rect 6210 19610 6234 19612
rect 6290 19610 6314 19612
rect 6370 19610 6394 19612
rect 6450 19610 6456 19612
rect 6210 19558 6212 19610
rect 6392 19558 6394 19610
rect 6148 19556 6154 19558
rect 6210 19556 6234 19558
rect 6290 19556 6314 19558
rect 6370 19556 6394 19558
rect 6450 19556 6456 19558
rect 6148 19547 6456 19556
rect 6148 18524 6456 18533
rect 6148 18522 6154 18524
rect 6210 18522 6234 18524
rect 6290 18522 6314 18524
rect 6370 18522 6394 18524
rect 6450 18522 6456 18524
rect 6210 18470 6212 18522
rect 6392 18470 6394 18522
rect 6148 18468 6154 18470
rect 6210 18468 6234 18470
rect 6290 18468 6314 18470
rect 6370 18468 6394 18470
rect 6450 18468 6456 18470
rect 6148 18459 6456 18468
rect 6092 18216 6144 18222
rect 6092 18158 6144 18164
rect 6104 18086 6132 18158
rect 6092 18080 6144 18086
rect 6656 18057 6684 22200
rect 6736 19712 6788 19718
rect 6736 19654 6788 19660
rect 6092 18022 6144 18028
rect 6642 18048 6698 18057
rect 6104 17746 6132 18022
rect 6642 17983 6698 17992
rect 6092 17740 6144 17746
rect 6092 17682 6144 17688
rect 6644 17672 6696 17678
rect 6644 17614 6696 17620
rect 6552 17536 6604 17542
rect 6552 17478 6604 17484
rect 6148 17436 6456 17445
rect 6148 17434 6154 17436
rect 6210 17434 6234 17436
rect 6290 17434 6314 17436
rect 6370 17434 6394 17436
rect 6450 17434 6456 17436
rect 6210 17382 6212 17434
rect 6392 17382 6394 17434
rect 6148 17380 6154 17382
rect 6210 17380 6234 17382
rect 6290 17380 6314 17382
rect 6370 17380 6394 17382
rect 6450 17380 6456 17382
rect 6148 17371 6456 17380
rect 6182 17096 6238 17105
rect 6182 17031 6238 17040
rect 5998 16688 6054 16697
rect 6196 16658 6224 17031
rect 6564 16998 6592 17478
rect 6552 16992 6604 16998
rect 6552 16934 6604 16940
rect 6552 16788 6604 16794
rect 6552 16730 6604 16736
rect 5998 16623 6054 16632
rect 6184 16652 6236 16658
rect 6184 16594 6236 16600
rect 5724 16584 5776 16590
rect 5724 16526 5776 16532
rect 5736 15994 5764 16526
rect 5908 16448 5960 16454
rect 5908 16390 5960 16396
rect 6000 16448 6052 16454
rect 6000 16390 6052 16396
rect 5920 16250 5948 16390
rect 5908 16244 5960 16250
rect 5908 16186 5960 16192
rect 6012 16130 6040 16390
rect 6148 16348 6456 16357
rect 6148 16346 6154 16348
rect 6210 16346 6234 16348
rect 6290 16346 6314 16348
rect 6370 16346 6394 16348
rect 6450 16346 6456 16348
rect 6210 16294 6212 16346
rect 6392 16294 6394 16346
rect 6148 16292 6154 16294
rect 6210 16292 6234 16294
rect 6290 16292 6314 16294
rect 6370 16292 6394 16294
rect 6450 16292 6456 16294
rect 6148 16283 6456 16292
rect 6564 16182 6592 16730
rect 6552 16176 6604 16182
rect 6012 16102 6132 16130
rect 6552 16118 6604 16124
rect 6000 16040 6052 16046
rect 5736 15978 5856 15994
rect 6000 15982 6052 15988
rect 5736 15972 5868 15978
rect 5736 15966 5816 15972
rect 5816 15914 5868 15920
rect 5632 15564 5684 15570
rect 5632 15506 5684 15512
rect 5540 15496 5592 15502
rect 5540 15438 5592 15444
rect 5552 14890 5580 15438
rect 5644 15162 5672 15506
rect 5828 15434 5856 15914
rect 6012 15706 6040 15982
rect 6104 15706 6132 16102
rect 6368 16108 6420 16114
rect 6368 16050 6420 16056
rect 6380 15910 6408 16050
rect 6368 15904 6420 15910
rect 6368 15846 6420 15852
rect 6000 15700 6052 15706
rect 6000 15642 6052 15648
rect 6092 15700 6144 15706
rect 6092 15642 6144 15648
rect 5816 15428 5868 15434
rect 5816 15370 5868 15376
rect 5632 15156 5684 15162
rect 5632 15098 5684 15104
rect 5724 15020 5776 15026
rect 5724 14962 5776 14968
rect 5540 14884 5592 14890
rect 5540 14826 5592 14832
rect 5448 13796 5500 13802
rect 5448 13738 5500 13744
rect 5552 13530 5580 14826
rect 5632 14816 5684 14822
rect 5632 14758 5684 14764
rect 5644 14550 5672 14758
rect 5632 14544 5684 14550
rect 5632 14486 5684 14492
rect 5736 14074 5764 14962
rect 5724 14068 5776 14074
rect 5724 14010 5776 14016
rect 5828 13954 5856 15370
rect 6380 15366 6408 15846
rect 6368 15360 6420 15366
rect 6368 15302 6420 15308
rect 6148 15260 6456 15269
rect 6148 15258 6154 15260
rect 6210 15258 6234 15260
rect 6290 15258 6314 15260
rect 6370 15258 6394 15260
rect 6450 15258 6456 15260
rect 6210 15206 6212 15258
rect 6392 15206 6394 15258
rect 6148 15204 6154 15206
rect 6210 15204 6234 15206
rect 6290 15204 6314 15206
rect 6370 15204 6394 15206
rect 6450 15204 6456 15206
rect 6148 15195 6456 15204
rect 6552 14272 6604 14278
rect 6552 14214 6604 14220
rect 6148 14172 6456 14181
rect 6148 14170 6154 14172
rect 6210 14170 6234 14172
rect 6290 14170 6314 14172
rect 6370 14170 6394 14172
rect 6450 14170 6456 14172
rect 6210 14118 6212 14170
rect 6392 14118 6394 14170
rect 6148 14116 6154 14118
rect 6210 14116 6234 14118
rect 6290 14116 6314 14118
rect 6370 14116 6394 14118
rect 6450 14116 6456 14118
rect 6148 14107 6456 14116
rect 6564 14074 6592 14214
rect 6552 14068 6604 14074
rect 6552 14010 6604 14016
rect 5736 13926 5856 13954
rect 6550 13968 6606 13977
rect 5540 13524 5592 13530
rect 5540 13466 5592 13472
rect 5448 13456 5500 13462
rect 5448 13398 5500 13404
rect 5356 13252 5408 13258
rect 5356 13194 5408 13200
rect 5262 12880 5318 12889
rect 5262 12815 5318 12824
rect 5276 12782 5304 12815
rect 5264 12776 5316 12782
rect 5264 12718 5316 12724
rect 5172 10804 5224 10810
rect 5172 10746 5224 10752
rect 5170 10160 5226 10169
rect 5170 10095 5226 10104
rect 5080 10056 5132 10062
rect 5080 9998 5132 10004
rect 4988 9988 5040 9994
rect 4988 9930 5040 9936
rect 4894 9480 4950 9489
rect 4894 9415 4950 9424
rect 4908 4826 4936 9415
rect 5000 9382 5028 9930
rect 4988 9376 5040 9382
rect 4988 9318 5040 9324
rect 5078 9208 5134 9217
rect 5078 9143 5134 9152
rect 5092 9110 5120 9143
rect 5080 9104 5132 9110
rect 5080 9046 5132 9052
rect 5080 8900 5132 8906
rect 5080 8842 5132 8848
rect 5092 8809 5120 8842
rect 5078 8800 5134 8809
rect 5078 8735 5134 8744
rect 5184 8566 5212 10095
rect 5264 10056 5316 10062
rect 5262 10024 5264 10033
rect 5316 10024 5318 10033
rect 5262 9959 5318 9968
rect 5264 9580 5316 9586
rect 5264 9522 5316 9528
rect 5276 9330 5304 9522
rect 5368 9450 5396 13194
rect 5460 12782 5488 13398
rect 5632 12844 5684 12850
rect 5632 12786 5684 12792
rect 5448 12776 5500 12782
rect 5448 12718 5500 12724
rect 5540 12708 5592 12714
rect 5540 12650 5592 12656
rect 5448 12164 5500 12170
rect 5448 12106 5500 12112
rect 5460 11898 5488 12106
rect 5448 11892 5500 11898
rect 5448 11834 5500 11840
rect 5460 11218 5488 11834
rect 5552 11354 5580 12650
rect 5644 12442 5672 12786
rect 5632 12436 5684 12442
rect 5632 12378 5684 12384
rect 5632 11620 5684 11626
rect 5632 11562 5684 11568
rect 5540 11348 5592 11354
rect 5540 11290 5592 11296
rect 5644 11218 5672 11562
rect 5448 11212 5500 11218
rect 5448 11154 5500 11160
rect 5632 11212 5684 11218
rect 5632 11154 5684 11160
rect 5630 11112 5686 11121
rect 5630 11047 5686 11056
rect 5540 10668 5592 10674
rect 5540 10610 5592 10616
rect 5448 10600 5500 10606
rect 5448 10542 5500 10548
rect 5460 10266 5488 10542
rect 5448 10260 5500 10266
rect 5448 10202 5500 10208
rect 5552 10130 5580 10610
rect 5540 10124 5592 10130
rect 5540 10066 5592 10072
rect 5540 9920 5592 9926
rect 5540 9862 5592 9868
rect 5446 9616 5502 9625
rect 5552 9586 5580 9862
rect 5446 9551 5502 9560
rect 5540 9580 5592 9586
rect 5356 9444 5408 9450
rect 5356 9386 5408 9392
rect 5276 9302 5396 9330
rect 5262 9072 5318 9081
rect 5262 9007 5318 9016
rect 5172 8560 5224 8566
rect 5172 8502 5224 8508
rect 5080 8424 5132 8430
rect 5080 8366 5132 8372
rect 5092 8294 5120 8366
rect 5080 8288 5132 8294
rect 5080 8230 5132 8236
rect 4988 8084 5040 8090
rect 4988 8026 5040 8032
rect 5000 7750 5028 8026
rect 5092 7954 5120 8230
rect 5080 7948 5132 7954
rect 5080 7890 5132 7896
rect 5092 7750 5120 7890
rect 5276 7818 5304 9007
rect 5264 7812 5316 7818
rect 5264 7754 5316 7760
rect 4988 7744 5040 7750
rect 4988 7686 5040 7692
rect 5080 7744 5132 7750
rect 5080 7686 5132 7692
rect 5000 7546 5028 7686
rect 4988 7540 5040 7546
rect 4988 7482 5040 7488
rect 5172 7336 5224 7342
rect 5172 7278 5224 7284
rect 5184 6662 5212 7278
rect 4988 6656 5040 6662
rect 4988 6598 5040 6604
rect 5172 6656 5224 6662
rect 5172 6598 5224 6604
rect 5000 6254 5028 6598
rect 4988 6248 5040 6254
rect 4988 6190 5040 6196
rect 5000 5574 5028 6190
rect 5184 5574 5212 6598
rect 5264 5772 5316 5778
rect 5264 5714 5316 5720
rect 4988 5568 5040 5574
rect 4988 5510 5040 5516
rect 5172 5568 5224 5574
rect 5172 5510 5224 5516
rect 4896 4820 4948 4826
rect 4896 4762 4948 4768
rect 4908 4622 4936 4762
rect 4896 4616 4948 4622
rect 4896 4558 4948 4564
rect 4802 4312 4858 4321
rect 4802 4247 4858 4256
rect 4620 3936 4672 3942
rect 5000 3913 5028 5510
rect 5080 5364 5132 5370
rect 5080 5306 5132 5312
rect 5092 5273 5120 5306
rect 5078 5264 5134 5273
rect 5184 5234 5212 5510
rect 5078 5199 5134 5208
rect 5172 5228 5224 5234
rect 5172 5170 5224 5176
rect 5170 5128 5226 5137
rect 5170 5063 5172 5072
rect 5224 5063 5226 5072
rect 5172 5034 5224 5040
rect 5276 4690 5304 5714
rect 5264 4684 5316 4690
rect 5264 4626 5316 4632
rect 5276 4282 5304 4626
rect 5264 4276 5316 4282
rect 5264 4218 5316 4224
rect 4620 3878 4672 3884
rect 4986 3904 5042 3913
rect 4986 3839 5042 3848
rect 5080 3392 5132 3398
rect 5080 3334 5132 3340
rect 5092 3194 5120 3334
rect 5080 3188 5132 3194
rect 5080 3130 5132 3136
rect 4988 2984 5040 2990
rect 4988 2926 5040 2932
rect 5000 2650 5028 2926
rect 4988 2644 5040 2650
rect 4988 2586 5040 2592
rect 5000 870 5120 898
rect 5000 800 5028 870
rect 3712 734 3924 762
rect 4066 0 4122 800
rect 4526 0 4582 800
rect 4986 0 5042 800
rect 5092 762 5120 870
rect 5368 762 5396 9302
rect 5460 8430 5488 9551
rect 5540 9522 5592 9528
rect 5644 9518 5672 11047
rect 5736 10674 5764 13926
rect 6550 13903 6606 13912
rect 6092 13864 6144 13870
rect 6092 13806 6144 13812
rect 6104 13705 6132 13806
rect 6090 13696 6146 13705
rect 6090 13631 6146 13640
rect 6564 13394 6592 13903
rect 6552 13388 6604 13394
rect 6552 13330 6604 13336
rect 6148 13084 6456 13093
rect 6148 13082 6154 13084
rect 6210 13082 6234 13084
rect 6290 13082 6314 13084
rect 6370 13082 6394 13084
rect 6450 13082 6456 13084
rect 6210 13030 6212 13082
rect 6392 13030 6394 13082
rect 6148 13028 6154 13030
rect 6210 13028 6234 13030
rect 6290 13028 6314 13030
rect 6370 13028 6394 13030
rect 6450 13028 6456 13030
rect 6148 13019 6456 13028
rect 5816 12844 5868 12850
rect 5816 12786 5868 12792
rect 5724 10668 5776 10674
rect 5724 10610 5776 10616
rect 5632 9512 5684 9518
rect 5632 9454 5684 9460
rect 5632 9376 5684 9382
rect 5630 9344 5632 9353
rect 5684 9344 5686 9353
rect 5736 9330 5764 10610
rect 5828 10266 5856 12786
rect 6552 12776 6604 12782
rect 6552 12718 6604 12724
rect 6564 12646 6592 12718
rect 6552 12640 6604 12646
rect 6552 12582 6604 12588
rect 6564 12306 6592 12582
rect 6656 12434 6684 17614
rect 6748 13938 6776 19654
rect 6828 18148 6880 18154
rect 6828 18090 6880 18096
rect 7012 18148 7064 18154
rect 7012 18090 7064 18096
rect 6736 13932 6788 13938
rect 6736 13874 6788 13880
rect 6840 13530 6868 18090
rect 7024 17882 7052 18090
rect 7012 17876 7064 17882
rect 7012 17818 7064 17824
rect 6920 17808 6972 17814
rect 6920 17750 6972 17756
rect 6932 17134 6960 17750
rect 6920 17128 6972 17134
rect 6920 17070 6972 17076
rect 6918 16416 6974 16425
rect 6918 16351 6974 16360
rect 6932 15978 6960 16351
rect 6920 15972 6972 15978
rect 6920 15914 6972 15920
rect 6920 15564 6972 15570
rect 6920 15506 6972 15512
rect 6932 15473 6960 15506
rect 6918 15464 6974 15473
rect 6918 15399 6974 15408
rect 7012 15360 7064 15366
rect 7012 15302 7064 15308
rect 6918 14784 6974 14793
rect 6918 14719 6974 14728
rect 6828 13524 6880 13530
rect 6828 13466 6880 13472
rect 6736 13184 6788 13190
rect 6736 13126 6788 13132
rect 6748 12714 6776 13126
rect 6840 12986 6868 13466
rect 6932 13258 6960 14719
rect 6920 13252 6972 13258
rect 6920 13194 6972 13200
rect 6828 12980 6880 12986
rect 6828 12922 6880 12928
rect 6840 12753 6868 12922
rect 6826 12744 6882 12753
rect 6736 12708 6788 12714
rect 6826 12679 6882 12688
rect 6736 12650 6788 12656
rect 6828 12436 6880 12442
rect 6656 12406 6776 12434
rect 6552 12300 6604 12306
rect 6552 12242 6604 12248
rect 6644 12300 6696 12306
rect 6644 12242 6696 12248
rect 6000 12096 6052 12102
rect 6000 12038 6052 12044
rect 6552 12096 6604 12102
rect 6552 12038 6604 12044
rect 6012 11354 6040 12038
rect 6148 11996 6456 12005
rect 6148 11994 6154 11996
rect 6210 11994 6234 11996
rect 6290 11994 6314 11996
rect 6370 11994 6394 11996
rect 6450 11994 6456 11996
rect 6210 11942 6212 11994
rect 6392 11942 6394 11994
rect 6148 11940 6154 11942
rect 6210 11940 6234 11942
rect 6290 11940 6314 11942
rect 6370 11940 6394 11942
rect 6450 11940 6456 11942
rect 6148 11931 6456 11940
rect 6564 11898 6592 12038
rect 6552 11892 6604 11898
rect 6552 11834 6604 11840
rect 6656 11778 6684 12242
rect 6564 11750 6684 11778
rect 6368 11552 6420 11558
rect 6368 11494 6420 11500
rect 6000 11348 6052 11354
rect 6000 11290 6052 11296
rect 6000 11212 6052 11218
rect 6000 11154 6052 11160
rect 5908 10532 5960 10538
rect 5908 10474 5960 10480
rect 5816 10260 5868 10266
rect 5816 10202 5868 10208
rect 5814 9480 5870 9489
rect 5814 9415 5816 9424
rect 5868 9415 5870 9424
rect 5816 9386 5868 9392
rect 5736 9302 5856 9330
rect 5630 9279 5686 9288
rect 5644 8922 5672 9279
rect 5552 8894 5672 8922
rect 5724 8900 5776 8906
rect 5448 8424 5500 8430
rect 5552 8401 5580 8894
rect 5724 8842 5776 8848
rect 5736 8514 5764 8842
rect 5828 8809 5856 9302
rect 5920 9178 5948 10474
rect 6012 10130 6040 11154
rect 6380 11014 6408 11494
rect 6564 11150 6592 11750
rect 6644 11688 6696 11694
rect 6644 11630 6696 11636
rect 6656 11150 6684 11630
rect 6552 11144 6604 11150
rect 6552 11086 6604 11092
rect 6644 11144 6696 11150
rect 6644 11086 6696 11092
rect 6368 11008 6420 11014
rect 6368 10950 6420 10956
rect 6552 11008 6604 11014
rect 6552 10950 6604 10956
rect 6644 11008 6696 11014
rect 6644 10950 6696 10956
rect 6148 10908 6456 10917
rect 6148 10906 6154 10908
rect 6210 10906 6234 10908
rect 6290 10906 6314 10908
rect 6370 10906 6394 10908
rect 6450 10906 6456 10908
rect 6210 10854 6212 10906
rect 6392 10854 6394 10906
rect 6148 10852 6154 10854
rect 6210 10852 6234 10854
rect 6290 10852 6314 10854
rect 6370 10852 6394 10854
rect 6450 10852 6456 10854
rect 6148 10843 6456 10852
rect 6090 10432 6146 10441
rect 6090 10367 6146 10376
rect 6000 10124 6052 10130
rect 6000 10066 6052 10072
rect 6012 9602 6040 10066
rect 6104 9926 6132 10367
rect 6564 10266 6592 10950
rect 6656 10810 6684 10950
rect 6644 10804 6696 10810
rect 6644 10746 6696 10752
rect 6642 10568 6698 10577
rect 6642 10503 6698 10512
rect 6552 10260 6604 10266
rect 6552 10202 6604 10208
rect 6274 10160 6330 10169
rect 6656 10130 6684 10503
rect 6748 10248 6776 12406
rect 6828 12378 6880 12384
rect 6840 10606 6868 12378
rect 6918 11928 6974 11937
rect 6918 11863 6920 11872
rect 6972 11863 6974 11872
rect 6920 11834 6972 11840
rect 7024 11354 7052 15302
rect 7116 15162 7144 22200
rect 7380 19712 7432 19718
rect 7380 19654 7432 19660
rect 7392 18193 7420 19654
rect 7378 18184 7434 18193
rect 7378 18119 7434 18128
rect 7576 18057 7604 22200
rect 7748 20596 7800 20602
rect 7748 20538 7800 20544
rect 7760 20058 7788 20538
rect 7748 20052 7800 20058
rect 7748 19994 7800 20000
rect 7656 19848 7708 19854
rect 7656 19790 7708 19796
rect 7562 18048 7618 18057
rect 7562 17983 7618 17992
rect 7472 17672 7524 17678
rect 7472 17614 7524 17620
rect 7380 17604 7432 17610
rect 7380 17546 7432 17552
rect 7392 17338 7420 17546
rect 7380 17332 7432 17338
rect 7380 17274 7432 17280
rect 7196 17128 7248 17134
rect 7196 17070 7248 17076
rect 7104 15156 7156 15162
rect 7104 15098 7156 15104
rect 7208 14890 7236 17070
rect 7286 16144 7342 16153
rect 7286 16079 7342 16088
rect 7300 15042 7328 16079
rect 7484 15162 7512 17614
rect 7564 16652 7616 16658
rect 7564 16594 7616 16600
rect 7576 15162 7604 16594
rect 7472 15156 7524 15162
rect 7472 15098 7524 15104
rect 7564 15156 7616 15162
rect 7564 15098 7616 15104
rect 7300 15014 7604 15042
rect 7288 14952 7340 14958
rect 7288 14894 7340 14900
rect 7196 14884 7248 14890
rect 7196 14826 7248 14832
rect 7104 14408 7156 14414
rect 7104 14350 7156 14356
rect 7116 13530 7144 14350
rect 7300 14074 7328 14894
rect 7380 14476 7432 14482
rect 7380 14418 7432 14424
rect 7288 14068 7340 14074
rect 7288 14010 7340 14016
rect 7196 14000 7248 14006
rect 7196 13942 7248 13948
rect 7104 13524 7156 13530
rect 7104 13466 7156 13472
rect 7104 12776 7156 12782
rect 7104 12718 7156 12724
rect 7116 11898 7144 12718
rect 7208 12170 7236 13942
rect 7392 13870 7420 14418
rect 7472 14340 7524 14346
rect 7472 14282 7524 14288
rect 7380 13864 7432 13870
rect 7380 13806 7432 13812
rect 7288 13728 7340 13734
rect 7288 13670 7340 13676
rect 7300 12442 7328 13670
rect 7392 13274 7420 13806
rect 7484 13394 7512 14282
rect 7576 13734 7604 15014
rect 7668 14482 7696 19790
rect 8036 18601 8064 22200
rect 8116 20256 8168 20262
rect 8116 20198 8168 20204
rect 8128 19786 8156 20198
rect 8392 19848 8444 19854
rect 8392 19790 8444 19796
rect 8116 19780 8168 19786
rect 8116 19722 8168 19728
rect 8022 18592 8078 18601
rect 8022 18527 8078 18536
rect 8024 18284 8076 18290
rect 8024 18226 8076 18232
rect 8036 18086 8064 18226
rect 8024 18080 8076 18086
rect 8024 18022 8076 18028
rect 7746 17776 7802 17785
rect 7746 17711 7802 17720
rect 7760 17134 7788 17711
rect 7932 17536 7984 17542
rect 7932 17478 7984 17484
rect 7944 17338 7972 17478
rect 7932 17332 7984 17338
rect 7932 17274 7984 17280
rect 7748 17128 7800 17134
rect 7748 17070 7800 17076
rect 7840 16108 7892 16114
rect 7840 16050 7892 16056
rect 7852 15706 7880 16050
rect 7932 15904 7984 15910
rect 7932 15846 7984 15852
rect 7840 15700 7892 15706
rect 7840 15642 7892 15648
rect 7746 15600 7802 15609
rect 7944 15570 7972 15846
rect 7746 15535 7748 15544
rect 7800 15535 7802 15544
rect 7932 15564 7984 15570
rect 7748 15506 7800 15512
rect 7932 15506 7984 15512
rect 8036 15450 8064 18022
rect 8128 17116 8156 19722
rect 8300 19508 8352 19514
rect 8300 19450 8352 19456
rect 8312 19281 8340 19450
rect 8298 19272 8354 19281
rect 8298 19207 8354 19216
rect 8298 18728 8354 18737
rect 8298 18663 8354 18672
rect 8312 18630 8340 18663
rect 8300 18624 8352 18630
rect 8300 18566 8352 18572
rect 8208 18080 8260 18086
rect 8208 18022 8260 18028
rect 8220 17270 8248 18022
rect 8404 17338 8432 19790
rect 8496 18465 8524 22200
rect 8956 22114 8984 22200
rect 9048 22114 9076 22222
rect 8956 22086 9076 22114
rect 9218 20360 9274 20369
rect 9218 20295 9220 20304
rect 9272 20295 9274 20304
rect 9220 20266 9272 20272
rect 8747 20156 9055 20165
rect 8747 20154 8753 20156
rect 8809 20154 8833 20156
rect 8889 20154 8913 20156
rect 8969 20154 8993 20156
rect 9049 20154 9055 20156
rect 8809 20102 8811 20154
rect 8991 20102 8993 20154
rect 8747 20100 8753 20102
rect 8809 20100 8833 20102
rect 8889 20100 8913 20102
rect 8969 20100 8993 20102
rect 9049 20100 9055 20102
rect 8747 20091 9055 20100
rect 8668 19372 8720 19378
rect 8668 19314 8720 19320
rect 8576 19168 8628 19174
rect 8576 19110 8628 19116
rect 8588 18873 8616 19110
rect 8574 18864 8630 18873
rect 8574 18799 8630 18808
rect 8576 18760 8628 18766
rect 8576 18702 8628 18708
rect 8482 18456 8538 18465
rect 8482 18391 8538 18400
rect 8484 18080 8536 18086
rect 8484 18022 8536 18028
rect 8392 17332 8444 17338
rect 8392 17274 8444 17280
rect 8208 17264 8260 17270
rect 8208 17206 8260 17212
rect 8392 17196 8444 17202
rect 8392 17138 8444 17144
rect 8128 17088 8340 17116
rect 8116 16652 8168 16658
rect 8116 16594 8168 16600
rect 8128 15638 8156 16594
rect 8312 16522 8340 17088
rect 8404 16998 8432 17138
rect 8392 16992 8444 16998
rect 8392 16934 8444 16940
rect 8300 16516 8352 16522
rect 8300 16458 8352 16464
rect 8312 15910 8340 16458
rect 8300 15904 8352 15910
rect 8298 15872 8300 15881
rect 8352 15872 8354 15881
rect 8298 15807 8354 15816
rect 8116 15632 8168 15638
rect 8168 15580 8340 15586
rect 8116 15574 8340 15580
rect 8128 15558 8340 15574
rect 7944 15422 8064 15450
rect 8208 15428 8260 15434
rect 7748 14952 7800 14958
rect 7748 14894 7800 14900
rect 7760 14550 7788 14894
rect 7748 14544 7800 14550
rect 7748 14486 7800 14492
rect 7656 14476 7708 14482
rect 7656 14418 7708 14424
rect 7840 14476 7892 14482
rect 7840 14418 7892 14424
rect 7852 14278 7880 14418
rect 7748 14272 7800 14278
rect 7840 14272 7892 14278
rect 7748 14214 7800 14220
rect 7838 14240 7840 14249
rect 7892 14240 7894 14249
rect 7760 14074 7788 14214
rect 7838 14175 7894 14184
rect 7748 14068 7800 14074
rect 7748 14010 7800 14016
rect 7656 13932 7708 13938
rect 7656 13874 7708 13880
rect 7564 13728 7616 13734
rect 7564 13670 7616 13676
rect 7472 13388 7524 13394
rect 7472 13330 7524 13336
rect 7392 13246 7512 13274
rect 7288 12436 7340 12442
rect 7288 12378 7340 12384
rect 7196 12164 7248 12170
rect 7196 12106 7248 12112
rect 7288 12096 7340 12102
rect 7288 12038 7340 12044
rect 7104 11892 7156 11898
rect 7104 11834 7156 11840
rect 7116 11694 7144 11834
rect 7104 11688 7156 11694
rect 7104 11630 7156 11636
rect 7116 11354 7144 11630
rect 7012 11348 7064 11354
rect 7012 11290 7064 11296
rect 7104 11348 7156 11354
rect 7104 11290 7156 11296
rect 6918 10704 6974 10713
rect 6918 10639 6920 10648
rect 6972 10639 6974 10648
rect 7196 10668 7248 10674
rect 6920 10610 6972 10616
rect 7196 10610 7248 10616
rect 6828 10600 6880 10606
rect 6828 10542 6880 10548
rect 7208 10470 7236 10610
rect 7196 10464 7248 10470
rect 7196 10406 7248 10412
rect 7104 10260 7156 10266
rect 6748 10220 6960 10248
rect 6826 10160 6882 10169
rect 6274 10095 6330 10104
rect 6644 10124 6696 10130
rect 6288 9994 6316 10095
rect 6644 10066 6696 10072
rect 6736 10124 6788 10130
rect 6826 10095 6882 10104
rect 6736 10066 6788 10072
rect 6276 9988 6328 9994
rect 6276 9930 6328 9936
rect 6092 9920 6144 9926
rect 6092 9862 6144 9868
rect 6148 9820 6456 9829
rect 6148 9818 6154 9820
rect 6210 9818 6234 9820
rect 6290 9818 6314 9820
rect 6370 9818 6394 9820
rect 6450 9818 6456 9820
rect 6210 9766 6212 9818
rect 6392 9766 6394 9818
rect 6148 9764 6154 9766
rect 6210 9764 6234 9766
rect 6290 9764 6314 9766
rect 6370 9764 6394 9766
rect 6450 9764 6456 9766
rect 6148 9755 6456 9764
rect 6550 9752 6606 9761
rect 6550 9687 6606 9696
rect 6184 9648 6236 9654
rect 6012 9586 6132 9602
rect 6184 9590 6236 9596
rect 6368 9648 6420 9654
rect 6368 9590 6420 9596
rect 6012 9580 6144 9586
rect 6012 9574 6092 9580
rect 6092 9522 6144 9528
rect 5908 9172 5960 9178
rect 5908 9114 5960 9120
rect 6090 9072 6146 9081
rect 6090 9007 6092 9016
rect 6144 9007 6146 9016
rect 6092 8978 6144 8984
rect 6196 8838 6224 9590
rect 6276 9580 6328 9586
rect 6276 9522 6328 9528
rect 6288 9353 6316 9522
rect 6380 9450 6408 9590
rect 6368 9444 6420 9450
rect 6368 9386 6420 9392
rect 6274 9344 6330 9353
rect 6274 9279 6330 9288
rect 6564 9178 6592 9687
rect 6748 9450 6776 10066
rect 6840 9625 6868 10095
rect 6826 9616 6882 9625
rect 6826 9551 6882 9560
rect 6736 9444 6788 9450
rect 6736 9386 6788 9392
rect 6552 9172 6604 9178
rect 6552 9114 6604 9120
rect 6826 9072 6882 9081
rect 6826 9007 6828 9016
rect 6880 9007 6882 9016
rect 6828 8978 6880 8984
rect 6184 8832 6236 8838
rect 5814 8800 5870 8809
rect 6184 8774 6236 8780
rect 6552 8832 6604 8838
rect 6552 8774 6604 8780
rect 6644 8832 6696 8838
rect 6932 8786 6960 10220
rect 7104 10202 7156 10208
rect 7012 9920 7064 9926
rect 7012 9862 7064 9868
rect 7024 9382 7052 9862
rect 7116 9761 7144 10202
rect 7102 9752 7158 9761
rect 7102 9687 7158 9696
rect 7012 9376 7064 9382
rect 7012 9318 7064 9324
rect 6644 8774 6696 8780
rect 5814 8735 5870 8744
rect 5644 8486 5764 8514
rect 5448 8366 5500 8372
rect 5538 8392 5594 8401
rect 5460 7342 5488 8366
rect 5538 8327 5594 8336
rect 5448 7336 5500 7342
rect 5448 7278 5500 7284
rect 5448 7200 5500 7206
rect 5448 7142 5500 7148
rect 5460 5817 5488 7142
rect 5552 5914 5580 8327
rect 5644 8090 5672 8486
rect 5724 8424 5776 8430
rect 5724 8366 5776 8372
rect 5736 8090 5764 8366
rect 5828 8294 5856 8735
rect 6148 8732 6456 8741
rect 6148 8730 6154 8732
rect 6210 8730 6234 8732
rect 6290 8730 6314 8732
rect 6370 8730 6394 8732
rect 6450 8730 6456 8732
rect 6210 8678 6212 8730
rect 6392 8678 6394 8730
rect 6148 8676 6154 8678
rect 6210 8676 6234 8678
rect 6290 8676 6314 8678
rect 6370 8676 6394 8678
rect 6450 8676 6456 8678
rect 6148 8667 6456 8676
rect 6564 8634 6592 8774
rect 6552 8628 6604 8634
rect 6552 8570 6604 8576
rect 6000 8492 6052 8498
rect 6000 8434 6052 8440
rect 5816 8288 5868 8294
rect 5816 8230 5868 8236
rect 5632 8084 5684 8090
rect 5632 8026 5684 8032
rect 5724 8084 5776 8090
rect 5724 8026 5776 8032
rect 5816 7404 5868 7410
rect 5816 7346 5868 7352
rect 5828 7002 5856 7346
rect 5908 7336 5960 7342
rect 5908 7278 5960 7284
rect 5816 6996 5868 7002
rect 5816 6938 5868 6944
rect 5632 6928 5684 6934
rect 5632 6870 5684 6876
rect 5644 6474 5672 6870
rect 5724 6792 5776 6798
rect 5724 6734 5776 6740
rect 5814 6760 5870 6769
rect 5736 6662 5764 6734
rect 5814 6695 5870 6704
rect 5828 6662 5856 6695
rect 5724 6656 5776 6662
rect 5722 6624 5724 6633
rect 5816 6656 5868 6662
rect 5776 6624 5778 6633
rect 5816 6598 5868 6604
rect 5722 6559 5778 6568
rect 5644 6446 5764 6474
rect 5632 6316 5684 6322
rect 5632 6258 5684 6264
rect 5540 5908 5592 5914
rect 5540 5850 5592 5856
rect 5446 5808 5502 5817
rect 5446 5743 5502 5752
rect 5448 5704 5500 5710
rect 5448 5646 5500 5652
rect 5460 5574 5488 5646
rect 5448 5568 5500 5574
rect 5446 5536 5448 5545
rect 5500 5536 5502 5545
rect 5446 5471 5502 5480
rect 5644 5409 5672 6258
rect 5630 5400 5686 5409
rect 5630 5335 5686 5344
rect 5632 5024 5684 5030
rect 5632 4966 5684 4972
rect 5644 4554 5672 4966
rect 5736 4706 5764 6446
rect 5816 5908 5868 5914
rect 5816 5850 5868 5856
rect 5828 5574 5856 5850
rect 5816 5568 5868 5574
rect 5816 5510 5868 5516
rect 5816 5228 5868 5234
rect 5816 5170 5868 5176
rect 5828 4826 5856 5170
rect 5920 4826 5948 7278
rect 6012 7274 6040 8434
rect 6368 7880 6420 7886
rect 6366 7848 6368 7857
rect 6420 7848 6422 7857
rect 6366 7783 6422 7792
rect 6148 7644 6456 7653
rect 6148 7642 6154 7644
rect 6210 7642 6234 7644
rect 6290 7642 6314 7644
rect 6370 7642 6394 7644
rect 6450 7642 6456 7644
rect 6210 7590 6212 7642
rect 6392 7590 6394 7642
rect 6148 7588 6154 7590
rect 6210 7588 6234 7590
rect 6290 7588 6314 7590
rect 6370 7588 6394 7590
rect 6450 7588 6456 7590
rect 6148 7579 6456 7588
rect 6656 7546 6684 8774
rect 6748 8758 6960 8786
rect 6644 7540 6696 7546
rect 6644 7482 6696 7488
rect 6092 7336 6144 7342
rect 6092 7278 6144 7284
rect 6000 7268 6052 7274
rect 6000 7210 6052 7216
rect 6000 6656 6052 6662
rect 6104 6644 6132 7278
rect 6366 6896 6422 6905
rect 6366 6831 6422 6840
rect 6380 6662 6408 6831
rect 6052 6616 6132 6644
rect 6368 6656 6420 6662
rect 6000 6598 6052 6604
rect 6368 6598 6420 6604
rect 6012 6322 6040 6598
rect 6148 6556 6456 6565
rect 6148 6554 6154 6556
rect 6210 6554 6234 6556
rect 6290 6554 6314 6556
rect 6370 6554 6394 6556
rect 6450 6554 6456 6556
rect 6210 6502 6212 6554
rect 6392 6502 6394 6554
rect 6148 6500 6154 6502
rect 6210 6500 6234 6502
rect 6290 6500 6314 6502
rect 6370 6500 6394 6502
rect 6450 6500 6456 6502
rect 6148 6491 6456 6500
rect 6000 6316 6052 6322
rect 6000 6258 6052 6264
rect 6276 6112 6328 6118
rect 6276 6054 6328 6060
rect 6550 6080 6606 6089
rect 6288 5642 6316 6054
rect 6748 6066 6776 8758
rect 6828 8628 6880 8634
rect 6828 8570 6880 8576
rect 6840 8294 6868 8570
rect 6920 8492 6972 8498
rect 6920 8434 6972 8440
rect 6828 8288 6880 8294
rect 6828 8230 6880 8236
rect 6840 7750 6868 8230
rect 6932 7886 6960 8434
rect 6920 7880 6972 7886
rect 6920 7822 6972 7828
rect 6828 7744 6880 7750
rect 6828 7686 6880 7692
rect 6840 6934 6868 7686
rect 6932 7449 6960 7822
rect 6918 7440 6974 7449
rect 6918 7375 6974 7384
rect 6918 7304 6974 7313
rect 6918 7239 6974 7248
rect 6828 6928 6880 6934
rect 6828 6870 6880 6876
rect 6826 6760 6882 6769
rect 6826 6695 6882 6704
rect 6840 6662 6868 6695
rect 6828 6656 6880 6662
rect 6828 6598 6880 6604
rect 6932 6322 6960 7239
rect 6920 6316 6972 6322
rect 6920 6258 6972 6264
rect 6550 6015 6606 6024
rect 6656 6038 6776 6066
rect 6564 5778 6592 6015
rect 6552 5772 6604 5778
rect 6552 5714 6604 5720
rect 6656 5658 6684 6038
rect 6734 5944 6790 5953
rect 6734 5879 6790 5888
rect 6276 5636 6328 5642
rect 6276 5578 6328 5584
rect 6564 5630 6684 5658
rect 6148 5468 6456 5477
rect 6148 5466 6154 5468
rect 6210 5466 6234 5468
rect 6290 5466 6314 5468
rect 6370 5466 6394 5468
rect 6450 5466 6456 5468
rect 6210 5414 6212 5466
rect 6392 5414 6394 5466
rect 6148 5412 6154 5414
rect 6210 5412 6234 5414
rect 6290 5412 6314 5414
rect 6370 5412 6394 5414
rect 6450 5412 6456 5414
rect 6148 5403 6456 5412
rect 6000 5160 6052 5166
rect 6000 5102 6052 5108
rect 5816 4820 5868 4826
rect 5816 4762 5868 4768
rect 5908 4820 5960 4826
rect 5908 4762 5960 4768
rect 5736 4678 5856 4706
rect 5632 4548 5684 4554
rect 5632 4490 5684 4496
rect 5540 4072 5592 4078
rect 5540 4014 5592 4020
rect 5448 3936 5500 3942
rect 5448 3878 5500 3884
rect 5460 3602 5488 3878
rect 5448 3596 5500 3602
rect 5448 3538 5500 3544
rect 5448 3460 5500 3466
rect 5448 3402 5500 3408
rect 5460 3194 5488 3402
rect 5448 3188 5500 3194
rect 5448 3130 5500 3136
rect 5448 3052 5500 3058
rect 5448 2994 5500 3000
rect 5460 800 5488 2994
rect 5552 2990 5580 4014
rect 5644 3602 5672 4490
rect 5724 4072 5776 4078
rect 5722 4040 5724 4049
rect 5776 4040 5778 4049
rect 5828 4010 5856 4678
rect 6012 4622 6040 5102
rect 6564 4690 6592 5630
rect 6644 5568 6696 5574
rect 6644 5510 6696 5516
rect 6656 5370 6684 5510
rect 6644 5364 6696 5370
rect 6644 5306 6696 5312
rect 6748 5250 6776 5879
rect 6932 5574 6960 6258
rect 7024 5914 7052 9318
rect 7208 7993 7236 10406
rect 7300 8906 7328 12038
rect 7484 11694 7512 13246
rect 7564 13184 7616 13190
rect 7564 13126 7616 13132
rect 7472 11688 7524 11694
rect 7472 11630 7524 11636
rect 7576 10266 7604 13126
rect 7668 12442 7696 13874
rect 7748 13456 7800 13462
rect 7748 13398 7800 13404
rect 7760 12782 7788 13398
rect 7748 12776 7800 12782
rect 7746 12744 7748 12753
rect 7840 12776 7892 12782
rect 7800 12744 7802 12753
rect 7840 12718 7892 12724
rect 7746 12679 7802 12688
rect 7656 12436 7708 12442
rect 7656 12378 7708 12384
rect 7748 12436 7800 12442
rect 7748 12378 7800 12384
rect 7656 12164 7708 12170
rect 7656 12106 7708 12112
rect 7564 10260 7616 10266
rect 7564 10202 7616 10208
rect 7562 9480 7618 9489
rect 7562 9415 7618 9424
rect 7470 9208 7526 9217
rect 7470 9143 7526 9152
rect 7484 8974 7512 9143
rect 7472 8968 7524 8974
rect 7472 8910 7524 8916
rect 7288 8900 7340 8906
rect 7288 8842 7340 8848
rect 7472 8832 7524 8838
rect 7472 8774 7524 8780
rect 7288 8492 7340 8498
rect 7288 8434 7340 8440
rect 7194 7984 7250 7993
rect 7104 7948 7156 7954
rect 7194 7919 7250 7928
rect 7104 7890 7156 7896
rect 7116 7750 7144 7890
rect 7104 7744 7156 7750
rect 7104 7686 7156 7692
rect 7116 7342 7144 7686
rect 7104 7336 7156 7342
rect 7104 7278 7156 7284
rect 7116 7002 7144 7278
rect 7208 7206 7236 7919
rect 7300 7546 7328 8434
rect 7380 8424 7432 8430
rect 7380 8366 7432 8372
rect 7288 7540 7340 7546
rect 7288 7482 7340 7488
rect 7196 7200 7248 7206
rect 7196 7142 7248 7148
rect 7104 6996 7156 7002
rect 7104 6938 7156 6944
rect 7116 6322 7144 6938
rect 7194 6760 7250 6769
rect 7194 6695 7250 6704
rect 7208 6662 7236 6695
rect 7196 6656 7248 6662
rect 7196 6598 7248 6604
rect 7104 6316 7156 6322
rect 7104 6258 7156 6264
rect 7012 5908 7064 5914
rect 7012 5850 7064 5856
rect 6920 5568 6972 5574
rect 6826 5536 6882 5545
rect 6920 5510 6972 5516
rect 6826 5471 6882 5480
rect 6656 5222 6776 5250
rect 6552 4684 6604 4690
rect 6552 4626 6604 4632
rect 6000 4616 6052 4622
rect 6000 4558 6052 4564
rect 6000 4480 6052 4486
rect 6000 4422 6052 4428
rect 6012 4146 6040 4422
rect 6148 4380 6456 4389
rect 6148 4378 6154 4380
rect 6210 4378 6234 4380
rect 6290 4378 6314 4380
rect 6370 4378 6394 4380
rect 6450 4378 6456 4380
rect 6210 4326 6212 4378
rect 6392 4326 6394 4378
rect 6148 4324 6154 4326
rect 6210 4324 6234 4326
rect 6290 4324 6314 4326
rect 6370 4324 6394 4326
rect 6450 4324 6456 4326
rect 6148 4315 6456 4324
rect 6552 4208 6604 4214
rect 6552 4150 6604 4156
rect 6000 4140 6052 4146
rect 6000 4082 6052 4088
rect 5722 3975 5778 3984
rect 5816 4004 5868 4010
rect 5816 3946 5868 3952
rect 6184 3936 6236 3942
rect 6184 3878 6236 3884
rect 6460 3936 6512 3942
rect 6460 3878 6512 3884
rect 5632 3596 5684 3602
rect 5632 3538 5684 3544
rect 5908 3596 5960 3602
rect 5908 3538 5960 3544
rect 5816 3528 5868 3534
rect 5816 3470 5868 3476
rect 5540 2984 5592 2990
rect 5540 2926 5592 2932
rect 5828 2650 5856 3470
rect 5920 3398 5948 3538
rect 6196 3534 6224 3878
rect 6472 3670 6500 3878
rect 6564 3738 6592 4150
rect 6552 3732 6604 3738
rect 6552 3674 6604 3680
rect 6460 3664 6512 3670
rect 6366 3632 6422 3641
rect 6460 3606 6512 3612
rect 6564 3602 6592 3674
rect 6366 3567 6368 3576
rect 6420 3567 6422 3576
rect 6552 3596 6604 3602
rect 6368 3538 6420 3544
rect 6552 3538 6604 3544
rect 6184 3528 6236 3534
rect 6184 3470 6236 3476
rect 5908 3392 5960 3398
rect 5908 3334 5960 3340
rect 6148 3292 6456 3301
rect 6148 3290 6154 3292
rect 6210 3290 6234 3292
rect 6290 3290 6314 3292
rect 6370 3290 6394 3292
rect 6450 3290 6456 3292
rect 6210 3238 6212 3290
rect 6392 3238 6394 3290
rect 6148 3236 6154 3238
rect 6210 3236 6234 3238
rect 6290 3236 6314 3238
rect 6370 3236 6394 3238
rect 6450 3236 6456 3238
rect 5906 3224 5962 3233
rect 6148 3227 6456 3236
rect 5906 3159 5962 3168
rect 5816 2644 5868 2650
rect 5816 2586 5868 2592
rect 5828 2514 5856 2586
rect 5816 2508 5868 2514
rect 5816 2450 5868 2456
rect 5920 800 5948 3159
rect 6550 3088 6606 3097
rect 6550 3023 6606 3032
rect 6564 2990 6592 3023
rect 6552 2984 6604 2990
rect 6552 2926 6604 2932
rect 6148 2204 6456 2213
rect 6148 2202 6154 2204
rect 6210 2202 6234 2204
rect 6290 2202 6314 2204
rect 6370 2202 6394 2204
rect 6450 2202 6456 2204
rect 6210 2150 6212 2202
rect 6392 2150 6394 2202
rect 6148 2148 6154 2150
rect 6210 2148 6234 2150
rect 6290 2148 6314 2150
rect 6370 2148 6394 2150
rect 6450 2148 6456 2150
rect 6148 2139 6456 2148
rect 6380 870 6500 898
rect 6380 800 6408 870
rect 5092 734 5396 762
rect 5446 0 5502 800
rect 5906 0 5962 800
rect 6366 0 6422 800
rect 6472 762 6500 870
rect 6656 762 6684 5222
rect 6736 4684 6788 4690
rect 6736 4626 6788 4632
rect 6748 4486 6776 4626
rect 6736 4480 6788 4486
rect 6736 4422 6788 4428
rect 6736 3664 6788 3670
rect 6734 3632 6736 3641
rect 6788 3632 6790 3641
rect 6734 3567 6790 3576
rect 6736 3392 6788 3398
rect 6736 3334 6788 3340
rect 6748 3194 6776 3334
rect 6736 3188 6788 3194
rect 6736 3130 6788 3136
rect 6840 800 6868 5471
rect 6932 3233 6960 5510
rect 7116 4826 7144 6258
rect 7104 4820 7156 4826
rect 7104 4762 7156 4768
rect 7116 4690 7144 4762
rect 7104 4684 7156 4690
rect 7104 4626 7156 4632
rect 7208 4570 7236 6598
rect 7392 6458 7420 8366
rect 7484 8090 7512 8774
rect 7576 8430 7604 9415
rect 7668 9042 7696 12106
rect 7760 11558 7788 12378
rect 7748 11552 7800 11558
rect 7748 11494 7800 11500
rect 7746 11112 7802 11121
rect 7746 11047 7802 11056
rect 7760 9926 7788 11047
rect 7748 9920 7800 9926
rect 7748 9862 7800 9868
rect 7760 9382 7788 9862
rect 7852 9450 7880 12718
rect 7944 11830 7972 15422
rect 8208 15370 8260 15376
rect 8220 15162 8248 15370
rect 8208 15156 8260 15162
rect 8128 15116 8208 15144
rect 8022 15056 8078 15065
rect 8022 14991 8078 15000
rect 8036 14278 8064 14991
rect 8024 14272 8076 14278
rect 8024 14214 8076 14220
rect 8036 12306 8064 14214
rect 8024 12300 8076 12306
rect 8024 12242 8076 12248
rect 7932 11824 7984 11830
rect 7932 11766 7984 11772
rect 8024 11756 8076 11762
rect 8024 11698 8076 11704
rect 7932 11688 7984 11694
rect 7932 11630 7984 11636
rect 7944 10810 7972 11630
rect 7932 10804 7984 10810
rect 7932 10746 7984 10752
rect 8036 10266 8064 11698
rect 8024 10260 8076 10266
rect 8024 10202 8076 10208
rect 8128 10130 8156 15116
rect 8208 15098 8260 15104
rect 8206 15056 8262 15065
rect 8206 14991 8262 15000
rect 8220 14890 8248 14991
rect 8208 14884 8260 14890
rect 8208 14826 8260 14832
rect 8312 14482 8340 15558
rect 8404 15450 8432 16934
rect 8496 15638 8524 18022
rect 8484 15632 8536 15638
rect 8484 15574 8536 15580
rect 8404 15422 8524 15450
rect 8392 15088 8444 15094
rect 8392 15030 8444 15036
rect 8404 14550 8432 15030
rect 8392 14544 8444 14550
rect 8392 14486 8444 14492
rect 8208 14476 8260 14482
rect 8208 14418 8260 14424
rect 8300 14476 8352 14482
rect 8300 14418 8352 14424
rect 8220 14278 8248 14418
rect 8208 14272 8260 14278
rect 8208 14214 8260 14220
rect 8208 13320 8260 13326
rect 8208 13262 8260 13268
rect 8220 12986 8248 13262
rect 8392 13184 8444 13190
rect 8392 13126 8444 13132
rect 8404 12986 8432 13126
rect 8208 12980 8260 12986
rect 8208 12922 8260 12928
rect 8392 12980 8444 12986
rect 8392 12922 8444 12928
rect 8392 12844 8444 12850
rect 8392 12786 8444 12792
rect 8300 12776 8352 12782
rect 8300 12718 8352 12724
rect 8312 12442 8340 12718
rect 8300 12436 8352 12442
rect 8300 12378 8352 12384
rect 8404 12356 8432 12786
rect 8496 12434 8524 15422
rect 8588 13274 8616 18702
rect 8680 16590 8708 19314
rect 9128 19304 9180 19310
rect 9128 19246 9180 19252
rect 9140 19145 9168 19246
rect 9126 19136 9182 19145
rect 8747 19068 9055 19077
rect 9126 19071 9182 19080
rect 8747 19066 8753 19068
rect 8809 19066 8833 19068
rect 8889 19066 8913 19068
rect 8969 19066 8993 19068
rect 9049 19066 9055 19068
rect 8809 19014 8811 19066
rect 8991 19014 8993 19066
rect 8747 19012 8753 19014
rect 8809 19012 8833 19014
rect 8889 19012 8913 19014
rect 8969 19012 8993 19014
rect 9049 19012 9055 19014
rect 8747 19003 9055 19012
rect 8944 18964 8996 18970
rect 8944 18906 8996 18912
rect 8850 18320 8906 18329
rect 8850 18255 8906 18264
rect 8864 18222 8892 18255
rect 8852 18216 8904 18222
rect 8852 18158 8904 18164
rect 8956 18154 8984 18906
rect 9128 18760 9180 18766
rect 9128 18702 9180 18708
rect 9220 18760 9272 18766
rect 9220 18702 9272 18708
rect 9036 18420 9088 18426
rect 9036 18362 9088 18368
rect 9048 18290 9076 18362
rect 9036 18284 9088 18290
rect 9036 18226 9088 18232
rect 8944 18148 8996 18154
rect 8944 18090 8996 18096
rect 8747 17980 9055 17989
rect 8747 17978 8753 17980
rect 8809 17978 8833 17980
rect 8889 17978 8913 17980
rect 8969 17978 8993 17980
rect 9049 17978 9055 17980
rect 8809 17926 8811 17978
rect 8991 17926 8993 17978
rect 8747 17924 8753 17926
rect 8809 17924 8833 17926
rect 8889 17924 8913 17926
rect 8969 17924 8993 17926
rect 9049 17924 9055 17926
rect 8747 17915 9055 17924
rect 9140 17678 9168 18702
rect 9232 17882 9260 18702
rect 9220 17876 9272 17882
rect 9220 17818 9272 17824
rect 9128 17672 9180 17678
rect 9128 17614 9180 17620
rect 9220 17604 9272 17610
rect 9220 17546 9272 17552
rect 9128 17536 9180 17542
rect 9128 17478 9180 17484
rect 9140 17338 9168 17478
rect 9128 17332 9180 17338
rect 9128 17274 9180 17280
rect 9128 16992 9180 16998
rect 9128 16934 9180 16940
rect 8747 16892 9055 16901
rect 8747 16890 8753 16892
rect 8809 16890 8833 16892
rect 8889 16890 8913 16892
rect 8969 16890 8993 16892
rect 9049 16890 9055 16892
rect 8809 16838 8811 16890
rect 8991 16838 8993 16890
rect 8747 16836 8753 16838
rect 8809 16836 8833 16838
rect 8889 16836 8913 16838
rect 8969 16836 8993 16838
rect 9049 16836 9055 16838
rect 8747 16827 9055 16836
rect 9140 16726 9168 16934
rect 9128 16720 9180 16726
rect 9128 16662 9180 16668
rect 8668 16584 8720 16590
rect 9232 16538 9260 17546
rect 9324 17270 9352 22222
rect 9402 22200 9458 23000
rect 9862 22200 9918 23000
rect 10322 22200 10378 23000
rect 10782 22200 10838 23000
rect 11242 22200 11298 23000
rect 11348 22222 11652 22250
rect 9416 19938 9444 22200
rect 9680 20392 9732 20398
rect 9680 20334 9732 20340
rect 9692 20058 9720 20334
rect 9680 20052 9732 20058
rect 9680 19994 9732 20000
rect 9416 19910 9628 19938
rect 9404 19848 9456 19854
rect 9404 19790 9456 19796
rect 9416 18834 9444 19790
rect 9496 19168 9548 19174
rect 9496 19110 9548 19116
rect 9404 18828 9456 18834
rect 9404 18770 9456 18776
rect 9402 18456 9458 18465
rect 9402 18391 9458 18400
rect 9416 18222 9444 18391
rect 9404 18216 9456 18222
rect 9404 18158 9456 18164
rect 9312 17264 9364 17270
rect 9312 17206 9364 17212
rect 9508 17082 9536 19110
rect 9600 18986 9628 19910
rect 9772 19848 9824 19854
rect 9772 19790 9824 19796
rect 9678 19000 9734 19009
rect 9600 18958 9678 18986
rect 9678 18935 9734 18944
rect 9784 18834 9812 19790
rect 9876 18902 9904 22200
rect 9956 19848 10008 19854
rect 9956 19790 10008 19796
rect 10048 19848 10100 19854
rect 10048 19790 10100 19796
rect 9968 19689 9996 19790
rect 9954 19680 10010 19689
rect 9954 19615 10010 19624
rect 10060 19378 10088 19790
rect 10140 19712 10192 19718
rect 10140 19654 10192 19660
rect 10048 19372 10100 19378
rect 10048 19314 10100 19320
rect 10060 19145 10088 19314
rect 10152 19242 10180 19654
rect 10140 19236 10192 19242
rect 10140 19178 10192 19184
rect 10046 19136 10102 19145
rect 10046 19071 10102 19080
rect 9956 18964 10008 18970
rect 9956 18906 10008 18912
rect 9864 18896 9916 18902
rect 9864 18838 9916 18844
rect 9772 18828 9824 18834
rect 9772 18770 9824 18776
rect 9634 18284 9686 18290
rect 9686 18244 9812 18272
rect 9634 18226 9686 18232
rect 9784 18136 9812 18244
rect 9968 18154 9996 18906
rect 10048 18896 10100 18902
rect 10048 18838 10100 18844
rect 9692 18108 9812 18136
rect 9956 18148 10008 18154
rect 9586 18048 9642 18057
rect 9586 17983 9642 17992
rect 8668 16526 8720 16532
rect 9140 16522 9260 16538
rect 9324 17054 9536 17082
rect 9324 16522 9352 17054
rect 9496 16584 9548 16590
rect 9496 16526 9548 16532
rect 9128 16516 9260 16522
rect 9180 16510 9260 16516
rect 9312 16516 9364 16522
rect 9128 16458 9180 16464
rect 9312 16458 9364 16464
rect 9140 15978 9168 16458
rect 9324 16402 9352 16458
rect 9232 16374 9352 16402
rect 9404 16448 9456 16454
rect 9404 16390 9456 16396
rect 8668 15972 8720 15978
rect 8668 15914 8720 15920
rect 9128 15972 9180 15978
rect 9128 15914 9180 15920
rect 8680 15162 8708 15914
rect 8747 15804 9055 15813
rect 8747 15802 8753 15804
rect 8809 15802 8833 15804
rect 8889 15802 8913 15804
rect 8969 15802 8993 15804
rect 9049 15802 9055 15804
rect 8809 15750 8811 15802
rect 8991 15750 8993 15802
rect 8747 15748 8753 15750
rect 8809 15748 8833 15750
rect 8889 15748 8913 15750
rect 8969 15748 8993 15750
rect 9049 15748 9055 15750
rect 8747 15739 9055 15748
rect 9140 15706 9168 15914
rect 9232 15910 9260 16374
rect 9312 16244 9364 16250
rect 9312 16186 9364 16192
rect 9324 15910 9352 16186
rect 9220 15904 9272 15910
rect 9220 15846 9272 15852
rect 9312 15904 9364 15910
rect 9312 15846 9364 15852
rect 9128 15700 9180 15706
rect 9128 15642 9180 15648
rect 8760 15428 8812 15434
rect 8760 15370 8812 15376
rect 8668 15156 8720 15162
rect 8668 15098 8720 15104
rect 8772 15042 8800 15370
rect 9140 15162 9168 15642
rect 9128 15156 9180 15162
rect 9128 15098 9180 15104
rect 8680 15014 8800 15042
rect 8680 14958 8708 15014
rect 8668 14952 8720 14958
rect 8668 14894 8720 14900
rect 9128 14952 9180 14958
rect 9128 14894 9180 14900
rect 8680 14006 8708 14894
rect 8747 14716 9055 14725
rect 8747 14714 8753 14716
rect 8809 14714 8833 14716
rect 8889 14714 8913 14716
rect 8969 14714 8993 14716
rect 9049 14714 9055 14716
rect 8809 14662 8811 14714
rect 8991 14662 8993 14714
rect 8747 14660 8753 14662
rect 8809 14660 8833 14662
rect 8889 14660 8913 14662
rect 8969 14660 8993 14662
rect 9049 14660 9055 14662
rect 8747 14651 9055 14660
rect 9140 14618 9168 14894
rect 9128 14612 9180 14618
rect 9128 14554 9180 14560
rect 9126 14512 9182 14521
rect 9126 14447 9128 14456
rect 9180 14447 9182 14456
rect 9128 14418 9180 14424
rect 9128 14272 9180 14278
rect 9128 14214 9180 14220
rect 8668 14000 8720 14006
rect 8668 13942 8720 13948
rect 8747 13628 9055 13637
rect 8747 13626 8753 13628
rect 8809 13626 8833 13628
rect 8889 13626 8913 13628
rect 8969 13626 8993 13628
rect 9049 13626 9055 13628
rect 8809 13574 8811 13626
rect 8991 13574 8993 13626
rect 8747 13572 8753 13574
rect 8809 13572 8833 13574
rect 8889 13572 8913 13574
rect 8969 13572 8993 13574
rect 9049 13572 9055 13574
rect 8747 13563 9055 13572
rect 8666 13424 8722 13433
rect 8666 13359 8668 13368
rect 8720 13359 8722 13368
rect 8668 13330 8720 13336
rect 8588 13246 8708 13274
rect 8496 12406 8616 12434
rect 8404 12328 8524 12356
rect 8300 12096 8352 12102
rect 8300 12038 8352 12044
rect 8208 11824 8260 11830
rect 8208 11766 8260 11772
rect 8116 10124 8168 10130
rect 7944 10084 8116 10112
rect 7840 9444 7892 9450
rect 7840 9386 7892 9392
rect 7748 9376 7800 9382
rect 7748 9318 7800 9324
rect 7840 9104 7892 9110
rect 7840 9046 7892 9052
rect 7656 9036 7708 9042
rect 7656 8978 7708 8984
rect 7852 8566 7880 9046
rect 7944 8634 7972 10084
rect 8116 10066 8168 10072
rect 8024 9988 8076 9994
rect 8024 9930 8076 9936
rect 8036 9178 8064 9930
rect 8220 9926 8248 11766
rect 8312 11558 8340 12038
rect 8300 11552 8352 11558
rect 8300 11494 8352 11500
rect 8300 11144 8352 11150
rect 8300 11086 8352 11092
rect 8208 9920 8260 9926
rect 8312 9908 8340 11086
rect 8496 10810 8524 12328
rect 8588 11150 8616 12406
rect 8576 11144 8628 11150
rect 8576 11086 8628 11092
rect 8576 11008 8628 11014
rect 8576 10950 8628 10956
rect 8588 10810 8616 10950
rect 8484 10804 8536 10810
rect 8484 10746 8536 10752
rect 8576 10804 8628 10810
rect 8576 10746 8628 10752
rect 8680 10690 8708 13246
rect 8747 12540 9055 12549
rect 8747 12538 8753 12540
rect 8809 12538 8833 12540
rect 8889 12538 8913 12540
rect 8969 12538 8993 12540
rect 9049 12538 9055 12540
rect 8809 12486 8811 12538
rect 8991 12486 8993 12538
rect 8747 12484 8753 12486
rect 8809 12484 8833 12486
rect 8889 12484 8913 12486
rect 8969 12484 8993 12486
rect 9049 12484 9055 12486
rect 8747 12475 9055 12484
rect 9140 12434 9168 14214
rect 9048 12406 9168 12434
rect 9048 11558 9076 12406
rect 9128 12096 9180 12102
rect 9128 12038 9180 12044
rect 9036 11552 9088 11558
rect 9036 11494 9088 11500
rect 8747 11452 9055 11461
rect 8747 11450 8753 11452
rect 8809 11450 8833 11452
rect 8889 11450 8913 11452
rect 8969 11450 8993 11452
rect 9049 11450 9055 11452
rect 8809 11398 8811 11450
rect 8991 11398 8993 11450
rect 8747 11396 8753 11398
rect 8809 11396 8833 11398
rect 8889 11396 8913 11398
rect 8969 11396 8993 11398
rect 9049 11396 9055 11398
rect 8747 11387 9055 11396
rect 9140 10996 9168 12038
rect 9048 10968 9168 10996
rect 9048 10810 9076 10968
rect 9036 10804 9088 10810
rect 9036 10746 9088 10752
rect 8496 10662 8708 10690
rect 8392 10600 8444 10606
rect 8496 10554 8524 10662
rect 8444 10548 8524 10554
rect 8392 10542 8524 10548
rect 8576 10600 8628 10606
rect 8576 10542 8628 10548
rect 8404 10526 8524 10542
rect 8404 10062 8432 10526
rect 8588 10130 8616 10542
rect 9128 10532 9180 10538
rect 9128 10474 9180 10480
rect 8747 10364 9055 10373
rect 8747 10362 8753 10364
rect 8809 10362 8833 10364
rect 8889 10362 8913 10364
rect 8969 10362 8993 10364
rect 9049 10362 9055 10364
rect 8809 10310 8811 10362
rect 8991 10310 8993 10362
rect 8747 10308 8753 10310
rect 8809 10308 8833 10310
rect 8889 10308 8913 10310
rect 8969 10308 8993 10310
rect 9049 10308 9055 10310
rect 8747 10299 9055 10308
rect 8576 10124 8628 10130
rect 8576 10066 8628 10072
rect 8392 10056 8444 10062
rect 8392 9998 8444 10004
rect 8312 9880 8524 9908
rect 8208 9862 8260 9868
rect 8024 9172 8076 9178
rect 8024 9114 8076 9120
rect 7932 8628 7984 8634
rect 7932 8570 7984 8576
rect 7656 8560 7708 8566
rect 7656 8502 7708 8508
rect 7840 8560 7892 8566
rect 7840 8502 7892 8508
rect 7564 8424 7616 8430
rect 7564 8366 7616 8372
rect 7472 8084 7524 8090
rect 7472 8026 7524 8032
rect 7564 7744 7616 7750
rect 7668 7732 7696 8502
rect 7748 8288 7800 8294
rect 7748 8230 7800 8236
rect 7616 7704 7696 7732
rect 7564 7686 7616 7692
rect 7576 7274 7604 7686
rect 7564 7268 7616 7274
rect 7564 7210 7616 7216
rect 7654 6896 7710 6905
rect 7760 6866 7788 8230
rect 7840 7812 7892 7818
rect 7840 7754 7892 7760
rect 7654 6831 7710 6840
rect 7748 6860 7800 6866
rect 7668 6662 7696 6831
rect 7748 6802 7800 6808
rect 7656 6656 7708 6662
rect 7656 6598 7708 6604
rect 7380 6452 7432 6458
rect 7380 6394 7432 6400
rect 7380 6316 7432 6322
rect 7380 6258 7432 6264
rect 7288 6112 7340 6118
rect 7288 6054 7340 6060
rect 7116 4542 7236 4570
rect 6918 3224 6974 3233
rect 6918 3159 6974 3168
rect 6920 3120 6972 3126
rect 6920 3062 6972 3068
rect 6932 2310 6960 3062
rect 7116 3058 7144 4542
rect 7104 3052 7156 3058
rect 7104 2994 7156 3000
rect 6920 2304 6972 2310
rect 6920 2246 6972 2252
rect 6932 2038 6960 2246
rect 6920 2032 6972 2038
rect 6920 1974 6972 1980
rect 7300 800 7328 6054
rect 7392 5778 7420 6258
rect 7564 6248 7616 6254
rect 7668 6225 7696 6598
rect 7564 6190 7616 6196
rect 7654 6216 7710 6225
rect 7576 5914 7604 6190
rect 7654 6151 7710 6160
rect 7746 5944 7802 5953
rect 7564 5908 7616 5914
rect 7746 5879 7748 5888
rect 7564 5850 7616 5856
rect 7800 5879 7802 5888
rect 7748 5850 7800 5856
rect 7472 5840 7524 5846
rect 7472 5782 7524 5788
rect 7380 5772 7432 5778
rect 7380 5714 7432 5720
rect 7380 5568 7432 5574
rect 7380 5510 7432 5516
rect 7392 5098 7420 5510
rect 7380 5092 7432 5098
rect 7380 5034 7432 5040
rect 7484 2774 7512 5782
rect 7748 5296 7800 5302
rect 7748 5238 7800 5244
rect 7564 5160 7616 5166
rect 7564 5102 7616 5108
rect 7576 4457 7604 5102
rect 7760 5098 7788 5238
rect 7748 5092 7800 5098
rect 7748 5034 7800 5040
rect 7656 4616 7708 4622
rect 7760 4593 7788 5034
rect 7852 4808 7880 7754
rect 7932 7404 7984 7410
rect 7932 7346 7984 7352
rect 7944 5370 7972 7346
rect 8036 6322 8064 9114
rect 8220 9110 8248 9862
rect 8496 9382 8524 9880
rect 9140 9518 9168 10474
rect 9128 9512 9180 9518
rect 9128 9454 9180 9460
rect 8392 9376 8444 9382
rect 8392 9318 8444 9324
rect 8484 9376 8536 9382
rect 8484 9318 8536 9324
rect 8208 9104 8260 9110
rect 8404 9058 8432 9318
rect 8208 9046 8260 9052
rect 8116 9036 8168 9042
rect 8116 8978 8168 8984
rect 8312 9030 8432 9058
rect 8128 7954 8156 8978
rect 8208 8832 8260 8838
rect 8208 8774 8260 8780
rect 8220 8362 8248 8774
rect 8208 8356 8260 8362
rect 8208 8298 8260 8304
rect 8208 8084 8260 8090
rect 8208 8026 8260 8032
rect 8116 7948 8168 7954
rect 8116 7890 8168 7896
rect 8220 7342 8248 8026
rect 8208 7336 8260 7342
rect 8208 7278 8260 7284
rect 8114 6760 8170 6769
rect 8114 6695 8170 6704
rect 8128 6662 8156 6695
rect 8116 6656 8168 6662
rect 8116 6598 8168 6604
rect 8116 6452 8168 6458
rect 8116 6394 8168 6400
rect 8024 6316 8076 6322
rect 8024 6258 8076 6264
rect 8036 5846 8064 6258
rect 8128 5914 8156 6394
rect 8220 6254 8248 7278
rect 8312 6905 8340 9030
rect 8392 7744 8444 7750
rect 8392 7686 8444 7692
rect 8404 7002 8432 7686
rect 8392 6996 8444 7002
rect 8392 6938 8444 6944
rect 8298 6896 8354 6905
rect 8298 6831 8354 6840
rect 8208 6248 8260 6254
rect 8208 6190 8260 6196
rect 8116 5908 8168 5914
rect 8116 5850 8168 5856
rect 8024 5840 8076 5846
rect 8024 5782 8076 5788
rect 8312 5658 8340 6831
rect 8390 6624 8446 6633
rect 8496 6610 8524 9318
rect 8747 9276 9055 9285
rect 8747 9274 8753 9276
rect 8809 9274 8833 9276
rect 8889 9274 8913 9276
rect 8969 9274 8993 9276
rect 9049 9274 9055 9276
rect 8809 9222 8811 9274
rect 8991 9222 8993 9274
rect 8747 9220 8753 9222
rect 8809 9220 8833 9222
rect 8889 9220 8913 9222
rect 8969 9220 8993 9222
rect 9049 9220 9055 9222
rect 8747 9211 9055 9220
rect 9128 8900 9180 8906
rect 9128 8842 9180 8848
rect 8576 8832 8628 8838
rect 8576 8774 8628 8780
rect 8668 8832 8720 8838
rect 8668 8774 8720 8780
rect 8588 8294 8616 8774
rect 8680 8634 8708 8774
rect 8668 8628 8720 8634
rect 8668 8570 8720 8576
rect 9140 8430 9168 8842
rect 8668 8424 8720 8430
rect 8668 8366 8720 8372
rect 9128 8424 9180 8430
rect 9128 8366 9180 8372
rect 8576 8288 8628 8294
rect 8576 8230 8628 8236
rect 8576 7744 8628 7750
rect 8680 7732 8708 8366
rect 8747 8188 9055 8197
rect 8747 8186 8753 8188
rect 8809 8186 8833 8188
rect 8889 8186 8913 8188
rect 8969 8186 8993 8188
rect 9049 8186 9055 8188
rect 8809 8134 8811 8186
rect 8991 8134 8993 8186
rect 8747 8132 8753 8134
rect 8809 8132 8833 8134
rect 8889 8132 8913 8134
rect 8969 8132 8993 8134
rect 9049 8132 9055 8134
rect 8747 8123 9055 8132
rect 9140 8129 9168 8366
rect 9126 8120 9182 8129
rect 9126 8055 9182 8064
rect 9232 7834 9260 15846
rect 9324 13308 9352 15846
rect 9416 15570 9444 16390
rect 9404 15564 9456 15570
rect 9404 15506 9456 15512
rect 9404 15360 9456 15366
rect 9402 15328 9404 15337
rect 9456 15328 9458 15337
rect 9402 15263 9458 15272
rect 9404 14816 9456 14822
rect 9404 14758 9456 14764
rect 9416 14482 9444 14758
rect 9404 14476 9456 14482
rect 9404 14418 9456 14424
rect 9508 13462 9536 16526
rect 9600 14278 9628 17983
rect 9692 15162 9720 18108
rect 9956 18090 10008 18096
rect 9770 18048 9826 18057
rect 9770 17983 9826 17992
rect 9784 16998 9812 17983
rect 9956 17876 10008 17882
rect 9956 17818 10008 17824
rect 9864 17672 9916 17678
rect 9864 17614 9916 17620
rect 9772 16992 9824 16998
rect 9772 16934 9824 16940
rect 9770 16552 9826 16561
rect 9770 16487 9772 16496
rect 9824 16487 9826 16496
rect 9772 16458 9824 16464
rect 9772 15972 9824 15978
rect 9772 15914 9824 15920
rect 9680 15156 9732 15162
rect 9680 15098 9732 15104
rect 9588 14272 9640 14278
rect 9784 14260 9812 15914
rect 9876 15144 9904 17614
rect 9968 16182 9996 17818
rect 10060 16232 10088 18838
rect 10140 18692 10192 18698
rect 10140 18634 10192 18640
rect 10152 18426 10180 18634
rect 10140 18420 10192 18426
rect 10140 18362 10192 18368
rect 10232 18352 10284 18358
rect 10232 18294 10284 18300
rect 10060 16204 10180 16232
rect 9956 16176 10008 16182
rect 9956 16118 10008 16124
rect 10048 16108 10100 16114
rect 10048 16050 10100 16056
rect 9956 15904 10008 15910
rect 9956 15846 10008 15852
rect 9968 15570 9996 15846
rect 9956 15564 10008 15570
rect 9956 15506 10008 15512
rect 9876 15116 9996 15144
rect 9864 15020 9916 15026
rect 9864 14962 9916 14968
rect 9588 14214 9640 14220
rect 9692 14232 9812 14260
rect 9692 14090 9720 14232
rect 9600 14062 9720 14090
rect 9770 14104 9826 14113
rect 9496 13456 9548 13462
rect 9496 13398 9548 13404
rect 9324 13280 9536 13308
rect 9312 13184 9364 13190
rect 9312 13126 9364 13132
rect 9404 13184 9456 13190
rect 9404 13126 9456 13132
rect 9324 12442 9352 13126
rect 9312 12436 9364 12442
rect 9312 12378 9364 12384
rect 9312 12232 9364 12238
rect 9312 12174 9364 12180
rect 9324 11898 9352 12174
rect 9312 11892 9364 11898
rect 9312 11834 9364 11840
rect 9312 11280 9364 11286
rect 9312 11222 9364 11228
rect 9324 10674 9352 11222
rect 9416 11218 9444 13126
rect 9508 12481 9536 13280
rect 9600 13190 9628 14062
rect 9770 14039 9772 14048
rect 9824 14039 9826 14048
rect 9772 14010 9824 14016
rect 9772 13932 9824 13938
rect 9772 13874 9824 13880
rect 9680 13796 9732 13802
rect 9680 13738 9732 13744
rect 9692 13530 9720 13738
rect 9680 13524 9732 13530
rect 9680 13466 9732 13472
rect 9588 13184 9640 13190
rect 9588 13126 9640 13132
rect 9680 13184 9732 13190
rect 9680 13126 9732 13132
rect 9588 12844 9640 12850
rect 9588 12786 9640 12792
rect 9494 12472 9550 12481
rect 9494 12407 9550 12416
rect 9600 12306 9628 12786
rect 9692 12434 9720 13126
rect 9784 12714 9812 13874
rect 9772 12708 9824 12714
rect 9772 12650 9824 12656
rect 9692 12406 9812 12434
rect 9496 12300 9548 12306
rect 9496 12242 9548 12248
rect 9588 12300 9640 12306
rect 9588 12242 9640 12248
rect 9508 12209 9536 12242
rect 9494 12200 9550 12209
rect 9494 12135 9550 12144
rect 9494 12064 9550 12073
rect 9494 11999 9550 12008
rect 9404 11212 9456 11218
rect 9404 11154 9456 11160
rect 9404 11008 9456 11014
rect 9404 10950 9456 10956
rect 9416 10810 9444 10950
rect 9404 10804 9456 10810
rect 9404 10746 9456 10752
rect 9312 10668 9364 10674
rect 9312 10610 9364 10616
rect 9312 10464 9364 10470
rect 9312 10406 9364 10412
rect 9324 10198 9352 10406
rect 9312 10192 9364 10198
rect 9312 10134 9364 10140
rect 9404 10124 9456 10130
rect 9404 10066 9456 10072
rect 9416 9722 9444 10066
rect 9404 9716 9456 9722
rect 9404 9658 9456 9664
rect 9508 8906 9536 11999
rect 9680 11756 9732 11762
rect 9680 11698 9732 11704
rect 9692 10810 9720 11698
rect 9784 11234 9812 12406
rect 9876 11626 9904 14962
rect 9968 12986 9996 15116
rect 10060 14618 10088 16050
rect 10048 14612 10100 14618
rect 10048 14554 10100 14560
rect 10048 14272 10100 14278
rect 10048 14214 10100 14220
rect 10060 13802 10088 14214
rect 10048 13796 10100 13802
rect 10048 13738 10100 13744
rect 9956 12980 10008 12986
rect 9956 12922 10008 12928
rect 9954 12336 10010 12345
rect 9954 12271 10010 12280
rect 9968 11694 9996 12271
rect 10048 12096 10100 12102
rect 10048 12038 10100 12044
rect 9956 11688 10008 11694
rect 9956 11630 10008 11636
rect 9864 11620 9916 11626
rect 9864 11562 9916 11568
rect 10060 11354 10088 12038
rect 10048 11348 10100 11354
rect 10048 11290 10100 11296
rect 9784 11206 9904 11234
rect 9772 11076 9824 11082
rect 9772 11018 9824 11024
rect 9680 10804 9732 10810
rect 9680 10746 9732 10752
rect 9588 10600 9640 10606
rect 9588 10542 9640 10548
rect 9600 10130 9628 10542
rect 9784 10146 9812 11018
rect 9876 10470 9904 11206
rect 9956 11076 10008 11082
rect 9956 11018 10008 11024
rect 9864 10464 9916 10470
rect 9864 10406 9916 10412
rect 9588 10124 9640 10130
rect 9588 10066 9640 10072
rect 9692 10118 9812 10146
rect 9692 9450 9720 10118
rect 9862 10024 9918 10033
rect 9862 9959 9918 9968
rect 9772 9920 9824 9926
rect 9772 9862 9824 9868
rect 9784 9654 9812 9862
rect 9772 9648 9824 9654
rect 9772 9590 9824 9596
rect 9680 9444 9732 9450
rect 9680 9386 9732 9392
rect 9876 9178 9904 9959
rect 9588 9172 9640 9178
rect 9588 9114 9640 9120
rect 9864 9172 9916 9178
rect 9864 9114 9916 9120
rect 9600 9042 9628 9114
rect 9968 9058 9996 11018
rect 10152 10742 10180 16204
rect 10244 16153 10272 18294
rect 10336 17354 10364 22200
rect 10692 20460 10744 20466
rect 10692 20402 10744 20408
rect 10600 19848 10652 19854
rect 10600 19790 10652 19796
rect 10416 19712 10468 19718
rect 10416 19654 10468 19660
rect 10428 18970 10456 19654
rect 10416 18964 10468 18970
rect 10416 18906 10468 18912
rect 10508 18828 10560 18834
rect 10508 18770 10560 18776
rect 10416 18624 10468 18630
rect 10416 18566 10468 18572
rect 10428 18358 10456 18566
rect 10416 18352 10468 18358
rect 10416 18294 10468 18300
rect 10520 18222 10548 18770
rect 10612 18465 10640 19790
rect 10598 18456 10654 18465
rect 10598 18391 10654 18400
rect 10508 18216 10560 18222
rect 10508 18158 10560 18164
rect 10336 17326 10640 17354
rect 10416 17196 10468 17202
rect 10416 17138 10468 17144
rect 10324 16448 10376 16454
rect 10324 16390 10376 16396
rect 10230 16144 10286 16153
rect 10230 16079 10286 16088
rect 10230 16008 10286 16017
rect 10230 15943 10286 15952
rect 10244 15706 10272 15943
rect 10232 15700 10284 15706
rect 10232 15642 10284 15648
rect 10232 14816 10284 14822
rect 10230 14784 10232 14793
rect 10284 14784 10286 14793
rect 10230 14719 10286 14728
rect 10336 14414 10364 16390
rect 10324 14408 10376 14414
rect 10324 14350 10376 14356
rect 10324 14272 10376 14278
rect 10428 14260 10456 17138
rect 10506 16144 10562 16153
rect 10506 16079 10562 16088
rect 10520 16046 10548 16079
rect 10508 16040 10560 16046
rect 10508 15982 10560 15988
rect 10612 15042 10640 17326
rect 10704 17270 10732 20402
rect 10692 17264 10744 17270
rect 10692 17206 10744 17212
rect 10692 16992 10744 16998
rect 10692 16934 10744 16940
rect 10704 16726 10732 16934
rect 10692 16720 10744 16726
rect 10692 16662 10744 16668
rect 10704 15570 10732 16662
rect 10796 16250 10824 22200
rect 11256 22114 11284 22200
rect 11348 22114 11376 22222
rect 11256 22086 11376 22114
rect 11244 21004 11296 21010
rect 11244 20946 11296 20952
rect 11060 20528 11112 20534
rect 11060 20470 11112 20476
rect 11072 19922 11100 20470
rect 11152 20324 11204 20330
rect 11152 20266 11204 20272
rect 11060 19916 11112 19922
rect 11060 19858 11112 19864
rect 11060 19712 11112 19718
rect 11060 19654 11112 19660
rect 10876 19168 10928 19174
rect 10876 19110 10928 19116
rect 10784 16244 10836 16250
rect 10784 16186 10836 16192
rect 10784 15972 10836 15978
rect 10784 15914 10836 15920
rect 10692 15564 10744 15570
rect 10692 15506 10744 15512
rect 10692 15360 10744 15366
rect 10692 15302 10744 15308
rect 10704 15162 10732 15302
rect 10692 15156 10744 15162
rect 10692 15098 10744 15104
rect 10612 15014 10732 15042
rect 10508 14884 10560 14890
rect 10508 14826 10560 14832
rect 10520 14618 10548 14826
rect 10508 14612 10560 14618
rect 10508 14554 10560 14560
rect 10508 14408 10560 14414
rect 10508 14350 10560 14356
rect 10376 14232 10456 14260
rect 10324 14214 10376 14220
rect 10416 14068 10468 14074
rect 10416 14010 10468 14016
rect 10324 14000 10376 14006
rect 10324 13942 10376 13948
rect 10232 13864 10284 13870
rect 10336 13852 10364 13942
rect 10284 13824 10364 13852
rect 10428 13852 10456 14010
rect 10520 13977 10548 14350
rect 10506 13968 10562 13977
rect 10506 13903 10562 13912
rect 10508 13864 10560 13870
rect 10428 13824 10508 13852
rect 10232 13806 10284 13812
rect 10508 13806 10560 13812
rect 10416 13184 10468 13190
rect 10416 13126 10468 13132
rect 10428 12986 10456 13126
rect 10416 12980 10468 12986
rect 10416 12922 10468 12928
rect 10520 12866 10548 13806
rect 10600 13728 10652 13734
rect 10600 13670 10652 13676
rect 10428 12838 10548 12866
rect 10232 11552 10284 11558
rect 10232 11494 10284 11500
rect 10244 11014 10272 11494
rect 10232 11008 10284 11014
rect 10232 10950 10284 10956
rect 10140 10736 10192 10742
rect 10140 10678 10192 10684
rect 10048 10668 10100 10674
rect 10048 10610 10100 10616
rect 10060 10062 10088 10610
rect 10152 10266 10180 10678
rect 10140 10260 10192 10266
rect 10140 10202 10192 10208
rect 10048 10056 10100 10062
rect 10048 9998 10100 10004
rect 10060 9450 10088 9998
rect 10152 9625 10180 10202
rect 10138 9616 10194 9625
rect 10138 9551 10194 9560
rect 10048 9444 10100 9450
rect 10048 9386 10100 9392
rect 9588 9036 9640 9042
rect 9588 8978 9640 8984
rect 9784 9030 9996 9058
rect 9496 8900 9548 8906
rect 9496 8842 9548 8848
rect 9588 8900 9640 8906
rect 9588 8842 9640 8848
rect 9600 8786 9628 8842
rect 8628 7704 8708 7732
rect 9140 7806 9260 7834
rect 9508 8758 9628 8786
rect 9312 7812 9364 7818
rect 8576 7686 8628 7692
rect 8588 7449 8616 7686
rect 8574 7440 8630 7449
rect 8574 7375 8630 7384
rect 8668 7404 8720 7410
rect 8668 7346 8720 7352
rect 8576 6860 8628 6866
rect 8576 6802 8628 6808
rect 8588 6769 8616 6802
rect 8574 6760 8630 6769
rect 8574 6695 8630 6704
rect 8446 6582 8524 6610
rect 8390 6559 8446 6568
rect 8404 6322 8432 6559
rect 8588 6338 8616 6695
rect 8680 6458 8708 7346
rect 8747 7100 9055 7109
rect 8747 7098 8753 7100
rect 8809 7098 8833 7100
rect 8889 7098 8913 7100
rect 8969 7098 8993 7100
rect 9049 7098 9055 7100
rect 8809 7046 8811 7098
rect 8991 7046 8993 7098
rect 8747 7044 8753 7046
rect 8809 7044 8833 7046
rect 8889 7044 8913 7046
rect 8969 7044 8993 7046
rect 9049 7044 9055 7046
rect 8747 7035 9055 7044
rect 9036 6860 9088 6866
rect 9036 6802 9088 6808
rect 9048 6633 9076 6802
rect 9140 6662 9168 7806
rect 9312 7754 9364 7760
rect 9324 7002 9352 7754
rect 9404 7744 9456 7750
rect 9404 7686 9456 7692
rect 9312 6996 9364 7002
rect 9312 6938 9364 6944
rect 9128 6656 9180 6662
rect 9034 6624 9090 6633
rect 9128 6598 9180 6604
rect 9034 6559 9090 6568
rect 9048 6458 9076 6559
rect 8668 6452 8720 6458
rect 8668 6394 8720 6400
rect 9036 6452 9088 6458
rect 9036 6394 9088 6400
rect 8392 6316 8444 6322
rect 8588 6310 8708 6338
rect 8392 6258 8444 6264
rect 8404 5846 8432 6258
rect 8484 6248 8536 6254
rect 8484 6190 8536 6196
rect 8496 6089 8524 6190
rect 8482 6080 8538 6089
rect 8482 6015 8538 6024
rect 8392 5840 8444 5846
rect 8392 5782 8444 5788
rect 8312 5630 8432 5658
rect 7932 5364 7984 5370
rect 7932 5306 7984 5312
rect 8300 5092 8352 5098
rect 8300 5034 8352 5040
rect 7932 4820 7984 4826
rect 7852 4780 7932 4808
rect 7932 4762 7984 4768
rect 7944 4690 7972 4762
rect 7932 4684 7984 4690
rect 7932 4626 7984 4632
rect 7656 4558 7708 4564
rect 7746 4584 7802 4593
rect 7562 4448 7618 4457
rect 7562 4383 7618 4392
rect 7564 4072 7616 4078
rect 7564 4014 7616 4020
rect 7576 3913 7604 4014
rect 7562 3904 7618 3913
rect 7562 3839 7618 3848
rect 7668 3126 7696 4558
rect 8312 4554 8340 5034
rect 7746 4519 7802 4528
rect 8300 4548 8352 4554
rect 8300 4490 8352 4496
rect 7840 4276 7892 4282
rect 7840 4218 7892 4224
rect 7852 4078 7880 4218
rect 7932 4208 7984 4214
rect 7932 4150 7984 4156
rect 8208 4208 8260 4214
rect 8208 4150 8260 4156
rect 7840 4072 7892 4078
rect 7840 4014 7892 4020
rect 7748 3732 7800 3738
rect 7748 3674 7800 3680
rect 7656 3120 7708 3126
rect 7656 3062 7708 3068
rect 7656 2984 7708 2990
rect 7656 2926 7708 2932
rect 7484 2746 7604 2774
rect 7576 2106 7604 2746
rect 7668 2446 7696 2926
rect 7656 2440 7708 2446
rect 7656 2382 7708 2388
rect 7564 2100 7616 2106
rect 7564 2042 7616 2048
rect 7760 800 7788 3674
rect 7840 3664 7892 3670
rect 7840 3606 7892 3612
rect 7852 2990 7880 3606
rect 7840 2984 7892 2990
rect 7840 2926 7892 2932
rect 7944 2446 7972 4150
rect 8114 4040 8170 4049
rect 8114 3975 8116 3984
rect 8168 3975 8170 3984
rect 8116 3946 8168 3952
rect 8024 3936 8076 3942
rect 8024 3878 8076 3884
rect 8036 3670 8064 3878
rect 8220 3720 8248 4150
rect 8404 4026 8432 5630
rect 8496 5166 8524 6015
rect 8576 5772 8628 5778
rect 8576 5714 8628 5720
rect 8484 5160 8536 5166
rect 8484 5102 8536 5108
rect 8484 5024 8536 5030
rect 8588 5001 8616 5714
rect 8484 4966 8536 4972
rect 8574 4992 8630 5001
rect 8496 4593 8524 4966
rect 8574 4927 8630 4936
rect 8680 4842 8708 6310
rect 8747 6012 9055 6021
rect 8747 6010 8753 6012
rect 8809 6010 8833 6012
rect 8889 6010 8913 6012
rect 8969 6010 8993 6012
rect 9049 6010 9055 6012
rect 8809 5958 8811 6010
rect 8991 5958 8993 6010
rect 8747 5956 8753 5958
rect 8809 5956 8833 5958
rect 8889 5956 8913 5958
rect 8969 5956 8993 5958
rect 9049 5956 9055 5958
rect 8747 5947 9055 5956
rect 9036 5840 9088 5846
rect 8956 5800 9036 5828
rect 8956 5642 8984 5800
rect 9036 5782 9088 5788
rect 9140 5681 9168 6598
rect 9416 6497 9444 7686
rect 9402 6488 9458 6497
rect 9402 6423 9458 6432
rect 9218 5944 9274 5953
rect 9218 5879 9274 5888
rect 9232 5760 9260 5879
rect 9508 5778 9536 8758
rect 9784 8430 9812 9030
rect 9956 8968 10008 8974
rect 9956 8910 10008 8916
rect 9968 8634 9996 8910
rect 9956 8628 10008 8634
rect 9956 8570 10008 8576
rect 9772 8424 9824 8430
rect 9864 8424 9916 8430
rect 9772 8366 9824 8372
rect 9862 8392 9864 8401
rect 9916 8392 9918 8401
rect 9588 7744 9640 7750
rect 9588 7686 9640 7692
rect 9600 7546 9628 7686
rect 9588 7540 9640 7546
rect 9588 7482 9640 7488
rect 9588 7336 9640 7342
rect 9586 7304 9588 7313
rect 9640 7304 9642 7313
rect 9586 7239 9642 7248
rect 9784 6866 9812 8366
rect 9862 8327 9918 8336
rect 9864 8288 9916 8294
rect 9864 8230 9916 8236
rect 9876 7206 9904 8230
rect 9864 7200 9916 7206
rect 9864 7142 9916 7148
rect 9772 6860 9824 6866
rect 9772 6802 9824 6808
rect 9586 6760 9642 6769
rect 9876 6746 9904 7142
rect 9586 6695 9642 6704
rect 9784 6718 9904 6746
rect 9600 6254 9628 6695
rect 9588 6248 9640 6254
rect 9588 6190 9640 6196
rect 9496 5772 9548 5778
rect 9232 5732 9444 5760
rect 9126 5672 9182 5681
rect 8944 5636 8996 5642
rect 9126 5607 9182 5616
rect 8944 5578 8996 5584
rect 8852 5568 8904 5574
rect 9232 5522 9260 5732
rect 9312 5636 9364 5642
rect 9312 5578 9364 5584
rect 8852 5510 8904 5516
rect 8864 5098 8892 5510
rect 8956 5494 9260 5522
rect 8956 5370 8984 5494
rect 9324 5386 9352 5578
rect 9416 5545 9444 5732
rect 9496 5714 9548 5720
rect 9402 5536 9458 5545
rect 9402 5471 9458 5480
rect 8944 5364 8996 5370
rect 8944 5306 8996 5312
rect 9048 5358 9352 5386
rect 9416 5370 9444 5471
rect 9404 5364 9456 5370
rect 8852 5092 8904 5098
rect 9048 5080 9076 5358
rect 9404 5306 9456 5312
rect 9312 5160 9364 5166
rect 9312 5102 9364 5108
rect 9494 5128 9550 5137
rect 9048 5052 9260 5080
rect 8852 5034 8904 5040
rect 8747 4924 9055 4933
rect 8747 4922 8753 4924
rect 8809 4922 8833 4924
rect 8889 4922 8913 4924
rect 8969 4922 8993 4924
rect 9049 4922 9055 4924
rect 8809 4870 8811 4922
rect 8991 4870 8993 4922
rect 8747 4868 8753 4870
rect 8809 4868 8833 4870
rect 8889 4868 8913 4870
rect 8969 4868 8993 4870
rect 9049 4868 9055 4870
rect 8747 4859 9055 4868
rect 8588 4814 8708 4842
rect 9126 4856 9182 4865
rect 8760 4820 8812 4826
rect 8588 4604 8616 4814
rect 8760 4762 8812 4768
rect 9036 4820 9088 4826
rect 9126 4791 9182 4800
rect 9036 4762 9088 4768
rect 8772 4729 8800 4762
rect 8758 4720 8814 4729
rect 8758 4655 8814 4664
rect 8482 4584 8538 4593
rect 8588 4576 8708 4604
rect 8482 4519 8538 4528
rect 8576 4140 8628 4146
rect 8128 3692 8248 3720
rect 8312 3998 8432 4026
rect 8496 4100 8576 4128
rect 8024 3664 8076 3670
rect 8024 3606 8076 3612
rect 8128 2650 8156 3692
rect 8206 3632 8262 3641
rect 8206 3567 8262 3576
rect 8116 2644 8168 2650
rect 8116 2586 8168 2592
rect 7932 2440 7984 2446
rect 7932 2382 7984 2388
rect 8220 800 8248 3567
rect 6472 734 6684 762
rect 6826 0 6882 800
rect 7286 0 7342 800
rect 7746 0 7802 800
rect 8206 0 8262 800
rect 8312 762 8340 3998
rect 8392 3936 8444 3942
rect 8496 3924 8524 4100
rect 8576 4082 8628 4088
rect 8444 3896 8524 3924
rect 8576 3936 8628 3942
rect 8574 3904 8576 3913
rect 8628 3904 8630 3913
rect 8392 3878 8444 3884
rect 8574 3839 8630 3848
rect 8576 3120 8628 3126
rect 8576 3062 8628 3068
rect 8588 2378 8616 3062
rect 8680 2582 8708 4576
rect 9048 4554 9076 4762
rect 9036 4548 9088 4554
rect 9036 4490 9088 4496
rect 9140 4282 9168 4791
rect 9128 4276 9180 4282
rect 9128 4218 9180 4224
rect 9232 4010 9260 5052
rect 9324 5030 9352 5102
rect 9416 5072 9494 5080
rect 9416 5063 9550 5072
rect 9416 5052 9536 5063
rect 9312 5024 9364 5030
rect 9312 4966 9364 4972
rect 9324 4622 9352 4966
rect 9312 4616 9364 4622
rect 9312 4558 9364 4564
rect 9416 4457 9444 5052
rect 9496 4480 9548 4486
rect 9402 4448 9458 4457
rect 9496 4422 9548 4428
rect 9402 4383 9458 4392
rect 9508 4282 9536 4422
rect 9496 4276 9548 4282
rect 9496 4218 9548 4224
rect 9508 4078 9536 4218
rect 9678 4176 9734 4185
rect 9678 4111 9680 4120
rect 9732 4111 9734 4120
rect 9680 4082 9732 4088
rect 9496 4072 9548 4078
rect 9496 4014 9548 4020
rect 9220 4004 9272 4010
rect 9220 3946 9272 3952
rect 9586 3904 9642 3913
rect 8747 3836 9055 3845
rect 9586 3839 9642 3848
rect 8747 3834 8753 3836
rect 8809 3834 8833 3836
rect 8889 3834 8913 3836
rect 8969 3834 8993 3836
rect 9049 3834 9055 3836
rect 8809 3782 8811 3834
rect 8991 3782 8993 3834
rect 8747 3780 8753 3782
rect 8809 3780 8833 3782
rect 8889 3780 8913 3782
rect 8969 3780 8993 3782
rect 9049 3780 9055 3782
rect 8747 3771 9055 3780
rect 9126 3360 9182 3369
rect 9126 3295 9182 3304
rect 9140 2990 9168 3295
rect 9312 3052 9364 3058
rect 9312 2994 9364 3000
rect 9128 2984 9180 2990
rect 9128 2926 9180 2932
rect 8747 2748 9055 2757
rect 8747 2746 8753 2748
rect 8809 2746 8833 2748
rect 8889 2746 8913 2748
rect 8969 2746 8993 2748
rect 9049 2746 9055 2748
rect 8809 2694 8811 2746
rect 8991 2694 8993 2746
rect 8747 2692 8753 2694
rect 8809 2692 8833 2694
rect 8889 2692 8913 2694
rect 8969 2692 8993 2694
rect 9049 2692 9055 2694
rect 8747 2683 9055 2692
rect 8668 2576 8720 2582
rect 8668 2518 8720 2524
rect 9126 2544 9182 2553
rect 9126 2479 9182 2488
rect 8576 2372 8628 2378
rect 8576 2314 8628 2320
rect 8588 870 8708 898
rect 8588 762 8616 870
rect 8680 800 8708 870
rect 9140 800 9168 2479
rect 9324 2378 9352 2994
rect 9312 2372 9364 2378
rect 9312 2314 9364 2320
rect 9600 800 9628 3839
rect 9784 3738 9812 6718
rect 9876 6662 9904 6718
rect 9956 6724 10008 6730
rect 9956 6666 10008 6672
rect 9864 6656 9916 6662
rect 9864 6598 9916 6604
rect 9968 6458 9996 6666
rect 9956 6452 10008 6458
rect 9956 6394 10008 6400
rect 9864 6248 9916 6254
rect 9864 6190 9916 6196
rect 9876 5846 9904 6190
rect 9864 5840 9916 5846
rect 9864 5782 9916 5788
rect 9956 5228 10008 5234
rect 9956 5170 10008 5176
rect 9968 5001 9996 5170
rect 9954 4992 10010 5001
rect 9954 4927 10010 4936
rect 9772 3732 9824 3738
rect 9772 3674 9824 3680
rect 9954 3632 10010 3641
rect 9954 3567 9956 3576
rect 10008 3567 10010 3576
rect 9956 3538 10008 3544
rect 9772 3460 9824 3466
rect 9772 3402 9824 3408
rect 9784 3194 9812 3402
rect 9956 3392 10008 3398
rect 9956 3334 10008 3340
rect 9772 3188 9824 3194
rect 9772 3130 9824 3136
rect 9968 3058 9996 3334
rect 9956 3052 10008 3058
rect 9956 2994 10008 3000
rect 9678 2952 9734 2961
rect 9678 2887 9680 2896
rect 9732 2887 9734 2896
rect 9680 2858 9732 2864
rect 10060 800 10088 9386
rect 10140 9376 10192 9382
rect 10140 9318 10192 9324
rect 10152 9042 10180 9318
rect 10140 9036 10192 9042
rect 10140 8978 10192 8984
rect 10138 8528 10194 8537
rect 10138 8463 10194 8472
rect 10152 5642 10180 8463
rect 10140 5636 10192 5642
rect 10140 5578 10192 5584
rect 10140 4684 10192 4690
rect 10140 4626 10192 4632
rect 10152 3126 10180 4626
rect 10140 3120 10192 3126
rect 10140 3062 10192 3068
rect 10152 2650 10180 3062
rect 10140 2644 10192 2650
rect 10140 2586 10192 2592
rect 8312 734 8616 762
rect 8666 0 8722 800
rect 9126 0 9182 800
rect 9586 0 9642 800
rect 10046 0 10102 800
rect 10244 762 10272 10950
rect 10322 9616 10378 9625
rect 10322 9551 10378 9560
rect 10336 9042 10364 9551
rect 10324 9036 10376 9042
rect 10324 8978 10376 8984
rect 10324 8288 10376 8294
rect 10428 8276 10456 12838
rect 10612 12442 10640 13670
rect 10600 12436 10652 12442
rect 10600 12378 10652 12384
rect 10704 12050 10732 15014
rect 10796 14113 10824 15914
rect 10782 14104 10838 14113
rect 10782 14039 10838 14048
rect 10888 13870 10916 19110
rect 11072 18766 11100 19654
rect 10968 18760 11020 18766
rect 10968 18702 11020 18708
rect 11060 18760 11112 18766
rect 11060 18702 11112 18708
rect 10980 17882 11008 18702
rect 10968 17876 11020 17882
rect 10968 17818 11020 17824
rect 10968 17264 11020 17270
rect 10968 17206 11020 17212
rect 10980 16998 11008 17206
rect 10968 16992 11020 16998
rect 10968 16934 11020 16940
rect 11072 16538 11100 18702
rect 11164 16590 11192 20266
rect 10980 16510 11100 16538
rect 11152 16584 11204 16590
rect 11152 16526 11204 16532
rect 10980 15162 11008 16510
rect 11060 16448 11112 16454
rect 11060 16390 11112 16396
rect 11072 16250 11100 16390
rect 11060 16244 11112 16250
rect 11060 16186 11112 16192
rect 11152 16244 11204 16250
rect 11152 16186 11204 16192
rect 11164 16130 11192 16186
rect 11072 16102 11192 16130
rect 11072 15366 11100 16102
rect 11152 16040 11204 16046
rect 11152 15982 11204 15988
rect 11164 15502 11192 15982
rect 11152 15496 11204 15502
rect 11152 15438 11204 15444
rect 11060 15360 11112 15366
rect 11058 15328 11060 15337
rect 11256 15348 11284 20946
rect 11624 20890 11652 22222
rect 11702 22200 11758 23000
rect 12162 22200 12218 23000
rect 12622 22200 12678 23000
rect 13082 22200 13138 23000
rect 13542 22200 13598 23000
rect 14002 22200 14058 23000
rect 14462 22200 14518 23000
rect 14568 22222 14872 22250
rect 11716 21010 11744 22200
rect 11704 21004 11756 21010
rect 11704 20946 11756 20952
rect 11624 20862 11744 20890
rect 11346 20700 11654 20709
rect 11346 20698 11352 20700
rect 11408 20698 11432 20700
rect 11488 20698 11512 20700
rect 11568 20698 11592 20700
rect 11648 20698 11654 20700
rect 11408 20646 11410 20698
rect 11590 20646 11592 20698
rect 11346 20644 11352 20646
rect 11408 20644 11432 20646
rect 11488 20644 11512 20646
rect 11568 20644 11592 20646
rect 11648 20644 11654 20646
rect 11346 20635 11654 20644
rect 11346 19612 11654 19621
rect 11346 19610 11352 19612
rect 11408 19610 11432 19612
rect 11488 19610 11512 19612
rect 11568 19610 11592 19612
rect 11648 19610 11654 19612
rect 11408 19558 11410 19610
rect 11590 19558 11592 19610
rect 11346 19556 11352 19558
rect 11408 19556 11432 19558
rect 11488 19556 11512 19558
rect 11568 19556 11592 19558
rect 11648 19556 11654 19558
rect 11346 19547 11654 19556
rect 11346 18524 11654 18533
rect 11346 18522 11352 18524
rect 11408 18522 11432 18524
rect 11488 18522 11512 18524
rect 11568 18522 11592 18524
rect 11648 18522 11654 18524
rect 11408 18470 11410 18522
rect 11590 18470 11592 18522
rect 11346 18468 11352 18470
rect 11408 18468 11432 18470
rect 11488 18468 11512 18470
rect 11568 18468 11592 18470
rect 11648 18468 11654 18470
rect 11346 18459 11654 18468
rect 11336 18080 11388 18086
rect 11336 18022 11388 18028
rect 11348 17882 11376 18022
rect 11610 17912 11666 17921
rect 11336 17876 11388 17882
rect 11610 17847 11666 17856
rect 11336 17818 11388 17824
rect 11624 17814 11652 17847
rect 11612 17808 11664 17814
rect 11612 17750 11664 17756
rect 11346 17436 11654 17445
rect 11346 17434 11352 17436
rect 11408 17434 11432 17436
rect 11488 17434 11512 17436
rect 11568 17434 11592 17436
rect 11648 17434 11654 17436
rect 11408 17382 11410 17434
rect 11590 17382 11592 17434
rect 11346 17380 11352 17382
rect 11408 17380 11432 17382
rect 11488 17380 11512 17382
rect 11568 17380 11592 17382
rect 11648 17380 11654 17382
rect 11346 17371 11654 17380
rect 11520 16992 11572 16998
rect 11520 16934 11572 16940
rect 11532 16833 11560 16934
rect 11518 16824 11574 16833
rect 11518 16759 11574 16768
rect 11346 16348 11654 16357
rect 11346 16346 11352 16348
rect 11408 16346 11432 16348
rect 11488 16346 11512 16348
rect 11568 16346 11592 16348
rect 11648 16346 11654 16348
rect 11408 16294 11410 16346
rect 11590 16294 11592 16346
rect 11346 16292 11352 16294
rect 11408 16292 11432 16294
rect 11488 16292 11512 16294
rect 11568 16292 11592 16294
rect 11648 16292 11654 16294
rect 11346 16283 11654 16292
rect 11612 16176 11664 16182
rect 11612 16118 11664 16124
rect 11624 15910 11652 16118
rect 11612 15904 11664 15910
rect 11612 15846 11664 15852
rect 11112 15328 11114 15337
rect 11058 15263 11114 15272
rect 11164 15320 11284 15348
rect 10968 15156 11020 15162
rect 10968 15098 11020 15104
rect 11060 14612 11112 14618
rect 11060 14554 11112 14560
rect 11072 14074 11100 14554
rect 11060 14068 11112 14074
rect 11060 14010 11112 14016
rect 10876 13864 10928 13870
rect 10876 13806 10928 13812
rect 10876 13728 10928 13734
rect 10876 13670 10928 13676
rect 10888 13190 10916 13670
rect 10968 13388 11020 13394
rect 10968 13330 11020 13336
rect 10876 13184 10928 13190
rect 10876 13126 10928 13132
rect 10980 13002 11008 13330
rect 10520 12022 10732 12050
rect 10796 12974 11008 13002
rect 10520 11218 10548 12022
rect 10796 11914 10824 12974
rect 10876 12708 10928 12714
rect 10876 12650 10928 12656
rect 10888 12306 10916 12650
rect 10968 12368 11020 12374
rect 10968 12310 11020 12316
rect 10876 12300 10928 12306
rect 10876 12242 10928 12248
rect 10612 11886 10824 11914
rect 10980 11898 11008 12310
rect 10968 11892 11020 11898
rect 10508 11212 10560 11218
rect 10508 11154 10560 11160
rect 10520 10742 10548 11154
rect 10508 10736 10560 10742
rect 10612 10713 10640 11886
rect 10968 11834 11020 11840
rect 10782 11792 10838 11801
rect 10692 11756 10744 11762
rect 10782 11727 10838 11736
rect 10692 11698 10744 11704
rect 10704 11286 10732 11698
rect 10796 11694 10824 11727
rect 10784 11688 10836 11694
rect 10784 11630 10836 11636
rect 10692 11280 10744 11286
rect 10692 11222 10744 11228
rect 10796 10996 10824 11630
rect 10980 11626 11008 11834
rect 11072 11830 11100 14010
rect 11164 12374 11192 15320
rect 11346 15260 11654 15269
rect 11346 15258 11352 15260
rect 11408 15258 11432 15260
rect 11488 15258 11512 15260
rect 11568 15258 11592 15260
rect 11648 15258 11654 15260
rect 11408 15206 11410 15258
rect 11590 15206 11592 15258
rect 11346 15204 11352 15206
rect 11408 15204 11432 15206
rect 11488 15204 11512 15206
rect 11568 15204 11592 15206
rect 11648 15204 11654 15206
rect 11346 15195 11654 15204
rect 11244 14544 11296 14550
rect 11244 14486 11296 14492
rect 11256 14074 11284 14486
rect 11346 14172 11654 14181
rect 11346 14170 11352 14172
rect 11408 14170 11432 14172
rect 11488 14170 11512 14172
rect 11568 14170 11592 14172
rect 11648 14170 11654 14172
rect 11408 14118 11410 14170
rect 11590 14118 11592 14170
rect 11346 14116 11352 14118
rect 11408 14116 11432 14118
rect 11488 14116 11512 14118
rect 11568 14116 11592 14118
rect 11648 14116 11654 14118
rect 11346 14107 11654 14116
rect 11244 14068 11296 14074
rect 11244 14010 11296 14016
rect 11520 13320 11572 13326
rect 11518 13288 11520 13297
rect 11572 13288 11574 13297
rect 11518 13223 11574 13232
rect 11244 13184 11296 13190
rect 11244 13126 11296 13132
rect 11152 12368 11204 12374
rect 11152 12310 11204 12316
rect 11152 12232 11204 12238
rect 11152 12174 11204 12180
rect 11060 11824 11112 11830
rect 11060 11766 11112 11772
rect 10968 11620 11020 11626
rect 10968 11562 11020 11568
rect 10980 11354 11008 11562
rect 10968 11348 11020 11354
rect 10968 11290 11020 11296
rect 11072 11082 11100 11766
rect 11164 11558 11192 12174
rect 11256 11898 11284 13126
rect 11346 13084 11654 13093
rect 11346 13082 11352 13084
rect 11408 13082 11432 13084
rect 11488 13082 11512 13084
rect 11568 13082 11592 13084
rect 11648 13082 11654 13084
rect 11408 13030 11410 13082
rect 11590 13030 11592 13082
rect 11346 13028 11352 13030
rect 11408 13028 11432 13030
rect 11488 13028 11512 13030
rect 11568 13028 11592 13030
rect 11648 13028 11654 13030
rect 11346 13019 11654 13028
rect 11716 12170 11744 20862
rect 11888 19712 11940 19718
rect 11888 19654 11940 19660
rect 11900 19514 11928 19654
rect 11888 19508 11940 19514
rect 11888 19450 11940 19456
rect 11794 16824 11850 16833
rect 11794 16759 11850 16768
rect 11808 14414 11836 16759
rect 11900 15473 11928 19450
rect 11980 18692 12032 18698
rect 11980 18634 12032 18640
rect 11992 18086 12020 18634
rect 11980 18080 12032 18086
rect 11980 18022 12032 18028
rect 11980 16448 12032 16454
rect 11980 16390 12032 16396
rect 12072 16448 12124 16454
rect 12072 16390 12124 16396
rect 11886 15464 11942 15473
rect 11886 15399 11942 15408
rect 11796 14408 11848 14414
rect 11796 14350 11848 14356
rect 11888 14272 11940 14278
rect 11888 14214 11940 14220
rect 11796 13864 11848 13870
rect 11796 13806 11848 13812
rect 11808 12628 11836 13806
rect 11900 12782 11928 14214
rect 11992 13870 12020 16390
rect 12084 16114 12112 16390
rect 12072 16108 12124 16114
rect 12072 16050 12124 16056
rect 12072 14816 12124 14822
rect 12072 14758 12124 14764
rect 11980 13864 12032 13870
rect 11980 13806 12032 13812
rect 11980 13388 12032 13394
rect 11980 13330 12032 13336
rect 11992 13190 12020 13330
rect 11980 13184 12032 13190
rect 11980 13126 12032 13132
rect 11992 13025 12020 13126
rect 11978 13016 12034 13025
rect 11978 12951 12034 12960
rect 12084 12850 12112 14758
rect 12072 12844 12124 12850
rect 12072 12786 12124 12792
rect 11888 12776 11940 12782
rect 11888 12718 11940 12724
rect 11808 12600 11928 12628
rect 11794 12472 11850 12481
rect 11794 12407 11850 12416
rect 11900 12434 11928 12600
rect 11808 12238 11836 12407
rect 11900 12406 12020 12434
rect 11796 12232 11848 12238
rect 11796 12174 11848 12180
rect 11888 12232 11940 12238
rect 11888 12174 11940 12180
rect 11704 12164 11756 12170
rect 11704 12106 11756 12112
rect 11346 11996 11654 12005
rect 11346 11994 11352 11996
rect 11408 11994 11432 11996
rect 11488 11994 11512 11996
rect 11568 11994 11592 11996
rect 11648 11994 11654 11996
rect 11408 11942 11410 11994
rect 11590 11942 11592 11994
rect 11346 11940 11352 11942
rect 11408 11940 11432 11942
rect 11488 11940 11512 11942
rect 11568 11940 11592 11942
rect 11648 11940 11654 11942
rect 11346 11931 11654 11940
rect 11244 11892 11296 11898
rect 11244 11834 11296 11840
rect 11716 11830 11744 12106
rect 11900 12050 11928 12174
rect 11992 12170 12020 12406
rect 11980 12164 12032 12170
rect 11980 12106 12032 12112
rect 11808 12022 11928 12050
rect 11704 11824 11756 11830
rect 11704 11766 11756 11772
rect 11336 11688 11388 11694
rect 11336 11630 11388 11636
rect 11152 11552 11204 11558
rect 11152 11494 11204 11500
rect 11060 11076 11112 11082
rect 11060 11018 11112 11024
rect 10796 10968 10916 10996
rect 10692 10804 10744 10810
rect 10692 10746 10744 10752
rect 10508 10678 10560 10684
rect 10598 10704 10654 10713
rect 10598 10639 10654 10648
rect 10600 9920 10652 9926
rect 10600 9862 10652 9868
rect 10612 9217 10640 9862
rect 10598 9208 10654 9217
rect 10598 9143 10654 9152
rect 10704 9042 10732 10746
rect 10888 10606 10916 10968
rect 10784 10600 10836 10606
rect 10784 10542 10836 10548
rect 10876 10600 10928 10606
rect 10876 10542 10928 10548
rect 10796 9994 10824 10542
rect 10784 9988 10836 9994
rect 10784 9930 10836 9936
rect 10784 9716 10836 9722
rect 10784 9658 10836 9664
rect 10692 9036 10744 9042
rect 10692 8978 10744 8984
rect 10600 8968 10652 8974
rect 10600 8910 10652 8916
rect 10508 8832 10560 8838
rect 10508 8774 10560 8780
rect 10520 8634 10548 8774
rect 10612 8634 10640 8910
rect 10508 8628 10560 8634
rect 10508 8570 10560 8576
rect 10600 8628 10652 8634
rect 10600 8570 10652 8576
rect 10376 8248 10456 8276
rect 10324 8230 10376 8236
rect 10612 8106 10640 8570
rect 10428 8078 10640 8106
rect 10428 7818 10456 8078
rect 10506 7984 10562 7993
rect 10506 7919 10562 7928
rect 10520 7818 10548 7919
rect 10598 7848 10654 7857
rect 10416 7812 10468 7818
rect 10416 7754 10468 7760
rect 10508 7812 10560 7818
rect 10598 7783 10654 7792
rect 10508 7754 10560 7760
rect 10612 7478 10640 7783
rect 10600 7472 10652 7478
rect 10600 7414 10652 7420
rect 10324 7200 10376 7206
rect 10324 7142 10376 7148
rect 10336 6798 10364 7142
rect 10508 6996 10560 7002
rect 10508 6938 10560 6944
rect 10324 6792 10376 6798
rect 10324 6734 10376 6740
rect 10416 6656 10468 6662
rect 10416 6598 10468 6604
rect 10428 6458 10456 6598
rect 10416 6452 10468 6458
rect 10416 6394 10468 6400
rect 10520 6338 10548 6938
rect 10704 6866 10732 8978
rect 10692 6860 10744 6866
rect 10692 6802 10744 6808
rect 10692 6724 10744 6730
rect 10692 6666 10744 6672
rect 10336 6310 10548 6338
rect 10600 6384 10652 6390
rect 10600 6326 10652 6332
rect 10336 5166 10364 6310
rect 10612 5953 10640 6326
rect 10704 6254 10732 6666
rect 10692 6248 10744 6254
rect 10692 6190 10744 6196
rect 10598 5944 10654 5953
rect 10598 5879 10654 5888
rect 10796 5710 10824 9658
rect 10968 9648 11020 9654
rect 10968 9590 11020 9596
rect 10876 9512 10928 9518
rect 10876 9454 10928 9460
rect 10888 8838 10916 9454
rect 10876 8832 10928 8838
rect 10876 8774 10928 8780
rect 10876 7948 10928 7954
rect 10876 7890 10928 7896
rect 10888 7857 10916 7890
rect 10874 7848 10930 7857
rect 10980 7818 11008 9590
rect 11060 9444 11112 9450
rect 11060 9386 11112 9392
rect 11072 8430 11100 9386
rect 11060 8424 11112 8430
rect 11060 8366 11112 8372
rect 10874 7783 10930 7792
rect 10968 7812 11020 7818
rect 10888 7274 10916 7783
rect 10968 7754 11020 7760
rect 10876 7268 10928 7274
rect 10876 7210 10928 7216
rect 11060 7200 11112 7206
rect 10888 7148 11060 7154
rect 10888 7142 11112 7148
rect 10888 7126 11100 7142
rect 10888 6633 10916 7126
rect 11058 6896 11114 6905
rect 11058 6831 11114 6840
rect 10968 6656 11020 6662
rect 10874 6624 10930 6633
rect 10968 6598 11020 6604
rect 10874 6559 10930 6568
rect 10876 6248 10928 6254
rect 10876 6190 10928 6196
rect 10888 5914 10916 6190
rect 10876 5908 10928 5914
rect 10876 5850 10928 5856
rect 10784 5704 10836 5710
rect 10784 5646 10836 5652
rect 10600 5636 10652 5642
rect 10600 5578 10652 5584
rect 10324 5160 10376 5166
rect 10322 5128 10324 5137
rect 10508 5160 10560 5166
rect 10376 5128 10378 5137
rect 10508 5102 10560 5108
rect 10322 5063 10378 5072
rect 10414 4992 10470 5001
rect 10414 4927 10470 4936
rect 10428 4826 10456 4927
rect 10416 4820 10468 4826
rect 10416 4762 10468 4768
rect 10324 4616 10376 4622
rect 10324 4558 10376 4564
rect 10336 4078 10364 4558
rect 10428 4214 10456 4762
rect 10520 4282 10548 5102
rect 10508 4276 10560 4282
rect 10508 4218 10560 4224
rect 10416 4208 10468 4214
rect 10416 4150 10468 4156
rect 10324 4072 10376 4078
rect 10324 4014 10376 4020
rect 10508 4004 10560 4010
rect 10508 3946 10560 3952
rect 10324 3596 10376 3602
rect 10324 3538 10376 3544
rect 10416 3596 10468 3602
rect 10416 3538 10468 3544
rect 10336 2582 10364 3538
rect 10428 3194 10456 3538
rect 10416 3188 10468 3194
rect 10416 3130 10468 3136
rect 10428 2650 10456 3130
rect 10520 3058 10548 3946
rect 10612 3097 10640 5578
rect 10692 5568 10744 5574
rect 10692 5510 10744 5516
rect 10784 5568 10836 5574
rect 10784 5510 10836 5516
rect 10704 5370 10732 5510
rect 10692 5364 10744 5370
rect 10692 5306 10744 5312
rect 10796 5273 10824 5510
rect 10782 5264 10838 5273
rect 10782 5199 10838 5208
rect 10876 4276 10928 4282
rect 10876 4218 10928 4224
rect 10888 3738 10916 4218
rect 10876 3732 10928 3738
rect 10876 3674 10928 3680
rect 10598 3088 10654 3097
rect 10508 3052 10560 3058
rect 10598 3023 10654 3032
rect 10508 2994 10560 3000
rect 10612 2990 10640 3023
rect 10600 2984 10652 2990
rect 10600 2926 10652 2932
rect 10876 2848 10928 2854
rect 10876 2790 10928 2796
rect 10888 2650 10916 2790
rect 10416 2644 10468 2650
rect 10416 2586 10468 2592
rect 10876 2644 10928 2650
rect 10876 2586 10928 2592
rect 10324 2576 10376 2582
rect 10324 2518 10376 2524
rect 10428 870 10548 898
rect 10428 762 10456 870
rect 10520 800 10548 870
rect 10980 800 11008 6598
rect 11072 5409 11100 6831
rect 11058 5400 11114 5409
rect 11058 5335 11114 5344
rect 11058 4176 11114 4185
rect 11058 4111 11114 4120
rect 11072 4078 11100 4111
rect 11060 4072 11112 4078
rect 11060 4014 11112 4020
rect 11060 3732 11112 3738
rect 11060 3674 11112 3680
rect 11072 3602 11100 3674
rect 11060 3596 11112 3602
rect 11060 3538 11112 3544
rect 11058 3496 11114 3505
rect 11058 3431 11114 3440
rect 11072 3398 11100 3431
rect 11060 3392 11112 3398
rect 11060 3334 11112 3340
rect 11058 3224 11114 3233
rect 11058 3159 11114 3168
rect 11072 3126 11100 3159
rect 11060 3120 11112 3126
rect 11060 3062 11112 3068
rect 10244 734 10456 762
rect 10506 0 10562 800
rect 10966 0 11022 800
rect 11164 762 11192 11494
rect 11348 11393 11376 11630
rect 11334 11384 11390 11393
rect 11334 11319 11336 11328
rect 11388 11319 11390 11328
rect 11336 11290 11388 11296
rect 11244 11076 11296 11082
rect 11244 11018 11296 11024
rect 11256 4162 11284 11018
rect 11346 10908 11654 10917
rect 11346 10906 11352 10908
rect 11408 10906 11432 10908
rect 11488 10906 11512 10908
rect 11568 10906 11592 10908
rect 11648 10906 11654 10908
rect 11408 10854 11410 10906
rect 11590 10854 11592 10906
rect 11346 10852 11352 10854
rect 11408 10852 11432 10854
rect 11488 10852 11512 10854
rect 11568 10852 11592 10854
rect 11648 10852 11654 10854
rect 11346 10843 11654 10852
rect 11716 10713 11744 11766
rect 11808 11626 11836 12022
rect 11980 11824 12032 11830
rect 11980 11766 12032 11772
rect 11888 11756 11940 11762
rect 11888 11698 11940 11704
rect 11796 11620 11848 11626
rect 11796 11562 11848 11568
rect 11702 10704 11758 10713
rect 11702 10639 11758 10648
rect 11704 10600 11756 10606
rect 11704 10542 11756 10548
rect 11612 10464 11664 10470
rect 11612 10406 11664 10412
rect 11624 10266 11652 10406
rect 11612 10260 11664 10266
rect 11612 10202 11664 10208
rect 11346 9820 11654 9829
rect 11346 9818 11352 9820
rect 11408 9818 11432 9820
rect 11488 9818 11512 9820
rect 11568 9818 11592 9820
rect 11648 9818 11654 9820
rect 11408 9766 11410 9818
rect 11590 9766 11592 9818
rect 11346 9764 11352 9766
rect 11408 9764 11432 9766
rect 11488 9764 11512 9766
rect 11568 9764 11592 9766
rect 11648 9764 11654 9766
rect 11346 9755 11654 9764
rect 11612 9376 11664 9382
rect 11612 9318 11664 9324
rect 11518 9208 11574 9217
rect 11518 9143 11574 9152
rect 11532 8945 11560 9143
rect 11624 8956 11652 9318
rect 11716 9024 11744 10542
rect 11808 9178 11836 11562
rect 11900 9450 11928 11698
rect 11992 11014 12020 11766
rect 12084 11665 12112 12786
rect 12070 11656 12126 11665
rect 12070 11591 12126 11600
rect 12072 11552 12124 11558
rect 12072 11494 12124 11500
rect 11980 11008 12032 11014
rect 11980 10950 12032 10956
rect 12084 10146 12112 11494
rect 12176 10198 12204 22200
rect 12532 20324 12584 20330
rect 12532 20266 12584 20272
rect 12440 19780 12492 19786
rect 12440 19722 12492 19728
rect 12452 19514 12480 19722
rect 12440 19508 12492 19514
rect 12440 19450 12492 19456
rect 12348 17604 12400 17610
rect 12348 17546 12400 17552
rect 12256 16652 12308 16658
rect 12256 16594 12308 16600
rect 12268 13818 12296 16594
rect 12360 15978 12388 17546
rect 12348 15972 12400 15978
rect 12348 15914 12400 15920
rect 12452 15609 12480 19450
rect 12544 19446 12572 20266
rect 12532 19440 12584 19446
rect 12532 19382 12584 19388
rect 12532 18624 12584 18630
rect 12532 18566 12584 18572
rect 12544 17921 12572 18566
rect 12530 17912 12586 17921
rect 12530 17847 12586 17856
rect 12532 17672 12584 17678
rect 12532 17614 12584 17620
rect 12544 17542 12572 17614
rect 12532 17536 12584 17542
rect 12532 17478 12584 17484
rect 12530 16960 12586 16969
rect 12530 16895 12586 16904
rect 12544 16794 12572 16895
rect 12532 16788 12584 16794
rect 12532 16730 12584 16736
rect 12532 16108 12584 16114
rect 12532 16050 12584 16056
rect 12544 16017 12572 16050
rect 12530 16008 12586 16017
rect 12530 15943 12586 15952
rect 12438 15600 12494 15609
rect 12438 15535 12494 15544
rect 12532 15360 12584 15366
rect 12532 15302 12584 15308
rect 12544 14906 12572 15302
rect 12636 15162 12664 22200
rect 13096 20482 13124 22200
rect 12912 20454 13124 20482
rect 12912 19854 12940 20454
rect 13556 20058 13584 22200
rect 14016 20534 14044 22200
rect 14004 20528 14056 20534
rect 14004 20470 14056 20476
rect 14476 20398 14504 22200
rect 14464 20392 14516 20398
rect 14464 20334 14516 20340
rect 13945 20156 14253 20165
rect 13945 20154 13951 20156
rect 14007 20154 14031 20156
rect 14087 20154 14111 20156
rect 14167 20154 14191 20156
rect 14247 20154 14253 20156
rect 14007 20102 14009 20154
rect 14189 20102 14191 20154
rect 13945 20100 13951 20102
rect 14007 20100 14031 20102
rect 14087 20100 14111 20102
rect 14167 20100 14191 20102
rect 14247 20100 14253 20102
rect 13945 20091 14253 20100
rect 13544 20052 13596 20058
rect 13544 19994 13596 20000
rect 14568 19938 14596 22222
rect 14844 22114 14872 22222
rect 14922 22200 14978 23000
rect 15382 22200 15438 23000
rect 15842 22200 15898 23000
rect 16302 22200 16358 23000
rect 16762 22200 16818 23000
rect 16868 22222 17080 22250
rect 14936 22114 14964 22200
rect 14844 22086 14964 22114
rect 14292 19910 14596 19938
rect 12900 19848 12952 19854
rect 12900 19790 12952 19796
rect 13084 19848 13136 19854
rect 13084 19790 13136 19796
rect 13636 19848 13688 19854
rect 13636 19790 13688 19796
rect 13096 19718 13124 19790
rect 13084 19712 13136 19718
rect 13084 19654 13136 19660
rect 12808 19440 12860 19446
rect 12808 19382 12860 19388
rect 12714 19000 12770 19009
rect 12714 18935 12770 18944
rect 12624 15156 12676 15162
rect 12624 15098 12676 15104
rect 12544 14878 12664 14906
rect 12532 14816 12584 14822
rect 12532 14758 12584 14764
rect 12544 14618 12572 14758
rect 12532 14612 12584 14618
rect 12532 14554 12584 14560
rect 12532 14408 12584 14414
rect 12452 14368 12532 14396
rect 12348 14272 12400 14278
rect 12348 14214 12400 14220
rect 12360 14006 12388 14214
rect 12348 14000 12400 14006
rect 12348 13942 12400 13948
rect 12268 13790 12388 13818
rect 12256 13728 12308 13734
rect 12256 13670 12308 13676
rect 12268 12646 12296 13670
rect 12256 12640 12308 12646
rect 12360 12617 12388 13790
rect 12452 13462 12480 14368
rect 12532 14350 12584 14356
rect 12532 14068 12584 14074
rect 12532 14010 12584 14016
rect 12440 13456 12492 13462
rect 12440 13398 12492 13404
rect 12544 13326 12572 14010
rect 12636 13376 12664 14878
rect 12728 14278 12756 18935
rect 12820 18057 12848 19382
rect 13096 19378 13124 19654
rect 13084 19372 13136 19378
rect 13136 19320 13216 19334
rect 13084 19314 13216 19320
rect 13096 19306 13216 19314
rect 13096 19249 13124 19306
rect 12900 19168 12952 19174
rect 12900 19110 12952 19116
rect 12912 18970 12940 19110
rect 12900 18964 12952 18970
rect 12900 18906 12952 18912
rect 13188 18766 13216 19306
rect 13360 18828 13412 18834
rect 13360 18770 13412 18776
rect 13176 18760 13228 18766
rect 13176 18702 13228 18708
rect 13372 18358 13400 18770
rect 13544 18624 13596 18630
rect 13544 18566 13596 18572
rect 13360 18352 13412 18358
rect 13360 18294 13412 18300
rect 13084 18080 13136 18086
rect 12806 18048 12862 18057
rect 12806 17983 12862 17992
rect 13082 18048 13084 18057
rect 13176 18080 13228 18086
rect 13136 18048 13138 18057
rect 13176 18022 13228 18028
rect 13082 17983 13138 17992
rect 12808 17740 12860 17746
rect 12808 17682 12860 17688
rect 12820 17270 12848 17682
rect 12992 17536 13044 17542
rect 12912 17496 12992 17524
rect 12808 17264 12860 17270
rect 12912 17241 12940 17496
rect 12992 17478 13044 17484
rect 13188 17338 13216 18022
rect 13452 17876 13504 17882
rect 13452 17818 13504 17824
rect 13464 17762 13492 17818
rect 13556 17814 13584 18566
rect 13280 17746 13492 17762
rect 13544 17808 13596 17814
rect 13544 17750 13596 17756
rect 13268 17740 13492 17746
rect 13320 17734 13492 17740
rect 13268 17682 13320 17688
rect 13176 17332 13228 17338
rect 13176 17274 13228 17280
rect 13360 17332 13412 17338
rect 13360 17274 13412 17280
rect 12808 17206 12860 17212
rect 12898 17232 12954 17241
rect 12898 17167 12954 17176
rect 12912 15094 12940 17167
rect 13372 16969 13400 17274
rect 13358 16960 13414 16969
rect 13358 16895 13414 16904
rect 13358 16824 13414 16833
rect 13358 16759 13414 16768
rect 13372 16590 13400 16759
rect 13360 16584 13412 16590
rect 13360 16526 13412 16532
rect 12992 16516 13044 16522
rect 12992 16458 13044 16464
rect 12900 15088 12952 15094
rect 12900 15030 12952 15036
rect 13004 14770 13032 16458
rect 13544 15088 13596 15094
rect 13544 15030 13596 15036
rect 13360 15020 13412 15026
rect 13360 14962 13412 14968
rect 12912 14742 13032 14770
rect 12716 14272 12768 14278
rect 12716 14214 12768 14220
rect 12636 13348 12848 13376
rect 12532 13320 12584 13326
rect 12532 13262 12584 13268
rect 12544 12646 12572 13262
rect 12820 13258 12848 13348
rect 12808 13252 12860 13258
rect 12808 13194 12860 13200
rect 12532 12640 12584 12646
rect 12256 12582 12308 12588
rect 12346 12608 12402 12617
rect 12532 12582 12584 12588
rect 12716 12640 12768 12646
rect 12716 12582 12768 12588
rect 12346 12543 12402 12552
rect 12544 12306 12572 12582
rect 12728 12434 12756 12582
rect 12636 12406 12756 12434
rect 12532 12300 12584 12306
rect 12532 12242 12584 12248
rect 12636 12170 12664 12406
rect 12256 12164 12308 12170
rect 12624 12164 12676 12170
rect 12308 12124 12388 12152
rect 12256 12106 12308 12112
rect 12256 11688 12308 11694
rect 12256 11630 12308 11636
rect 12268 11257 12296 11630
rect 12254 11248 12310 11257
rect 12254 11183 12310 11192
rect 12256 11076 12308 11082
rect 12256 11018 12308 11024
rect 11992 10118 12112 10146
rect 12164 10192 12216 10198
rect 12164 10134 12216 10140
rect 11888 9444 11940 9450
rect 11888 9386 11940 9392
rect 11796 9172 11848 9178
rect 11796 9114 11848 9120
rect 11716 8996 11928 9024
rect 11334 8936 11390 8945
rect 11334 8871 11390 8880
rect 11518 8936 11574 8945
rect 11624 8928 11744 8956
rect 11518 8871 11574 8880
rect 11348 8838 11376 8871
rect 11336 8832 11388 8838
rect 11336 8774 11388 8780
rect 11346 8732 11654 8741
rect 11346 8730 11352 8732
rect 11408 8730 11432 8732
rect 11488 8730 11512 8732
rect 11568 8730 11592 8732
rect 11648 8730 11654 8732
rect 11408 8678 11410 8730
rect 11590 8678 11592 8730
rect 11346 8676 11352 8678
rect 11408 8676 11432 8678
rect 11488 8676 11512 8678
rect 11568 8676 11592 8678
rect 11648 8676 11654 8678
rect 11346 8667 11654 8676
rect 11334 8256 11390 8265
rect 11334 8191 11390 8200
rect 11348 7993 11376 8191
rect 11334 7984 11390 7993
rect 11334 7919 11336 7928
rect 11388 7919 11390 7928
rect 11336 7890 11388 7896
rect 11346 7644 11654 7653
rect 11346 7642 11352 7644
rect 11408 7642 11432 7644
rect 11488 7642 11512 7644
rect 11568 7642 11592 7644
rect 11648 7642 11654 7644
rect 11408 7590 11410 7642
rect 11590 7590 11592 7642
rect 11346 7588 11352 7590
rect 11408 7588 11432 7590
rect 11488 7588 11512 7590
rect 11568 7588 11592 7590
rect 11648 7588 11654 7590
rect 11346 7579 11654 7588
rect 11716 7002 11744 8928
rect 11796 8832 11848 8838
rect 11796 8774 11848 8780
rect 11704 6996 11756 7002
rect 11704 6938 11756 6944
rect 11808 6730 11836 8774
rect 11796 6724 11848 6730
rect 11796 6666 11848 6672
rect 11346 6556 11654 6565
rect 11346 6554 11352 6556
rect 11408 6554 11432 6556
rect 11488 6554 11512 6556
rect 11568 6554 11592 6556
rect 11648 6554 11654 6556
rect 11408 6502 11410 6554
rect 11590 6502 11592 6554
rect 11346 6500 11352 6502
rect 11408 6500 11432 6502
rect 11488 6500 11512 6502
rect 11568 6500 11592 6502
rect 11648 6500 11654 6502
rect 11346 6491 11654 6500
rect 11336 6384 11388 6390
rect 11336 6326 11388 6332
rect 11518 6352 11574 6361
rect 11348 5953 11376 6326
rect 11518 6287 11574 6296
rect 11532 6254 11560 6287
rect 11520 6248 11572 6254
rect 11520 6190 11572 6196
rect 11796 6248 11848 6254
rect 11796 6190 11848 6196
rect 11532 5953 11560 6190
rect 11334 5944 11390 5953
rect 11334 5879 11390 5888
rect 11518 5944 11574 5953
rect 11518 5879 11574 5888
rect 11702 5808 11758 5817
rect 11702 5743 11758 5752
rect 11716 5574 11744 5743
rect 11808 5710 11836 6190
rect 11796 5704 11848 5710
rect 11796 5646 11848 5652
rect 11704 5568 11756 5574
rect 11704 5510 11756 5516
rect 11346 5468 11654 5477
rect 11346 5466 11352 5468
rect 11408 5466 11432 5468
rect 11488 5466 11512 5468
rect 11568 5466 11592 5468
rect 11648 5466 11654 5468
rect 11408 5414 11410 5466
rect 11590 5414 11592 5466
rect 11346 5412 11352 5414
rect 11408 5412 11432 5414
rect 11488 5412 11512 5414
rect 11568 5412 11592 5414
rect 11648 5412 11654 5414
rect 11346 5403 11654 5412
rect 11794 5264 11850 5273
rect 11794 5199 11850 5208
rect 11808 5166 11836 5199
rect 11796 5160 11848 5166
rect 11796 5102 11848 5108
rect 11900 4842 11928 8996
rect 11992 5250 12020 10118
rect 12072 10056 12124 10062
rect 12268 10044 12296 11018
rect 12360 10305 12388 12124
rect 12624 12106 12676 12112
rect 12532 12096 12584 12102
rect 12532 12038 12584 12044
rect 12440 11348 12492 11354
rect 12440 11290 12492 11296
rect 12452 11014 12480 11290
rect 12544 11218 12572 12038
rect 12532 11212 12584 11218
rect 12532 11154 12584 11160
rect 12440 11008 12492 11014
rect 12440 10950 12492 10956
rect 12452 10742 12480 10950
rect 12440 10736 12492 10742
rect 12440 10678 12492 10684
rect 12346 10296 12402 10305
rect 12346 10231 12402 10240
rect 12348 10192 12400 10198
rect 12348 10134 12400 10140
rect 12072 9998 12124 10004
rect 12176 10016 12296 10044
rect 12084 9722 12112 9998
rect 12072 9716 12124 9722
rect 12072 9658 12124 9664
rect 12176 9382 12204 10016
rect 12360 9704 12388 10134
rect 12452 10062 12480 10678
rect 12532 10260 12584 10266
rect 12532 10202 12584 10208
rect 12440 10056 12492 10062
rect 12440 9998 12492 10004
rect 12360 9676 12480 9704
rect 12452 9586 12480 9676
rect 12440 9580 12492 9586
rect 12440 9522 12492 9528
rect 12256 9444 12308 9450
rect 12256 9386 12308 9392
rect 12164 9376 12216 9382
rect 12164 9318 12216 9324
rect 12268 8072 12296 9386
rect 12452 8838 12480 9522
rect 12440 8832 12492 8838
rect 12440 8774 12492 8780
rect 12544 8401 12572 10202
rect 12530 8392 12586 8401
rect 12530 8327 12586 8336
rect 12544 8294 12572 8327
rect 12532 8288 12584 8294
rect 12532 8230 12584 8236
rect 12636 8090 12664 12106
rect 12716 11756 12768 11762
rect 12716 11698 12768 11704
rect 12728 11082 12756 11698
rect 12820 11150 12848 13194
rect 12808 11144 12860 11150
rect 12808 11086 12860 11092
rect 12716 11076 12768 11082
rect 12716 11018 12768 11024
rect 12808 10736 12860 10742
rect 12808 10678 12860 10684
rect 12820 10305 12848 10678
rect 12806 10296 12862 10305
rect 12806 10231 12862 10240
rect 12716 9920 12768 9926
rect 12716 9862 12768 9868
rect 12728 9586 12756 9862
rect 12716 9580 12768 9586
rect 12716 9522 12768 9528
rect 12624 8084 12676 8090
rect 12268 8044 12480 8072
rect 12452 7868 12480 8044
rect 12624 8026 12676 8032
rect 12530 7984 12586 7993
rect 12530 7919 12532 7928
rect 12584 7919 12586 7928
rect 12532 7890 12584 7896
rect 12360 7840 12480 7868
rect 12072 7744 12124 7750
rect 12072 7686 12124 7692
rect 12084 7546 12112 7686
rect 12072 7540 12124 7546
rect 12072 7482 12124 7488
rect 12256 7268 12308 7274
rect 12256 7210 12308 7216
rect 12070 7032 12126 7041
rect 12070 6967 12126 6976
rect 12084 5817 12112 6967
rect 12268 6934 12296 7210
rect 12256 6928 12308 6934
rect 12256 6870 12308 6876
rect 12164 6180 12216 6186
rect 12164 6122 12216 6128
rect 12070 5808 12126 5817
rect 12070 5743 12126 5752
rect 11992 5234 12112 5250
rect 11992 5228 12124 5234
rect 11992 5222 12072 5228
rect 12072 5170 12124 5176
rect 12176 5098 12204 6122
rect 12256 5228 12308 5234
rect 12256 5170 12308 5176
rect 12164 5092 12216 5098
rect 12164 5034 12216 5040
rect 11900 4814 12020 4842
rect 12268 4826 12296 5170
rect 11888 4752 11940 4758
rect 11888 4694 11940 4700
rect 11346 4380 11654 4389
rect 11346 4378 11352 4380
rect 11408 4378 11432 4380
rect 11488 4378 11512 4380
rect 11568 4378 11592 4380
rect 11648 4378 11654 4380
rect 11408 4326 11410 4378
rect 11590 4326 11592 4378
rect 11346 4324 11352 4326
rect 11408 4324 11432 4326
rect 11488 4324 11512 4326
rect 11568 4324 11592 4326
rect 11648 4324 11654 4326
rect 11346 4315 11654 4324
rect 11900 4282 11928 4694
rect 11888 4276 11940 4282
rect 11888 4218 11940 4224
rect 11256 4134 11928 4162
rect 11428 4072 11480 4078
rect 11428 4014 11480 4020
rect 11242 3632 11298 3641
rect 11242 3567 11244 3576
rect 11296 3567 11298 3576
rect 11244 3538 11296 3544
rect 11440 3398 11468 4014
rect 11428 3392 11480 3398
rect 11428 3334 11480 3340
rect 11704 3392 11756 3398
rect 11704 3334 11756 3340
rect 11346 3292 11654 3301
rect 11346 3290 11352 3292
rect 11408 3290 11432 3292
rect 11488 3290 11512 3292
rect 11568 3290 11592 3292
rect 11648 3290 11654 3292
rect 11408 3238 11410 3290
rect 11590 3238 11592 3290
rect 11346 3236 11352 3238
rect 11408 3236 11432 3238
rect 11488 3236 11512 3238
rect 11568 3236 11592 3238
rect 11648 3236 11654 3238
rect 11346 3227 11654 3236
rect 11716 3194 11744 3334
rect 11704 3188 11756 3194
rect 11704 3130 11756 3136
rect 11796 3052 11848 3058
rect 11796 2994 11848 3000
rect 11808 2650 11836 2994
rect 11796 2644 11848 2650
rect 11796 2586 11848 2592
rect 11346 2204 11654 2213
rect 11346 2202 11352 2204
rect 11408 2202 11432 2204
rect 11488 2202 11512 2204
rect 11568 2202 11592 2204
rect 11648 2202 11654 2204
rect 11408 2150 11410 2202
rect 11590 2150 11592 2202
rect 11346 2148 11352 2150
rect 11408 2148 11432 2150
rect 11488 2148 11512 2150
rect 11568 2148 11592 2150
rect 11648 2148 11654 2150
rect 11346 2139 11654 2148
rect 11348 870 11468 898
rect 11348 762 11376 870
rect 11440 800 11468 870
rect 11900 800 11928 4134
rect 11992 3194 12020 4814
rect 12256 4820 12308 4826
rect 12256 4762 12308 4768
rect 12268 4554 12296 4762
rect 12256 4548 12308 4554
rect 12256 4490 12308 4496
rect 12072 4276 12124 4282
rect 12072 4218 12124 4224
rect 12084 4078 12112 4218
rect 12072 4072 12124 4078
rect 12072 4014 12124 4020
rect 12084 3670 12112 4014
rect 12072 3664 12124 3670
rect 12072 3606 12124 3612
rect 11980 3188 12032 3194
rect 11980 3130 12032 3136
rect 11992 3058 12020 3130
rect 11980 3052 12032 3058
rect 11980 2994 12032 3000
rect 12360 800 12388 7840
rect 12440 7744 12492 7750
rect 12440 7686 12492 7692
rect 12452 6662 12480 7686
rect 12440 6656 12492 6662
rect 12440 6598 12492 6604
rect 12624 6452 12676 6458
rect 12624 6394 12676 6400
rect 12440 6248 12492 6254
rect 12440 6190 12492 6196
rect 12532 6248 12584 6254
rect 12532 6190 12584 6196
rect 12452 5710 12480 6190
rect 12544 6118 12572 6190
rect 12532 6112 12584 6118
rect 12532 6054 12584 6060
rect 12636 5953 12664 6394
rect 12622 5944 12678 5953
rect 12622 5879 12678 5888
rect 12532 5772 12584 5778
rect 12532 5714 12584 5720
rect 12440 5704 12492 5710
rect 12440 5646 12492 5652
rect 12440 5568 12492 5574
rect 12438 5536 12440 5545
rect 12492 5536 12494 5545
rect 12438 5471 12494 5480
rect 12544 5302 12572 5714
rect 12532 5296 12584 5302
rect 12532 5238 12584 5244
rect 12636 5166 12664 5879
rect 12532 5160 12584 5166
rect 12532 5102 12584 5108
rect 12624 5160 12676 5166
rect 12624 5102 12676 5108
rect 12544 5030 12572 5102
rect 12532 5024 12584 5030
rect 12530 4992 12532 5001
rect 12584 4992 12586 5001
rect 12530 4927 12586 4936
rect 12636 4622 12664 5102
rect 12624 4616 12676 4622
rect 12624 4558 12676 4564
rect 12728 4185 12756 9522
rect 12808 8288 12860 8294
rect 12808 8230 12860 8236
rect 12820 5778 12848 8230
rect 12912 7274 12940 14742
rect 13176 14272 13228 14278
rect 13176 14214 13228 14220
rect 12992 12096 13044 12102
rect 12992 12038 13044 12044
rect 13004 10470 13032 12038
rect 13188 11370 13216 14214
rect 13372 13870 13400 14962
rect 13452 14884 13504 14890
rect 13452 14826 13504 14832
rect 13464 14346 13492 14826
rect 13556 14532 13584 15030
rect 13648 14822 13676 19790
rect 13820 19372 13872 19378
rect 13820 19314 13872 19320
rect 13728 18760 13780 18766
rect 13728 18702 13780 18708
rect 13740 18290 13768 18702
rect 13728 18284 13780 18290
rect 13728 18226 13780 18232
rect 13740 17746 13768 18226
rect 13728 17740 13780 17746
rect 13728 17682 13780 17688
rect 13832 16794 13860 19314
rect 13945 19068 14253 19077
rect 13945 19066 13951 19068
rect 14007 19066 14031 19068
rect 14087 19066 14111 19068
rect 14167 19066 14191 19068
rect 14247 19066 14253 19068
rect 14007 19014 14009 19066
rect 14189 19014 14191 19066
rect 13945 19012 13951 19014
rect 14007 19012 14031 19014
rect 14087 19012 14111 19014
rect 14167 19012 14191 19014
rect 14247 19012 14253 19014
rect 13945 19003 14253 19012
rect 14188 18828 14240 18834
rect 14188 18770 14240 18776
rect 14200 18426 14228 18770
rect 14292 18698 14320 19910
rect 14832 19848 14884 19854
rect 14832 19790 14884 19796
rect 14372 19780 14424 19786
rect 14372 19722 14424 19728
rect 14464 19780 14516 19786
rect 14464 19722 14516 19728
rect 14384 18698 14412 19722
rect 14280 18692 14332 18698
rect 14280 18634 14332 18640
rect 14372 18692 14424 18698
rect 14372 18634 14424 18640
rect 14188 18420 14240 18426
rect 14188 18362 14240 18368
rect 14372 18352 14424 18358
rect 14372 18294 14424 18300
rect 14188 18284 14240 18290
rect 14188 18226 14240 18232
rect 14200 18170 14228 18226
rect 14200 18142 14320 18170
rect 13945 17980 14253 17989
rect 13945 17978 13951 17980
rect 14007 17978 14031 17980
rect 14087 17978 14111 17980
rect 14167 17978 14191 17980
rect 14247 17978 14253 17980
rect 14007 17926 14009 17978
rect 14189 17926 14191 17978
rect 13945 17924 13951 17926
rect 14007 17924 14031 17926
rect 14087 17924 14111 17926
rect 14167 17924 14191 17926
rect 14247 17924 14253 17926
rect 13945 17915 14253 17924
rect 13945 16892 14253 16901
rect 13945 16890 13951 16892
rect 14007 16890 14031 16892
rect 14087 16890 14111 16892
rect 14167 16890 14191 16892
rect 14247 16890 14253 16892
rect 14007 16838 14009 16890
rect 14189 16838 14191 16890
rect 13945 16836 13951 16838
rect 14007 16836 14031 16838
rect 14087 16836 14111 16838
rect 14167 16836 14191 16838
rect 14247 16836 14253 16838
rect 13945 16827 14253 16836
rect 13820 16788 13872 16794
rect 13820 16730 13872 16736
rect 13728 16516 13780 16522
rect 13728 16458 13780 16464
rect 13740 15910 13768 16458
rect 13832 16454 13860 16730
rect 13820 16448 13872 16454
rect 13820 16390 13872 16396
rect 13728 15904 13780 15910
rect 13728 15846 13780 15852
rect 13740 15502 13768 15846
rect 13945 15804 14253 15813
rect 13945 15802 13951 15804
rect 14007 15802 14031 15804
rect 14087 15802 14111 15804
rect 14167 15802 14191 15804
rect 14247 15802 14253 15804
rect 14007 15750 14009 15802
rect 14189 15750 14191 15802
rect 13945 15748 13951 15750
rect 14007 15748 14031 15750
rect 14087 15748 14111 15750
rect 14167 15748 14191 15750
rect 14247 15748 14253 15750
rect 13945 15739 14253 15748
rect 13728 15496 13780 15502
rect 13728 15438 13780 15444
rect 13740 15366 13768 15438
rect 13728 15360 13780 15366
rect 13728 15302 13780 15308
rect 13820 15360 13872 15366
rect 13820 15302 13872 15308
rect 13740 14958 13768 15302
rect 13728 14952 13780 14958
rect 13728 14894 13780 14900
rect 13636 14816 13688 14822
rect 13636 14758 13688 14764
rect 13636 14544 13688 14550
rect 13556 14504 13636 14532
rect 13636 14486 13688 14492
rect 13740 14482 13768 14894
rect 13728 14476 13780 14482
rect 13728 14418 13780 14424
rect 13452 14340 13504 14346
rect 13452 14282 13504 14288
rect 13544 14340 13596 14346
rect 13544 14282 13596 14288
rect 13556 13938 13584 14282
rect 13636 14272 13688 14278
rect 13740 14260 13768 14418
rect 13832 14414 13860 15302
rect 14292 15065 14320 18142
rect 14384 17746 14412 18294
rect 14372 17740 14424 17746
rect 14372 17682 14424 17688
rect 14372 17196 14424 17202
rect 14372 17138 14424 17144
rect 14278 15056 14334 15065
rect 14278 14991 14334 15000
rect 13945 14716 14253 14725
rect 13945 14714 13951 14716
rect 14007 14714 14031 14716
rect 14087 14714 14111 14716
rect 14167 14714 14191 14716
rect 14247 14714 14253 14716
rect 14007 14662 14009 14714
rect 14189 14662 14191 14714
rect 13945 14660 13951 14662
rect 14007 14660 14031 14662
rect 14087 14660 14111 14662
rect 14167 14660 14191 14662
rect 14247 14660 14253 14662
rect 13945 14651 14253 14660
rect 13820 14408 13872 14414
rect 13820 14350 13872 14356
rect 13688 14232 13768 14260
rect 13636 14214 13688 14220
rect 13648 14074 13676 14214
rect 13636 14068 13688 14074
rect 13636 14010 13688 14016
rect 13544 13932 13596 13938
rect 13544 13874 13596 13880
rect 13360 13864 13412 13870
rect 13360 13806 13412 13812
rect 13372 12434 13400 13806
rect 13556 13734 13584 13874
rect 13544 13728 13596 13734
rect 13544 13670 13596 13676
rect 14280 13728 14332 13734
rect 14280 13670 14332 13676
rect 13945 13628 14253 13637
rect 13945 13626 13951 13628
rect 14007 13626 14031 13628
rect 14087 13626 14111 13628
rect 14167 13626 14191 13628
rect 14247 13626 14253 13628
rect 14007 13574 14009 13626
rect 14189 13574 14191 13626
rect 13945 13572 13951 13574
rect 14007 13572 14031 13574
rect 14087 13572 14111 13574
rect 14167 13572 14191 13574
rect 14247 13572 14253 13574
rect 13945 13563 14253 13572
rect 13820 13524 13872 13530
rect 13820 13466 13872 13472
rect 13096 11342 13216 11370
rect 13280 12406 13400 12434
rect 12992 10464 13044 10470
rect 12992 10406 13044 10412
rect 13096 8922 13124 11342
rect 13176 11280 13228 11286
rect 13176 11222 13228 11228
rect 13004 8894 13124 8922
rect 13004 8072 13032 8894
rect 13188 8537 13216 11222
rect 13280 9353 13308 12406
rect 13832 11898 13860 13466
rect 14292 13190 14320 13670
rect 14384 13530 14412 17138
rect 14372 13524 14424 13530
rect 14372 13466 14424 13472
rect 14096 13184 14148 13190
rect 14096 13126 14148 13132
rect 14280 13184 14332 13190
rect 14280 13126 14332 13132
rect 14108 12986 14136 13126
rect 14096 12980 14148 12986
rect 14096 12922 14148 12928
rect 14292 12918 14320 13126
rect 14280 12912 14332 12918
rect 14280 12854 14332 12860
rect 14292 12782 14320 12854
rect 14372 12844 14424 12850
rect 14372 12786 14424 12792
rect 14280 12776 14332 12782
rect 14280 12718 14332 12724
rect 13945 12540 14253 12549
rect 13945 12538 13951 12540
rect 14007 12538 14031 12540
rect 14087 12538 14111 12540
rect 14167 12538 14191 12540
rect 14247 12538 14253 12540
rect 14007 12486 14009 12538
rect 14189 12486 14191 12538
rect 13945 12484 13951 12486
rect 14007 12484 14031 12486
rect 14087 12484 14111 12486
rect 14167 12484 14191 12486
rect 14247 12484 14253 12486
rect 13945 12475 14253 12484
rect 13912 12232 13964 12238
rect 13912 12174 13964 12180
rect 13924 12102 13952 12174
rect 13912 12096 13964 12102
rect 13912 12038 13964 12044
rect 14188 12096 14240 12102
rect 14292 12084 14320 12718
rect 14384 12238 14412 12786
rect 14372 12232 14424 12238
rect 14372 12174 14424 12180
rect 14240 12056 14320 12084
rect 14188 12038 14240 12044
rect 13820 11892 13872 11898
rect 13820 11834 13872 11840
rect 13728 11552 13780 11558
rect 13924 11540 13952 12038
rect 14200 11694 14228 12038
rect 14188 11688 14240 11694
rect 14188 11630 14240 11636
rect 13728 11494 13780 11500
rect 13832 11512 13952 11540
rect 13544 11280 13596 11286
rect 13544 11222 13596 11228
rect 13450 10296 13506 10305
rect 13450 10231 13506 10240
rect 13464 10198 13492 10231
rect 13452 10192 13504 10198
rect 13452 10134 13504 10140
rect 13360 9988 13412 9994
rect 13360 9930 13412 9936
rect 13372 9674 13400 9930
rect 13556 9674 13584 11222
rect 13740 10742 13768 11494
rect 13728 10736 13780 10742
rect 13728 10678 13780 10684
rect 13636 10668 13688 10674
rect 13636 10610 13688 10616
rect 13648 9722 13676 10610
rect 13728 10464 13780 10470
rect 13728 10406 13780 10412
rect 13740 10266 13768 10406
rect 13728 10260 13780 10266
rect 13728 10202 13780 10208
rect 13728 10124 13780 10130
rect 13728 10066 13780 10072
rect 13372 9646 13584 9674
rect 13636 9716 13688 9722
rect 13636 9658 13688 9664
rect 13266 9344 13322 9353
rect 13266 9279 13322 9288
rect 13268 8900 13320 8906
rect 13268 8842 13320 8848
rect 13174 8528 13230 8537
rect 13174 8463 13230 8472
rect 13280 8362 13308 8842
rect 13268 8356 13320 8362
rect 13188 8316 13268 8344
rect 13004 8044 13124 8072
rect 12992 7948 13044 7954
rect 12992 7890 13044 7896
rect 13004 7342 13032 7890
rect 12992 7336 13044 7342
rect 12992 7278 13044 7284
rect 12900 7268 12952 7274
rect 12900 7210 12952 7216
rect 13004 6934 13032 7278
rect 12992 6928 13044 6934
rect 12992 6870 13044 6876
rect 12808 5772 12860 5778
rect 12808 5714 12860 5720
rect 12808 5568 12860 5574
rect 12808 5510 12860 5516
rect 12900 5568 12952 5574
rect 12900 5510 12952 5516
rect 12820 5370 12848 5510
rect 12808 5364 12860 5370
rect 12808 5306 12860 5312
rect 12912 4690 12940 5510
rect 13096 5137 13124 8044
rect 13082 5128 13138 5137
rect 13082 5063 13138 5072
rect 13096 4758 13124 5063
rect 13084 4752 13136 4758
rect 13084 4694 13136 4700
rect 12900 4684 12952 4690
rect 12900 4626 12952 4632
rect 13188 4486 13216 8316
rect 13268 8298 13320 8304
rect 13268 6452 13320 6458
rect 13268 6394 13320 6400
rect 13280 5914 13308 6394
rect 13268 5908 13320 5914
rect 13268 5850 13320 5856
rect 13372 5352 13400 9646
rect 13636 9580 13688 9586
rect 13636 9522 13688 9528
rect 13648 9178 13676 9522
rect 13636 9172 13688 9178
rect 13636 9114 13688 9120
rect 13542 8936 13598 8945
rect 13542 8871 13544 8880
rect 13596 8871 13598 8880
rect 13544 8842 13596 8848
rect 13542 8528 13598 8537
rect 13542 8463 13598 8472
rect 13452 8288 13504 8294
rect 13452 8230 13504 8236
rect 13464 5370 13492 8230
rect 13280 5324 13400 5352
rect 13452 5364 13504 5370
rect 13176 4480 13228 4486
rect 13176 4422 13228 4428
rect 13280 4282 13308 5324
rect 13452 5306 13504 5312
rect 13464 5250 13492 5306
rect 13556 5273 13584 8463
rect 13740 8294 13768 10066
rect 13832 9625 13860 11512
rect 13945 11452 14253 11461
rect 13945 11450 13951 11452
rect 14007 11450 14031 11452
rect 14087 11450 14111 11452
rect 14167 11450 14191 11452
rect 14247 11450 14253 11452
rect 14007 11398 14009 11450
rect 14189 11398 14191 11450
rect 13945 11396 13951 11398
rect 14007 11396 14031 11398
rect 14087 11396 14111 11398
rect 14167 11396 14191 11398
rect 14247 11396 14253 11398
rect 13945 11387 14253 11396
rect 14280 11348 14332 11354
rect 14280 11290 14332 11296
rect 13945 10364 14253 10373
rect 13945 10362 13951 10364
rect 14007 10362 14031 10364
rect 14087 10362 14111 10364
rect 14167 10362 14191 10364
rect 14247 10362 14253 10364
rect 14007 10310 14009 10362
rect 14189 10310 14191 10362
rect 13945 10308 13951 10310
rect 14007 10308 14031 10310
rect 14087 10308 14111 10310
rect 14167 10308 14191 10310
rect 14247 10308 14253 10310
rect 13945 10299 14253 10308
rect 13912 9920 13964 9926
rect 13912 9862 13964 9868
rect 13818 9616 13874 9625
rect 13818 9551 13874 9560
rect 13820 9512 13872 9518
rect 13820 9454 13872 9460
rect 13832 9042 13860 9454
rect 13924 9382 13952 9862
rect 14002 9480 14058 9489
rect 14002 9415 14004 9424
rect 14056 9415 14058 9424
rect 14004 9386 14056 9392
rect 13912 9376 13964 9382
rect 13912 9318 13964 9324
rect 13945 9276 14253 9285
rect 13945 9274 13951 9276
rect 14007 9274 14031 9276
rect 14087 9274 14111 9276
rect 14167 9274 14191 9276
rect 14247 9274 14253 9276
rect 14007 9222 14009 9274
rect 14189 9222 14191 9274
rect 13945 9220 13951 9222
rect 14007 9220 14031 9222
rect 14087 9220 14111 9222
rect 14167 9220 14191 9222
rect 14247 9220 14253 9222
rect 13945 9211 14253 9220
rect 13820 9036 13872 9042
rect 13820 8978 13872 8984
rect 13832 8634 13860 8978
rect 13820 8628 13872 8634
rect 13820 8570 13872 8576
rect 13728 8288 13780 8294
rect 13728 8230 13780 8236
rect 13945 8188 14253 8197
rect 13945 8186 13951 8188
rect 14007 8186 14031 8188
rect 14087 8186 14111 8188
rect 14167 8186 14191 8188
rect 14247 8186 14253 8188
rect 14007 8134 14009 8186
rect 14189 8134 14191 8186
rect 13945 8132 13951 8134
rect 14007 8132 14031 8134
rect 14087 8132 14111 8134
rect 14167 8132 14191 8134
rect 14247 8132 14253 8134
rect 13726 8120 13782 8129
rect 13945 8123 14253 8132
rect 13726 8055 13728 8064
rect 13780 8055 13782 8064
rect 13728 8026 13780 8032
rect 13740 7478 13768 8026
rect 14292 7993 14320 11290
rect 14372 11212 14424 11218
rect 14372 11154 14424 11160
rect 14384 10044 14412 11154
rect 14476 11082 14504 19722
rect 14648 19304 14700 19310
rect 14568 19252 14648 19258
rect 14568 19246 14700 19252
rect 14568 19230 14688 19246
rect 14568 18834 14596 19230
rect 14740 19168 14792 19174
rect 14740 19110 14792 19116
rect 14752 18902 14780 19110
rect 14740 18896 14792 18902
rect 14740 18838 14792 18844
rect 14556 18828 14608 18834
rect 14556 18770 14608 18776
rect 14648 18760 14700 18766
rect 14648 18702 14700 18708
rect 14660 18426 14688 18702
rect 14648 18420 14700 18426
rect 14648 18362 14700 18368
rect 14740 16652 14792 16658
rect 14740 16594 14792 16600
rect 14752 16454 14780 16594
rect 14740 16448 14792 16454
rect 14740 16390 14792 16396
rect 14844 16250 14872 19790
rect 15396 18193 15424 22200
rect 15856 20602 15884 22200
rect 15844 20596 15896 20602
rect 15844 20538 15896 20544
rect 16316 19242 16344 22200
rect 16776 22114 16804 22200
rect 16868 22114 16896 22222
rect 16776 22086 16896 22114
rect 16544 20700 16852 20709
rect 16544 20698 16550 20700
rect 16606 20698 16630 20700
rect 16686 20698 16710 20700
rect 16766 20698 16790 20700
rect 16846 20698 16852 20700
rect 16606 20646 16608 20698
rect 16788 20646 16790 20698
rect 16544 20644 16550 20646
rect 16606 20644 16630 20646
rect 16686 20644 16710 20646
rect 16766 20644 16790 20646
rect 16846 20644 16852 20646
rect 16544 20635 16852 20644
rect 16948 19712 17000 19718
rect 16948 19654 17000 19660
rect 16544 19612 16852 19621
rect 16544 19610 16550 19612
rect 16606 19610 16630 19612
rect 16686 19610 16710 19612
rect 16766 19610 16790 19612
rect 16846 19610 16852 19612
rect 16606 19558 16608 19610
rect 16788 19558 16790 19610
rect 16544 19556 16550 19558
rect 16606 19556 16630 19558
rect 16686 19556 16710 19558
rect 16766 19556 16790 19558
rect 16846 19556 16852 19558
rect 16544 19547 16852 19556
rect 16960 19242 16988 19654
rect 17052 19310 17080 22222
rect 17222 22200 17278 23000
rect 17682 22200 17738 23000
rect 18142 22200 18198 23000
rect 18602 22200 18658 23000
rect 19062 22200 19118 23000
rect 19522 22200 19578 23000
rect 19982 22200 20038 23000
rect 20442 22200 20498 23000
rect 20902 22200 20958 23000
rect 21362 22200 21418 23000
rect 21822 22200 21878 23000
rect 22282 22200 22338 23000
rect 22742 22200 22798 23000
rect 17236 20330 17264 22200
rect 17224 20324 17276 20330
rect 17224 20266 17276 20272
rect 17040 19304 17092 19310
rect 17040 19246 17092 19252
rect 16304 19236 16356 19242
rect 16304 19178 16356 19184
rect 16948 19236 17000 19242
rect 16948 19178 17000 19184
rect 17696 18986 17724 22200
rect 18156 19174 18184 22200
rect 18144 19168 18196 19174
rect 18144 19110 18196 19116
rect 17512 18970 17724 18986
rect 17500 18964 17724 18970
rect 17552 18958 17724 18964
rect 17500 18906 17552 18912
rect 18616 18873 18644 22200
rect 19076 20058 19104 22200
rect 19143 20156 19451 20165
rect 19143 20154 19149 20156
rect 19205 20154 19229 20156
rect 19285 20154 19309 20156
rect 19365 20154 19389 20156
rect 19445 20154 19451 20156
rect 19205 20102 19207 20154
rect 19387 20102 19389 20154
rect 19143 20100 19149 20102
rect 19205 20100 19229 20102
rect 19285 20100 19309 20102
rect 19365 20100 19389 20102
rect 19445 20100 19451 20102
rect 19143 20091 19451 20100
rect 19064 20052 19116 20058
rect 19064 19994 19116 20000
rect 19143 19068 19451 19077
rect 19143 19066 19149 19068
rect 19205 19066 19229 19068
rect 19285 19066 19309 19068
rect 19365 19066 19389 19068
rect 19445 19066 19451 19068
rect 19205 19014 19207 19066
rect 19387 19014 19389 19066
rect 19143 19012 19149 19014
rect 19205 19012 19229 19014
rect 19285 19012 19309 19014
rect 19365 19012 19389 19014
rect 19445 19012 19451 19014
rect 19143 19003 19451 19012
rect 18602 18864 18658 18873
rect 18602 18799 18658 18808
rect 16396 18760 16448 18766
rect 19536 18737 19564 22200
rect 19616 19508 19668 19514
rect 19616 19450 19668 19456
rect 16396 18702 16448 18708
rect 19522 18728 19578 18737
rect 16120 18624 16172 18630
rect 16120 18566 16172 18572
rect 15382 18184 15438 18193
rect 15382 18119 15438 18128
rect 16132 18086 16160 18566
rect 16408 18290 16436 18702
rect 17868 18692 17920 18698
rect 19522 18663 19578 18672
rect 17868 18634 17920 18640
rect 16948 18624 17000 18630
rect 16948 18566 17000 18572
rect 16544 18524 16852 18533
rect 16544 18522 16550 18524
rect 16606 18522 16630 18524
rect 16686 18522 16710 18524
rect 16766 18522 16790 18524
rect 16846 18522 16852 18524
rect 16606 18470 16608 18522
rect 16788 18470 16790 18522
rect 16544 18468 16550 18470
rect 16606 18468 16630 18470
rect 16686 18468 16710 18470
rect 16766 18468 16790 18470
rect 16846 18468 16852 18470
rect 16544 18459 16852 18468
rect 16396 18284 16448 18290
rect 16396 18226 16448 18232
rect 16120 18080 16172 18086
rect 16120 18022 16172 18028
rect 15108 17740 15160 17746
rect 15108 17682 15160 17688
rect 15120 17066 15148 17682
rect 15844 17264 15896 17270
rect 15844 17206 15896 17212
rect 15108 17060 15160 17066
rect 15108 17002 15160 17008
rect 15476 16992 15528 16998
rect 15476 16934 15528 16940
rect 15200 16516 15252 16522
rect 15200 16458 15252 16464
rect 15384 16516 15436 16522
rect 15384 16458 15436 16464
rect 14832 16244 14884 16250
rect 14832 16186 14884 16192
rect 15108 16108 15160 16114
rect 15108 16050 15160 16056
rect 14832 15904 14884 15910
rect 14832 15846 14884 15852
rect 14648 15428 14700 15434
rect 14648 15370 14700 15376
rect 14556 15156 14608 15162
rect 14556 15098 14608 15104
rect 14568 12753 14596 15098
rect 14554 12744 14610 12753
rect 14554 12679 14610 12688
rect 14556 12640 14608 12646
rect 14556 12582 14608 12588
rect 14568 11830 14596 12582
rect 14660 12374 14688 15370
rect 14740 15360 14792 15366
rect 14740 15302 14792 15308
rect 14648 12368 14700 12374
rect 14648 12310 14700 12316
rect 14660 12170 14688 12310
rect 14752 12209 14780 15302
rect 14844 12986 14872 15846
rect 14924 15496 14976 15502
rect 14924 15438 14976 15444
rect 14936 14618 14964 15438
rect 15016 15020 15068 15026
rect 15016 14962 15068 14968
rect 15028 14929 15056 14962
rect 15014 14920 15070 14929
rect 15014 14855 15070 14864
rect 14924 14612 14976 14618
rect 14924 14554 14976 14560
rect 15028 13530 15056 14855
rect 15120 14074 15148 16050
rect 15212 16046 15240 16458
rect 15396 16182 15424 16458
rect 15384 16176 15436 16182
rect 15384 16118 15436 16124
rect 15200 16040 15252 16046
rect 15200 15982 15252 15988
rect 15212 15416 15240 15982
rect 15488 15450 15516 16934
rect 15856 16794 15884 17206
rect 16132 17105 16160 18022
rect 16960 17898 16988 18566
rect 17880 18426 17908 18634
rect 18236 18624 18288 18630
rect 18236 18566 18288 18572
rect 17868 18420 17920 18426
rect 17868 18362 17920 18368
rect 17776 18284 17828 18290
rect 17776 18226 17828 18232
rect 16868 17882 16988 17898
rect 16856 17876 16988 17882
rect 16908 17870 16988 17876
rect 16856 17818 16908 17824
rect 16396 17740 16448 17746
rect 16396 17682 16448 17688
rect 16408 17270 16436 17682
rect 16544 17436 16852 17445
rect 16544 17434 16550 17436
rect 16606 17434 16630 17436
rect 16686 17434 16710 17436
rect 16766 17434 16790 17436
rect 16846 17434 16852 17436
rect 16606 17382 16608 17434
rect 16788 17382 16790 17434
rect 16544 17380 16550 17382
rect 16606 17380 16630 17382
rect 16686 17380 16710 17382
rect 16766 17380 16790 17382
rect 16846 17380 16852 17382
rect 16544 17371 16852 17380
rect 16396 17264 16448 17270
rect 16210 17232 16266 17241
rect 16396 17206 16448 17212
rect 16210 17167 16212 17176
rect 16264 17167 16266 17176
rect 16212 17138 16264 17144
rect 16118 17096 16174 17105
rect 16118 17031 16174 17040
rect 17788 16998 17816 18226
rect 17776 16992 17828 16998
rect 17776 16934 17828 16940
rect 15844 16788 15896 16794
rect 15844 16730 15896 16736
rect 17880 16561 17908 18362
rect 18248 18358 18276 18566
rect 18236 18352 18288 18358
rect 18236 18294 18288 18300
rect 18972 18284 19024 18290
rect 18972 18226 19024 18232
rect 18984 17542 19012 18226
rect 19143 17980 19451 17989
rect 19143 17978 19149 17980
rect 19205 17978 19229 17980
rect 19285 17978 19309 17980
rect 19365 17978 19389 17980
rect 19445 17978 19451 17980
rect 19205 17926 19207 17978
rect 19387 17926 19389 17978
rect 19143 17924 19149 17926
rect 19205 17924 19229 17926
rect 19285 17924 19309 17926
rect 19365 17924 19389 17926
rect 19445 17924 19451 17926
rect 19143 17915 19451 17924
rect 19628 17785 19656 19450
rect 19996 19281 20024 22200
rect 20456 20262 20484 22200
rect 20916 20369 20944 22200
rect 20902 20360 20958 20369
rect 20902 20295 20958 20304
rect 20444 20256 20496 20262
rect 20444 20198 20496 20204
rect 21376 20058 21404 22200
rect 21836 20890 21864 22200
rect 21652 20862 21864 20890
rect 21548 20392 21600 20398
rect 21548 20334 21600 20340
rect 21364 20052 21416 20058
rect 21364 19994 21416 20000
rect 21560 19922 21588 20334
rect 21548 19916 21600 19922
rect 21548 19858 21600 19864
rect 21088 19780 21140 19786
rect 21088 19722 21140 19728
rect 20168 19712 20220 19718
rect 20168 19654 20220 19660
rect 19982 19272 20038 19281
rect 19982 19207 20038 19216
rect 19708 18760 19760 18766
rect 19708 18702 19760 18708
rect 19614 17776 19670 17785
rect 19614 17711 19670 17720
rect 18972 17536 19024 17542
rect 18972 17478 19024 17484
rect 19628 17241 19656 17711
rect 19720 17610 19748 18702
rect 19892 18624 19944 18630
rect 19892 18566 19944 18572
rect 19904 17678 19932 18566
rect 19892 17672 19944 17678
rect 19892 17614 19944 17620
rect 19708 17604 19760 17610
rect 19708 17546 19760 17552
rect 19614 17232 19670 17241
rect 19064 17196 19116 17202
rect 19614 17167 19670 17176
rect 19064 17138 19116 17144
rect 18052 17128 18104 17134
rect 18052 17070 18104 17076
rect 18064 16794 18092 17070
rect 18052 16788 18104 16794
rect 18052 16730 18104 16736
rect 17866 16552 17922 16561
rect 16396 16516 16448 16522
rect 17866 16487 17922 16496
rect 17960 16516 18012 16522
rect 16396 16458 16448 16464
rect 17960 16458 18012 16464
rect 15844 15904 15896 15910
rect 15844 15846 15896 15852
rect 15856 15638 15884 15846
rect 15844 15632 15896 15638
rect 15844 15574 15896 15580
rect 15488 15434 15608 15450
rect 15384 15428 15436 15434
rect 15212 15388 15384 15416
rect 15212 15026 15240 15388
rect 15488 15428 15620 15434
rect 15488 15422 15568 15428
rect 15384 15370 15436 15376
rect 15568 15370 15620 15376
rect 16408 15162 16436 16458
rect 16544 16348 16852 16357
rect 16544 16346 16550 16348
rect 16606 16346 16630 16348
rect 16686 16346 16710 16348
rect 16766 16346 16790 16348
rect 16846 16346 16852 16348
rect 16606 16294 16608 16346
rect 16788 16294 16790 16346
rect 16544 16292 16550 16294
rect 16606 16292 16630 16294
rect 16686 16292 16710 16294
rect 16766 16292 16790 16294
rect 16846 16292 16852 16294
rect 16544 16283 16852 16292
rect 17500 15360 17552 15366
rect 17500 15302 17552 15308
rect 16544 15260 16852 15269
rect 16544 15258 16550 15260
rect 16606 15258 16630 15260
rect 16686 15258 16710 15260
rect 16766 15258 16790 15260
rect 16846 15258 16852 15260
rect 16606 15206 16608 15258
rect 16788 15206 16790 15258
rect 16544 15204 16550 15206
rect 16606 15204 16630 15206
rect 16686 15204 16710 15206
rect 16766 15204 16790 15206
rect 16846 15204 16852 15206
rect 16544 15195 16852 15204
rect 16396 15156 16448 15162
rect 16396 15098 16448 15104
rect 15200 15020 15252 15026
rect 15200 14962 15252 14968
rect 15212 14618 15240 14962
rect 16212 14884 16264 14890
rect 16212 14826 16264 14832
rect 15200 14612 15252 14618
rect 15200 14554 15252 14560
rect 16224 14414 16252 14826
rect 16396 14476 16448 14482
rect 16396 14418 16448 14424
rect 15568 14408 15620 14414
rect 15568 14350 15620 14356
rect 16212 14408 16264 14414
rect 16212 14350 16264 14356
rect 15108 14068 15160 14074
rect 15108 14010 15160 14016
rect 15016 13524 15068 13530
rect 15016 13466 15068 13472
rect 14832 12980 14884 12986
rect 14832 12922 14884 12928
rect 14924 12232 14976 12238
rect 14738 12200 14794 12209
rect 14648 12164 14700 12170
rect 14924 12174 14976 12180
rect 14738 12135 14794 12144
rect 14648 12106 14700 12112
rect 14740 12096 14792 12102
rect 14740 12038 14792 12044
rect 14556 11824 14608 11830
rect 14556 11766 14608 11772
rect 14752 11286 14780 12038
rect 14740 11280 14792 11286
rect 14740 11222 14792 11228
rect 14464 11076 14516 11082
rect 14464 11018 14516 11024
rect 14464 10736 14516 10742
rect 14464 10678 14516 10684
rect 14476 10266 14504 10678
rect 14648 10464 14700 10470
rect 14648 10406 14700 10412
rect 14464 10260 14516 10266
rect 14464 10202 14516 10208
rect 14554 10160 14610 10169
rect 14554 10095 14610 10104
rect 14464 10056 14516 10062
rect 14384 10016 14464 10044
rect 14464 9998 14516 10004
rect 14568 8634 14596 10095
rect 14660 9654 14688 10406
rect 14936 10266 14964 12174
rect 15120 11762 15148 14010
rect 15580 13462 15608 14350
rect 16212 14272 16264 14278
rect 16212 14214 16264 14220
rect 15568 13456 15620 13462
rect 15568 13398 15620 13404
rect 15936 13184 15988 13190
rect 15936 13126 15988 13132
rect 15948 12850 15976 13126
rect 15936 12844 15988 12850
rect 15936 12786 15988 12792
rect 15108 11756 15160 11762
rect 15108 11698 15160 11704
rect 15108 11144 15160 11150
rect 15108 11086 15160 11092
rect 15120 10674 15148 11086
rect 15200 11008 15252 11014
rect 15200 10950 15252 10956
rect 15108 10668 15160 10674
rect 15108 10610 15160 10616
rect 14924 10260 14976 10266
rect 14924 10202 14976 10208
rect 14738 10024 14794 10033
rect 14738 9959 14794 9968
rect 14648 9648 14700 9654
rect 14648 9590 14700 9596
rect 14556 8628 14608 8634
rect 14556 8570 14608 8576
rect 14464 8424 14516 8430
rect 14464 8366 14516 8372
rect 14278 7984 14334 7993
rect 14278 7919 14334 7928
rect 14188 7812 14240 7818
rect 14188 7754 14240 7760
rect 14372 7812 14424 7818
rect 14372 7754 14424 7760
rect 13728 7472 13780 7478
rect 13634 7440 13690 7449
rect 13728 7414 13780 7420
rect 13634 7375 13690 7384
rect 13648 6089 13676 7375
rect 14200 7290 14228 7754
rect 14280 7744 14332 7750
rect 14280 7686 14332 7692
rect 14292 7546 14320 7686
rect 14280 7540 14332 7546
rect 14280 7482 14332 7488
rect 13820 7268 13872 7274
rect 14200 7262 14320 7290
rect 13820 7210 13872 7216
rect 13832 7002 13860 7210
rect 13945 7100 14253 7109
rect 13945 7098 13951 7100
rect 14007 7098 14031 7100
rect 14087 7098 14111 7100
rect 14167 7098 14191 7100
rect 14247 7098 14253 7100
rect 14007 7046 14009 7098
rect 14189 7046 14191 7098
rect 13945 7044 13951 7046
rect 14007 7044 14031 7046
rect 14087 7044 14111 7046
rect 14167 7044 14191 7046
rect 14247 7044 14253 7046
rect 13945 7035 14253 7044
rect 13820 6996 13872 7002
rect 13820 6938 13872 6944
rect 13820 6656 13872 6662
rect 13820 6598 13872 6604
rect 13634 6080 13690 6089
rect 13634 6015 13690 6024
rect 13372 5222 13492 5250
rect 13542 5264 13598 5273
rect 13372 5030 13400 5222
rect 13542 5199 13598 5208
rect 13452 5160 13504 5166
rect 13452 5102 13504 5108
rect 13360 5024 13412 5030
rect 13360 4966 13412 4972
rect 13268 4276 13320 4282
rect 13268 4218 13320 4224
rect 12714 4176 12770 4185
rect 12714 4111 12770 4120
rect 12808 4140 12860 4146
rect 12808 4082 12860 4088
rect 12820 800 12848 4082
rect 13464 3058 13492 5102
rect 13636 4616 13688 4622
rect 13636 4558 13688 4564
rect 13544 3528 13596 3534
rect 13544 3470 13596 3476
rect 13556 3058 13584 3470
rect 13648 3466 13676 4558
rect 13832 4146 13860 6598
rect 13945 6012 14253 6021
rect 13945 6010 13951 6012
rect 14007 6010 14031 6012
rect 14087 6010 14111 6012
rect 14167 6010 14191 6012
rect 14247 6010 14253 6012
rect 14007 5958 14009 6010
rect 14189 5958 14191 6010
rect 13945 5956 13951 5958
rect 14007 5956 14031 5958
rect 14087 5956 14111 5958
rect 14167 5956 14191 5958
rect 14247 5956 14253 5958
rect 13945 5947 14253 5956
rect 14292 5794 14320 7262
rect 14384 6798 14412 7754
rect 14372 6792 14424 6798
rect 14372 6734 14424 6740
rect 14476 6458 14504 8366
rect 14556 8016 14608 8022
rect 14556 7958 14608 7964
rect 14568 6866 14596 7958
rect 14556 6860 14608 6866
rect 14556 6802 14608 6808
rect 14660 6730 14688 9590
rect 14752 6866 14780 9959
rect 14832 9376 14884 9382
rect 14832 9318 14884 9324
rect 14740 6860 14792 6866
rect 14740 6802 14792 6808
rect 14648 6724 14700 6730
rect 14648 6666 14700 6672
rect 14752 6474 14780 6802
rect 14464 6452 14516 6458
rect 14464 6394 14516 6400
rect 14660 6446 14780 6474
rect 14292 5766 14412 5794
rect 14384 5642 14412 5766
rect 14280 5636 14332 5642
rect 14280 5578 14332 5584
rect 14372 5636 14424 5642
rect 14372 5578 14424 5584
rect 13945 4924 14253 4933
rect 13945 4922 13951 4924
rect 14007 4922 14031 4924
rect 14087 4922 14111 4924
rect 14167 4922 14191 4924
rect 14247 4922 14253 4924
rect 14007 4870 14009 4922
rect 14189 4870 14191 4922
rect 13945 4868 13951 4870
rect 14007 4868 14031 4870
rect 14087 4868 14111 4870
rect 14167 4868 14191 4870
rect 14247 4868 14253 4870
rect 13945 4859 14253 4868
rect 13820 4140 13872 4146
rect 13820 4082 13872 4088
rect 13945 3836 14253 3845
rect 13945 3834 13951 3836
rect 14007 3834 14031 3836
rect 14087 3834 14111 3836
rect 14167 3834 14191 3836
rect 14247 3834 14253 3836
rect 14007 3782 14009 3834
rect 14189 3782 14191 3834
rect 13945 3780 13951 3782
rect 14007 3780 14031 3782
rect 14087 3780 14111 3782
rect 14167 3780 14191 3782
rect 14247 3780 14253 3782
rect 13945 3771 14253 3780
rect 13636 3460 13688 3466
rect 13636 3402 13688 3408
rect 13728 3392 13780 3398
rect 13728 3334 13780 3340
rect 13740 3058 13768 3334
rect 14292 3058 14320 5578
rect 14660 4729 14688 6446
rect 14740 6384 14792 6390
rect 14740 6326 14792 6332
rect 14646 4720 14702 4729
rect 14646 4655 14702 4664
rect 14752 4622 14780 6326
rect 14844 5114 14872 9318
rect 14936 7206 14964 10202
rect 15016 9716 15068 9722
rect 15016 9658 15068 9664
rect 15028 7342 15056 9658
rect 15120 9586 15148 10610
rect 15108 9580 15160 9586
rect 15108 9522 15160 9528
rect 15108 8628 15160 8634
rect 15108 8570 15160 8576
rect 15120 8090 15148 8570
rect 15108 8084 15160 8090
rect 15108 8026 15160 8032
rect 15212 7954 15240 10950
rect 15568 10736 15620 10742
rect 15568 10678 15620 10684
rect 15292 10056 15344 10062
rect 15292 9998 15344 10004
rect 15304 8838 15332 9998
rect 15580 9926 15608 10678
rect 15568 9920 15620 9926
rect 15568 9862 15620 9868
rect 15660 9920 15712 9926
rect 15660 9862 15712 9868
rect 15292 8832 15344 8838
rect 15292 8774 15344 8780
rect 15200 7948 15252 7954
rect 15200 7890 15252 7896
rect 15108 7880 15160 7886
rect 15108 7822 15160 7828
rect 15120 7546 15148 7822
rect 15108 7540 15160 7546
rect 15108 7482 15160 7488
rect 15016 7336 15068 7342
rect 15016 7278 15068 7284
rect 14924 7200 14976 7206
rect 14924 7142 14976 7148
rect 15028 6934 15056 7278
rect 15016 6928 15068 6934
rect 15016 6870 15068 6876
rect 15200 5228 15252 5234
rect 15200 5170 15252 5176
rect 14844 5086 14964 5114
rect 14832 5024 14884 5030
rect 14832 4966 14884 4972
rect 14844 4690 14872 4966
rect 14832 4684 14884 4690
rect 14832 4626 14884 4632
rect 14740 4616 14792 4622
rect 14740 4558 14792 4564
rect 14372 4480 14424 4486
rect 14372 4422 14424 4428
rect 14384 4146 14412 4422
rect 14372 4140 14424 4146
rect 14372 4082 14424 4088
rect 14556 4004 14608 4010
rect 14556 3946 14608 3952
rect 14568 3058 14596 3946
rect 14936 3534 14964 5086
rect 15212 4049 15240 5170
rect 15198 4040 15254 4049
rect 15198 3975 15254 3984
rect 14924 3528 14976 3534
rect 15304 3505 15332 8774
rect 15382 8528 15438 8537
rect 15382 8463 15384 8472
rect 15436 8463 15438 8472
rect 15384 8434 15436 8440
rect 15476 8084 15528 8090
rect 15476 8026 15528 8032
rect 15488 7546 15516 8026
rect 15476 7540 15528 7546
rect 15476 7482 15528 7488
rect 15476 7404 15528 7410
rect 15476 7346 15528 7352
rect 15488 6866 15516 7346
rect 15476 6860 15528 6866
rect 15476 6802 15528 6808
rect 15580 6322 15608 9862
rect 15672 9586 15700 9862
rect 16224 9625 16252 14214
rect 16408 13938 16436 14418
rect 17224 14340 17276 14346
rect 17224 14282 17276 14288
rect 16544 14172 16852 14181
rect 16544 14170 16550 14172
rect 16606 14170 16630 14172
rect 16686 14170 16710 14172
rect 16766 14170 16790 14172
rect 16846 14170 16852 14172
rect 16606 14118 16608 14170
rect 16788 14118 16790 14170
rect 16544 14116 16550 14118
rect 16606 14116 16630 14118
rect 16686 14116 16710 14118
rect 16766 14116 16790 14118
rect 16846 14116 16852 14118
rect 16544 14107 16852 14116
rect 17236 14074 17264 14282
rect 17224 14068 17276 14074
rect 17224 14010 17276 14016
rect 16396 13932 16448 13938
rect 16396 13874 16448 13880
rect 16544 13084 16852 13093
rect 16544 13082 16550 13084
rect 16606 13082 16630 13084
rect 16686 13082 16710 13084
rect 16766 13082 16790 13084
rect 16846 13082 16852 13084
rect 16606 13030 16608 13082
rect 16788 13030 16790 13082
rect 16544 13028 16550 13030
rect 16606 13028 16630 13030
rect 16686 13028 16710 13030
rect 16766 13028 16790 13030
rect 16846 13028 16852 13030
rect 16544 13019 16852 13028
rect 16672 12844 16724 12850
rect 16672 12786 16724 12792
rect 16578 12744 16634 12753
rect 16578 12679 16634 12688
rect 16592 12170 16620 12679
rect 16684 12306 16712 12786
rect 16672 12300 16724 12306
rect 16672 12242 16724 12248
rect 16580 12164 16632 12170
rect 16580 12106 16632 12112
rect 16544 11996 16852 12005
rect 16544 11994 16550 11996
rect 16606 11994 16630 11996
rect 16686 11994 16710 11996
rect 16766 11994 16790 11996
rect 16846 11994 16852 11996
rect 16606 11942 16608 11994
rect 16788 11942 16790 11994
rect 16544 11940 16550 11942
rect 16606 11940 16630 11942
rect 16686 11940 16710 11942
rect 16766 11940 16790 11942
rect 16846 11940 16852 11942
rect 16544 11931 16852 11940
rect 16396 11756 16448 11762
rect 16396 11698 16448 11704
rect 16304 11552 16356 11558
rect 16304 11494 16356 11500
rect 16316 11150 16344 11494
rect 16304 11144 16356 11150
rect 16304 11086 16356 11092
rect 16316 10674 16344 11086
rect 16408 10810 16436 11698
rect 16764 11280 16816 11286
rect 16816 11228 17080 11234
rect 16764 11222 17080 11228
rect 16776 11206 17080 11222
rect 16544 10908 16852 10917
rect 16544 10906 16550 10908
rect 16606 10906 16630 10908
rect 16686 10906 16710 10908
rect 16766 10906 16790 10908
rect 16846 10906 16852 10908
rect 16606 10854 16608 10906
rect 16788 10854 16790 10906
rect 16544 10852 16550 10854
rect 16606 10852 16630 10854
rect 16686 10852 16710 10854
rect 16766 10852 16790 10854
rect 16846 10852 16852 10854
rect 16544 10843 16852 10852
rect 16396 10804 16448 10810
rect 16396 10746 16448 10752
rect 16948 10804 17000 10810
rect 16948 10746 17000 10752
rect 16304 10668 16356 10674
rect 16304 10610 16356 10616
rect 16960 10062 16988 10746
rect 16948 10056 17000 10062
rect 16948 9998 17000 10004
rect 16304 9988 16356 9994
rect 16304 9930 16356 9936
rect 16210 9616 16266 9625
rect 15660 9580 15712 9586
rect 16210 9551 16266 9560
rect 15660 9522 15712 9528
rect 15568 6316 15620 6322
rect 15568 6258 15620 6264
rect 15672 5574 15700 9522
rect 15752 9172 15804 9178
rect 15752 9114 15804 9120
rect 15764 8634 15792 9114
rect 16212 8900 16264 8906
rect 16212 8842 16264 8848
rect 15752 8628 15804 8634
rect 15752 8570 15804 8576
rect 15752 7880 15804 7886
rect 15752 7822 15804 7828
rect 15764 7750 15792 7822
rect 15752 7744 15804 7750
rect 15752 7686 15804 7692
rect 15764 5817 15792 7686
rect 15844 6112 15896 6118
rect 15844 6054 15896 6060
rect 15750 5808 15806 5817
rect 15750 5743 15806 5752
rect 15660 5568 15712 5574
rect 15660 5510 15712 5516
rect 15856 5234 15884 6054
rect 15844 5228 15896 5234
rect 15844 5170 15896 5176
rect 15476 5160 15528 5166
rect 15476 5102 15528 5108
rect 15488 4826 15516 5102
rect 15476 4820 15528 4826
rect 15476 4762 15528 4768
rect 16028 4684 16080 4690
rect 16028 4626 16080 4632
rect 15844 4616 15896 4622
rect 15844 4558 15896 4564
rect 15752 4208 15804 4214
rect 15752 4150 15804 4156
rect 15384 4072 15436 4078
rect 15384 4014 15436 4020
rect 14924 3470 14976 3476
rect 15290 3496 15346 3505
rect 15290 3431 15346 3440
rect 15396 3058 15424 4014
rect 15568 3188 15620 3194
rect 15568 3130 15620 3136
rect 13452 3052 13504 3058
rect 13452 2994 13504 3000
rect 13544 3052 13596 3058
rect 13544 2994 13596 3000
rect 13728 3052 13780 3058
rect 13728 2994 13780 3000
rect 14280 3052 14332 3058
rect 14280 2994 14332 3000
rect 14556 3052 14608 3058
rect 14556 2994 14608 3000
rect 14924 3052 14976 3058
rect 14924 2994 14976 3000
rect 15384 3052 15436 3058
rect 15384 2994 15436 3000
rect 13176 2984 13228 2990
rect 13556 2938 13584 2994
rect 13228 2932 13584 2938
rect 13176 2926 13584 2932
rect 13820 2984 13872 2990
rect 13820 2926 13872 2932
rect 13188 2910 13584 2926
rect 13268 2848 13320 2854
rect 13268 2790 13320 2796
rect 13728 2848 13780 2854
rect 13728 2790 13780 2796
rect 13280 800 13308 2790
rect 13740 800 13768 2790
rect 13832 2446 13860 2926
rect 13945 2748 14253 2757
rect 13945 2746 13951 2748
rect 14007 2746 14031 2748
rect 14087 2746 14111 2748
rect 14167 2746 14191 2748
rect 14247 2746 14253 2748
rect 14007 2694 14009 2746
rect 14189 2694 14191 2746
rect 13945 2692 13951 2694
rect 14007 2692 14031 2694
rect 14087 2692 14111 2694
rect 14167 2692 14191 2694
rect 14247 2692 14253 2694
rect 13945 2683 14253 2692
rect 14568 2650 14596 2994
rect 14648 2848 14700 2854
rect 14648 2790 14700 2796
rect 14556 2644 14608 2650
rect 14556 2586 14608 2592
rect 13820 2440 13872 2446
rect 13820 2382 13872 2388
rect 14188 2304 14240 2310
rect 14188 2246 14240 2252
rect 14200 800 14228 2246
rect 14660 800 14688 2790
rect 14936 2650 14964 2994
rect 15108 2916 15160 2922
rect 15108 2858 15160 2864
rect 14924 2644 14976 2650
rect 14924 2586 14976 2592
rect 15120 800 15148 2858
rect 15580 800 15608 3130
rect 15764 3058 15792 4150
rect 15856 3738 15884 4558
rect 15936 4480 15988 4486
rect 15936 4422 15988 4428
rect 15948 4010 15976 4422
rect 15936 4004 15988 4010
rect 15936 3946 15988 3952
rect 16040 3942 16068 4626
rect 16028 3936 16080 3942
rect 16028 3878 16080 3884
rect 16224 3738 16252 8842
rect 16316 6186 16344 9930
rect 16544 9820 16852 9829
rect 16544 9818 16550 9820
rect 16606 9818 16630 9820
rect 16686 9818 16710 9820
rect 16766 9818 16790 9820
rect 16846 9818 16852 9820
rect 16606 9766 16608 9818
rect 16788 9766 16790 9818
rect 16544 9764 16550 9766
rect 16606 9764 16630 9766
rect 16686 9764 16710 9766
rect 16766 9764 16790 9766
rect 16846 9764 16852 9766
rect 16544 9755 16852 9764
rect 16488 9580 16540 9586
rect 16488 9522 16540 9528
rect 16500 9178 16528 9522
rect 16948 9376 17000 9382
rect 16948 9318 17000 9324
rect 16488 9172 16540 9178
rect 16488 9114 16540 9120
rect 16960 8906 16988 9318
rect 16948 8900 17000 8906
rect 16948 8842 17000 8848
rect 16544 8732 16852 8741
rect 16544 8730 16550 8732
rect 16606 8730 16630 8732
rect 16686 8730 16710 8732
rect 16766 8730 16790 8732
rect 16846 8730 16852 8732
rect 16606 8678 16608 8730
rect 16788 8678 16790 8730
rect 16544 8676 16550 8678
rect 16606 8676 16630 8678
rect 16686 8676 16710 8678
rect 16766 8676 16790 8678
rect 16846 8676 16852 8678
rect 16544 8667 16852 8676
rect 16488 8288 16540 8294
rect 16488 8230 16540 8236
rect 16500 8090 16528 8230
rect 16396 8084 16448 8090
rect 16396 8026 16448 8032
rect 16488 8084 16540 8090
rect 16488 8026 16540 8032
rect 16408 7750 16436 8026
rect 16396 7744 16448 7750
rect 16396 7686 16448 7692
rect 16408 7177 16436 7686
rect 16544 7644 16852 7653
rect 16544 7642 16550 7644
rect 16606 7642 16630 7644
rect 16686 7642 16710 7644
rect 16766 7642 16790 7644
rect 16846 7642 16852 7644
rect 16606 7590 16608 7642
rect 16788 7590 16790 7642
rect 16544 7588 16550 7590
rect 16606 7588 16630 7590
rect 16686 7588 16710 7590
rect 16766 7588 16790 7590
rect 16846 7588 16852 7590
rect 16544 7579 16852 7588
rect 16960 7313 16988 8842
rect 17052 8838 17080 11206
rect 17130 10704 17186 10713
rect 17130 10639 17186 10648
rect 17040 8832 17092 8838
rect 17040 8774 17092 8780
rect 16946 7304 17002 7313
rect 16946 7239 17002 7248
rect 16394 7168 16450 7177
rect 16394 7103 16450 7112
rect 16946 6760 17002 6769
rect 16946 6695 17002 6704
rect 16544 6556 16852 6565
rect 16544 6554 16550 6556
rect 16606 6554 16630 6556
rect 16686 6554 16710 6556
rect 16766 6554 16790 6556
rect 16846 6554 16852 6556
rect 16606 6502 16608 6554
rect 16788 6502 16790 6554
rect 16544 6500 16550 6502
rect 16606 6500 16630 6502
rect 16686 6500 16710 6502
rect 16766 6500 16790 6502
rect 16846 6500 16852 6502
rect 16544 6491 16852 6500
rect 16304 6180 16356 6186
rect 16304 6122 16356 6128
rect 16396 5568 16448 5574
rect 16394 5536 16396 5545
rect 16448 5536 16450 5545
rect 16394 5471 16450 5480
rect 16544 5468 16852 5477
rect 16544 5466 16550 5468
rect 16606 5466 16630 5468
rect 16686 5466 16710 5468
rect 16766 5466 16790 5468
rect 16846 5466 16852 5468
rect 16606 5414 16608 5466
rect 16788 5414 16790 5466
rect 16544 5412 16550 5414
rect 16606 5412 16630 5414
rect 16686 5412 16710 5414
rect 16766 5412 16790 5414
rect 16846 5412 16852 5414
rect 16544 5403 16852 5412
rect 16960 4826 16988 6695
rect 17052 5302 17080 8774
rect 17040 5296 17092 5302
rect 17040 5238 17092 5244
rect 17040 5160 17092 5166
rect 17040 5102 17092 5108
rect 16948 4820 17000 4826
rect 16948 4762 17000 4768
rect 16960 4622 16988 4762
rect 16948 4616 17000 4622
rect 16948 4558 17000 4564
rect 16396 4480 16448 4486
rect 16396 4422 16448 4428
rect 15844 3732 15896 3738
rect 15844 3674 15896 3680
rect 16212 3732 16264 3738
rect 16212 3674 16264 3680
rect 16304 3460 16356 3466
rect 16304 3402 16356 3408
rect 16212 3392 16264 3398
rect 16212 3334 16264 3340
rect 16224 3058 16252 3334
rect 16316 3194 16344 3402
rect 16304 3188 16356 3194
rect 16304 3130 16356 3136
rect 15752 3052 15804 3058
rect 15752 2994 15804 3000
rect 16212 3052 16264 3058
rect 16212 2994 16264 3000
rect 15764 2650 15792 2994
rect 15936 2984 15988 2990
rect 15936 2926 15988 2932
rect 15948 2650 15976 2926
rect 16028 2916 16080 2922
rect 16028 2858 16080 2864
rect 15752 2644 15804 2650
rect 15752 2586 15804 2592
rect 15936 2644 15988 2650
rect 15936 2586 15988 2592
rect 16040 800 16068 2858
rect 16408 1986 16436 4422
rect 16544 4380 16852 4389
rect 16544 4378 16550 4380
rect 16606 4378 16630 4380
rect 16686 4378 16710 4380
rect 16766 4378 16790 4380
rect 16846 4378 16852 4380
rect 16606 4326 16608 4378
rect 16788 4326 16790 4378
rect 16544 4324 16550 4326
rect 16606 4324 16630 4326
rect 16686 4324 16710 4326
rect 16766 4324 16790 4326
rect 16846 4324 16852 4326
rect 16544 4315 16852 4324
rect 16960 4146 16988 4558
rect 16948 4140 17000 4146
rect 16948 4082 17000 4088
rect 16544 3292 16852 3301
rect 16544 3290 16550 3292
rect 16606 3290 16630 3292
rect 16686 3290 16710 3292
rect 16766 3290 16790 3292
rect 16846 3290 16852 3292
rect 16606 3238 16608 3290
rect 16788 3238 16790 3290
rect 16544 3236 16550 3238
rect 16606 3236 16630 3238
rect 16686 3236 16710 3238
rect 16766 3236 16790 3238
rect 16846 3236 16852 3238
rect 16544 3227 16852 3236
rect 17052 3058 17080 5102
rect 17144 4078 17172 10639
rect 17236 9489 17264 14010
rect 17408 13320 17460 13326
rect 17408 13262 17460 13268
rect 17420 13190 17448 13262
rect 17408 13184 17460 13190
rect 17408 13126 17460 13132
rect 17512 12850 17540 15302
rect 17972 13870 18000 16458
rect 18972 16448 19024 16454
rect 18972 16390 19024 16396
rect 18984 16114 19012 16390
rect 18972 16108 19024 16114
rect 18972 16050 19024 16056
rect 18052 14952 18104 14958
rect 18052 14894 18104 14900
rect 18064 14618 18092 14894
rect 18696 14816 18748 14822
rect 18696 14758 18748 14764
rect 18052 14612 18104 14618
rect 18052 14554 18104 14560
rect 18708 14006 18736 14758
rect 18984 14521 19012 16050
rect 18970 14512 19026 14521
rect 18970 14447 19026 14456
rect 19076 14278 19104 17138
rect 19143 16892 19451 16901
rect 19143 16890 19149 16892
rect 19205 16890 19229 16892
rect 19285 16890 19309 16892
rect 19365 16890 19389 16892
rect 19445 16890 19451 16892
rect 19205 16838 19207 16890
rect 19387 16838 19389 16890
rect 19143 16836 19149 16838
rect 19205 16836 19229 16838
rect 19285 16836 19309 16838
rect 19365 16836 19389 16838
rect 19445 16836 19451 16838
rect 19143 16827 19451 16836
rect 19143 15804 19451 15813
rect 19143 15802 19149 15804
rect 19205 15802 19229 15804
rect 19285 15802 19309 15804
rect 19365 15802 19389 15804
rect 19445 15802 19451 15804
rect 19205 15750 19207 15802
rect 19387 15750 19389 15802
rect 19143 15748 19149 15750
rect 19205 15748 19229 15750
rect 19285 15748 19309 15750
rect 19365 15748 19389 15750
rect 19445 15748 19451 15750
rect 19143 15739 19451 15748
rect 19904 15706 19932 17614
rect 20180 17338 20208 19654
rect 20996 19372 21048 19378
rect 20996 19314 21048 19320
rect 20904 19304 20956 19310
rect 20904 19246 20956 19252
rect 20352 18692 20404 18698
rect 20352 18634 20404 18640
rect 20168 17332 20220 17338
rect 20168 17274 20220 17280
rect 20364 16998 20392 18634
rect 20916 18329 20944 19246
rect 21008 18970 21036 19314
rect 20996 18964 21048 18970
rect 20996 18906 21048 18912
rect 21008 18426 21036 18906
rect 20996 18420 21048 18426
rect 20996 18362 21048 18368
rect 20902 18320 20958 18329
rect 20902 18255 20958 18264
rect 20916 18154 20944 18255
rect 20904 18148 20956 18154
rect 20904 18090 20956 18096
rect 21008 17882 21036 18362
rect 20996 17876 21048 17882
rect 20996 17818 21048 17824
rect 21008 17338 21036 17818
rect 21100 17542 21128 19722
rect 21560 19514 21588 19858
rect 21548 19508 21600 19514
rect 21548 19450 21600 19456
rect 21652 19174 21680 20862
rect 21742 20700 22050 20709
rect 21742 20698 21748 20700
rect 21804 20698 21828 20700
rect 21884 20698 21908 20700
rect 21964 20698 21988 20700
rect 22044 20698 22050 20700
rect 21804 20646 21806 20698
rect 21986 20646 21988 20698
rect 21742 20644 21748 20646
rect 21804 20644 21828 20646
rect 21884 20644 21908 20646
rect 21964 20644 21988 20646
rect 22044 20644 22050 20646
rect 21742 20635 22050 20644
rect 22296 20466 22324 22200
rect 22284 20460 22336 20466
rect 22284 20402 22336 20408
rect 21742 19612 22050 19621
rect 21742 19610 21748 19612
rect 21804 19610 21828 19612
rect 21884 19610 21908 19612
rect 21964 19610 21988 19612
rect 22044 19610 22050 19612
rect 21804 19558 21806 19610
rect 21986 19558 21988 19610
rect 21742 19556 21748 19558
rect 21804 19556 21828 19558
rect 21884 19556 21908 19558
rect 21964 19556 21988 19558
rect 22044 19556 22050 19558
rect 21742 19547 22050 19556
rect 21640 19168 21692 19174
rect 21640 19110 21692 19116
rect 22756 18766 22784 22200
rect 22744 18760 22796 18766
rect 22744 18702 22796 18708
rect 21742 18524 22050 18533
rect 21742 18522 21748 18524
rect 21804 18522 21828 18524
rect 21884 18522 21908 18524
rect 21964 18522 21988 18524
rect 22044 18522 22050 18524
rect 21804 18470 21806 18522
rect 21986 18470 21988 18522
rect 21742 18468 21748 18470
rect 21804 18468 21828 18470
rect 21884 18468 21908 18470
rect 21964 18468 21988 18470
rect 22044 18468 22050 18470
rect 21742 18459 22050 18468
rect 21088 17536 21140 17542
rect 21088 17478 21140 17484
rect 20996 17332 21048 17338
rect 20996 17274 21048 17280
rect 20352 16992 20404 16998
rect 20352 16934 20404 16940
rect 20076 15904 20128 15910
rect 20076 15846 20128 15852
rect 19892 15700 19944 15706
rect 19892 15642 19944 15648
rect 20088 15162 20116 15846
rect 20076 15156 20128 15162
rect 20076 15098 20128 15104
rect 20168 15088 20220 15094
rect 20168 15030 20220 15036
rect 19800 15020 19852 15026
rect 19800 14962 19852 14968
rect 19143 14716 19451 14725
rect 19143 14714 19149 14716
rect 19205 14714 19229 14716
rect 19285 14714 19309 14716
rect 19365 14714 19389 14716
rect 19445 14714 19451 14716
rect 19205 14662 19207 14714
rect 19387 14662 19389 14714
rect 19143 14660 19149 14662
rect 19205 14660 19229 14662
rect 19285 14660 19309 14662
rect 19365 14660 19389 14662
rect 19445 14660 19451 14662
rect 19143 14651 19451 14660
rect 19812 14278 19840 14962
rect 19064 14272 19116 14278
rect 19064 14214 19116 14220
rect 19800 14272 19852 14278
rect 19800 14214 19852 14220
rect 18696 14000 18748 14006
rect 18696 13942 18748 13948
rect 18972 14000 19024 14006
rect 18972 13942 19024 13948
rect 17960 13864 18012 13870
rect 17960 13806 18012 13812
rect 17972 12889 18000 13806
rect 18052 13252 18104 13258
rect 18052 13194 18104 13200
rect 18064 12986 18092 13194
rect 18144 13184 18196 13190
rect 18144 13126 18196 13132
rect 18052 12980 18104 12986
rect 18052 12922 18104 12928
rect 17958 12880 18014 12889
rect 17500 12844 17552 12850
rect 17958 12815 18014 12824
rect 17500 12786 17552 12792
rect 18156 12782 18184 13126
rect 18144 12776 18196 12782
rect 18144 12718 18196 12724
rect 18156 12424 18184 12718
rect 18236 12436 18288 12442
rect 18156 12396 18236 12424
rect 18236 12378 18288 12384
rect 18248 11898 18276 12378
rect 18984 12345 19012 13942
rect 19143 13628 19451 13637
rect 19143 13626 19149 13628
rect 19205 13626 19229 13628
rect 19285 13626 19309 13628
rect 19365 13626 19389 13628
rect 19445 13626 19451 13628
rect 19205 13574 19207 13626
rect 19387 13574 19389 13626
rect 19143 13572 19149 13574
rect 19205 13572 19229 13574
rect 19285 13572 19309 13574
rect 19365 13572 19389 13574
rect 19445 13572 19451 13574
rect 19143 13563 19451 13572
rect 19522 13424 19578 13433
rect 19522 13359 19578 13368
rect 19536 12986 19564 13359
rect 19708 13320 19760 13326
rect 19708 13262 19760 13268
rect 19524 12980 19576 12986
rect 19524 12922 19576 12928
rect 19616 12640 19668 12646
rect 19616 12582 19668 12588
rect 19143 12540 19451 12549
rect 19143 12538 19149 12540
rect 19205 12538 19229 12540
rect 19285 12538 19309 12540
rect 19365 12538 19389 12540
rect 19445 12538 19451 12540
rect 19205 12486 19207 12538
rect 19387 12486 19389 12538
rect 19143 12484 19149 12486
rect 19205 12484 19229 12486
rect 19285 12484 19309 12486
rect 19365 12484 19389 12486
rect 19445 12484 19451 12486
rect 19143 12475 19451 12484
rect 18970 12336 19026 12345
rect 18970 12271 19026 12280
rect 18236 11892 18288 11898
rect 18236 11834 18288 11840
rect 18880 11552 18932 11558
rect 18880 11494 18932 11500
rect 18972 11552 19024 11558
rect 18972 11494 19024 11500
rect 17972 11082 18184 11098
rect 17684 11076 17736 11082
rect 17972 11076 18196 11082
rect 17972 11070 18144 11076
rect 17972 11064 18000 11070
rect 17736 11036 18000 11064
rect 17684 11018 17736 11024
rect 18144 11018 18196 11024
rect 17960 10600 18012 10606
rect 17960 10542 18012 10548
rect 17972 10062 18000 10542
rect 17960 10056 18012 10062
rect 17960 9998 18012 10004
rect 17972 9674 18000 9998
rect 17972 9646 18092 9674
rect 17776 9580 17828 9586
rect 17776 9522 17828 9528
rect 17222 9480 17278 9489
rect 17222 9415 17278 9424
rect 17592 8832 17644 8838
rect 17592 8774 17644 8780
rect 17316 8492 17368 8498
rect 17316 8434 17368 8440
rect 17224 7744 17276 7750
rect 17224 7686 17276 7692
rect 17236 5137 17264 7686
rect 17222 5128 17278 5137
rect 17222 5063 17278 5072
rect 17224 4480 17276 4486
rect 17224 4422 17276 4428
rect 17132 4072 17184 4078
rect 17132 4014 17184 4020
rect 17144 3670 17172 4014
rect 17236 3942 17264 4422
rect 17328 4078 17356 8434
rect 17408 8288 17460 8294
rect 17408 8230 17460 8236
rect 17420 4486 17448 8230
rect 17604 7818 17632 8774
rect 17788 7857 17816 9522
rect 18064 9518 18092 9646
rect 18052 9512 18104 9518
rect 18052 9454 18104 9460
rect 18064 9178 18092 9454
rect 18052 9172 18104 9178
rect 18052 9114 18104 9120
rect 18156 8362 18184 11018
rect 18512 9920 18564 9926
rect 18512 9862 18564 9868
rect 18144 8356 18196 8362
rect 18144 8298 18196 8304
rect 18142 8256 18198 8265
rect 18142 8191 18198 8200
rect 17774 7848 17830 7857
rect 17592 7812 17644 7818
rect 17774 7783 17830 7792
rect 17592 7754 17644 7760
rect 17500 5772 17552 5778
rect 17500 5714 17552 5720
rect 17512 4690 17540 5714
rect 17604 4758 17632 7754
rect 17684 7744 17736 7750
rect 17684 7686 17736 7692
rect 17696 7449 17724 7686
rect 17788 7546 17816 7783
rect 17776 7540 17828 7546
rect 17776 7482 17828 7488
rect 17868 7472 17920 7478
rect 17682 7440 17738 7449
rect 17868 7414 17920 7420
rect 17682 7375 17738 7384
rect 17776 5568 17828 5574
rect 17776 5510 17828 5516
rect 17788 5370 17816 5510
rect 17776 5364 17828 5370
rect 17776 5306 17828 5312
rect 17592 4752 17644 4758
rect 17592 4694 17644 4700
rect 17500 4684 17552 4690
rect 17500 4626 17552 4632
rect 17776 4548 17828 4554
rect 17776 4490 17828 4496
rect 17408 4480 17460 4486
rect 17408 4422 17460 4428
rect 17592 4480 17644 4486
rect 17592 4422 17644 4428
rect 17684 4480 17736 4486
rect 17684 4422 17736 4428
rect 17604 4282 17632 4422
rect 17592 4276 17644 4282
rect 17592 4218 17644 4224
rect 17408 4208 17460 4214
rect 17408 4150 17460 4156
rect 17316 4072 17368 4078
rect 17316 4014 17368 4020
rect 17224 3936 17276 3942
rect 17224 3878 17276 3884
rect 17420 3738 17448 4150
rect 17408 3732 17460 3738
rect 17408 3674 17460 3680
rect 17132 3664 17184 3670
rect 17132 3606 17184 3612
rect 17040 3052 17092 3058
rect 17040 2994 17092 3000
rect 17696 2961 17724 4422
rect 17788 3058 17816 4490
rect 17880 4146 17908 7414
rect 17958 7168 18014 7177
rect 17958 7103 18014 7112
rect 17868 4140 17920 4146
rect 17868 4082 17920 4088
rect 17880 3534 17908 4082
rect 17868 3528 17920 3534
rect 17868 3470 17920 3476
rect 17868 3188 17920 3194
rect 17868 3130 17920 3136
rect 17776 3052 17828 3058
rect 17776 2994 17828 3000
rect 17682 2952 17738 2961
rect 17408 2916 17460 2922
rect 17682 2887 17738 2896
rect 17408 2858 17460 2864
rect 16948 2848 17000 2854
rect 16948 2790 17000 2796
rect 16544 2204 16852 2213
rect 16544 2202 16550 2204
rect 16606 2202 16630 2204
rect 16686 2202 16710 2204
rect 16766 2202 16790 2204
rect 16846 2202 16852 2204
rect 16606 2150 16608 2202
rect 16788 2150 16790 2202
rect 16544 2148 16550 2150
rect 16606 2148 16630 2150
rect 16686 2148 16710 2150
rect 16766 2148 16790 2150
rect 16846 2148 16852 2150
rect 16544 2139 16852 2148
rect 16408 1958 16528 1986
rect 16500 800 16528 1958
rect 16960 800 16988 2790
rect 17420 800 17448 2858
rect 17880 800 17908 3130
rect 17972 2650 18000 7103
rect 18156 4078 18184 8191
rect 18144 4072 18196 4078
rect 18144 4014 18196 4020
rect 18524 3602 18552 9862
rect 18892 9586 18920 11494
rect 18880 9580 18932 9586
rect 18880 9522 18932 9528
rect 18892 8974 18920 9522
rect 18880 8968 18932 8974
rect 18880 8910 18932 8916
rect 18880 8832 18932 8838
rect 18880 8774 18932 8780
rect 18892 8634 18920 8774
rect 18880 8628 18932 8634
rect 18880 8570 18932 8576
rect 18892 8265 18920 8570
rect 18984 8566 19012 11494
rect 19143 11452 19451 11461
rect 19143 11450 19149 11452
rect 19205 11450 19229 11452
rect 19285 11450 19309 11452
rect 19365 11450 19389 11452
rect 19445 11450 19451 11452
rect 19205 11398 19207 11450
rect 19387 11398 19389 11450
rect 19143 11396 19149 11398
rect 19205 11396 19229 11398
rect 19285 11396 19309 11398
rect 19365 11396 19389 11398
rect 19445 11396 19451 11398
rect 19143 11387 19451 11396
rect 19524 11076 19576 11082
rect 19524 11018 19576 11024
rect 19536 10470 19564 11018
rect 19524 10464 19576 10470
rect 19524 10406 19576 10412
rect 19143 10364 19451 10373
rect 19143 10362 19149 10364
rect 19205 10362 19229 10364
rect 19285 10362 19309 10364
rect 19365 10362 19389 10364
rect 19445 10362 19451 10364
rect 19205 10310 19207 10362
rect 19387 10310 19389 10362
rect 19143 10308 19149 10310
rect 19205 10308 19229 10310
rect 19285 10308 19309 10310
rect 19365 10308 19389 10310
rect 19445 10308 19451 10310
rect 19143 10299 19451 10308
rect 19340 9988 19392 9994
rect 19340 9930 19392 9936
rect 19156 9920 19208 9926
rect 19156 9862 19208 9868
rect 19168 9518 19196 9862
rect 19352 9722 19380 9930
rect 19340 9716 19392 9722
rect 19340 9658 19392 9664
rect 19156 9512 19208 9518
rect 19076 9472 19156 9500
rect 19076 9178 19104 9472
rect 19156 9454 19208 9460
rect 19143 9276 19451 9285
rect 19143 9274 19149 9276
rect 19205 9274 19229 9276
rect 19285 9274 19309 9276
rect 19365 9274 19389 9276
rect 19445 9274 19451 9276
rect 19205 9222 19207 9274
rect 19387 9222 19389 9274
rect 19143 9220 19149 9222
rect 19205 9220 19229 9222
rect 19285 9220 19309 9222
rect 19365 9220 19389 9222
rect 19445 9220 19451 9222
rect 19143 9211 19451 9220
rect 19064 9172 19116 9178
rect 19064 9114 19116 9120
rect 18972 8560 19024 8566
rect 18972 8502 19024 8508
rect 18878 8256 18934 8265
rect 18878 8191 18934 8200
rect 19143 8188 19451 8197
rect 19143 8186 19149 8188
rect 19205 8186 19229 8188
rect 19285 8186 19309 8188
rect 19365 8186 19389 8188
rect 19445 8186 19451 8188
rect 19205 8134 19207 8186
rect 19387 8134 19389 8186
rect 19143 8132 19149 8134
rect 19205 8132 19229 8134
rect 19285 8132 19309 8134
rect 19365 8132 19389 8134
rect 19445 8132 19451 8134
rect 19143 8123 19451 8132
rect 19536 8022 19564 10406
rect 19628 10130 19656 12582
rect 19720 12442 19748 13262
rect 19708 12436 19760 12442
rect 19708 12378 19760 12384
rect 19812 11801 19840 14214
rect 19798 11792 19854 11801
rect 19798 11727 19854 11736
rect 19892 11756 19944 11762
rect 19892 11698 19944 11704
rect 19708 10532 19760 10538
rect 19708 10474 19760 10480
rect 19616 10124 19668 10130
rect 19616 10066 19668 10072
rect 19616 9648 19668 9654
rect 19616 9590 19668 9596
rect 19524 8016 19576 8022
rect 19524 7958 19576 7964
rect 19143 7100 19451 7109
rect 19143 7098 19149 7100
rect 19205 7098 19229 7100
rect 19285 7098 19309 7100
rect 19365 7098 19389 7100
rect 19445 7098 19451 7100
rect 19205 7046 19207 7098
rect 19387 7046 19389 7098
rect 19143 7044 19149 7046
rect 19205 7044 19229 7046
rect 19285 7044 19309 7046
rect 19365 7044 19389 7046
rect 19445 7044 19451 7046
rect 19143 7035 19451 7044
rect 19143 6012 19451 6021
rect 19143 6010 19149 6012
rect 19205 6010 19229 6012
rect 19285 6010 19309 6012
rect 19365 6010 19389 6012
rect 19445 6010 19451 6012
rect 19205 5958 19207 6010
rect 19387 5958 19389 6010
rect 19143 5956 19149 5958
rect 19205 5956 19229 5958
rect 19285 5956 19309 5958
rect 19365 5956 19389 5958
rect 19445 5956 19451 5958
rect 19143 5947 19451 5956
rect 19628 5914 19656 9590
rect 19720 8906 19748 10474
rect 19904 10062 19932 11698
rect 20076 10668 20128 10674
rect 20076 10610 20128 10616
rect 19892 10056 19944 10062
rect 19892 9998 19944 10004
rect 20088 8974 20116 10610
rect 20180 9654 20208 15030
rect 20364 14414 20392 16934
rect 21008 16794 21036 17274
rect 20996 16788 21048 16794
rect 20996 16730 21048 16736
rect 21100 16153 21128 17478
rect 21742 17436 22050 17445
rect 21742 17434 21748 17436
rect 21804 17434 21828 17436
rect 21884 17434 21908 17436
rect 21964 17434 21988 17436
rect 22044 17434 22050 17436
rect 21804 17382 21806 17434
rect 21986 17382 21988 17434
rect 21742 17380 21748 17382
rect 21804 17380 21828 17382
rect 21884 17380 21908 17382
rect 21964 17380 21988 17382
rect 22044 17380 22050 17382
rect 21742 17371 22050 17380
rect 21456 16788 21508 16794
rect 21456 16730 21508 16736
rect 21364 16448 21416 16454
rect 21364 16390 21416 16396
rect 21086 16144 21142 16153
rect 21086 16079 21142 16088
rect 21180 16108 21232 16114
rect 21376 16096 21404 16390
rect 21468 16114 21496 16730
rect 21742 16348 22050 16357
rect 21742 16346 21748 16348
rect 21804 16346 21828 16348
rect 21884 16346 21908 16348
rect 21964 16346 21988 16348
rect 22044 16346 22050 16348
rect 21804 16294 21806 16346
rect 21986 16294 21988 16346
rect 21742 16292 21748 16294
rect 21804 16292 21828 16294
rect 21884 16292 21908 16294
rect 21964 16292 21988 16294
rect 22044 16292 22050 16294
rect 21742 16283 22050 16292
rect 21232 16068 21404 16096
rect 21180 16050 21232 16056
rect 20720 15496 20772 15502
rect 20720 15438 20772 15444
rect 20536 15360 20588 15366
rect 20536 15302 20588 15308
rect 20352 14408 20404 14414
rect 20352 14350 20404 14356
rect 20260 13932 20312 13938
rect 20260 13874 20312 13880
rect 20272 11354 20300 13874
rect 20260 11348 20312 11354
rect 20260 11290 20312 11296
rect 20548 9994 20576 15302
rect 20732 15026 20760 15438
rect 21272 15428 21324 15434
rect 21272 15370 21324 15376
rect 20720 15020 20772 15026
rect 20720 14962 20772 14968
rect 20732 14618 20760 14962
rect 20720 14612 20772 14618
rect 20720 14554 20772 14560
rect 20732 14074 20760 14554
rect 20812 14340 20864 14346
rect 20812 14282 20864 14288
rect 20720 14068 20772 14074
rect 20720 14010 20772 14016
rect 20732 13326 20760 14010
rect 20824 13433 20852 14282
rect 21284 14074 21312 15370
rect 21272 14068 21324 14074
rect 21272 14010 21324 14016
rect 20810 13424 20866 13433
rect 20810 13359 20866 13368
rect 20720 13320 20772 13326
rect 20720 13262 20772 13268
rect 20628 13252 20680 13258
rect 20628 13194 20680 13200
rect 20536 9988 20588 9994
rect 20536 9930 20588 9936
rect 20168 9648 20220 9654
rect 20168 9590 20220 9596
rect 20076 8968 20128 8974
rect 20076 8910 20128 8916
rect 19708 8900 19760 8906
rect 19708 8842 19760 8848
rect 19720 6254 19748 8842
rect 20640 8634 20668 13194
rect 20732 12986 20760 13262
rect 20904 13184 20956 13190
rect 20904 13126 20956 13132
rect 21180 13184 21232 13190
rect 21180 13126 21232 13132
rect 20720 12980 20772 12986
rect 20720 12922 20772 12928
rect 20916 12850 20944 13126
rect 20904 12844 20956 12850
rect 20904 12786 20956 12792
rect 20996 11212 21048 11218
rect 20996 11154 21048 11160
rect 21008 10810 21036 11154
rect 20996 10804 21048 10810
rect 20996 10746 21048 10752
rect 21008 10266 21036 10746
rect 20996 10260 21048 10266
rect 20996 10202 21048 10208
rect 20812 9376 20864 9382
rect 20812 9318 20864 9324
rect 20628 8628 20680 8634
rect 20628 8570 20680 8576
rect 19708 6248 19760 6254
rect 19708 6190 19760 6196
rect 19616 5908 19668 5914
rect 19616 5850 19668 5856
rect 20640 5846 20668 8570
rect 20824 7478 20852 9318
rect 20812 7472 20864 7478
rect 20812 7414 20864 7420
rect 19064 5840 19116 5846
rect 19064 5782 19116 5788
rect 20628 5840 20680 5846
rect 20628 5782 20680 5788
rect 19076 4622 19104 5782
rect 21192 5778 21220 13126
rect 21272 12980 21324 12986
rect 21272 12922 21324 12928
rect 21284 12442 21312 12922
rect 21272 12436 21324 12442
rect 21272 12378 21324 12384
rect 21284 11898 21312 12378
rect 21272 11892 21324 11898
rect 21272 11834 21324 11840
rect 21284 11354 21312 11834
rect 21272 11348 21324 11354
rect 21272 11290 21324 11296
rect 21272 9376 21324 9382
rect 21272 9318 21324 9324
rect 21284 8838 21312 9318
rect 21272 8832 21324 8838
rect 21272 8774 21324 8780
rect 21284 8294 21312 8774
rect 21272 8288 21324 8294
rect 21272 8230 21324 8236
rect 21284 7954 21312 8230
rect 21272 7948 21324 7954
rect 21272 7890 21324 7896
rect 21284 7546 21312 7890
rect 21272 7540 21324 7546
rect 21272 7482 21324 7488
rect 21376 5817 21404 16068
rect 21456 16108 21508 16114
rect 21456 16050 21508 16056
rect 21468 15502 21496 16050
rect 21456 15496 21508 15502
rect 21456 15438 21508 15444
rect 21742 15260 22050 15269
rect 21742 15258 21748 15260
rect 21804 15258 21828 15260
rect 21884 15258 21908 15260
rect 21964 15258 21988 15260
rect 22044 15258 22050 15260
rect 21804 15206 21806 15258
rect 21986 15206 21988 15258
rect 21742 15204 21748 15206
rect 21804 15204 21828 15206
rect 21884 15204 21908 15206
rect 21964 15204 21988 15206
rect 22044 15204 22050 15206
rect 21742 15195 22050 15204
rect 21456 14612 21508 14618
rect 21456 14554 21508 14560
rect 21468 13530 21496 14554
rect 21742 14172 22050 14181
rect 21742 14170 21748 14172
rect 21804 14170 21828 14172
rect 21884 14170 21908 14172
rect 21964 14170 21988 14172
rect 22044 14170 22050 14172
rect 21804 14118 21806 14170
rect 21986 14118 21988 14170
rect 21742 14116 21748 14118
rect 21804 14116 21828 14118
rect 21884 14116 21908 14118
rect 21964 14116 21988 14118
rect 22044 14116 22050 14118
rect 21742 14107 22050 14116
rect 21548 14068 21600 14074
rect 21548 14010 21600 14016
rect 21456 13524 21508 13530
rect 21456 13466 21508 13472
rect 21560 8090 21588 14010
rect 21742 13084 22050 13093
rect 21742 13082 21748 13084
rect 21804 13082 21828 13084
rect 21884 13082 21908 13084
rect 21964 13082 21988 13084
rect 22044 13082 22050 13084
rect 21804 13030 21806 13082
rect 21986 13030 21988 13082
rect 21742 13028 21748 13030
rect 21804 13028 21828 13030
rect 21884 13028 21908 13030
rect 21964 13028 21988 13030
rect 22044 13028 22050 13030
rect 21742 13019 22050 13028
rect 21742 11996 22050 12005
rect 21742 11994 21748 11996
rect 21804 11994 21828 11996
rect 21884 11994 21908 11996
rect 21964 11994 21988 11996
rect 22044 11994 22050 11996
rect 21804 11942 21806 11994
rect 21986 11942 21988 11994
rect 21742 11940 21748 11942
rect 21804 11940 21828 11942
rect 21884 11940 21908 11942
rect 21964 11940 21988 11942
rect 22044 11940 22050 11942
rect 21742 11931 22050 11940
rect 21742 10908 22050 10917
rect 21742 10906 21748 10908
rect 21804 10906 21828 10908
rect 21884 10906 21908 10908
rect 21964 10906 21988 10908
rect 22044 10906 22050 10908
rect 21804 10854 21806 10906
rect 21986 10854 21988 10906
rect 21742 10852 21748 10854
rect 21804 10852 21828 10854
rect 21884 10852 21908 10854
rect 21964 10852 21988 10854
rect 22044 10852 22050 10854
rect 21742 10843 22050 10852
rect 21742 9820 22050 9829
rect 21742 9818 21748 9820
rect 21804 9818 21828 9820
rect 21884 9818 21908 9820
rect 21964 9818 21988 9820
rect 22044 9818 22050 9820
rect 21804 9766 21806 9818
rect 21986 9766 21988 9818
rect 21742 9764 21748 9766
rect 21804 9764 21828 9766
rect 21884 9764 21908 9766
rect 21964 9764 21988 9766
rect 22044 9764 22050 9766
rect 21742 9755 22050 9764
rect 21742 8732 22050 8741
rect 21742 8730 21748 8732
rect 21804 8730 21828 8732
rect 21884 8730 21908 8732
rect 21964 8730 21988 8732
rect 22044 8730 22050 8732
rect 21804 8678 21806 8730
rect 21986 8678 21988 8730
rect 21742 8676 21748 8678
rect 21804 8676 21828 8678
rect 21884 8676 21908 8678
rect 21964 8676 21988 8678
rect 22044 8676 22050 8678
rect 21742 8667 22050 8676
rect 21548 8084 21600 8090
rect 21548 8026 21600 8032
rect 21742 7644 22050 7653
rect 21742 7642 21748 7644
rect 21804 7642 21828 7644
rect 21884 7642 21908 7644
rect 21964 7642 21988 7644
rect 22044 7642 22050 7644
rect 21804 7590 21806 7642
rect 21986 7590 21988 7642
rect 21742 7588 21748 7590
rect 21804 7588 21828 7590
rect 21884 7588 21908 7590
rect 21964 7588 21988 7590
rect 22044 7588 22050 7590
rect 21742 7579 22050 7588
rect 21742 6556 22050 6565
rect 21742 6554 21748 6556
rect 21804 6554 21828 6556
rect 21884 6554 21908 6556
rect 21964 6554 21988 6556
rect 22044 6554 22050 6556
rect 21804 6502 21806 6554
rect 21986 6502 21988 6554
rect 21742 6500 21748 6502
rect 21804 6500 21828 6502
rect 21884 6500 21908 6502
rect 21964 6500 21988 6502
rect 22044 6500 22050 6502
rect 21742 6491 22050 6500
rect 21362 5808 21418 5817
rect 21180 5772 21232 5778
rect 21362 5743 21418 5752
rect 21180 5714 21232 5720
rect 20260 5568 20312 5574
rect 20260 5510 20312 5516
rect 20628 5568 20680 5574
rect 20628 5510 20680 5516
rect 19614 5128 19670 5137
rect 19614 5063 19670 5072
rect 19143 4924 19451 4933
rect 19143 4922 19149 4924
rect 19205 4922 19229 4924
rect 19285 4922 19309 4924
rect 19365 4922 19389 4924
rect 19445 4922 19451 4924
rect 19205 4870 19207 4922
rect 19387 4870 19389 4922
rect 19143 4868 19149 4870
rect 19205 4868 19229 4870
rect 19285 4868 19309 4870
rect 19365 4868 19389 4870
rect 19445 4868 19451 4870
rect 19143 4859 19451 4868
rect 19064 4616 19116 4622
rect 19064 4558 19116 4564
rect 19064 4208 19116 4214
rect 19064 4150 19116 4156
rect 18604 3664 18656 3670
rect 18604 3606 18656 3612
rect 18512 3596 18564 3602
rect 18512 3538 18564 3544
rect 18420 3528 18472 3534
rect 18420 3470 18472 3476
rect 18236 3392 18288 3398
rect 18236 3334 18288 3340
rect 18248 2922 18276 3334
rect 18432 3058 18460 3470
rect 18616 3058 18644 3606
rect 18788 3188 18840 3194
rect 18788 3130 18840 3136
rect 18420 3052 18472 3058
rect 18420 2994 18472 3000
rect 18604 3052 18656 3058
rect 18604 2994 18656 3000
rect 18236 2916 18288 2922
rect 18236 2858 18288 2864
rect 17960 2644 18012 2650
rect 17960 2586 18012 2592
rect 18328 2576 18380 2582
rect 18328 2518 18380 2524
rect 18340 800 18368 2518
rect 18432 2378 18460 2994
rect 18420 2372 18472 2378
rect 18420 2314 18472 2320
rect 18800 800 18828 3130
rect 19076 3058 19104 4150
rect 19143 3836 19451 3845
rect 19143 3834 19149 3836
rect 19205 3834 19229 3836
rect 19285 3834 19309 3836
rect 19365 3834 19389 3836
rect 19445 3834 19451 3836
rect 19205 3782 19207 3834
rect 19387 3782 19389 3834
rect 19143 3780 19149 3782
rect 19205 3780 19229 3782
rect 19285 3780 19309 3782
rect 19365 3780 19389 3782
rect 19445 3780 19451 3782
rect 19143 3771 19451 3780
rect 19248 3188 19300 3194
rect 19432 3188 19484 3194
rect 19300 3148 19432 3176
rect 19248 3130 19300 3136
rect 19432 3130 19484 3136
rect 19628 3058 19656 5063
rect 20272 4826 20300 5510
rect 20640 5234 20668 5510
rect 21742 5468 22050 5477
rect 21742 5466 21748 5468
rect 21804 5466 21828 5468
rect 21884 5466 21908 5468
rect 21964 5466 21988 5468
rect 22044 5466 22050 5468
rect 21804 5414 21806 5466
rect 21986 5414 21988 5466
rect 21742 5412 21748 5414
rect 21804 5412 21828 5414
rect 21884 5412 21908 5414
rect 21964 5412 21988 5414
rect 22044 5412 22050 5414
rect 21742 5403 22050 5412
rect 20628 5228 20680 5234
rect 20628 5170 20680 5176
rect 20904 5160 20956 5166
rect 20904 5102 20956 5108
rect 20260 4820 20312 4826
rect 20260 4762 20312 4768
rect 19892 4548 19944 4554
rect 19892 4490 19944 4496
rect 19904 3058 19932 4490
rect 20168 3460 20220 3466
rect 20168 3402 20220 3408
rect 19064 3052 19116 3058
rect 19524 3052 19576 3058
rect 19116 3012 19196 3040
rect 19064 2994 19116 3000
rect 19064 2916 19116 2922
rect 19064 2858 19116 2864
rect 19076 1442 19104 2858
rect 19168 2854 19196 3012
rect 19524 2994 19576 3000
rect 19616 3052 19668 3058
rect 19892 3052 19944 3058
rect 19668 3012 19840 3040
rect 19616 2994 19668 3000
rect 19156 2848 19208 2854
rect 19156 2790 19208 2796
rect 19143 2748 19451 2757
rect 19143 2746 19149 2748
rect 19205 2746 19229 2748
rect 19285 2746 19309 2748
rect 19365 2746 19389 2748
rect 19445 2746 19451 2748
rect 19205 2694 19207 2746
rect 19387 2694 19389 2746
rect 19143 2692 19149 2694
rect 19205 2692 19229 2694
rect 19285 2692 19309 2694
rect 19365 2692 19389 2694
rect 19445 2692 19451 2694
rect 19143 2683 19451 2692
rect 19536 1578 19564 2994
rect 19812 2938 19840 3012
rect 19892 2994 19944 3000
rect 19984 3052 20036 3058
rect 19984 2994 20036 3000
rect 19996 2938 20024 2994
rect 19812 2910 20024 2938
rect 19536 1550 19748 1578
rect 19076 1414 19288 1442
rect 19260 800 19288 1414
rect 19720 800 19748 1550
rect 20180 800 20208 3402
rect 20916 3058 20944 5102
rect 22468 4684 22520 4690
rect 22468 4626 22520 4632
rect 21742 4380 22050 4389
rect 21742 4378 21748 4380
rect 21804 4378 21828 4380
rect 21884 4378 21908 4380
rect 21964 4378 21988 4380
rect 22044 4378 22050 4380
rect 21804 4326 21806 4378
rect 21986 4326 21988 4378
rect 21742 4324 21748 4326
rect 21804 4324 21828 4326
rect 21884 4324 21908 4326
rect 21964 4324 21988 4326
rect 22044 4324 22050 4326
rect 21742 4315 22050 4324
rect 21548 3392 21600 3398
rect 21548 3334 21600 3340
rect 20904 3052 20956 3058
rect 20904 2994 20956 3000
rect 21088 2984 21140 2990
rect 21088 2926 21140 2932
rect 20628 2916 20680 2922
rect 20628 2858 20680 2864
rect 20640 800 20668 2858
rect 21100 800 21128 2926
rect 21560 800 21588 3334
rect 21742 3292 22050 3301
rect 21742 3290 21748 3292
rect 21804 3290 21828 3292
rect 21884 3290 21908 3292
rect 21964 3290 21988 3292
rect 22044 3290 22050 3292
rect 21804 3238 21806 3290
rect 21986 3238 21988 3290
rect 21742 3236 21748 3238
rect 21804 3236 21828 3238
rect 21884 3236 21908 3238
rect 21964 3236 21988 3238
rect 22044 3236 22050 3238
rect 21742 3227 22050 3236
rect 22100 3120 22152 3126
rect 22100 3062 22152 3068
rect 21742 2204 22050 2213
rect 21742 2202 21748 2204
rect 21804 2202 21828 2204
rect 21884 2202 21908 2204
rect 21964 2202 21988 2204
rect 22044 2202 22050 2204
rect 21804 2150 21806 2202
rect 21986 2150 21988 2202
rect 21742 2148 21748 2150
rect 21804 2148 21828 2150
rect 21884 2148 21908 2150
rect 21964 2148 21988 2150
rect 22044 2148 22050 2150
rect 21742 2139 22050 2148
rect 22112 1442 22140 3062
rect 22020 1414 22140 1442
rect 22020 800 22048 1414
rect 22480 800 22508 4626
rect 11164 734 11376 762
rect 11426 0 11482 800
rect 11886 0 11942 800
rect 12346 0 12402 800
rect 12806 0 12862 800
rect 13266 0 13322 800
rect 13726 0 13782 800
rect 14186 0 14242 800
rect 14646 0 14702 800
rect 15106 0 15162 800
rect 15566 0 15622 800
rect 16026 0 16082 800
rect 16486 0 16542 800
rect 16946 0 17002 800
rect 17406 0 17462 800
rect 17866 0 17922 800
rect 18326 0 18382 800
rect 18786 0 18842 800
rect 19246 0 19302 800
rect 19706 0 19762 800
rect 20166 0 20222 800
rect 20626 0 20682 800
rect 21086 0 21142 800
rect 21546 0 21602 800
rect 22006 0 22062 800
rect 22466 0 22522 800
<< via2 >>
rect 2778 20984 2834 21040
rect 2870 20576 2926 20632
rect 2778 19352 2834 19408
rect 2594 18128 2650 18184
rect 2318 17720 2374 17776
rect 1950 16904 2006 16960
rect 1858 16496 1914 16552
rect 2686 17312 2742 17368
rect 2962 20168 3018 20224
rect 3054 19760 3110 19816
rect 3238 18944 3294 19000
rect 3555 20154 3611 20156
rect 3635 20154 3691 20156
rect 3715 20154 3771 20156
rect 3795 20154 3851 20156
rect 3555 20102 3601 20154
rect 3601 20102 3611 20154
rect 3635 20102 3665 20154
rect 3665 20102 3677 20154
rect 3677 20102 3691 20154
rect 3715 20102 3729 20154
rect 3729 20102 3741 20154
rect 3741 20102 3771 20154
rect 3795 20102 3805 20154
rect 3805 20102 3851 20154
rect 3555 20100 3611 20102
rect 3635 20100 3691 20102
rect 3715 20100 3771 20102
rect 3795 20100 3851 20102
rect 3555 19066 3611 19068
rect 3635 19066 3691 19068
rect 3715 19066 3771 19068
rect 3795 19066 3851 19068
rect 3555 19014 3601 19066
rect 3601 19014 3611 19066
rect 3635 19014 3665 19066
rect 3665 19014 3677 19066
rect 3677 19014 3691 19066
rect 3715 19014 3729 19066
rect 3729 19014 3741 19066
rect 3741 19014 3771 19066
rect 3795 19014 3805 19066
rect 3805 19014 3851 19066
rect 3555 19012 3611 19014
rect 3635 19012 3691 19014
rect 3715 19012 3771 19014
rect 3795 19012 3851 19014
rect 3555 17978 3611 17980
rect 3635 17978 3691 17980
rect 3715 17978 3771 17980
rect 3795 17978 3851 17980
rect 3555 17926 3601 17978
rect 3601 17926 3611 17978
rect 3635 17926 3665 17978
rect 3665 17926 3677 17978
rect 3677 17926 3691 17978
rect 3715 17926 3729 17978
rect 3729 17926 3741 17978
rect 3741 17926 3771 17978
rect 3795 17926 3805 17978
rect 3805 17926 3851 17978
rect 3555 17924 3611 17926
rect 3635 17924 3691 17926
rect 3715 17924 3771 17926
rect 3795 17924 3851 17926
rect 3555 16890 3611 16892
rect 3635 16890 3691 16892
rect 3715 16890 3771 16892
rect 3795 16890 3851 16892
rect 3555 16838 3601 16890
rect 3601 16838 3611 16890
rect 3635 16838 3665 16890
rect 3665 16838 3677 16890
rect 3677 16838 3691 16890
rect 3715 16838 3729 16890
rect 3729 16838 3741 16890
rect 3741 16838 3771 16890
rect 3795 16838 3805 16890
rect 3805 16838 3851 16890
rect 3555 16836 3611 16838
rect 3635 16836 3691 16838
rect 3715 16836 3771 16838
rect 3795 16836 3851 16838
rect 2870 16088 2926 16144
rect 1858 14048 1914 14104
rect 2778 14456 2834 14512
rect 1582 13640 1638 13696
rect 1766 12008 1822 12064
rect 1674 9172 1730 9208
rect 1674 9152 1676 9172
rect 1676 9152 1728 9172
rect 1728 9152 1730 9172
rect 1490 8744 1546 8800
rect 2226 13776 2282 13832
rect 1950 13232 2006 13288
rect 3054 15680 3110 15736
rect 2962 14864 3018 14920
rect 2870 11600 2926 11656
rect 3146 15272 3202 15328
rect 1674 6568 1730 6624
rect 1398 5888 1454 5944
rect 2042 5208 2098 5264
rect 2870 7384 2926 7440
rect 1674 2216 1730 2272
rect 2502 3984 2558 4040
rect 3606 16532 3608 16552
rect 3608 16532 3660 16552
rect 3660 16532 3662 16552
rect 3606 16496 3662 16532
rect 3882 15952 3938 16008
rect 3555 15802 3611 15804
rect 3635 15802 3691 15804
rect 3715 15802 3771 15804
rect 3795 15802 3851 15804
rect 3555 15750 3601 15802
rect 3601 15750 3611 15802
rect 3635 15750 3665 15802
rect 3665 15750 3677 15802
rect 3677 15750 3691 15802
rect 3715 15750 3729 15802
rect 3729 15750 3741 15802
rect 3741 15750 3771 15802
rect 3795 15750 3805 15802
rect 3805 15750 3851 15802
rect 3555 15748 3611 15750
rect 3635 15748 3691 15750
rect 3715 15748 3771 15750
rect 3795 15748 3851 15750
rect 3555 14714 3611 14716
rect 3635 14714 3691 14716
rect 3715 14714 3771 14716
rect 3795 14714 3851 14716
rect 3555 14662 3601 14714
rect 3601 14662 3611 14714
rect 3635 14662 3665 14714
rect 3665 14662 3677 14714
rect 3677 14662 3691 14714
rect 3715 14662 3729 14714
rect 3729 14662 3741 14714
rect 3741 14662 3771 14714
rect 3795 14662 3805 14714
rect 3805 14662 3851 14714
rect 3555 14660 3611 14662
rect 3635 14660 3691 14662
rect 3715 14660 3771 14662
rect 3795 14660 3851 14662
rect 3555 13626 3611 13628
rect 3635 13626 3691 13628
rect 3715 13626 3771 13628
rect 3795 13626 3851 13628
rect 3555 13574 3601 13626
rect 3601 13574 3611 13626
rect 3635 13574 3665 13626
rect 3665 13574 3677 13626
rect 3677 13574 3691 13626
rect 3715 13574 3729 13626
rect 3729 13574 3741 13626
rect 3741 13574 3771 13626
rect 3795 13574 3805 13626
rect 3805 13574 3851 13626
rect 3555 13572 3611 13574
rect 3635 13572 3691 13574
rect 3715 13572 3771 13574
rect 3795 13572 3851 13574
rect 3422 12824 3478 12880
rect 3330 12416 3386 12472
rect 3238 11600 3294 11656
rect 3555 12538 3611 12540
rect 3635 12538 3691 12540
rect 3715 12538 3771 12540
rect 3795 12538 3851 12540
rect 3555 12486 3601 12538
rect 3601 12486 3611 12538
rect 3635 12486 3665 12538
rect 3665 12486 3677 12538
rect 3677 12486 3691 12538
rect 3715 12486 3729 12538
rect 3729 12486 3741 12538
rect 3741 12486 3771 12538
rect 3795 12486 3805 12538
rect 3805 12486 3851 12538
rect 3555 12484 3611 12486
rect 3635 12484 3691 12486
rect 3715 12484 3771 12486
rect 3795 12484 3851 12486
rect 3555 11450 3611 11452
rect 3635 11450 3691 11452
rect 3715 11450 3771 11452
rect 3795 11450 3851 11452
rect 3555 11398 3601 11450
rect 3601 11398 3611 11450
rect 3635 11398 3665 11450
rect 3665 11398 3677 11450
rect 3677 11398 3691 11450
rect 3715 11398 3729 11450
rect 3729 11398 3741 11450
rect 3741 11398 3771 11450
rect 3795 11398 3805 11450
rect 3805 11398 3851 11450
rect 3555 11396 3611 11398
rect 3635 11396 3691 11398
rect 3715 11396 3771 11398
rect 3795 11396 3851 11398
rect 3555 10362 3611 10364
rect 3635 10362 3691 10364
rect 3715 10362 3771 10364
rect 3795 10362 3851 10364
rect 3555 10310 3601 10362
rect 3601 10310 3611 10362
rect 3635 10310 3665 10362
rect 3665 10310 3677 10362
rect 3677 10310 3691 10362
rect 3715 10310 3729 10362
rect 3729 10310 3741 10362
rect 3741 10310 3771 10362
rect 3795 10310 3805 10362
rect 3805 10310 3851 10362
rect 3555 10308 3611 10310
rect 3635 10308 3691 10310
rect 3715 10308 3771 10310
rect 3795 10308 3851 10310
rect 4066 13232 4122 13288
rect 4618 14728 4674 14784
rect 4066 10784 4122 10840
rect 3974 9968 4030 10024
rect 3882 9832 3938 9888
rect 3790 9560 3846 9616
rect 3555 9274 3611 9276
rect 3635 9274 3691 9276
rect 3715 9274 3771 9276
rect 3795 9274 3851 9276
rect 3555 9222 3601 9274
rect 3601 9222 3611 9274
rect 3635 9222 3665 9274
rect 3665 9222 3677 9274
rect 3677 9222 3691 9274
rect 3715 9222 3729 9274
rect 3729 9222 3741 9274
rect 3741 9222 3771 9274
rect 3795 9222 3805 9274
rect 3805 9222 3851 9274
rect 3555 9220 3611 9222
rect 3635 9220 3691 9222
rect 3715 9220 3771 9222
rect 3795 9220 3851 9222
rect 3555 8186 3611 8188
rect 3635 8186 3691 8188
rect 3715 8186 3771 8188
rect 3795 8186 3851 8188
rect 3555 8134 3601 8186
rect 3601 8134 3611 8186
rect 3635 8134 3665 8186
rect 3665 8134 3677 8186
rect 3677 8134 3691 8186
rect 3715 8134 3729 8186
rect 3729 8134 3741 8186
rect 3741 8134 3771 8186
rect 3795 8134 3805 8186
rect 3805 8134 3851 8186
rect 3555 8132 3611 8134
rect 3635 8132 3691 8134
rect 3715 8132 3771 8134
rect 3795 8132 3851 8134
rect 3974 7520 4030 7576
rect 3422 7112 3478 7168
rect 3555 7098 3611 7100
rect 3635 7098 3691 7100
rect 3715 7098 3771 7100
rect 3795 7098 3851 7100
rect 3555 7046 3601 7098
rect 3601 7046 3611 7098
rect 3635 7046 3665 7098
rect 3665 7046 3677 7098
rect 3677 7046 3691 7098
rect 3715 7046 3729 7098
rect 3729 7046 3741 7098
rect 3741 7046 3771 7098
rect 3795 7046 3805 7098
rect 3805 7046 3851 7098
rect 3555 7044 3611 7046
rect 3635 7044 3691 7046
rect 3715 7044 3771 7046
rect 3795 7044 3851 7046
rect 4342 8916 4344 8936
rect 4344 8916 4396 8936
rect 4396 8916 4398 8936
rect 4342 8880 4398 8916
rect 4250 7928 4306 7984
rect 3422 6740 3424 6760
rect 3424 6740 3476 6760
rect 3476 6740 3478 6760
rect 3422 6704 3478 6740
rect 3146 6296 3202 6352
rect 3330 6296 3386 6352
rect 5354 15000 5410 15056
rect 5262 14864 5318 14920
rect 4894 11192 4950 11248
rect 3555 6010 3611 6012
rect 3635 6010 3691 6012
rect 3715 6010 3771 6012
rect 3795 6010 3851 6012
rect 3555 5958 3601 6010
rect 3601 5958 3611 6010
rect 3635 5958 3665 6010
rect 3665 5958 3677 6010
rect 3677 5958 3691 6010
rect 3715 5958 3729 6010
rect 3729 5958 3741 6010
rect 3741 5958 3771 6010
rect 3795 5958 3805 6010
rect 3805 5958 3851 6010
rect 3555 5956 3611 5958
rect 3635 5956 3691 5958
rect 3715 5956 3771 5958
rect 3795 5956 3851 5958
rect 3974 5344 4030 5400
rect 3790 5108 3792 5128
rect 3792 5108 3844 5128
rect 3844 5108 3846 5128
rect 3790 5072 3846 5108
rect 3555 4922 3611 4924
rect 3635 4922 3691 4924
rect 3715 4922 3771 4924
rect 3795 4922 3851 4924
rect 3555 4870 3601 4922
rect 3601 4870 3611 4922
rect 3635 4870 3665 4922
rect 3665 4870 3677 4922
rect 3677 4870 3691 4922
rect 3715 4870 3729 4922
rect 3729 4870 3741 4922
rect 3741 4870 3771 4922
rect 3795 4870 3805 4922
rect 3805 4870 3851 4922
rect 3555 4868 3611 4870
rect 3635 4868 3691 4870
rect 3715 4868 3771 4870
rect 3795 4868 3851 4870
rect 3330 3848 3386 3904
rect 3238 3440 3294 3496
rect 2870 3032 2926 3088
rect 3974 4664 4030 4720
rect 3555 3834 3611 3836
rect 3635 3834 3691 3836
rect 3715 3834 3771 3836
rect 3795 3834 3851 3836
rect 3555 3782 3601 3834
rect 3601 3782 3611 3834
rect 3635 3782 3665 3834
rect 3665 3782 3677 3834
rect 3677 3782 3691 3834
rect 3715 3782 3729 3834
rect 3729 3782 3741 3834
rect 3741 3782 3771 3834
rect 3795 3782 3805 3834
rect 3805 3782 3851 3834
rect 3555 3780 3611 3782
rect 3635 3780 3691 3782
rect 3715 3780 3771 3782
rect 3795 3780 3851 3782
rect 3555 2746 3611 2748
rect 3635 2746 3691 2748
rect 3715 2746 3771 2748
rect 3795 2746 3851 2748
rect 3555 2694 3601 2746
rect 3601 2694 3611 2746
rect 3635 2694 3665 2746
rect 3665 2694 3677 2746
rect 3677 2694 3691 2746
rect 3715 2694 3729 2746
rect 3729 2694 3741 2746
rect 3741 2694 3771 2746
rect 3795 2694 3805 2746
rect 3805 2694 3851 2746
rect 3555 2692 3611 2694
rect 3635 2692 3691 2694
rect 3715 2692 3771 2694
rect 3795 2692 3851 2694
rect 3422 2624 3478 2680
rect 3422 1808 3478 1864
rect 4710 4664 4766 4720
rect 5078 11600 5134 11656
rect 5078 11192 5134 11248
rect 6154 20698 6210 20700
rect 6234 20698 6290 20700
rect 6314 20698 6370 20700
rect 6394 20698 6450 20700
rect 6154 20646 6200 20698
rect 6200 20646 6210 20698
rect 6234 20646 6264 20698
rect 6264 20646 6276 20698
rect 6276 20646 6290 20698
rect 6314 20646 6328 20698
rect 6328 20646 6340 20698
rect 6340 20646 6370 20698
rect 6394 20646 6404 20698
rect 6404 20646 6450 20698
rect 6154 20644 6210 20646
rect 6234 20644 6290 20646
rect 6314 20644 6370 20646
rect 6394 20644 6450 20646
rect 6154 19610 6210 19612
rect 6234 19610 6290 19612
rect 6314 19610 6370 19612
rect 6394 19610 6450 19612
rect 6154 19558 6200 19610
rect 6200 19558 6210 19610
rect 6234 19558 6264 19610
rect 6264 19558 6276 19610
rect 6276 19558 6290 19610
rect 6314 19558 6328 19610
rect 6328 19558 6340 19610
rect 6340 19558 6370 19610
rect 6394 19558 6404 19610
rect 6404 19558 6450 19610
rect 6154 19556 6210 19558
rect 6234 19556 6290 19558
rect 6314 19556 6370 19558
rect 6394 19556 6450 19558
rect 6154 18522 6210 18524
rect 6234 18522 6290 18524
rect 6314 18522 6370 18524
rect 6394 18522 6450 18524
rect 6154 18470 6200 18522
rect 6200 18470 6210 18522
rect 6234 18470 6264 18522
rect 6264 18470 6276 18522
rect 6276 18470 6290 18522
rect 6314 18470 6328 18522
rect 6328 18470 6340 18522
rect 6340 18470 6370 18522
rect 6394 18470 6404 18522
rect 6404 18470 6450 18522
rect 6154 18468 6210 18470
rect 6234 18468 6290 18470
rect 6314 18468 6370 18470
rect 6394 18468 6450 18470
rect 6642 17992 6698 18048
rect 6154 17434 6210 17436
rect 6234 17434 6290 17436
rect 6314 17434 6370 17436
rect 6394 17434 6450 17436
rect 6154 17382 6200 17434
rect 6200 17382 6210 17434
rect 6234 17382 6264 17434
rect 6264 17382 6276 17434
rect 6276 17382 6290 17434
rect 6314 17382 6328 17434
rect 6328 17382 6340 17434
rect 6340 17382 6370 17434
rect 6394 17382 6404 17434
rect 6404 17382 6450 17434
rect 6154 17380 6210 17382
rect 6234 17380 6290 17382
rect 6314 17380 6370 17382
rect 6394 17380 6450 17382
rect 6182 17040 6238 17096
rect 5998 16632 6054 16688
rect 6154 16346 6210 16348
rect 6234 16346 6290 16348
rect 6314 16346 6370 16348
rect 6394 16346 6450 16348
rect 6154 16294 6200 16346
rect 6200 16294 6210 16346
rect 6234 16294 6264 16346
rect 6264 16294 6276 16346
rect 6276 16294 6290 16346
rect 6314 16294 6328 16346
rect 6328 16294 6340 16346
rect 6340 16294 6370 16346
rect 6394 16294 6404 16346
rect 6404 16294 6450 16346
rect 6154 16292 6210 16294
rect 6234 16292 6290 16294
rect 6314 16292 6370 16294
rect 6394 16292 6450 16294
rect 6154 15258 6210 15260
rect 6234 15258 6290 15260
rect 6314 15258 6370 15260
rect 6394 15258 6450 15260
rect 6154 15206 6200 15258
rect 6200 15206 6210 15258
rect 6234 15206 6264 15258
rect 6264 15206 6276 15258
rect 6276 15206 6290 15258
rect 6314 15206 6328 15258
rect 6328 15206 6340 15258
rect 6340 15206 6370 15258
rect 6394 15206 6404 15258
rect 6404 15206 6450 15258
rect 6154 15204 6210 15206
rect 6234 15204 6290 15206
rect 6314 15204 6370 15206
rect 6394 15204 6450 15206
rect 6154 14170 6210 14172
rect 6234 14170 6290 14172
rect 6314 14170 6370 14172
rect 6394 14170 6450 14172
rect 6154 14118 6200 14170
rect 6200 14118 6210 14170
rect 6234 14118 6264 14170
rect 6264 14118 6276 14170
rect 6276 14118 6290 14170
rect 6314 14118 6328 14170
rect 6328 14118 6340 14170
rect 6340 14118 6370 14170
rect 6394 14118 6404 14170
rect 6404 14118 6450 14170
rect 6154 14116 6210 14118
rect 6234 14116 6290 14118
rect 6314 14116 6370 14118
rect 6394 14116 6450 14118
rect 5262 12824 5318 12880
rect 5170 10104 5226 10160
rect 4894 9424 4950 9480
rect 5078 9152 5134 9208
rect 5078 8744 5134 8800
rect 5262 10004 5264 10024
rect 5264 10004 5316 10024
rect 5316 10004 5318 10024
rect 5262 9968 5318 10004
rect 5630 11056 5686 11112
rect 5446 9560 5502 9616
rect 5262 9016 5318 9072
rect 4802 4256 4858 4312
rect 5078 5208 5134 5264
rect 5170 5092 5226 5128
rect 5170 5072 5172 5092
rect 5172 5072 5224 5092
rect 5224 5072 5226 5092
rect 4986 3848 5042 3904
rect 6550 13912 6606 13968
rect 6090 13640 6146 13696
rect 6154 13082 6210 13084
rect 6234 13082 6290 13084
rect 6314 13082 6370 13084
rect 6394 13082 6450 13084
rect 6154 13030 6200 13082
rect 6200 13030 6210 13082
rect 6234 13030 6264 13082
rect 6264 13030 6276 13082
rect 6276 13030 6290 13082
rect 6314 13030 6328 13082
rect 6328 13030 6340 13082
rect 6340 13030 6370 13082
rect 6394 13030 6404 13082
rect 6404 13030 6450 13082
rect 6154 13028 6210 13030
rect 6234 13028 6290 13030
rect 6314 13028 6370 13030
rect 6394 13028 6450 13030
rect 5630 9324 5632 9344
rect 5632 9324 5684 9344
rect 5684 9324 5686 9344
rect 5630 9288 5686 9324
rect 6918 16360 6974 16416
rect 6918 15408 6974 15464
rect 6918 14728 6974 14784
rect 6826 12688 6882 12744
rect 6154 11994 6210 11996
rect 6234 11994 6290 11996
rect 6314 11994 6370 11996
rect 6394 11994 6450 11996
rect 6154 11942 6200 11994
rect 6200 11942 6210 11994
rect 6234 11942 6264 11994
rect 6264 11942 6276 11994
rect 6276 11942 6290 11994
rect 6314 11942 6328 11994
rect 6328 11942 6340 11994
rect 6340 11942 6370 11994
rect 6394 11942 6404 11994
rect 6404 11942 6450 11994
rect 6154 11940 6210 11942
rect 6234 11940 6290 11942
rect 6314 11940 6370 11942
rect 6394 11940 6450 11942
rect 5814 9444 5870 9480
rect 5814 9424 5816 9444
rect 5816 9424 5868 9444
rect 5868 9424 5870 9444
rect 6154 10906 6210 10908
rect 6234 10906 6290 10908
rect 6314 10906 6370 10908
rect 6394 10906 6450 10908
rect 6154 10854 6200 10906
rect 6200 10854 6210 10906
rect 6234 10854 6264 10906
rect 6264 10854 6276 10906
rect 6276 10854 6290 10906
rect 6314 10854 6328 10906
rect 6328 10854 6340 10906
rect 6340 10854 6370 10906
rect 6394 10854 6404 10906
rect 6404 10854 6450 10906
rect 6154 10852 6210 10854
rect 6234 10852 6290 10854
rect 6314 10852 6370 10854
rect 6394 10852 6450 10854
rect 6090 10376 6146 10432
rect 6642 10512 6698 10568
rect 6274 10104 6330 10160
rect 6918 11892 6974 11928
rect 6918 11872 6920 11892
rect 6920 11872 6972 11892
rect 6972 11872 6974 11892
rect 7378 18128 7434 18184
rect 7562 17992 7618 18048
rect 7286 16088 7342 16144
rect 8022 18536 8078 18592
rect 7746 17720 7802 17776
rect 7746 15564 7802 15600
rect 7746 15544 7748 15564
rect 7748 15544 7800 15564
rect 7800 15544 7802 15564
rect 8298 19216 8354 19272
rect 8298 18672 8354 18728
rect 9218 20324 9274 20360
rect 9218 20304 9220 20324
rect 9220 20304 9272 20324
rect 9272 20304 9274 20324
rect 8753 20154 8809 20156
rect 8833 20154 8889 20156
rect 8913 20154 8969 20156
rect 8993 20154 9049 20156
rect 8753 20102 8799 20154
rect 8799 20102 8809 20154
rect 8833 20102 8863 20154
rect 8863 20102 8875 20154
rect 8875 20102 8889 20154
rect 8913 20102 8927 20154
rect 8927 20102 8939 20154
rect 8939 20102 8969 20154
rect 8993 20102 9003 20154
rect 9003 20102 9049 20154
rect 8753 20100 8809 20102
rect 8833 20100 8889 20102
rect 8913 20100 8969 20102
rect 8993 20100 9049 20102
rect 8574 18808 8630 18864
rect 8482 18400 8538 18456
rect 8298 15852 8300 15872
rect 8300 15852 8352 15872
rect 8352 15852 8354 15872
rect 8298 15816 8354 15852
rect 7838 14220 7840 14240
rect 7840 14220 7892 14240
rect 7892 14220 7894 14240
rect 7838 14184 7894 14220
rect 6918 10668 6974 10704
rect 6918 10648 6920 10668
rect 6920 10648 6972 10668
rect 6972 10648 6974 10668
rect 6826 10104 6882 10160
rect 6154 9818 6210 9820
rect 6234 9818 6290 9820
rect 6314 9818 6370 9820
rect 6394 9818 6450 9820
rect 6154 9766 6200 9818
rect 6200 9766 6210 9818
rect 6234 9766 6264 9818
rect 6264 9766 6276 9818
rect 6276 9766 6290 9818
rect 6314 9766 6328 9818
rect 6328 9766 6340 9818
rect 6340 9766 6370 9818
rect 6394 9766 6404 9818
rect 6404 9766 6450 9818
rect 6154 9764 6210 9766
rect 6234 9764 6290 9766
rect 6314 9764 6370 9766
rect 6394 9764 6450 9766
rect 6550 9696 6606 9752
rect 6090 9036 6146 9072
rect 6090 9016 6092 9036
rect 6092 9016 6144 9036
rect 6144 9016 6146 9036
rect 6274 9288 6330 9344
rect 6826 9560 6882 9616
rect 6826 9036 6882 9072
rect 6826 9016 6828 9036
rect 6828 9016 6880 9036
rect 6880 9016 6882 9036
rect 5814 8744 5870 8800
rect 7102 9696 7158 9752
rect 5538 8336 5594 8392
rect 6154 8730 6210 8732
rect 6234 8730 6290 8732
rect 6314 8730 6370 8732
rect 6394 8730 6450 8732
rect 6154 8678 6200 8730
rect 6200 8678 6210 8730
rect 6234 8678 6264 8730
rect 6264 8678 6276 8730
rect 6276 8678 6290 8730
rect 6314 8678 6328 8730
rect 6328 8678 6340 8730
rect 6340 8678 6370 8730
rect 6394 8678 6404 8730
rect 6404 8678 6450 8730
rect 6154 8676 6210 8678
rect 6234 8676 6290 8678
rect 6314 8676 6370 8678
rect 6394 8676 6450 8678
rect 5814 6704 5870 6760
rect 5722 6604 5724 6624
rect 5724 6604 5776 6624
rect 5776 6604 5778 6624
rect 5722 6568 5778 6604
rect 5446 5752 5502 5808
rect 5446 5516 5448 5536
rect 5448 5516 5500 5536
rect 5500 5516 5502 5536
rect 5446 5480 5502 5516
rect 5630 5344 5686 5400
rect 6366 7828 6368 7848
rect 6368 7828 6420 7848
rect 6420 7828 6422 7848
rect 6366 7792 6422 7828
rect 6154 7642 6210 7644
rect 6234 7642 6290 7644
rect 6314 7642 6370 7644
rect 6394 7642 6450 7644
rect 6154 7590 6200 7642
rect 6200 7590 6210 7642
rect 6234 7590 6264 7642
rect 6264 7590 6276 7642
rect 6276 7590 6290 7642
rect 6314 7590 6328 7642
rect 6328 7590 6340 7642
rect 6340 7590 6370 7642
rect 6394 7590 6404 7642
rect 6404 7590 6450 7642
rect 6154 7588 6210 7590
rect 6234 7588 6290 7590
rect 6314 7588 6370 7590
rect 6394 7588 6450 7590
rect 6366 6840 6422 6896
rect 6154 6554 6210 6556
rect 6234 6554 6290 6556
rect 6314 6554 6370 6556
rect 6394 6554 6450 6556
rect 6154 6502 6200 6554
rect 6200 6502 6210 6554
rect 6234 6502 6264 6554
rect 6264 6502 6276 6554
rect 6276 6502 6290 6554
rect 6314 6502 6328 6554
rect 6328 6502 6340 6554
rect 6340 6502 6370 6554
rect 6394 6502 6404 6554
rect 6404 6502 6450 6554
rect 6154 6500 6210 6502
rect 6234 6500 6290 6502
rect 6314 6500 6370 6502
rect 6394 6500 6450 6502
rect 6550 6024 6606 6080
rect 6918 7384 6974 7440
rect 6918 7248 6974 7304
rect 6826 6704 6882 6760
rect 6734 5888 6790 5944
rect 6154 5466 6210 5468
rect 6234 5466 6290 5468
rect 6314 5466 6370 5468
rect 6394 5466 6450 5468
rect 6154 5414 6200 5466
rect 6200 5414 6210 5466
rect 6234 5414 6264 5466
rect 6264 5414 6276 5466
rect 6276 5414 6290 5466
rect 6314 5414 6328 5466
rect 6328 5414 6340 5466
rect 6340 5414 6370 5466
rect 6394 5414 6404 5466
rect 6404 5414 6450 5466
rect 6154 5412 6210 5414
rect 6234 5412 6290 5414
rect 6314 5412 6370 5414
rect 6394 5412 6450 5414
rect 5722 4020 5724 4040
rect 5724 4020 5776 4040
rect 5776 4020 5778 4040
rect 5722 3984 5778 4020
rect 7746 12724 7748 12744
rect 7748 12724 7800 12744
rect 7800 12724 7802 12744
rect 7746 12688 7802 12724
rect 7562 9424 7618 9480
rect 7470 9152 7526 9208
rect 7194 7928 7250 7984
rect 7194 6704 7250 6760
rect 6826 5480 6882 5536
rect 6154 4378 6210 4380
rect 6234 4378 6290 4380
rect 6314 4378 6370 4380
rect 6394 4378 6450 4380
rect 6154 4326 6200 4378
rect 6200 4326 6210 4378
rect 6234 4326 6264 4378
rect 6264 4326 6276 4378
rect 6276 4326 6290 4378
rect 6314 4326 6328 4378
rect 6328 4326 6340 4378
rect 6340 4326 6370 4378
rect 6394 4326 6404 4378
rect 6404 4326 6450 4378
rect 6154 4324 6210 4326
rect 6234 4324 6290 4326
rect 6314 4324 6370 4326
rect 6394 4324 6450 4326
rect 6366 3596 6422 3632
rect 6366 3576 6368 3596
rect 6368 3576 6420 3596
rect 6420 3576 6422 3596
rect 6154 3290 6210 3292
rect 6234 3290 6290 3292
rect 6314 3290 6370 3292
rect 6394 3290 6450 3292
rect 6154 3238 6200 3290
rect 6200 3238 6210 3290
rect 6234 3238 6264 3290
rect 6264 3238 6276 3290
rect 6276 3238 6290 3290
rect 6314 3238 6328 3290
rect 6328 3238 6340 3290
rect 6340 3238 6370 3290
rect 6394 3238 6404 3290
rect 6404 3238 6450 3290
rect 6154 3236 6210 3238
rect 6234 3236 6290 3238
rect 6314 3236 6370 3238
rect 6394 3236 6450 3238
rect 5906 3168 5962 3224
rect 6550 3032 6606 3088
rect 6154 2202 6210 2204
rect 6234 2202 6290 2204
rect 6314 2202 6370 2204
rect 6394 2202 6450 2204
rect 6154 2150 6200 2202
rect 6200 2150 6210 2202
rect 6234 2150 6264 2202
rect 6264 2150 6276 2202
rect 6276 2150 6290 2202
rect 6314 2150 6328 2202
rect 6328 2150 6340 2202
rect 6340 2150 6370 2202
rect 6394 2150 6404 2202
rect 6404 2150 6450 2202
rect 6154 2148 6210 2150
rect 6234 2148 6290 2150
rect 6314 2148 6370 2150
rect 6394 2148 6450 2150
rect 6734 3612 6736 3632
rect 6736 3612 6788 3632
rect 6788 3612 6790 3632
rect 6734 3576 6790 3612
rect 7746 11056 7802 11112
rect 8022 15000 8078 15056
rect 8206 15000 8262 15056
rect 9126 19080 9182 19136
rect 8753 19066 8809 19068
rect 8833 19066 8889 19068
rect 8913 19066 8969 19068
rect 8993 19066 9049 19068
rect 8753 19014 8799 19066
rect 8799 19014 8809 19066
rect 8833 19014 8863 19066
rect 8863 19014 8875 19066
rect 8875 19014 8889 19066
rect 8913 19014 8927 19066
rect 8927 19014 8939 19066
rect 8939 19014 8969 19066
rect 8993 19014 9003 19066
rect 9003 19014 9049 19066
rect 8753 19012 8809 19014
rect 8833 19012 8889 19014
rect 8913 19012 8969 19014
rect 8993 19012 9049 19014
rect 8850 18264 8906 18320
rect 8753 17978 8809 17980
rect 8833 17978 8889 17980
rect 8913 17978 8969 17980
rect 8993 17978 9049 17980
rect 8753 17926 8799 17978
rect 8799 17926 8809 17978
rect 8833 17926 8863 17978
rect 8863 17926 8875 17978
rect 8875 17926 8889 17978
rect 8913 17926 8927 17978
rect 8927 17926 8939 17978
rect 8939 17926 8969 17978
rect 8993 17926 9003 17978
rect 9003 17926 9049 17978
rect 8753 17924 8809 17926
rect 8833 17924 8889 17926
rect 8913 17924 8969 17926
rect 8993 17924 9049 17926
rect 8753 16890 8809 16892
rect 8833 16890 8889 16892
rect 8913 16890 8969 16892
rect 8993 16890 9049 16892
rect 8753 16838 8799 16890
rect 8799 16838 8809 16890
rect 8833 16838 8863 16890
rect 8863 16838 8875 16890
rect 8875 16838 8889 16890
rect 8913 16838 8927 16890
rect 8927 16838 8939 16890
rect 8939 16838 8969 16890
rect 8993 16838 9003 16890
rect 9003 16838 9049 16890
rect 8753 16836 8809 16838
rect 8833 16836 8889 16838
rect 8913 16836 8969 16838
rect 8993 16836 9049 16838
rect 9402 18400 9458 18456
rect 9678 18944 9734 19000
rect 9954 19624 10010 19680
rect 10046 19080 10102 19136
rect 9586 17992 9642 18048
rect 8753 15802 8809 15804
rect 8833 15802 8889 15804
rect 8913 15802 8969 15804
rect 8993 15802 9049 15804
rect 8753 15750 8799 15802
rect 8799 15750 8809 15802
rect 8833 15750 8863 15802
rect 8863 15750 8875 15802
rect 8875 15750 8889 15802
rect 8913 15750 8927 15802
rect 8927 15750 8939 15802
rect 8939 15750 8969 15802
rect 8993 15750 9003 15802
rect 9003 15750 9049 15802
rect 8753 15748 8809 15750
rect 8833 15748 8889 15750
rect 8913 15748 8969 15750
rect 8993 15748 9049 15750
rect 8753 14714 8809 14716
rect 8833 14714 8889 14716
rect 8913 14714 8969 14716
rect 8993 14714 9049 14716
rect 8753 14662 8799 14714
rect 8799 14662 8809 14714
rect 8833 14662 8863 14714
rect 8863 14662 8875 14714
rect 8875 14662 8889 14714
rect 8913 14662 8927 14714
rect 8927 14662 8939 14714
rect 8939 14662 8969 14714
rect 8993 14662 9003 14714
rect 9003 14662 9049 14714
rect 8753 14660 8809 14662
rect 8833 14660 8889 14662
rect 8913 14660 8969 14662
rect 8993 14660 9049 14662
rect 9126 14476 9182 14512
rect 9126 14456 9128 14476
rect 9128 14456 9180 14476
rect 9180 14456 9182 14476
rect 8753 13626 8809 13628
rect 8833 13626 8889 13628
rect 8913 13626 8969 13628
rect 8993 13626 9049 13628
rect 8753 13574 8799 13626
rect 8799 13574 8809 13626
rect 8833 13574 8863 13626
rect 8863 13574 8875 13626
rect 8875 13574 8889 13626
rect 8913 13574 8927 13626
rect 8927 13574 8939 13626
rect 8939 13574 8969 13626
rect 8993 13574 9003 13626
rect 9003 13574 9049 13626
rect 8753 13572 8809 13574
rect 8833 13572 8889 13574
rect 8913 13572 8969 13574
rect 8993 13572 9049 13574
rect 8666 13388 8722 13424
rect 8666 13368 8668 13388
rect 8668 13368 8720 13388
rect 8720 13368 8722 13388
rect 8753 12538 8809 12540
rect 8833 12538 8889 12540
rect 8913 12538 8969 12540
rect 8993 12538 9049 12540
rect 8753 12486 8799 12538
rect 8799 12486 8809 12538
rect 8833 12486 8863 12538
rect 8863 12486 8875 12538
rect 8875 12486 8889 12538
rect 8913 12486 8927 12538
rect 8927 12486 8939 12538
rect 8939 12486 8969 12538
rect 8993 12486 9003 12538
rect 9003 12486 9049 12538
rect 8753 12484 8809 12486
rect 8833 12484 8889 12486
rect 8913 12484 8969 12486
rect 8993 12484 9049 12486
rect 8753 11450 8809 11452
rect 8833 11450 8889 11452
rect 8913 11450 8969 11452
rect 8993 11450 9049 11452
rect 8753 11398 8799 11450
rect 8799 11398 8809 11450
rect 8833 11398 8863 11450
rect 8863 11398 8875 11450
rect 8875 11398 8889 11450
rect 8913 11398 8927 11450
rect 8927 11398 8939 11450
rect 8939 11398 8969 11450
rect 8993 11398 9003 11450
rect 9003 11398 9049 11450
rect 8753 11396 8809 11398
rect 8833 11396 8889 11398
rect 8913 11396 8969 11398
rect 8993 11396 9049 11398
rect 8753 10362 8809 10364
rect 8833 10362 8889 10364
rect 8913 10362 8969 10364
rect 8993 10362 9049 10364
rect 8753 10310 8799 10362
rect 8799 10310 8809 10362
rect 8833 10310 8863 10362
rect 8863 10310 8875 10362
rect 8875 10310 8889 10362
rect 8913 10310 8927 10362
rect 8927 10310 8939 10362
rect 8939 10310 8969 10362
rect 8993 10310 9003 10362
rect 9003 10310 9049 10362
rect 8753 10308 8809 10310
rect 8833 10308 8889 10310
rect 8913 10308 8969 10310
rect 8993 10308 9049 10310
rect 7654 6840 7710 6896
rect 6918 3168 6974 3224
rect 7654 6160 7710 6216
rect 7746 5908 7802 5944
rect 7746 5888 7748 5908
rect 7748 5888 7800 5908
rect 7800 5888 7802 5908
rect 8114 6704 8170 6760
rect 8298 6840 8354 6896
rect 8390 6568 8446 6624
rect 8753 9274 8809 9276
rect 8833 9274 8889 9276
rect 8913 9274 8969 9276
rect 8993 9274 9049 9276
rect 8753 9222 8799 9274
rect 8799 9222 8809 9274
rect 8833 9222 8863 9274
rect 8863 9222 8875 9274
rect 8875 9222 8889 9274
rect 8913 9222 8927 9274
rect 8927 9222 8939 9274
rect 8939 9222 8969 9274
rect 8993 9222 9003 9274
rect 9003 9222 9049 9274
rect 8753 9220 8809 9222
rect 8833 9220 8889 9222
rect 8913 9220 8969 9222
rect 8993 9220 9049 9222
rect 8753 8186 8809 8188
rect 8833 8186 8889 8188
rect 8913 8186 8969 8188
rect 8993 8186 9049 8188
rect 8753 8134 8799 8186
rect 8799 8134 8809 8186
rect 8833 8134 8863 8186
rect 8863 8134 8875 8186
rect 8875 8134 8889 8186
rect 8913 8134 8927 8186
rect 8927 8134 8939 8186
rect 8939 8134 8969 8186
rect 8993 8134 9003 8186
rect 9003 8134 9049 8186
rect 8753 8132 8809 8134
rect 8833 8132 8889 8134
rect 8913 8132 8969 8134
rect 8993 8132 9049 8134
rect 9126 8064 9182 8120
rect 9402 15308 9404 15328
rect 9404 15308 9456 15328
rect 9456 15308 9458 15328
rect 9402 15272 9458 15308
rect 9770 17992 9826 18048
rect 9770 16516 9826 16552
rect 9770 16496 9772 16516
rect 9772 16496 9824 16516
rect 9824 16496 9826 16516
rect 9770 14068 9826 14104
rect 9770 14048 9772 14068
rect 9772 14048 9824 14068
rect 9824 14048 9826 14068
rect 9494 12416 9550 12472
rect 9494 12144 9550 12200
rect 9494 12008 9550 12064
rect 9954 12280 10010 12336
rect 9862 9968 9918 10024
rect 10598 18400 10654 18456
rect 10230 16088 10286 16144
rect 10230 15952 10286 16008
rect 10230 14764 10232 14784
rect 10232 14764 10284 14784
rect 10284 14764 10286 14784
rect 10230 14728 10286 14764
rect 10506 16088 10562 16144
rect 10506 13912 10562 13968
rect 10138 9560 10194 9616
rect 8574 7384 8630 7440
rect 8574 6704 8630 6760
rect 8753 7098 8809 7100
rect 8833 7098 8889 7100
rect 8913 7098 8969 7100
rect 8993 7098 9049 7100
rect 8753 7046 8799 7098
rect 8799 7046 8809 7098
rect 8833 7046 8863 7098
rect 8863 7046 8875 7098
rect 8875 7046 8889 7098
rect 8913 7046 8927 7098
rect 8927 7046 8939 7098
rect 8939 7046 8969 7098
rect 8993 7046 9003 7098
rect 9003 7046 9049 7098
rect 8753 7044 8809 7046
rect 8833 7044 8889 7046
rect 8913 7044 8969 7046
rect 8993 7044 9049 7046
rect 9034 6568 9090 6624
rect 8482 6024 8538 6080
rect 7562 4392 7618 4448
rect 7562 3848 7618 3904
rect 7746 4528 7802 4584
rect 8114 4004 8170 4040
rect 8114 3984 8116 4004
rect 8116 3984 8168 4004
rect 8168 3984 8170 4004
rect 8574 4936 8630 4992
rect 8753 6010 8809 6012
rect 8833 6010 8889 6012
rect 8913 6010 8969 6012
rect 8993 6010 9049 6012
rect 8753 5958 8799 6010
rect 8799 5958 8809 6010
rect 8833 5958 8863 6010
rect 8863 5958 8875 6010
rect 8875 5958 8889 6010
rect 8913 5958 8927 6010
rect 8927 5958 8939 6010
rect 8939 5958 8969 6010
rect 8993 5958 9003 6010
rect 9003 5958 9049 6010
rect 8753 5956 8809 5958
rect 8833 5956 8889 5958
rect 8913 5956 8969 5958
rect 8993 5956 9049 5958
rect 9402 6432 9458 6488
rect 9218 5888 9274 5944
rect 9862 8372 9864 8392
rect 9864 8372 9916 8392
rect 9916 8372 9918 8392
rect 9586 7284 9588 7304
rect 9588 7284 9640 7304
rect 9640 7284 9642 7304
rect 9586 7248 9642 7284
rect 9862 8336 9918 8372
rect 9586 6704 9642 6760
rect 9126 5616 9182 5672
rect 9402 5480 9458 5536
rect 8753 4922 8809 4924
rect 8833 4922 8889 4924
rect 8913 4922 8969 4924
rect 8993 4922 9049 4924
rect 8753 4870 8799 4922
rect 8799 4870 8809 4922
rect 8833 4870 8863 4922
rect 8863 4870 8875 4922
rect 8875 4870 8889 4922
rect 8913 4870 8927 4922
rect 8927 4870 8939 4922
rect 8939 4870 8969 4922
rect 8993 4870 9003 4922
rect 9003 4870 9049 4922
rect 8753 4868 8809 4870
rect 8833 4868 8889 4870
rect 8913 4868 8969 4870
rect 8993 4868 9049 4870
rect 9126 4800 9182 4856
rect 8758 4664 8814 4720
rect 8482 4528 8538 4584
rect 8206 3576 8262 3632
rect 8574 3884 8576 3904
rect 8576 3884 8628 3904
rect 8628 3884 8630 3904
rect 8574 3848 8630 3884
rect 9494 5072 9550 5128
rect 9402 4392 9458 4448
rect 9678 4140 9734 4176
rect 9678 4120 9680 4140
rect 9680 4120 9732 4140
rect 9732 4120 9734 4140
rect 9586 3848 9642 3904
rect 8753 3834 8809 3836
rect 8833 3834 8889 3836
rect 8913 3834 8969 3836
rect 8993 3834 9049 3836
rect 8753 3782 8799 3834
rect 8799 3782 8809 3834
rect 8833 3782 8863 3834
rect 8863 3782 8875 3834
rect 8875 3782 8889 3834
rect 8913 3782 8927 3834
rect 8927 3782 8939 3834
rect 8939 3782 8969 3834
rect 8993 3782 9003 3834
rect 9003 3782 9049 3834
rect 8753 3780 8809 3782
rect 8833 3780 8889 3782
rect 8913 3780 8969 3782
rect 8993 3780 9049 3782
rect 9126 3304 9182 3360
rect 8753 2746 8809 2748
rect 8833 2746 8889 2748
rect 8913 2746 8969 2748
rect 8993 2746 9049 2748
rect 8753 2694 8799 2746
rect 8799 2694 8809 2746
rect 8833 2694 8863 2746
rect 8863 2694 8875 2746
rect 8875 2694 8889 2746
rect 8913 2694 8927 2746
rect 8927 2694 8939 2746
rect 8939 2694 8969 2746
rect 8993 2694 9003 2746
rect 9003 2694 9049 2746
rect 8753 2692 8809 2694
rect 8833 2692 8889 2694
rect 8913 2692 8969 2694
rect 8993 2692 9049 2694
rect 9126 2488 9182 2544
rect 9954 4936 10010 4992
rect 9954 3596 10010 3632
rect 9954 3576 9956 3596
rect 9956 3576 10008 3596
rect 10008 3576 10010 3596
rect 9678 2916 9734 2952
rect 9678 2896 9680 2916
rect 9680 2896 9732 2916
rect 9732 2896 9734 2916
rect 10138 8472 10194 8528
rect 10322 9560 10378 9616
rect 10782 14048 10838 14104
rect 11352 20698 11408 20700
rect 11432 20698 11488 20700
rect 11512 20698 11568 20700
rect 11592 20698 11648 20700
rect 11352 20646 11398 20698
rect 11398 20646 11408 20698
rect 11432 20646 11462 20698
rect 11462 20646 11474 20698
rect 11474 20646 11488 20698
rect 11512 20646 11526 20698
rect 11526 20646 11538 20698
rect 11538 20646 11568 20698
rect 11592 20646 11602 20698
rect 11602 20646 11648 20698
rect 11352 20644 11408 20646
rect 11432 20644 11488 20646
rect 11512 20644 11568 20646
rect 11592 20644 11648 20646
rect 11352 19610 11408 19612
rect 11432 19610 11488 19612
rect 11512 19610 11568 19612
rect 11592 19610 11648 19612
rect 11352 19558 11398 19610
rect 11398 19558 11408 19610
rect 11432 19558 11462 19610
rect 11462 19558 11474 19610
rect 11474 19558 11488 19610
rect 11512 19558 11526 19610
rect 11526 19558 11538 19610
rect 11538 19558 11568 19610
rect 11592 19558 11602 19610
rect 11602 19558 11648 19610
rect 11352 19556 11408 19558
rect 11432 19556 11488 19558
rect 11512 19556 11568 19558
rect 11592 19556 11648 19558
rect 11352 18522 11408 18524
rect 11432 18522 11488 18524
rect 11512 18522 11568 18524
rect 11592 18522 11648 18524
rect 11352 18470 11398 18522
rect 11398 18470 11408 18522
rect 11432 18470 11462 18522
rect 11462 18470 11474 18522
rect 11474 18470 11488 18522
rect 11512 18470 11526 18522
rect 11526 18470 11538 18522
rect 11538 18470 11568 18522
rect 11592 18470 11602 18522
rect 11602 18470 11648 18522
rect 11352 18468 11408 18470
rect 11432 18468 11488 18470
rect 11512 18468 11568 18470
rect 11592 18468 11648 18470
rect 11610 17856 11666 17912
rect 11352 17434 11408 17436
rect 11432 17434 11488 17436
rect 11512 17434 11568 17436
rect 11592 17434 11648 17436
rect 11352 17382 11398 17434
rect 11398 17382 11408 17434
rect 11432 17382 11462 17434
rect 11462 17382 11474 17434
rect 11474 17382 11488 17434
rect 11512 17382 11526 17434
rect 11526 17382 11538 17434
rect 11538 17382 11568 17434
rect 11592 17382 11602 17434
rect 11602 17382 11648 17434
rect 11352 17380 11408 17382
rect 11432 17380 11488 17382
rect 11512 17380 11568 17382
rect 11592 17380 11648 17382
rect 11518 16768 11574 16824
rect 11352 16346 11408 16348
rect 11432 16346 11488 16348
rect 11512 16346 11568 16348
rect 11592 16346 11648 16348
rect 11352 16294 11398 16346
rect 11398 16294 11408 16346
rect 11432 16294 11462 16346
rect 11462 16294 11474 16346
rect 11474 16294 11488 16346
rect 11512 16294 11526 16346
rect 11526 16294 11538 16346
rect 11538 16294 11568 16346
rect 11592 16294 11602 16346
rect 11602 16294 11648 16346
rect 11352 16292 11408 16294
rect 11432 16292 11488 16294
rect 11512 16292 11568 16294
rect 11592 16292 11648 16294
rect 11058 15308 11060 15328
rect 11060 15308 11112 15328
rect 11112 15308 11114 15328
rect 11058 15272 11114 15308
rect 10782 11736 10838 11792
rect 11352 15258 11408 15260
rect 11432 15258 11488 15260
rect 11512 15258 11568 15260
rect 11592 15258 11648 15260
rect 11352 15206 11398 15258
rect 11398 15206 11408 15258
rect 11432 15206 11462 15258
rect 11462 15206 11474 15258
rect 11474 15206 11488 15258
rect 11512 15206 11526 15258
rect 11526 15206 11538 15258
rect 11538 15206 11568 15258
rect 11592 15206 11602 15258
rect 11602 15206 11648 15258
rect 11352 15204 11408 15206
rect 11432 15204 11488 15206
rect 11512 15204 11568 15206
rect 11592 15204 11648 15206
rect 11352 14170 11408 14172
rect 11432 14170 11488 14172
rect 11512 14170 11568 14172
rect 11592 14170 11648 14172
rect 11352 14118 11398 14170
rect 11398 14118 11408 14170
rect 11432 14118 11462 14170
rect 11462 14118 11474 14170
rect 11474 14118 11488 14170
rect 11512 14118 11526 14170
rect 11526 14118 11538 14170
rect 11538 14118 11568 14170
rect 11592 14118 11602 14170
rect 11602 14118 11648 14170
rect 11352 14116 11408 14118
rect 11432 14116 11488 14118
rect 11512 14116 11568 14118
rect 11592 14116 11648 14118
rect 11518 13268 11520 13288
rect 11520 13268 11572 13288
rect 11572 13268 11574 13288
rect 11518 13232 11574 13268
rect 11352 13082 11408 13084
rect 11432 13082 11488 13084
rect 11512 13082 11568 13084
rect 11592 13082 11648 13084
rect 11352 13030 11398 13082
rect 11398 13030 11408 13082
rect 11432 13030 11462 13082
rect 11462 13030 11474 13082
rect 11474 13030 11488 13082
rect 11512 13030 11526 13082
rect 11526 13030 11538 13082
rect 11538 13030 11568 13082
rect 11592 13030 11602 13082
rect 11602 13030 11648 13082
rect 11352 13028 11408 13030
rect 11432 13028 11488 13030
rect 11512 13028 11568 13030
rect 11592 13028 11648 13030
rect 11794 16768 11850 16824
rect 11886 15408 11942 15464
rect 11978 12960 12034 13016
rect 11794 12416 11850 12472
rect 11352 11994 11408 11996
rect 11432 11994 11488 11996
rect 11512 11994 11568 11996
rect 11592 11994 11648 11996
rect 11352 11942 11398 11994
rect 11398 11942 11408 11994
rect 11432 11942 11462 11994
rect 11462 11942 11474 11994
rect 11474 11942 11488 11994
rect 11512 11942 11526 11994
rect 11526 11942 11538 11994
rect 11538 11942 11568 11994
rect 11592 11942 11602 11994
rect 11602 11942 11648 11994
rect 11352 11940 11408 11942
rect 11432 11940 11488 11942
rect 11512 11940 11568 11942
rect 11592 11940 11648 11942
rect 10598 10648 10654 10704
rect 10598 9152 10654 9208
rect 10506 7928 10562 7984
rect 10598 7792 10654 7848
rect 10598 5888 10654 5944
rect 10874 7792 10930 7848
rect 11058 6840 11114 6896
rect 10874 6568 10930 6624
rect 10322 5108 10324 5128
rect 10324 5108 10376 5128
rect 10376 5108 10378 5128
rect 10322 5072 10378 5108
rect 10414 4936 10470 4992
rect 10782 5208 10838 5264
rect 10598 3032 10654 3088
rect 11058 5344 11114 5400
rect 11058 4120 11114 4176
rect 11058 3440 11114 3496
rect 11058 3168 11114 3224
rect 11334 11348 11390 11384
rect 11334 11328 11336 11348
rect 11336 11328 11388 11348
rect 11388 11328 11390 11348
rect 11352 10906 11408 10908
rect 11432 10906 11488 10908
rect 11512 10906 11568 10908
rect 11592 10906 11648 10908
rect 11352 10854 11398 10906
rect 11398 10854 11408 10906
rect 11432 10854 11462 10906
rect 11462 10854 11474 10906
rect 11474 10854 11488 10906
rect 11512 10854 11526 10906
rect 11526 10854 11538 10906
rect 11538 10854 11568 10906
rect 11592 10854 11602 10906
rect 11602 10854 11648 10906
rect 11352 10852 11408 10854
rect 11432 10852 11488 10854
rect 11512 10852 11568 10854
rect 11592 10852 11648 10854
rect 11702 10648 11758 10704
rect 11352 9818 11408 9820
rect 11432 9818 11488 9820
rect 11512 9818 11568 9820
rect 11592 9818 11648 9820
rect 11352 9766 11398 9818
rect 11398 9766 11408 9818
rect 11432 9766 11462 9818
rect 11462 9766 11474 9818
rect 11474 9766 11488 9818
rect 11512 9766 11526 9818
rect 11526 9766 11538 9818
rect 11538 9766 11568 9818
rect 11592 9766 11602 9818
rect 11602 9766 11648 9818
rect 11352 9764 11408 9766
rect 11432 9764 11488 9766
rect 11512 9764 11568 9766
rect 11592 9764 11648 9766
rect 11518 9152 11574 9208
rect 12070 11600 12126 11656
rect 12530 17856 12586 17912
rect 12530 16904 12586 16960
rect 12530 15952 12586 16008
rect 12438 15544 12494 15600
rect 13951 20154 14007 20156
rect 14031 20154 14087 20156
rect 14111 20154 14167 20156
rect 14191 20154 14247 20156
rect 13951 20102 13997 20154
rect 13997 20102 14007 20154
rect 14031 20102 14061 20154
rect 14061 20102 14073 20154
rect 14073 20102 14087 20154
rect 14111 20102 14125 20154
rect 14125 20102 14137 20154
rect 14137 20102 14167 20154
rect 14191 20102 14201 20154
rect 14201 20102 14247 20154
rect 13951 20100 14007 20102
rect 14031 20100 14087 20102
rect 14111 20100 14167 20102
rect 14191 20100 14247 20102
rect 12714 18944 12770 19000
rect 12806 17992 12862 18048
rect 13082 18028 13084 18048
rect 13084 18028 13136 18048
rect 13136 18028 13138 18048
rect 13082 17992 13138 18028
rect 12898 17176 12954 17232
rect 13358 16904 13414 16960
rect 13358 16768 13414 16824
rect 12346 12552 12402 12608
rect 12254 11192 12310 11248
rect 11334 8880 11390 8936
rect 11518 8880 11574 8936
rect 11352 8730 11408 8732
rect 11432 8730 11488 8732
rect 11512 8730 11568 8732
rect 11592 8730 11648 8732
rect 11352 8678 11398 8730
rect 11398 8678 11408 8730
rect 11432 8678 11462 8730
rect 11462 8678 11474 8730
rect 11474 8678 11488 8730
rect 11512 8678 11526 8730
rect 11526 8678 11538 8730
rect 11538 8678 11568 8730
rect 11592 8678 11602 8730
rect 11602 8678 11648 8730
rect 11352 8676 11408 8678
rect 11432 8676 11488 8678
rect 11512 8676 11568 8678
rect 11592 8676 11648 8678
rect 11334 8200 11390 8256
rect 11334 7948 11390 7984
rect 11334 7928 11336 7948
rect 11336 7928 11388 7948
rect 11388 7928 11390 7948
rect 11352 7642 11408 7644
rect 11432 7642 11488 7644
rect 11512 7642 11568 7644
rect 11592 7642 11648 7644
rect 11352 7590 11398 7642
rect 11398 7590 11408 7642
rect 11432 7590 11462 7642
rect 11462 7590 11474 7642
rect 11474 7590 11488 7642
rect 11512 7590 11526 7642
rect 11526 7590 11538 7642
rect 11538 7590 11568 7642
rect 11592 7590 11602 7642
rect 11602 7590 11648 7642
rect 11352 7588 11408 7590
rect 11432 7588 11488 7590
rect 11512 7588 11568 7590
rect 11592 7588 11648 7590
rect 11352 6554 11408 6556
rect 11432 6554 11488 6556
rect 11512 6554 11568 6556
rect 11592 6554 11648 6556
rect 11352 6502 11398 6554
rect 11398 6502 11408 6554
rect 11432 6502 11462 6554
rect 11462 6502 11474 6554
rect 11474 6502 11488 6554
rect 11512 6502 11526 6554
rect 11526 6502 11538 6554
rect 11538 6502 11568 6554
rect 11592 6502 11602 6554
rect 11602 6502 11648 6554
rect 11352 6500 11408 6502
rect 11432 6500 11488 6502
rect 11512 6500 11568 6502
rect 11592 6500 11648 6502
rect 11518 6296 11574 6352
rect 11334 5888 11390 5944
rect 11518 5888 11574 5944
rect 11702 5752 11758 5808
rect 11352 5466 11408 5468
rect 11432 5466 11488 5468
rect 11512 5466 11568 5468
rect 11592 5466 11648 5468
rect 11352 5414 11398 5466
rect 11398 5414 11408 5466
rect 11432 5414 11462 5466
rect 11462 5414 11474 5466
rect 11474 5414 11488 5466
rect 11512 5414 11526 5466
rect 11526 5414 11538 5466
rect 11538 5414 11568 5466
rect 11592 5414 11602 5466
rect 11602 5414 11648 5466
rect 11352 5412 11408 5414
rect 11432 5412 11488 5414
rect 11512 5412 11568 5414
rect 11592 5412 11648 5414
rect 11794 5208 11850 5264
rect 12346 10240 12402 10296
rect 12530 8336 12586 8392
rect 12806 10240 12862 10296
rect 12530 7948 12586 7984
rect 12530 7928 12532 7948
rect 12532 7928 12584 7948
rect 12584 7928 12586 7948
rect 12070 6976 12126 7032
rect 12070 5752 12126 5808
rect 11352 4378 11408 4380
rect 11432 4378 11488 4380
rect 11512 4378 11568 4380
rect 11592 4378 11648 4380
rect 11352 4326 11398 4378
rect 11398 4326 11408 4378
rect 11432 4326 11462 4378
rect 11462 4326 11474 4378
rect 11474 4326 11488 4378
rect 11512 4326 11526 4378
rect 11526 4326 11538 4378
rect 11538 4326 11568 4378
rect 11592 4326 11602 4378
rect 11602 4326 11648 4378
rect 11352 4324 11408 4326
rect 11432 4324 11488 4326
rect 11512 4324 11568 4326
rect 11592 4324 11648 4326
rect 11242 3596 11298 3632
rect 11242 3576 11244 3596
rect 11244 3576 11296 3596
rect 11296 3576 11298 3596
rect 11352 3290 11408 3292
rect 11432 3290 11488 3292
rect 11512 3290 11568 3292
rect 11592 3290 11648 3292
rect 11352 3238 11398 3290
rect 11398 3238 11408 3290
rect 11432 3238 11462 3290
rect 11462 3238 11474 3290
rect 11474 3238 11488 3290
rect 11512 3238 11526 3290
rect 11526 3238 11538 3290
rect 11538 3238 11568 3290
rect 11592 3238 11602 3290
rect 11602 3238 11648 3290
rect 11352 3236 11408 3238
rect 11432 3236 11488 3238
rect 11512 3236 11568 3238
rect 11592 3236 11648 3238
rect 11352 2202 11408 2204
rect 11432 2202 11488 2204
rect 11512 2202 11568 2204
rect 11592 2202 11648 2204
rect 11352 2150 11398 2202
rect 11398 2150 11408 2202
rect 11432 2150 11462 2202
rect 11462 2150 11474 2202
rect 11474 2150 11488 2202
rect 11512 2150 11526 2202
rect 11526 2150 11538 2202
rect 11538 2150 11568 2202
rect 11592 2150 11602 2202
rect 11602 2150 11648 2202
rect 11352 2148 11408 2150
rect 11432 2148 11488 2150
rect 11512 2148 11568 2150
rect 11592 2148 11648 2150
rect 12622 5888 12678 5944
rect 12438 5516 12440 5536
rect 12440 5516 12492 5536
rect 12492 5516 12494 5536
rect 12438 5480 12494 5516
rect 12530 4972 12532 4992
rect 12532 4972 12584 4992
rect 12584 4972 12586 4992
rect 12530 4936 12586 4972
rect 13951 19066 14007 19068
rect 14031 19066 14087 19068
rect 14111 19066 14167 19068
rect 14191 19066 14247 19068
rect 13951 19014 13997 19066
rect 13997 19014 14007 19066
rect 14031 19014 14061 19066
rect 14061 19014 14073 19066
rect 14073 19014 14087 19066
rect 14111 19014 14125 19066
rect 14125 19014 14137 19066
rect 14137 19014 14167 19066
rect 14191 19014 14201 19066
rect 14201 19014 14247 19066
rect 13951 19012 14007 19014
rect 14031 19012 14087 19014
rect 14111 19012 14167 19014
rect 14191 19012 14247 19014
rect 13951 17978 14007 17980
rect 14031 17978 14087 17980
rect 14111 17978 14167 17980
rect 14191 17978 14247 17980
rect 13951 17926 13997 17978
rect 13997 17926 14007 17978
rect 14031 17926 14061 17978
rect 14061 17926 14073 17978
rect 14073 17926 14087 17978
rect 14111 17926 14125 17978
rect 14125 17926 14137 17978
rect 14137 17926 14167 17978
rect 14191 17926 14201 17978
rect 14201 17926 14247 17978
rect 13951 17924 14007 17926
rect 14031 17924 14087 17926
rect 14111 17924 14167 17926
rect 14191 17924 14247 17926
rect 13951 16890 14007 16892
rect 14031 16890 14087 16892
rect 14111 16890 14167 16892
rect 14191 16890 14247 16892
rect 13951 16838 13997 16890
rect 13997 16838 14007 16890
rect 14031 16838 14061 16890
rect 14061 16838 14073 16890
rect 14073 16838 14087 16890
rect 14111 16838 14125 16890
rect 14125 16838 14137 16890
rect 14137 16838 14167 16890
rect 14191 16838 14201 16890
rect 14201 16838 14247 16890
rect 13951 16836 14007 16838
rect 14031 16836 14087 16838
rect 14111 16836 14167 16838
rect 14191 16836 14247 16838
rect 13951 15802 14007 15804
rect 14031 15802 14087 15804
rect 14111 15802 14167 15804
rect 14191 15802 14247 15804
rect 13951 15750 13997 15802
rect 13997 15750 14007 15802
rect 14031 15750 14061 15802
rect 14061 15750 14073 15802
rect 14073 15750 14087 15802
rect 14111 15750 14125 15802
rect 14125 15750 14137 15802
rect 14137 15750 14167 15802
rect 14191 15750 14201 15802
rect 14201 15750 14247 15802
rect 13951 15748 14007 15750
rect 14031 15748 14087 15750
rect 14111 15748 14167 15750
rect 14191 15748 14247 15750
rect 14278 15000 14334 15056
rect 13951 14714 14007 14716
rect 14031 14714 14087 14716
rect 14111 14714 14167 14716
rect 14191 14714 14247 14716
rect 13951 14662 13997 14714
rect 13997 14662 14007 14714
rect 14031 14662 14061 14714
rect 14061 14662 14073 14714
rect 14073 14662 14087 14714
rect 14111 14662 14125 14714
rect 14125 14662 14137 14714
rect 14137 14662 14167 14714
rect 14191 14662 14201 14714
rect 14201 14662 14247 14714
rect 13951 14660 14007 14662
rect 14031 14660 14087 14662
rect 14111 14660 14167 14662
rect 14191 14660 14247 14662
rect 13951 13626 14007 13628
rect 14031 13626 14087 13628
rect 14111 13626 14167 13628
rect 14191 13626 14247 13628
rect 13951 13574 13997 13626
rect 13997 13574 14007 13626
rect 14031 13574 14061 13626
rect 14061 13574 14073 13626
rect 14073 13574 14087 13626
rect 14111 13574 14125 13626
rect 14125 13574 14137 13626
rect 14137 13574 14167 13626
rect 14191 13574 14201 13626
rect 14201 13574 14247 13626
rect 13951 13572 14007 13574
rect 14031 13572 14087 13574
rect 14111 13572 14167 13574
rect 14191 13572 14247 13574
rect 13951 12538 14007 12540
rect 14031 12538 14087 12540
rect 14111 12538 14167 12540
rect 14191 12538 14247 12540
rect 13951 12486 13997 12538
rect 13997 12486 14007 12538
rect 14031 12486 14061 12538
rect 14061 12486 14073 12538
rect 14073 12486 14087 12538
rect 14111 12486 14125 12538
rect 14125 12486 14137 12538
rect 14137 12486 14167 12538
rect 14191 12486 14201 12538
rect 14201 12486 14247 12538
rect 13951 12484 14007 12486
rect 14031 12484 14087 12486
rect 14111 12484 14167 12486
rect 14191 12484 14247 12486
rect 13450 10240 13506 10296
rect 13266 9288 13322 9344
rect 13174 8472 13230 8528
rect 13082 5072 13138 5128
rect 13542 8900 13598 8936
rect 13542 8880 13544 8900
rect 13544 8880 13596 8900
rect 13596 8880 13598 8900
rect 13542 8472 13598 8528
rect 13951 11450 14007 11452
rect 14031 11450 14087 11452
rect 14111 11450 14167 11452
rect 14191 11450 14247 11452
rect 13951 11398 13997 11450
rect 13997 11398 14007 11450
rect 14031 11398 14061 11450
rect 14061 11398 14073 11450
rect 14073 11398 14087 11450
rect 14111 11398 14125 11450
rect 14125 11398 14137 11450
rect 14137 11398 14167 11450
rect 14191 11398 14201 11450
rect 14201 11398 14247 11450
rect 13951 11396 14007 11398
rect 14031 11396 14087 11398
rect 14111 11396 14167 11398
rect 14191 11396 14247 11398
rect 13951 10362 14007 10364
rect 14031 10362 14087 10364
rect 14111 10362 14167 10364
rect 14191 10362 14247 10364
rect 13951 10310 13997 10362
rect 13997 10310 14007 10362
rect 14031 10310 14061 10362
rect 14061 10310 14073 10362
rect 14073 10310 14087 10362
rect 14111 10310 14125 10362
rect 14125 10310 14137 10362
rect 14137 10310 14167 10362
rect 14191 10310 14201 10362
rect 14201 10310 14247 10362
rect 13951 10308 14007 10310
rect 14031 10308 14087 10310
rect 14111 10308 14167 10310
rect 14191 10308 14247 10310
rect 13818 9560 13874 9616
rect 14002 9444 14058 9480
rect 14002 9424 14004 9444
rect 14004 9424 14056 9444
rect 14056 9424 14058 9444
rect 13951 9274 14007 9276
rect 14031 9274 14087 9276
rect 14111 9274 14167 9276
rect 14191 9274 14247 9276
rect 13951 9222 13997 9274
rect 13997 9222 14007 9274
rect 14031 9222 14061 9274
rect 14061 9222 14073 9274
rect 14073 9222 14087 9274
rect 14111 9222 14125 9274
rect 14125 9222 14137 9274
rect 14137 9222 14167 9274
rect 14191 9222 14201 9274
rect 14201 9222 14247 9274
rect 13951 9220 14007 9222
rect 14031 9220 14087 9222
rect 14111 9220 14167 9222
rect 14191 9220 14247 9222
rect 13951 8186 14007 8188
rect 14031 8186 14087 8188
rect 14111 8186 14167 8188
rect 14191 8186 14247 8188
rect 13951 8134 13997 8186
rect 13997 8134 14007 8186
rect 14031 8134 14061 8186
rect 14061 8134 14073 8186
rect 14073 8134 14087 8186
rect 14111 8134 14125 8186
rect 14125 8134 14137 8186
rect 14137 8134 14167 8186
rect 14191 8134 14201 8186
rect 14201 8134 14247 8186
rect 13951 8132 14007 8134
rect 14031 8132 14087 8134
rect 14111 8132 14167 8134
rect 14191 8132 14247 8134
rect 13726 8084 13782 8120
rect 13726 8064 13728 8084
rect 13728 8064 13780 8084
rect 13780 8064 13782 8084
rect 16550 20698 16606 20700
rect 16630 20698 16686 20700
rect 16710 20698 16766 20700
rect 16790 20698 16846 20700
rect 16550 20646 16596 20698
rect 16596 20646 16606 20698
rect 16630 20646 16660 20698
rect 16660 20646 16672 20698
rect 16672 20646 16686 20698
rect 16710 20646 16724 20698
rect 16724 20646 16736 20698
rect 16736 20646 16766 20698
rect 16790 20646 16800 20698
rect 16800 20646 16846 20698
rect 16550 20644 16606 20646
rect 16630 20644 16686 20646
rect 16710 20644 16766 20646
rect 16790 20644 16846 20646
rect 16550 19610 16606 19612
rect 16630 19610 16686 19612
rect 16710 19610 16766 19612
rect 16790 19610 16846 19612
rect 16550 19558 16596 19610
rect 16596 19558 16606 19610
rect 16630 19558 16660 19610
rect 16660 19558 16672 19610
rect 16672 19558 16686 19610
rect 16710 19558 16724 19610
rect 16724 19558 16736 19610
rect 16736 19558 16766 19610
rect 16790 19558 16800 19610
rect 16800 19558 16846 19610
rect 16550 19556 16606 19558
rect 16630 19556 16686 19558
rect 16710 19556 16766 19558
rect 16790 19556 16846 19558
rect 19149 20154 19205 20156
rect 19229 20154 19285 20156
rect 19309 20154 19365 20156
rect 19389 20154 19445 20156
rect 19149 20102 19195 20154
rect 19195 20102 19205 20154
rect 19229 20102 19259 20154
rect 19259 20102 19271 20154
rect 19271 20102 19285 20154
rect 19309 20102 19323 20154
rect 19323 20102 19335 20154
rect 19335 20102 19365 20154
rect 19389 20102 19399 20154
rect 19399 20102 19445 20154
rect 19149 20100 19205 20102
rect 19229 20100 19285 20102
rect 19309 20100 19365 20102
rect 19389 20100 19445 20102
rect 19149 19066 19205 19068
rect 19229 19066 19285 19068
rect 19309 19066 19365 19068
rect 19389 19066 19445 19068
rect 19149 19014 19195 19066
rect 19195 19014 19205 19066
rect 19229 19014 19259 19066
rect 19259 19014 19271 19066
rect 19271 19014 19285 19066
rect 19309 19014 19323 19066
rect 19323 19014 19335 19066
rect 19335 19014 19365 19066
rect 19389 19014 19399 19066
rect 19399 19014 19445 19066
rect 19149 19012 19205 19014
rect 19229 19012 19285 19014
rect 19309 19012 19365 19014
rect 19389 19012 19445 19014
rect 18602 18808 18658 18864
rect 15382 18128 15438 18184
rect 19522 18672 19578 18728
rect 16550 18522 16606 18524
rect 16630 18522 16686 18524
rect 16710 18522 16766 18524
rect 16790 18522 16846 18524
rect 16550 18470 16596 18522
rect 16596 18470 16606 18522
rect 16630 18470 16660 18522
rect 16660 18470 16672 18522
rect 16672 18470 16686 18522
rect 16710 18470 16724 18522
rect 16724 18470 16736 18522
rect 16736 18470 16766 18522
rect 16790 18470 16800 18522
rect 16800 18470 16846 18522
rect 16550 18468 16606 18470
rect 16630 18468 16686 18470
rect 16710 18468 16766 18470
rect 16790 18468 16846 18470
rect 14554 12688 14610 12744
rect 15014 14864 15070 14920
rect 16550 17434 16606 17436
rect 16630 17434 16686 17436
rect 16710 17434 16766 17436
rect 16790 17434 16846 17436
rect 16550 17382 16596 17434
rect 16596 17382 16606 17434
rect 16630 17382 16660 17434
rect 16660 17382 16672 17434
rect 16672 17382 16686 17434
rect 16710 17382 16724 17434
rect 16724 17382 16736 17434
rect 16736 17382 16766 17434
rect 16790 17382 16800 17434
rect 16800 17382 16846 17434
rect 16550 17380 16606 17382
rect 16630 17380 16686 17382
rect 16710 17380 16766 17382
rect 16790 17380 16846 17382
rect 16210 17196 16266 17232
rect 16210 17176 16212 17196
rect 16212 17176 16264 17196
rect 16264 17176 16266 17196
rect 16118 17040 16174 17096
rect 19149 17978 19205 17980
rect 19229 17978 19285 17980
rect 19309 17978 19365 17980
rect 19389 17978 19445 17980
rect 19149 17926 19195 17978
rect 19195 17926 19205 17978
rect 19229 17926 19259 17978
rect 19259 17926 19271 17978
rect 19271 17926 19285 17978
rect 19309 17926 19323 17978
rect 19323 17926 19335 17978
rect 19335 17926 19365 17978
rect 19389 17926 19399 17978
rect 19399 17926 19445 17978
rect 19149 17924 19205 17926
rect 19229 17924 19285 17926
rect 19309 17924 19365 17926
rect 19389 17924 19445 17926
rect 20902 20304 20958 20360
rect 19982 19216 20038 19272
rect 19614 17720 19670 17776
rect 19614 17176 19670 17232
rect 17866 16496 17922 16552
rect 16550 16346 16606 16348
rect 16630 16346 16686 16348
rect 16710 16346 16766 16348
rect 16790 16346 16846 16348
rect 16550 16294 16596 16346
rect 16596 16294 16606 16346
rect 16630 16294 16660 16346
rect 16660 16294 16672 16346
rect 16672 16294 16686 16346
rect 16710 16294 16724 16346
rect 16724 16294 16736 16346
rect 16736 16294 16766 16346
rect 16790 16294 16800 16346
rect 16800 16294 16846 16346
rect 16550 16292 16606 16294
rect 16630 16292 16686 16294
rect 16710 16292 16766 16294
rect 16790 16292 16846 16294
rect 16550 15258 16606 15260
rect 16630 15258 16686 15260
rect 16710 15258 16766 15260
rect 16790 15258 16846 15260
rect 16550 15206 16596 15258
rect 16596 15206 16606 15258
rect 16630 15206 16660 15258
rect 16660 15206 16672 15258
rect 16672 15206 16686 15258
rect 16710 15206 16724 15258
rect 16724 15206 16736 15258
rect 16736 15206 16766 15258
rect 16790 15206 16800 15258
rect 16800 15206 16846 15258
rect 16550 15204 16606 15206
rect 16630 15204 16686 15206
rect 16710 15204 16766 15206
rect 16790 15204 16846 15206
rect 14738 12144 14794 12200
rect 14554 10104 14610 10160
rect 14738 9968 14794 10024
rect 14278 7928 14334 7984
rect 13634 7384 13690 7440
rect 13951 7098 14007 7100
rect 14031 7098 14087 7100
rect 14111 7098 14167 7100
rect 14191 7098 14247 7100
rect 13951 7046 13997 7098
rect 13997 7046 14007 7098
rect 14031 7046 14061 7098
rect 14061 7046 14073 7098
rect 14073 7046 14087 7098
rect 14111 7046 14125 7098
rect 14125 7046 14137 7098
rect 14137 7046 14167 7098
rect 14191 7046 14201 7098
rect 14201 7046 14247 7098
rect 13951 7044 14007 7046
rect 14031 7044 14087 7046
rect 14111 7044 14167 7046
rect 14191 7044 14247 7046
rect 13634 6024 13690 6080
rect 13542 5208 13598 5264
rect 12714 4120 12770 4176
rect 13951 6010 14007 6012
rect 14031 6010 14087 6012
rect 14111 6010 14167 6012
rect 14191 6010 14247 6012
rect 13951 5958 13997 6010
rect 13997 5958 14007 6010
rect 14031 5958 14061 6010
rect 14061 5958 14073 6010
rect 14073 5958 14087 6010
rect 14111 5958 14125 6010
rect 14125 5958 14137 6010
rect 14137 5958 14167 6010
rect 14191 5958 14201 6010
rect 14201 5958 14247 6010
rect 13951 5956 14007 5958
rect 14031 5956 14087 5958
rect 14111 5956 14167 5958
rect 14191 5956 14247 5958
rect 13951 4922 14007 4924
rect 14031 4922 14087 4924
rect 14111 4922 14167 4924
rect 14191 4922 14247 4924
rect 13951 4870 13997 4922
rect 13997 4870 14007 4922
rect 14031 4870 14061 4922
rect 14061 4870 14073 4922
rect 14073 4870 14087 4922
rect 14111 4870 14125 4922
rect 14125 4870 14137 4922
rect 14137 4870 14167 4922
rect 14191 4870 14201 4922
rect 14201 4870 14247 4922
rect 13951 4868 14007 4870
rect 14031 4868 14087 4870
rect 14111 4868 14167 4870
rect 14191 4868 14247 4870
rect 13951 3834 14007 3836
rect 14031 3834 14087 3836
rect 14111 3834 14167 3836
rect 14191 3834 14247 3836
rect 13951 3782 13997 3834
rect 13997 3782 14007 3834
rect 14031 3782 14061 3834
rect 14061 3782 14073 3834
rect 14073 3782 14087 3834
rect 14111 3782 14125 3834
rect 14125 3782 14137 3834
rect 14137 3782 14167 3834
rect 14191 3782 14201 3834
rect 14201 3782 14247 3834
rect 13951 3780 14007 3782
rect 14031 3780 14087 3782
rect 14111 3780 14167 3782
rect 14191 3780 14247 3782
rect 14646 4664 14702 4720
rect 15198 3984 15254 4040
rect 15382 8492 15438 8528
rect 15382 8472 15384 8492
rect 15384 8472 15436 8492
rect 15436 8472 15438 8492
rect 16550 14170 16606 14172
rect 16630 14170 16686 14172
rect 16710 14170 16766 14172
rect 16790 14170 16846 14172
rect 16550 14118 16596 14170
rect 16596 14118 16606 14170
rect 16630 14118 16660 14170
rect 16660 14118 16672 14170
rect 16672 14118 16686 14170
rect 16710 14118 16724 14170
rect 16724 14118 16736 14170
rect 16736 14118 16766 14170
rect 16790 14118 16800 14170
rect 16800 14118 16846 14170
rect 16550 14116 16606 14118
rect 16630 14116 16686 14118
rect 16710 14116 16766 14118
rect 16790 14116 16846 14118
rect 16550 13082 16606 13084
rect 16630 13082 16686 13084
rect 16710 13082 16766 13084
rect 16790 13082 16846 13084
rect 16550 13030 16596 13082
rect 16596 13030 16606 13082
rect 16630 13030 16660 13082
rect 16660 13030 16672 13082
rect 16672 13030 16686 13082
rect 16710 13030 16724 13082
rect 16724 13030 16736 13082
rect 16736 13030 16766 13082
rect 16790 13030 16800 13082
rect 16800 13030 16846 13082
rect 16550 13028 16606 13030
rect 16630 13028 16686 13030
rect 16710 13028 16766 13030
rect 16790 13028 16846 13030
rect 16578 12688 16634 12744
rect 16550 11994 16606 11996
rect 16630 11994 16686 11996
rect 16710 11994 16766 11996
rect 16790 11994 16846 11996
rect 16550 11942 16596 11994
rect 16596 11942 16606 11994
rect 16630 11942 16660 11994
rect 16660 11942 16672 11994
rect 16672 11942 16686 11994
rect 16710 11942 16724 11994
rect 16724 11942 16736 11994
rect 16736 11942 16766 11994
rect 16790 11942 16800 11994
rect 16800 11942 16846 11994
rect 16550 11940 16606 11942
rect 16630 11940 16686 11942
rect 16710 11940 16766 11942
rect 16790 11940 16846 11942
rect 16550 10906 16606 10908
rect 16630 10906 16686 10908
rect 16710 10906 16766 10908
rect 16790 10906 16846 10908
rect 16550 10854 16596 10906
rect 16596 10854 16606 10906
rect 16630 10854 16660 10906
rect 16660 10854 16672 10906
rect 16672 10854 16686 10906
rect 16710 10854 16724 10906
rect 16724 10854 16736 10906
rect 16736 10854 16766 10906
rect 16790 10854 16800 10906
rect 16800 10854 16846 10906
rect 16550 10852 16606 10854
rect 16630 10852 16686 10854
rect 16710 10852 16766 10854
rect 16790 10852 16846 10854
rect 16210 9560 16266 9616
rect 15750 5752 15806 5808
rect 15290 3440 15346 3496
rect 13951 2746 14007 2748
rect 14031 2746 14087 2748
rect 14111 2746 14167 2748
rect 14191 2746 14247 2748
rect 13951 2694 13997 2746
rect 13997 2694 14007 2746
rect 14031 2694 14061 2746
rect 14061 2694 14073 2746
rect 14073 2694 14087 2746
rect 14111 2694 14125 2746
rect 14125 2694 14137 2746
rect 14137 2694 14167 2746
rect 14191 2694 14201 2746
rect 14201 2694 14247 2746
rect 13951 2692 14007 2694
rect 14031 2692 14087 2694
rect 14111 2692 14167 2694
rect 14191 2692 14247 2694
rect 16550 9818 16606 9820
rect 16630 9818 16686 9820
rect 16710 9818 16766 9820
rect 16790 9818 16846 9820
rect 16550 9766 16596 9818
rect 16596 9766 16606 9818
rect 16630 9766 16660 9818
rect 16660 9766 16672 9818
rect 16672 9766 16686 9818
rect 16710 9766 16724 9818
rect 16724 9766 16736 9818
rect 16736 9766 16766 9818
rect 16790 9766 16800 9818
rect 16800 9766 16846 9818
rect 16550 9764 16606 9766
rect 16630 9764 16686 9766
rect 16710 9764 16766 9766
rect 16790 9764 16846 9766
rect 16550 8730 16606 8732
rect 16630 8730 16686 8732
rect 16710 8730 16766 8732
rect 16790 8730 16846 8732
rect 16550 8678 16596 8730
rect 16596 8678 16606 8730
rect 16630 8678 16660 8730
rect 16660 8678 16672 8730
rect 16672 8678 16686 8730
rect 16710 8678 16724 8730
rect 16724 8678 16736 8730
rect 16736 8678 16766 8730
rect 16790 8678 16800 8730
rect 16800 8678 16846 8730
rect 16550 8676 16606 8678
rect 16630 8676 16686 8678
rect 16710 8676 16766 8678
rect 16790 8676 16846 8678
rect 16550 7642 16606 7644
rect 16630 7642 16686 7644
rect 16710 7642 16766 7644
rect 16790 7642 16846 7644
rect 16550 7590 16596 7642
rect 16596 7590 16606 7642
rect 16630 7590 16660 7642
rect 16660 7590 16672 7642
rect 16672 7590 16686 7642
rect 16710 7590 16724 7642
rect 16724 7590 16736 7642
rect 16736 7590 16766 7642
rect 16790 7590 16800 7642
rect 16800 7590 16846 7642
rect 16550 7588 16606 7590
rect 16630 7588 16686 7590
rect 16710 7588 16766 7590
rect 16790 7588 16846 7590
rect 17130 10648 17186 10704
rect 16946 7248 17002 7304
rect 16394 7112 16450 7168
rect 16946 6704 17002 6760
rect 16550 6554 16606 6556
rect 16630 6554 16686 6556
rect 16710 6554 16766 6556
rect 16790 6554 16846 6556
rect 16550 6502 16596 6554
rect 16596 6502 16606 6554
rect 16630 6502 16660 6554
rect 16660 6502 16672 6554
rect 16672 6502 16686 6554
rect 16710 6502 16724 6554
rect 16724 6502 16736 6554
rect 16736 6502 16766 6554
rect 16790 6502 16800 6554
rect 16800 6502 16846 6554
rect 16550 6500 16606 6502
rect 16630 6500 16686 6502
rect 16710 6500 16766 6502
rect 16790 6500 16846 6502
rect 16394 5516 16396 5536
rect 16396 5516 16448 5536
rect 16448 5516 16450 5536
rect 16394 5480 16450 5516
rect 16550 5466 16606 5468
rect 16630 5466 16686 5468
rect 16710 5466 16766 5468
rect 16790 5466 16846 5468
rect 16550 5414 16596 5466
rect 16596 5414 16606 5466
rect 16630 5414 16660 5466
rect 16660 5414 16672 5466
rect 16672 5414 16686 5466
rect 16710 5414 16724 5466
rect 16724 5414 16736 5466
rect 16736 5414 16766 5466
rect 16790 5414 16800 5466
rect 16800 5414 16846 5466
rect 16550 5412 16606 5414
rect 16630 5412 16686 5414
rect 16710 5412 16766 5414
rect 16790 5412 16846 5414
rect 16550 4378 16606 4380
rect 16630 4378 16686 4380
rect 16710 4378 16766 4380
rect 16790 4378 16846 4380
rect 16550 4326 16596 4378
rect 16596 4326 16606 4378
rect 16630 4326 16660 4378
rect 16660 4326 16672 4378
rect 16672 4326 16686 4378
rect 16710 4326 16724 4378
rect 16724 4326 16736 4378
rect 16736 4326 16766 4378
rect 16790 4326 16800 4378
rect 16800 4326 16846 4378
rect 16550 4324 16606 4326
rect 16630 4324 16686 4326
rect 16710 4324 16766 4326
rect 16790 4324 16846 4326
rect 16550 3290 16606 3292
rect 16630 3290 16686 3292
rect 16710 3290 16766 3292
rect 16790 3290 16846 3292
rect 16550 3238 16596 3290
rect 16596 3238 16606 3290
rect 16630 3238 16660 3290
rect 16660 3238 16672 3290
rect 16672 3238 16686 3290
rect 16710 3238 16724 3290
rect 16724 3238 16736 3290
rect 16736 3238 16766 3290
rect 16790 3238 16800 3290
rect 16800 3238 16846 3290
rect 16550 3236 16606 3238
rect 16630 3236 16686 3238
rect 16710 3236 16766 3238
rect 16790 3236 16846 3238
rect 18970 14456 19026 14512
rect 19149 16890 19205 16892
rect 19229 16890 19285 16892
rect 19309 16890 19365 16892
rect 19389 16890 19445 16892
rect 19149 16838 19195 16890
rect 19195 16838 19205 16890
rect 19229 16838 19259 16890
rect 19259 16838 19271 16890
rect 19271 16838 19285 16890
rect 19309 16838 19323 16890
rect 19323 16838 19335 16890
rect 19335 16838 19365 16890
rect 19389 16838 19399 16890
rect 19399 16838 19445 16890
rect 19149 16836 19205 16838
rect 19229 16836 19285 16838
rect 19309 16836 19365 16838
rect 19389 16836 19445 16838
rect 19149 15802 19205 15804
rect 19229 15802 19285 15804
rect 19309 15802 19365 15804
rect 19389 15802 19445 15804
rect 19149 15750 19195 15802
rect 19195 15750 19205 15802
rect 19229 15750 19259 15802
rect 19259 15750 19271 15802
rect 19271 15750 19285 15802
rect 19309 15750 19323 15802
rect 19323 15750 19335 15802
rect 19335 15750 19365 15802
rect 19389 15750 19399 15802
rect 19399 15750 19445 15802
rect 19149 15748 19205 15750
rect 19229 15748 19285 15750
rect 19309 15748 19365 15750
rect 19389 15748 19445 15750
rect 20902 18264 20958 18320
rect 21748 20698 21804 20700
rect 21828 20698 21884 20700
rect 21908 20698 21964 20700
rect 21988 20698 22044 20700
rect 21748 20646 21794 20698
rect 21794 20646 21804 20698
rect 21828 20646 21858 20698
rect 21858 20646 21870 20698
rect 21870 20646 21884 20698
rect 21908 20646 21922 20698
rect 21922 20646 21934 20698
rect 21934 20646 21964 20698
rect 21988 20646 21998 20698
rect 21998 20646 22044 20698
rect 21748 20644 21804 20646
rect 21828 20644 21884 20646
rect 21908 20644 21964 20646
rect 21988 20644 22044 20646
rect 21748 19610 21804 19612
rect 21828 19610 21884 19612
rect 21908 19610 21964 19612
rect 21988 19610 22044 19612
rect 21748 19558 21794 19610
rect 21794 19558 21804 19610
rect 21828 19558 21858 19610
rect 21858 19558 21870 19610
rect 21870 19558 21884 19610
rect 21908 19558 21922 19610
rect 21922 19558 21934 19610
rect 21934 19558 21964 19610
rect 21988 19558 21998 19610
rect 21998 19558 22044 19610
rect 21748 19556 21804 19558
rect 21828 19556 21884 19558
rect 21908 19556 21964 19558
rect 21988 19556 22044 19558
rect 21748 18522 21804 18524
rect 21828 18522 21884 18524
rect 21908 18522 21964 18524
rect 21988 18522 22044 18524
rect 21748 18470 21794 18522
rect 21794 18470 21804 18522
rect 21828 18470 21858 18522
rect 21858 18470 21870 18522
rect 21870 18470 21884 18522
rect 21908 18470 21922 18522
rect 21922 18470 21934 18522
rect 21934 18470 21964 18522
rect 21988 18470 21998 18522
rect 21998 18470 22044 18522
rect 21748 18468 21804 18470
rect 21828 18468 21884 18470
rect 21908 18468 21964 18470
rect 21988 18468 22044 18470
rect 19149 14714 19205 14716
rect 19229 14714 19285 14716
rect 19309 14714 19365 14716
rect 19389 14714 19445 14716
rect 19149 14662 19195 14714
rect 19195 14662 19205 14714
rect 19229 14662 19259 14714
rect 19259 14662 19271 14714
rect 19271 14662 19285 14714
rect 19309 14662 19323 14714
rect 19323 14662 19335 14714
rect 19335 14662 19365 14714
rect 19389 14662 19399 14714
rect 19399 14662 19445 14714
rect 19149 14660 19205 14662
rect 19229 14660 19285 14662
rect 19309 14660 19365 14662
rect 19389 14660 19445 14662
rect 17958 12824 18014 12880
rect 19149 13626 19205 13628
rect 19229 13626 19285 13628
rect 19309 13626 19365 13628
rect 19389 13626 19445 13628
rect 19149 13574 19195 13626
rect 19195 13574 19205 13626
rect 19229 13574 19259 13626
rect 19259 13574 19271 13626
rect 19271 13574 19285 13626
rect 19309 13574 19323 13626
rect 19323 13574 19335 13626
rect 19335 13574 19365 13626
rect 19389 13574 19399 13626
rect 19399 13574 19445 13626
rect 19149 13572 19205 13574
rect 19229 13572 19285 13574
rect 19309 13572 19365 13574
rect 19389 13572 19445 13574
rect 19522 13368 19578 13424
rect 19149 12538 19205 12540
rect 19229 12538 19285 12540
rect 19309 12538 19365 12540
rect 19389 12538 19445 12540
rect 19149 12486 19195 12538
rect 19195 12486 19205 12538
rect 19229 12486 19259 12538
rect 19259 12486 19271 12538
rect 19271 12486 19285 12538
rect 19309 12486 19323 12538
rect 19323 12486 19335 12538
rect 19335 12486 19365 12538
rect 19389 12486 19399 12538
rect 19399 12486 19445 12538
rect 19149 12484 19205 12486
rect 19229 12484 19285 12486
rect 19309 12484 19365 12486
rect 19389 12484 19445 12486
rect 18970 12280 19026 12336
rect 17222 9424 17278 9480
rect 17222 5072 17278 5128
rect 18142 8200 18198 8256
rect 17774 7792 17830 7848
rect 17682 7384 17738 7440
rect 17958 7112 18014 7168
rect 17682 2896 17738 2952
rect 16550 2202 16606 2204
rect 16630 2202 16686 2204
rect 16710 2202 16766 2204
rect 16790 2202 16846 2204
rect 16550 2150 16596 2202
rect 16596 2150 16606 2202
rect 16630 2150 16660 2202
rect 16660 2150 16672 2202
rect 16672 2150 16686 2202
rect 16710 2150 16724 2202
rect 16724 2150 16736 2202
rect 16736 2150 16766 2202
rect 16790 2150 16800 2202
rect 16800 2150 16846 2202
rect 16550 2148 16606 2150
rect 16630 2148 16686 2150
rect 16710 2148 16766 2150
rect 16790 2148 16846 2150
rect 19149 11450 19205 11452
rect 19229 11450 19285 11452
rect 19309 11450 19365 11452
rect 19389 11450 19445 11452
rect 19149 11398 19195 11450
rect 19195 11398 19205 11450
rect 19229 11398 19259 11450
rect 19259 11398 19271 11450
rect 19271 11398 19285 11450
rect 19309 11398 19323 11450
rect 19323 11398 19335 11450
rect 19335 11398 19365 11450
rect 19389 11398 19399 11450
rect 19399 11398 19445 11450
rect 19149 11396 19205 11398
rect 19229 11396 19285 11398
rect 19309 11396 19365 11398
rect 19389 11396 19445 11398
rect 19149 10362 19205 10364
rect 19229 10362 19285 10364
rect 19309 10362 19365 10364
rect 19389 10362 19445 10364
rect 19149 10310 19195 10362
rect 19195 10310 19205 10362
rect 19229 10310 19259 10362
rect 19259 10310 19271 10362
rect 19271 10310 19285 10362
rect 19309 10310 19323 10362
rect 19323 10310 19335 10362
rect 19335 10310 19365 10362
rect 19389 10310 19399 10362
rect 19399 10310 19445 10362
rect 19149 10308 19205 10310
rect 19229 10308 19285 10310
rect 19309 10308 19365 10310
rect 19389 10308 19445 10310
rect 19149 9274 19205 9276
rect 19229 9274 19285 9276
rect 19309 9274 19365 9276
rect 19389 9274 19445 9276
rect 19149 9222 19195 9274
rect 19195 9222 19205 9274
rect 19229 9222 19259 9274
rect 19259 9222 19271 9274
rect 19271 9222 19285 9274
rect 19309 9222 19323 9274
rect 19323 9222 19335 9274
rect 19335 9222 19365 9274
rect 19389 9222 19399 9274
rect 19399 9222 19445 9274
rect 19149 9220 19205 9222
rect 19229 9220 19285 9222
rect 19309 9220 19365 9222
rect 19389 9220 19445 9222
rect 18878 8200 18934 8256
rect 19149 8186 19205 8188
rect 19229 8186 19285 8188
rect 19309 8186 19365 8188
rect 19389 8186 19445 8188
rect 19149 8134 19195 8186
rect 19195 8134 19205 8186
rect 19229 8134 19259 8186
rect 19259 8134 19271 8186
rect 19271 8134 19285 8186
rect 19309 8134 19323 8186
rect 19323 8134 19335 8186
rect 19335 8134 19365 8186
rect 19389 8134 19399 8186
rect 19399 8134 19445 8186
rect 19149 8132 19205 8134
rect 19229 8132 19285 8134
rect 19309 8132 19365 8134
rect 19389 8132 19445 8134
rect 19798 11736 19854 11792
rect 19149 7098 19205 7100
rect 19229 7098 19285 7100
rect 19309 7098 19365 7100
rect 19389 7098 19445 7100
rect 19149 7046 19195 7098
rect 19195 7046 19205 7098
rect 19229 7046 19259 7098
rect 19259 7046 19271 7098
rect 19271 7046 19285 7098
rect 19309 7046 19323 7098
rect 19323 7046 19335 7098
rect 19335 7046 19365 7098
rect 19389 7046 19399 7098
rect 19399 7046 19445 7098
rect 19149 7044 19205 7046
rect 19229 7044 19285 7046
rect 19309 7044 19365 7046
rect 19389 7044 19445 7046
rect 19149 6010 19205 6012
rect 19229 6010 19285 6012
rect 19309 6010 19365 6012
rect 19389 6010 19445 6012
rect 19149 5958 19195 6010
rect 19195 5958 19205 6010
rect 19229 5958 19259 6010
rect 19259 5958 19271 6010
rect 19271 5958 19285 6010
rect 19309 5958 19323 6010
rect 19323 5958 19335 6010
rect 19335 5958 19365 6010
rect 19389 5958 19399 6010
rect 19399 5958 19445 6010
rect 19149 5956 19205 5958
rect 19229 5956 19285 5958
rect 19309 5956 19365 5958
rect 19389 5956 19445 5958
rect 21748 17434 21804 17436
rect 21828 17434 21884 17436
rect 21908 17434 21964 17436
rect 21988 17434 22044 17436
rect 21748 17382 21794 17434
rect 21794 17382 21804 17434
rect 21828 17382 21858 17434
rect 21858 17382 21870 17434
rect 21870 17382 21884 17434
rect 21908 17382 21922 17434
rect 21922 17382 21934 17434
rect 21934 17382 21964 17434
rect 21988 17382 21998 17434
rect 21998 17382 22044 17434
rect 21748 17380 21804 17382
rect 21828 17380 21884 17382
rect 21908 17380 21964 17382
rect 21988 17380 22044 17382
rect 21086 16088 21142 16144
rect 21748 16346 21804 16348
rect 21828 16346 21884 16348
rect 21908 16346 21964 16348
rect 21988 16346 22044 16348
rect 21748 16294 21794 16346
rect 21794 16294 21804 16346
rect 21828 16294 21858 16346
rect 21858 16294 21870 16346
rect 21870 16294 21884 16346
rect 21908 16294 21922 16346
rect 21922 16294 21934 16346
rect 21934 16294 21964 16346
rect 21988 16294 21998 16346
rect 21998 16294 22044 16346
rect 21748 16292 21804 16294
rect 21828 16292 21884 16294
rect 21908 16292 21964 16294
rect 21988 16292 22044 16294
rect 20810 13368 20866 13424
rect 21748 15258 21804 15260
rect 21828 15258 21884 15260
rect 21908 15258 21964 15260
rect 21988 15258 22044 15260
rect 21748 15206 21794 15258
rect 21794 15206 21804 15258
rect 21828 15206 21858 15258
rect 21858 15206 21870 15258
rect 21870 15206 21884 15258
rect 21908 15206 21922 15258
rect 21922 15206 21934 15258
rect 21934 15206 21964 15258
rect 21988 15206 21998 15258
rect 21998 15206 22044 15258
rect 21748 15204 21804 15206
rect 21828 15204 21884 15206
rect 21908 15204 21964 15206
rect 21988 15204 22044 15206
rect 21748 14170 21804 14172
rect 21828 14170 21884 14172
rect 21908 14170 21964 14172
rect 21988 14170 22044 14172
rect 21748 14118 21794 14170
rect 21794 14118 21804 14170
rect 21828 14118 21858 14170
rect 21858 14118 21870 14170
rect 21870 14118 21884 14170
rect 21908 14118 21922 14170
rect 21922 14118 21934 14170
rect 21934 14118 21964 14170
rect 21988 14118 21998 14170
rect 21998 14118 22044 14170
rect 21748 14116 21804 14118
rect 21828 14116 21884 14118
rect 21908 14116 21964 14118
rect 21988 14116 22044 14118
rect 21748 13082 21804 13084
rect 21828 13082 21884 13084
rect 21908 13082 21964 13084
rect 21988 13082 22044 13084
rect 21748 13030 21794 13082
rect 21794 13030 21804 13082
rect 21828 13030 21858 13082
rect 21858 13030 21870 13082
rect 21870 13030 21884 13082
rect 21908 13030 21922 13082
rect 21922 13030 21934 13082
rect 21934 13030 21964 13082
rect 21988 13030 21998 13082
rect 21998 13030 22044 13082
rect 21748 13028 21804 13030
rect 21828 13028 21884 13030
rect 21908 13028 21964 13030
rect 21988 13028 22044 13030
rect 21748 11994 21804 11996
rect 21828 11994 21884 11996
rect 21908 11994 21964 11996
rect 21988 11994 22044 11996
rect 21748 11942 21794 11994
rect 21794 11942 21804 11994
rect 21828 11942 21858 11994
rect 21858 11942 21870 11994
rect 21870 11942 21884 11994
rect 21908 11942 21922 11994
rect 21922 11942 21934 11994
rect 21934 11942 21964 11994
rect 21988 11942 21998 11994
rect 21998 11942 22044 11994
rect 21748 11940 21804 11942
rect 21828 11940 21884 11942
rect 21908 11940 21964 11942
rect 21988 11940 22044 11942
rect 21748 10906 21804 10908
rect 21828 10906 21884 10908
rect 21908 10906 21964 10908
rect 21988 10906 22044 10908
rect 21748 10854 21794 10906
rect 21794 10854 21804 10906
rect 21828 10854 21858 10906
rect 21858 10854 21870 10906
rect 21870 10854 21884 10906
rect 21908 10854 21922 10906
rect 21922 10854 21934 10906
rect 21934 10854 21964 10906
rect 21988 10854 21998 10906
rect 21998 10854 22044 10906
rect 21748 10852 21804 10854
rect 21828 10852 21884 10854
rect 21908 10852 21964 10854
rect 21988 10852 22044 10854
rect 21748 9818 21804 9820
rect 21828 9818 21884 9820
rect 21908 9818 21964 9820
rect 21988 9818 22044 9820
rect 21748 9766 21794 9818
rect 21794 9766 21804 9818
rect 21828 9766 21858 9818
rect 21858 9766 21870 9818
rect 21870 9766 21884 9818
rect 21908 9766 21922 9818
rect 21922 9766 21934 9818
rect 21934 9766 21964 9818
rect 21988 9766 21998 9818
rect 21998 9766 22044 9818
rect 21748 9764 21804 9766
rect 21828 9764 21884 9766
rect 21908 9764 21964 9766
rect 21988 9764 22044 9766
rect 21748 8730 21804 8732
rect 21828 8730 21884 8732
rect 21908 8730 21964 8732
rect 21988 8730 22044 8732
rect 21748 8678 21794 8730
rect 21794 8678 21804 8730
rect 21828 8678 21858 8730
rect 21858 8678 21870 8730
rect 21870 8678 21884 8730
rect 21908 8678 21922 8730
rect 21922 8678 21934 8730
rect 21934 8678 21964 8730
rect 21988 8678 21998 8730
rect 21998 8678 22044 8730
rect 21748 8676 21804 8678
rect 21828 8676 21884 8678
rect 21908 8676 21964 8678
rect 21988 8676 22044 8678
rect 21748 7642 21804 7644
rect 21828 7642 21884 7644
rect 21908 7642 21964 7644
rect 21988 7642 22044 7644
rect 21748 7590 21794 7642
rect 21794 7590 21804 7642
rect 21828 7590 21858 7642
rect 21858 7590 21870 7642
rect 21870 7590 21884 7642
rect 21908 7590 21922 7642
rect 21922 7590 21934 7642
rect 21934 7590 21964 7642
rect 21988 7590 21998 7642
rect 21998 7590 22044 7642
rect 21748 7588 21804 7590
rect 21828 7588 21884 7590
rect 21908 7588 21964 7590
rect 21988 7588 22044 7590
rect 21748 6554 21804 6556
rect 21828 6554 21884 6556
rect 21908 6554 21964 6556
rect 21988 6554 22044 6556
rect 21748 6502 21794 6554
rect 21794 6502 21804 6554
rect 21828 6502 21858 6554
rect 21858 6502 21870 6554
rect 21870 6502 21884 6554
rect 21908 6502 21922 6554
rect 21922 6502 21934 6554
rect 21934 6502 21964 6554
rect 21988 6502 21998 6554
rect 21998 6502 22044 6554
rect 21748 6500 21804 6502
rect 21828 6500 21884 6502
rect 21908 6500 21964 6502
rect 21988 6500 22044 6502
rect 21362 5752 21418 5808
rect 19614 5072 19670 5128
rect 19149 4922 19205 4924
rect 19229 4922 19285 4924
rect 19309 4922 19365 4924
rect 19389 4922 19445 4924
rect 19149 4870 19195 4922
rect 19195 4870 19205 4922
rect 19229 4870 19259 4922
rect 19259 4870 19271 4922
rect 19271 4870 19285 4922
rect 19309 4870 19323 4922
rect 19323 4870 19335 4922
rect 19335 4870 19365 4922
rect 19389 4870 19399 4922
rect 19399 4870 19445 4922
rect 19149 4868 19205 4870
rect 19229 4868 19285 4870
rect 19309 4868 19365 4870
rect 19389 4868 19445 4870
rect 19149 3834 19205 3836
rect 19229 3834 19285 3836
rect 19309 3834 19365 3836
rect 19389 3834 19445 3836
rect 19149 3782 19195 3834
rect 19195 3782 19205 3834
rect 19229 3782 19259 3834
rect 19259 3782 19271 3834
rect 19271 3782 19285 3834
rect 19309 3782 19323 3834
rect 19323 3782 19335 3834
rect 19335 3782 19365 3834
rect 19389 3782 19399 3834
rect 19399 3782 19445 3834
rect 19149 3780 19205 3782
rect 19229 3780 19285 3782
rect 19309 3780 19365 3782
rect 19389 3780 19445 3782
rect 21748 5466 21804 5468
rect 21828 5466 21884 5468
rect 21908 5466 21964 5468
rect 21988 5466 22044 5468
rect 21748 5414 21794 5466
rect 21794 5414 21804 5466
rect 21828 5414 21858 5466
rect 21858 5414 21870 5466
rect 21870 5414 21884 5466
rect 21908 5414 21922 5466
rect 21922 5414 21934 5466
rect 21934 5414 21964 5466
rect 21988 5414 21998 5466
rect 21998 5414 22044 5466
rect 21748 5412 21804 5414
rect 21828 5412 21884 5414
rect 21908 5412 21964 5414
rect 21988 5412 22044 5414
rect 19149 2746 19205 2748
rect 19229 2746 19285 2748
rect 19309 2746 19365 2748
rect 19389 2746 19445 2748
rect 19149 2694 19195 2746
rect 19195 2694 19205 2746
rect 19229 2694 19259 2746
rect 19259 2694 19271 2746
rect 19271 2694 19285 2746
rect 19309 2694 19323 2746
rect 19323 2694 19335 2746
rect 19335 2694 19365 2746
rect 19389 2694 19399 2746
rect 19399 2694 19445 2746
rect 19149 2692 19205 2694
rect 19229 2692 19285 2694
rect 19309 2692 19365 2694
rect 19389 2692 19445 2694
rect 21748 4378 21804 4380
rect 21828 4378 21884 4380
rect 21908 4378 21964 4380
rect 21988 4378 22044 4380
rect 21748 4326 21794 4378
rect 21794 4326 21804 4378
rect 21828 4326 21858 4378
rect 21858 4326 21870 4378
rect 21870 4326 21884 4378
rect 21908 4326 21922 4378
rect 21922 4326 21934 4378
rect 21934 4326 21964 4378
rect 21988 4326 21998 4378
rect 21998 4326 22044 4378
rect 21748 4324 21804 4326
rect 21828 4324 21884 4326
rect 21908 4324 21964 4326
rect 21988 4324 22044 4326
rect 21748 3290 21804 3292
rect 21828 3290 21884 3292
rect 21908 3290 21964 3292
rect 21988 3290 22044 3292
rect 21748 3238 21794 3290
rect 21794 3238 21804 3290
rect 21828 3238 21858 3290
rect 21858 3238 21870 3290
rect 21870 3238 21884 3290
rect 21908 3238 21922 3290
rect 21922 3238 21934 3290
rect 21934 3238 21964 3290
rect 21988 3238 21998 3290
rect 21998 3238 22044 3290
rect 21748 3236 21804 3238
rect 21828 3236 21884 3238
rect 21908 3236 21964 3238
rect 21988 3236 22044 3238
rect 21748 2202 21804 2204
rect 21828 2202 21884 2204
rect 21908 2202 21964 2204
rect 21988 2202 22044 2204
rect 21748 2150 21794 2202
rect 21794 2150 21804 2202
rect 21828 2150 21858 2202
rect 21858 2150 21870 2202
rect 21870 2150 21884 2202
rect 21908 2150 21922 2202
rect 21922 2150 21934 2202
rect 21934 2150 21964 2202
rect 21988 2150 21998 2202
rect 21998 2150 22044 2202
rect 21748 2148 21804 2150
rect 21828 2148 21884 2150
rect 21908 2148 21964 2150
rect 21988 2148 22044 2150
<< metal3 >>
rect 0 21042 800 21072
rect 2773 21042 2839 21045
rect 0 21040 2839 21042
rect 0 20984 2778 21040
rect 2834 20984 2839 21040
rect 0 20982 2839 20984
rect 0 20952 800 20982
rect 2773 20979 2839 20982
rect 6144 20704 6460 20705
rect 0 20634 800 20664
rect 6144 20640 6150 20704
rect 6214 20640 6230 20704
rect 6294 20640 6310 20704
rect 6374 20640 6390 20704
rect 6454 20640 6460 20704
rect 6144 20639 6460 20640
rect 11342 20704 11658 20705
rect 11342 20640 11348 20704
rect 11412 20640 11428 20704
rect 11492 20640 11508 20704
rect 11572 20640 11588 20704
rect 11652 20640 11658 20704
rect 11342 20639 11658 20640
rect 16540 20704 16856 20705
rect 16540 20640 16546 20704
rect 16610 20640 16626 20704
rect 16690 20640 16706 20704
rect 16770 20640 16786 20704
rect 16850 20640 16856 20704
rect 16540 20639 16856 20640
rect 21738 20704 22054 20705
rect 21738 20640 21744 20704
rect 21808 20640 21824 20704
rect 21888 20640 21904 20704
rect 21968 20640 21984 20704
rect 22048 20640 22054 20704
rect 21738 20639 22054 20640
rect 2865 20634 2931 20637
rect 0 20632 2931 20634
rect 0 20576 2870 20632
rect 2926 20576 2931 20632
rect 0 20574 2931 20576
rect 0 20544 800 20574
rect 2865 20571 2931 20574
rect 9213 20362 9279 20365
rect 20897 20362 20963 20365
rect 9213 20360 20963 20362
rect 9213 20304 9218 20360
rect 9274 20304 20902 20360
rect 20958 20304 20963 20360
rect 9213 20302 20963 20304
rect 9213 20299 9279 20302
rect 20897 20299 20963 20302
rect 0 20226 800 20256
rect 2957 20226 3023 20229
rect 0 20224 3023 20226
rect 0 20168 2962 20224
rect 3018 20168 3023 20224
rect 0 20166 3023 20168
rect 0 20136 800 20166
rect 2957 20163 3023 20166
rect 3545 20160 3861 20161
rect 3545 20096 3551 20160
rect 3615 20096 3631 20160
rect 3695 20096 3711 20160
rect 3775 20096 3791 20160
rect 3855 20096 3861 20160
rect 3545 20095 3861 20096
rect 8743 20160 9059 20161
rect 8743 20096 8749 20160
rect 8813 20096 8829 20160
rect 8893 20096 8909 20160
rect 8973 20096 8989 20160
rect 9053 20096 9059 20160
rect 8743 20095 9059 20096
rect 13941 20160 14257 20161
rect 13941 20096 13947 20160
rect 14011 20096 14027 20160
rect 14091 20096 14107 20160
rect 14171 20096 14187 20160
rect 14251 20096 14257 20160
rect 13941 20095 14257 20096
rect 19139 20160 19455 20161
rect 19139 20096 19145 20160
rect 19209 20096 19225 20160
rect 19289 20096 19305 20160
rect 19369 20096 19385 20160
rect 19449 20096 19455 20160
rect 19139 20095 19455 20096
rect 0 19818 800 19848
rect 3049 19818 3115 19821
rect 0 19816 3115 19818
rect 0 19760 3054 19816
rect 3110 19760 3115 19816
rect 0 19758 3115 19760
rect 0 19728 800 19758
rect 3049 19755 3115 19758
rect 9949 19682 10015 19685
rect 11094 19682 11100 19684
rect 9949 19680 11100 19682
rect 9949 19624 9954 19680
rect 10010 19624 11100 19680
rect 9949 19622 11100 19624
rect 9949 19619 10015 19622
rect 11094 19620 11100 19622
rect 11164 19620 11170 19684
rect 6144 19616 6460 19617
rect 6144 19552 6150 19616
rect 6214 19552 6230 19616
rect 6294 19552 6310 19616
rect 6374 19552 6390 19616
rect 6454 19552 6460 19616
rect 6144 19551 6460 19552
rect 11342 19616 11658 19617
rect 11342 19552 11348 19616
rect 11412 19552 11428 19616
rect 11492 19552 11508 19616
rect 11572 19552 11588 19616
rect 11652 19552 11658 19616
rect 11342 19551 11658 19552
rect 16540 19616 16856 19617
rect 16540 19552 16546 19616
rect 16610 19552 16626 19616
rect 16690 19552 16706 19616
rect 16770 19552 16786 19616
rect 16850 19552 16856 19616
rect 16540 19551 16856 19552
rect 21738 19616 22054 19617
rect 21738 19552 21744 19616
rect 21808 19552 21824 19616
rect 21888 19552 21904 19616
rect 21968 19552 21984 19616
rect 22048 19552 22054 19616
rect 21738 19551 22054 19552
rect 0 19410 800 19440
rect 2773 19410 2839 19413
rect 0 19408 2839 19410
rect 0 19352 2778 19408
rect 2834 19352 2839 19408
rect 0 19350 2839 19352
rect 0 19320 800 19350
rect 2773 19347 2839 19350
rect 8293 19274 8359 19277
rect 19977 19274 20043 19277
rect 8293 19272 20043 19274
rect 8293 19216 8298 19272
rect 8354 19216 19982 19272
rect 20038 19216 20043 19272
rect 8293 19214 20043 19216
rect 8293 19211 8359 19214
rect 19977 19211 20043 19214
rect 9121 19138 9187 19141
rect 9438 19138 9444 19140
rect 9121 19136 9444 19138
rect 9121 19080 9126 19136
rect 9182 19080 9444 19136
rect 9121 19078 9444 19080
rect 9121 19075 9187 19078
rect 9438 19076 9444 19078
rect 9508 19076 9514 19140
rect 9806 19076 9812 19140
rect 9876 19138 9882 19140
rect 10041 19138 10107 19141
rect 9876 19136 10107 19138
rect 9876 19080 10046 19136
rect 10102 19080 10107 19136
rect 9876 19078 10107 19080
rect 9876 19076 9882 19078
rect 10041 19075 10107 19078
rect 3545 19072 3861 19073
rect 0 19002 800 19032
rect 3545 19008 3551 19072
rect 3615 19008 3631 19072
rect 3695 19008 3711 19072
rect 3775 19008 3791 19072
rect 3855 19008 3861 19072
rect 3545 19007 3861 19008
rect 8743 19072 9059 19073
rect 8743 19008 8749 19072
rect 8813 19008 8829 19072
rect 8893 19008 8909 19072
rect 8973 19008 8989 19072
rect 9053 19008 9059 19072
rect 8743 19007 9059 19008
rect 13941 19072 14257 19073
rect 13941 19008 13947 19072
rect 14011 19008 14027 19072
rect 14091 19008 14107 19072
rect 14171 19008 14187 19072
rect 14251 19008 14257 19072
rect 13941 19007 14257 19008
rect 19139 19072 19455 19073
rect 19139 19008 19145 19072
rect 19209 19008 19225 19072
rect 19289 19008 19305 19072
rect 19369 19008 19385 19072
rect 19449 19008 19455 19072
rect 19139 19007 19455 19008
rect 3233 19002 3299 19005
rect 0 19000 3299 19002
rect 0 18944 3238 19000
rect 3294 18944 3299 19000
rect 0 18942 3299 18944
rect 0 18912 800 18942
rect 3233 18939 3299 18942
rect 9673 19002 9739 19005
rect 12709 19002 12775 19005
rect 9673 19000 12775 19002
rect 9673 18944 9678 19000
rect 9734 18944 12714 19000
rect 12770 18944 12775 19000
rect 9673 18942 12775 18944
rect 9673 18939 9739 18942
rect 12709 18939 12775 18942
rect 8569 18866 8635 18869
rect 18597 18866 18663 18869
rect 8569 18864 18663 18866
rect 8569 18808 8574 18864
rect 8630 18808 18602 18864
rect 18658 18808 18663 18864
rect 8569 18806 18663 18808
rect 8569 18803 8635 18806
rect 18597 18803 18663 18806
rect 8293 18730 8359 18733
rect 19517 18730 19583 18733
rect 8293 18728 19583 18730
rect 8293 18672 8298 18728
rect 8354 18672 19522 18728
rect 19578 18672 19583 18728
rect 8293 18670 19583 18672
rect 8293 18667 8359 18670
rect 19517 18667 19583 18670
rect 0 18594 800 18624
rect 2814 18594 2820 18596
rect 0 18534 2820 18594
rect 0 18504 800 18534
rect 2814 18532 2820 18534
rect 2884 18532 2890 18596
rect 8017 18594 8083 18597
rect 10910 18594 10916 18596
rect 8017 18592 10916 18594
rect 8017 18536 8022 18592
rect 8078 18536 10916 18592
rect 8017 18534 10916 18536
rect 8017 18531 8083 18534
rect 10910 18532 10916 18534
rect 10980 18532 10986 18596
rect 6144 18528 6460 18529
rect 6144 18464 6150 18528
rect 6214 18464 6230 18528
rect 6294 18464 6310 18528
rect 6374 18464 6390 18528
rect 6454 18464 6460 18528
rect 6144 18463 6460 18464
rect 11342 18528 11658 18529
rect 11342 18464 11348 18528
rect 11412 18464 11428 18528
rect 11492 18464 11508 18528
rect 11572 18464 11588 18528
rect 11652 18464 11658 18528
rect 11342 18463 11658 18464
rect 16540 18528 16856 18529
rect 16540 18464 16546 18528
rect 16610 18464 16626 18528
rect 16690 18464 16706 18528
rect 16770 18464 16786 18528
rect 16850 18464 16856 18528
rect 16540 18463 16856 18464
rect 21738 18528 22054 18529
rect 21738 18464 21744 18528
rect 21808 18464 21824 18528
rect 21888 18464 21904 18528
rect 21968 18464 21984 18528
rect 22048 18464 22054 18528
rect 21738 18463 22054 18464
rect 8477 18458 8543 18461
rect 9254 18458 9260 18460
rect 8477 18456 9260 18458
rect 8477 18400 8482 18456
rect 8538 18400 9260 18456
rect 8477 18398 9260 18400
rect 8477 18395 8543 18398
rect 9254 18396 9260 18398
rect 9324 18396 9330 18460
rect 9397 18458 9463 18461
rect 10593 18458 10659 18461
rect 9397 18456 10659 18458
rect 9397 18400 9402 18456
rect 9458 18400 10598 18456
rect 10654 18400 10659 18456
rect 9397 18398 10659 18400
rect 9397 18395 9463 18398
rect 10593 18395 10659 18398
rect 8845 18322 8911 18325
rect 20897 18322 20963 18325
rect 8845 18320 20963 18322
rect 8845 18264 8850 18320
rect 8906 18264 20902 18320
rect 20958 18264 20963 18320
rect 8845 18262 20963 18264
rect 8845 18259 8911 18262
rect 20897 18259 20963 18262
rect 0 18186 800 18216
rect 2589 18186 2655 18189
rect 0 18184 2655 18186
rect 0 18128 2594 18184
rect 2650 18128 2655 18184
rect 0 18126 2655 18128
rect 0 18096 800 18126
rect 2589 18123 2655 18126
rect 7373 18186 7439 18189
rect 15377 18186 15443 18189
rect 7373 18184 15443 18186
rect 7373 18128 7378 18184
rect 7434 18128 15382 18184
rect 15438 18128 15443 18184
rect 7373 18126 15443 18128
rect 7373 18123 7439 18126
rect 15377 18123 15443 18126
rect 6637 18052 6703 18053
rect 6637 18048 6684 18052
rect 6748 18050 6754 18052
rect 7557 18050 7623 18053
rect 8150 18050 8156 18052
rect 6637 17992 6642 18048
rect 6637 17988 6684 17992
rect 6748 17990 6794 18050
rect 7557 18048 8156 18050
rect 7557 17992 7562 18048
rect 7618 17992 8156 18048
rect 7557 17990 8156 17992
rect 6748 17988 6754 17990
rect 6637 17987 6703 17988
rect 7557 17987 7623 17990
rect 8150 17988 8156 17990
rect 8220 17988 8226 18052
rect 9438 17988 9444 18052
rect 9508 18050 9514 18052
rect 9581 18050 9647 18053
rect 9508 18048 9647 18050
rect 9508 17992 9586 18048
rect 9642 17992 9647 18048
rect 9508 17990 9647 17992
rect 9508 17988 9514 17990
rect 9581 17987 9647 17990
rect 9765 18050 9831 18053
rect 12801 18050 12867 18053
rect 13077 18050 13143 18053
rect 9765 18048 13143 18050
rect 9765 17992 9770 18048
rect 9826 17992 12806 18048
rect 12862 17992 13082 18048
rect 13138 17992 13143 18048
rect 9765 17990 13143 17992
rect 9765 17987 9831 17990
rect 12801 17987 12867 17990
rect 13077 17987 13143 17990
rect 3545 17984 3861 17985
rect 3545 17920 3551 17984
rect 3615 17920 3631 17984
rect 3695 17920 3711 17984
rect 3775 17920 3791 17984
rect 3855 17920 3861 17984
rect 3545 17919 3861 17920
rect 8743 17984 9059 17985
rect 8743 17920 8749 17984
rect 8813 17920 8829 17984
rect 8893 17920 8909 17984
rect 8973 17920 8989 17984
rect 9053 17920 9059 17984
rect 8743 17919 9059 17920
rect 13941 17984 14257 17985
rect 13941 17920 13947 17984
rect 14011 17920 14027 17984
rect 14091 17920 14107 17984
rect 14171 17920 14187 17984
rect 14251 17920 14257 17984
rect 13941 17919 14257 17920
rect 19139 17984 19455 17985
rect 19139 17920 19145 17984
rect 19209 17920 19225 17984
rect 19289 17920 19305 17984
rect 19369 17920 19385 17984
rect 19449 17920 19455 17984
rect 19139 17919 19455 17920
rect 11605 17914 11671 17917
rect 12525 17914 12591 17917
rect 11605 17912 12591 17914
rect 11605 17856 11610 17912
rect 11666 17856 12530 17912
rect 12586 17856 12591 17912
rect 11605 17854 12591 17856
rect 11605 17851 11671 17854
rect 12525 17851 12591 17854
rect 0 17778 800 17808
rect 2313 17778 2379 17781
rect 0 17776 2379 17778
rect 0 17720 2318 17776
rect 2374 17720 2379 17776
rect 0 17718 2379 17720
rect 0 17688 800 17718
rect 2313 17715 2379 17718
rect 7741 17778 7807 17781
rect 19609 17778 19675 17781
rect 7741 17776 19675 17778
rect 7741 17720 7746 17776
rect 7802 17720 19614 17776
rect 19670 17720 19675 17776
rect 7741 17718 19675 17720
rect 7741 17715 7807 17718
rect 19609 17715 19675 17718
rect 6144 17440 6460 17441
rect 0 17370 800 17400
rect 6144 17376 6150 17440
rect 6214 17376 6230 17440
rect 6294 17376 6310 17440
rect 6374 17376 6390 17440
rect 6454 17376 6460 17440
rect 6144 17375 6460 17376
rect 11342 17440 11658 17441
rect 11342 17376 11348 17440
rect 11412 17376 11428 17440
rect 11492 17376 11508 17440
rect 11572 17376 11588 17440
rect 11652 17376 11658 17440
rect 11342 17375 11658 17376
rect 16540 17440 16856 17441
rect 16540 17376 16546 17440
rect 16610 17376 16626 17440
rect 16690 17376 16706 17440
rect 16770 17376 16786 17440
rect 16850 17376 16856 17440
rect 16540 17375 16856 17376
rect 21738 17440 22054 17441
rect 21738 17376 21744 17440
rect 21808 17376 21824 17440
rect 21888 17376 21904 17440
rect 21968 17376 21984 17440
rect 22048 17376 22054 17440
rect 21738 17375 22054 17376
rect 2681 17370 2747 17373
rect 0 17368 2747 17370
rect 0 17312 2686 17368
rect 2742 17312 2747 17368
rect 0 17310 2747 17312
rect 0 17280 800 17310
rect 2681 17307 2747 17310
rect 12893 17234 12959 17237
rect 16205 17234 16271 17237
rect 12893 17232 16271 17234
rect 12893 17176 12898 17232
rect 12954 17176 16210 17232
rect 16266 17176 16271 17232
rect 12893 17174 16271 17176
rect 12893 17171 12959 17174
rect 16205 17171 16271 17174
rect 19609 17234 19675 17237
rect 22200 17234 23000 17264
rect 19609 17232 23000 17234
rect 19609 17176 19614 17232
rect 19670 17176 23000 17232
rect 19609 17174 23000 17176
rect 19609 17171 19675 17174
rect 22200 17144 23000 17174
rect 6177 17098 6243 17101
rect 16113 17098 16179 17101
rect 6177 17096 16179 17098
rect 6177 17040 6182 17096
rect 6238 17040 16118 17096
rect 16174 17040 16179 17096
rect 6177 17038 16179 17040
rect 6177 17035 6243 17038
rect 16113 17035 16179 17038
rect 0 16962 800 16992
rect 1945 16962 2011 16965
rect 0 16960 2011 16962
rect 0 16904 1950 16960
rect 2006 16904 2011 16960
rect 0 16902 2011 16904
rect 0 16872 800 16902
rect 1945 16899 2011 16902
rect 12525 16962 12591 16965
rect 13353 16962 13419 16965
rect 12525 16960 13419 16962
rect 12525 16904 12530 16960
rect 12586 16904 13358 16960
rect 13414 16904 13419 16960
rect 12525 16902 13419 16904
rect 12525 16899 12591 16902
rect 13353 16899 13419 16902
rect 3545 16896 3861 16897
rect 3545 16832 3551 16896
rect 3615 16832 3631 16896
rect 3695 16832 3711 16896
rect 3775 16832 3791 16896
rect 3855 16832 3861 16896
rect 3545 16831 3861 16832
rect 8743 16896 9059 16897
rect 8743 16832 8749 16896
rect 8813 16832 8829 16896
rect 8893 16832 8909 16896
rect 8973 16832 8989 16896
rect 9053 16832 9059 16896
rect 8743 16831 9059 16832
rect 13941 16896 14257 16897
rect 13941 16832 13947 16896
rect 14011 16832 14027 16896
rect 14091 16832 14107 16896
rect 14171 16832 14187 16896
rect 14251 16832 14257 16896
rect 13941 16831 14257 16832
rect 19139 16896 19455 16897
rect 19139 16832 19145 16896
rect 19209 16832 19225 16896
rect 19289 16832 19305 16896
rect 19369 16832 19385 16896
rect 19449 16832 19455 16896
rect 19139 16831 19455 16832
rect 11513 16826 11579 16829
rect 11789 16826 11855 16829
rect 13353 16826 13419 16829
rect 11513 16824 13419 16826
rect 11513 16768 11518 16824
rect 11574 16768 11794 16824
rect 11850 16768 13358 16824
rect 13414 16768 13419 16824
rect 11513 16766 13419 16768
rect 11513 16763 11579 16766
rect 11789 16763 11855 16766
rect 13353 16763 13419 16766
rect 5993 16690 6059 16693
rect 6862 16690 6868 16692
rect 5993 16688 6868 16690
rect 5993 16632 5998 16688
rect 6054 16632 6868 16688
rect 5993 16630 6868 16632
rect 5993 16627 6059 16630
rect 6862 16628 6868 16630
rect 6932 16628 6938 16692
rect 0 16554 800 16584
rect 1853 16554 1919 16557
rect 0 16552 1919 16554
rect 0 16496 1858 16552
rect 1914 16496 1919 16552
rect 0 16494 1919 16496
rect 0 16464 800 16494
rect 1853 16491 1919 16494
rect 3601 16554 3667 16557
rect 9765 16554 9831 16557
rect 17861 16554 17927 16557
rect 3601 16552 9831 16554
rect 3601 16496 3606 16552
rect 3662 16496 9770 16552
rect 9826 16496 9831 16552
rect 3601 16494 9831 16496
rect 3601 16491 3667 16494
rect 9765 16491 9831 16494
rect 9952 16552 17927 16554
rect 9952 16496 17866 16552
rect 17922 16496 17927 16552
rect 9952 16494 17927 16496
rect 6913 16418 6979 16421
rect 9952 16418 10012 16494
rect 17861 16491 17927 16494
rect 6913 16416 10012 16418
rect 6913 16360 6918 16416
rect 6974 16360 10012 16416
rect 6913 16358 10012 16360
rect 6913 16355 6979 16358
rect 6144 16352 6460 16353
rect 6144 16288 6150 16352
rect 6214 16288 6230 16352
rect 6294 16288 6310 16352
rect 6374 16288 6390 16352
rect 6454 16288 6460 16352
rect 6144 16287 6460 16288
rect 11342 16352 11658 16353
rect 11342 16288 11348 16352
rect 11412 16288 11428 16352
rect 11492 16288 11508 16352
rect 11572 16288 11588 16352
rect 11652 16288 11658 16352
rect 11342 16287 11658 16288
rect 16540 16352 16856 16353
rect 16540 16288 16546 16352
rect 16610 16288 16626 16352
rect 16690 16288 16706 16352
rect 16770 16288 16786 16352
rect 16850 16288 16856 16352
rect 16540 16287 16856 16288
rect 21738 16352 22054 16353
rect 21738 16288 21744 16352
rect 21808 16288 21824 16352
rect 21888 16288 21904 16352
rect 21968 16288 21984 16352
rect 22048 16288 22054 16352
rect 21738 16287 22054 16288
rect 0 16146 800 16176
rect 2865 16146 2931 16149
rect 0 16144 2931 16146
rect 0 16088 2870 16144
rect 2926 16088 2931 16144
rect 0 16086 2931 16088
rect 0 16056 800 16086
rect 2865 16083 2931 16086
rect 7281 16146 7347 16149
rect 10225 16146 10291 16149
rect 10501 16146 10567 16149
rect 21081 16146 21147 16149
rect 7281 16144 10426 16146
rect 7281 16088 7286 16144
rect 7342 16088 10230 16144
rect 10286 16088 10426 16144
rect 7281 16086 10426 16088
rect 7281 16083 7347 16086
rect 10225 16083 10291 16086
rect 3877 16010 3943 16013
rect 10225 16010 10291 16013
rect 3877 16008 10291 16010
rect 3877 15952 3882 16008
rect 3938 15952 10230 16008
rect 10286 15952 10291 16008
rect 3877 15950 10291 15952
rect 10366 16010 10426 16086
rect 10501 16144 21147 16146
rect 10501 16088 10506 16144
rect 10562 16088 21086 16144
rect 21142 16088 21147 16144
rect 10501 16086 21147 16088
rect 10501 16083 10567 16086
rect 21081 16083 21147 16086
rect 12525 16010 12591 16013
rect 10366 16008 12591 16010
rect 10366 15952 12530 16008
rect 12586 15952 12591 16008
rect 10366 15950 12591 15952
rect 3877 15947 3943 15950
rect 10225 15947 10291 15950
rect 12525 15947 12591 15950
rect 7230 15812 7236 15876
rect 7300 15874 7306 15876
rect 8293 15874 8359 15877
rect 7300 15872 8359 15874
rect 7300 15816 8298 15872
rect 8354 15816 8359 15872
rect 7300 15814 8359 15816
rect 7300 15812 7306 15814
rect 8293 15811 8359 15814
rect 3545 15808 3861 15809
rect 0 15738 800 15768
rect 3545 15744 3551 15808
rect 3615 15744 3631 15808
rect 3695 15744 3711 15808
rect 3775 15744 3791 15808
rect 3855 15744 3861 15808
rect 3545 15743 3861 15744
rect 8743 15808 9059 15809
rect 8743 15744 8749 15808
rect 8813 15744 8829 15808
rect 8893 15744 8909 15808
rect 8973 15744 8989 15808
rect 9053 15744 9059 15808
rect 8743 15743 9059 15744
rect 13941 15808 14257 15809
rect 13941 15744 13947 15808
rect 14011 15744 14027 15808
rect 14091 15744 14107 15808
rect 14171 15744 14187 15808
rect 14251 15744 14257 15808
rect 13941 15743 14257 15744
rect 19139 15808 19455 15809
rect 19139 15744 19145 15808
rect 19209 15744 19225 15808
rect 19289 15744 19305 15808
rect 19369 15744 19385 15808
rect 19449 15744 19455 15808
rect 19139 15743 19455 15744
rect 3049 15738 3115 15741
rect 0 15736 3115 15738
rect 0 15680 3054 15736
rect 3110 15680 3115 15736
rect 0 15678 3115 15680
rect 0 15648 800 15678
rect 3049 15675 3115 15678
rect 7741 15602 7807 15605
rect 12433 15602 12499 15605
rect 7741 15600 12499 15602
rect 7741 15544 7746 15600
rect 7802 15544 12438 15600
rect 12494 15544 12499 15600
rect 7741 15542 12499 15544
rect 7741 15539 7807 15542
rect 12433 15539 12499 15542
rect 6913 15466 6979 15469
rect 11881 15466 11947 15469
rect 6913 15464 11947 15466
rect 6913 15408 6918 15464
rect 6974 15408 11886 15464
rect 11942 15408 11947 15464
rect 6913 15406 11947 15408
rect 6913 15403 6979 15406
rect 11881 15403 11947 15406
rect 0 15330 800 15360
rect 3141 15330 3207 15333
rect 9397 15332 9463 15333
rect 9397 15330 9444 15332
rect 0 15328 3207 15330
rect 0 15272 3146 15328
rect 3202 15272 3207 15328
rect 0 15270 3207 15272
rect 9352 15328 9444 15330
rect 9508 15330 9514 15332
rect 11053 15330 11119 15333
rect 9508 15328 11119 15330
rect 9352 15272 9402 15328
rect 9508 15272 11058 15328
rect 11114 15272 11119 15328
rect 9352 15270 9444 15272
rect 0 15240 800 15270
rect 3141 15267 3207 15270
rect 9397 15268 9444 15270
rect 9508 15270 11119 15272
rect 9508 15268 9514 15270
rect 9397 15267 9463 15268
rect 11053 15267 11119 15270
rect 6144 15264 6460 15265
rect 6144 15200 6150 15264
rect 6214 15200 6230 15264
rect 6294 15200 6310 15264
rect 6374 15200 6390 15264
rect 6454 15200 6460 15264
rect 6144 15199 6460 15200
rect 11342 15264 11658 15265
rect 11342 15200 11348 15264
rect 11412 15200 11428 15264
rect 11492 15200 11508 15264
rect 11572 15200 11588 15264
rect 11652 15200 11658 15264
rect 11342 15199 11658 15200
rect 16540 15264 16856 15265
rect 16540 15200 16546 15264
rect 16610 15200 16626 15264
rect 16690 15200 16706 15264
rect 16770 15200 16786 15264
rect 16850 15200 16856 15264
rect 16540 15199 16856 15200
rect 21738 15264 22054 15265
rect 21738 15200 21744 15264
rect 21808 15200 21824 15264
rect 21888 15200 21904 15264
rect 21968 15200 21984 15264
rect 22048 15200 22054 15264
rect 21738 15199 22054 15200
rect 5349 15058 5415 15061
rect 8017 15058 8083 15061
rect 5349 15056 8083 15058
rect 5349 15000 5354 15056
rect 5410 15000 8022 15056
rect 8078 15000 8083 15056
rect 5349 14998 8083 15000
rect 5349 14995 5415 14998
rect 8017 14995 8083 14998
rect 8201 15058 8267 15061
rect 14273 15058 14339 15061
rect 8201 15056 14339 15058
rect 8201 15000 8206 15056
rect 8262 15000 14278 15056
rect 14334 15000 14339 15056
rect 8201 14998 14339 15000
rect 8201 14995 8267 14998
rect 14273 14995 14339 14998
rect 0 14922 800 14952
rect 2957 14922 3023 14925
rect 0 14920 3023 14922
rect 0 14864 2962 14920
rect 3018 14864 3023 14920
rect 0 14862 3023 14864
rect 0 14832 800 14862
rect 2957 14859 3023 14862
rect 5257 14922 5323 14925
rect 5574 14922 5580 14924
rect 5257 14920 5580 14922
rect 5257 14864 5262 14920
rect 5318 14864 5580 14920
rect 5257 14862 5580 14864
rect 5257 14859 5323 14862
rect 5574 14860 5580 14862
rect 5644 14922 5650 14924
rect 15009 14922 15075 14925
rect 5644 14920 15075 14922
rect 5644 14864 15014 14920
rect 15070 14864 15075 14920
rect 5644 14862 15075 14864
rect 5644 14860 5650 14862
rect 15009 14859 15075 14862
rect 4613 14786 4679 14789
rect 6913 14786 6979 14789
rect 10225 14788 10291 14789
rect 4613 14784 6979 14786
rect 4613 14728 4618 14784
rect 4674 14728 6918 14784
rect 6974 14728 6979 14784
rect 4613 14726 6979 14728
rect 4613 14723 4679 14726
rect 6913 14723 6979 14726
rect 10174 14724 10180 14788
rect 10244 14786 10291 14788
rect 10244 14784 10336 14786
rect 10286 14728 10336 14784
rect 10244 14726 10336 14728
rect 10244 14724 10291 14726
rect 10225 14723 10291 14724
rect 3545 14720 3861 14721
rect 3545 14656 3551 14720
rect 3615 14656 3631 14720
rect 3695 14656 3711 14720
rect 3775 14656 3791 14720
rect 3855 14656 3861 14720
rect 3545 14655 3861 14656
rect 8743 14720 9059 14721
rect 8743 14656 8749 14720
rect 8813 14656 8829 14720
rect 8893 14656 8909 14720
rect 8973 14656 8989 14720
rect 9053 14656 9059 14720
rect 8743 14655 9059 14656
rect 13941 14720 14257 14721
rect 13941 14656 13947 14720
rect 14011 14656 14027 14720
rect 14091 14656 14107 14720
rect 14171 14656 14187 14720
rect 14251 14656 14257 14720
rect 13941 14655 14257 14656
rect 19139 14720 19455 14721
rect 19139 14656 19145 14720
rect 19209 14656 19225 14720
rect 19289 14656 19305 14720
rect 19369 14656 19385 14720
rect 19449 14656 19455 14720
rect 19139 14655 19455 14656
rect 0 14514 800 14544
rect 2773 14514 2839 14517
rect 0 14512 2839 14514
rect 0 14456 2778 14512
rect 2834 14456 2839 14512
rect 0 14454 2839 14456
rect 0 14424 800 14454
rect 2773 14451 2839 14454
rect 9121 14514 9187 14517
rect 18965 14514 19031 14517
rect 9121 14512 19031 14514
rect 9121 14456 9126 14512
rect 9182 14456 18970 14512
rect 19026 14456 19031 14512
rect 9121 14454 19031 14456
rect 9121 14451 9187 14454
rect 18965 14451 19031 14454
rect 7833 14244 7899 14245
rect 7782 14180 7788 14244
rect 7852 14242 7899 14244
rect 7852 14240 7944 14242
rect 7894 14184 7944 14240
rect 7852 14182 7944 14184
rect 7852 14180 7899 14182
rect 7833 14179 7899 14180
rect 6144 14176 6460 14177
rect 0 14106 800 14136
rect 6144 14112 6150 14176
rect 6214 14112 6230 14176
rect 6294 14112 6310 14176
rect 6374 14112 6390 14176
rect 6454 14112 6460 14176
rect 6144 14111 6460 14112
rect 11342 14176 11658 14177
rect 11342 14112 11348 14176
rect 11412 14112 11428 14176
rect 11492 14112 11508 14176
rect 11572 14112 11588 14176
rect 11652 14112 11658 14176
rect 11342 14111 11658 14112
rect 16540 14176 16856 14177
rect 16540 14112 16546 14176
rect 16610 14112 16626 14176
rect 16690 14112 16706 14176
rect 16770 14112 16786 14176
rect 16850 14112 16856 14176
rect 16540 14111 16856 14112
rect 21738 14176 22054 14177
rect 21738 14112 21744 14176
rect 21808 14112 21824 14176
rect 21888 14112 21904 14176
rect 21968 14112 21984 14176
rect 22048 14112 22054 14176
rect 21738 14111 22054 14112
rect 1853 14106 1919 14109
rect 0 14104 1919 14106
rect 0 14048 1858 14104
rect 1914 14048 1919 14104
rect 0 14046 1919 14048
rect 0 14016 800 14046
rect 1853 14043 1919 14046
rect 9765 14106 9831 14109
rect 10777 14106 10843 14109
rect 9765 14104 10843 14106
rect 9765 14048 9770 14104
rect 9826 14048 10782 14104
rect 10838 14048 10843 14104
rect 9765 14046 10843 14048
rect 9765 14043 9831 14046
rect 10777 14043 10843 14046
rect 6545 13970 6611 13973
rect 10501 13970 10567 13973
rect 6545 13968 10567 13970
rect 6545 13912 6550 13968
rect 6606 13912 10506 13968
rect 10562 13912 10567 13968
rect 6545 13910 10567 13912
rect 6545 13907 6611 13910
rect 10501 13907 10567 13910
rect 2221 13834 2287 13837
rect 2814 13834 2820 13836
rect 2221 13832 2820 13834
rect 2221 13776 2226 13832
rect 2282 13776 2820 13832
rect 2221 13774 2820 13776
rect 2221 13771 2287 13774
rect 2814 13772 2820 13774
rect 2884 13772 2890 13836
rect 0 13698 800 13728
rect 1577 13698 1643 13701
rect 0 13696 1643 13698
rect 0 13640 1582 13696
rect 1638 13640 1643 13696
rect 0 13638 1643 13640
rect 0 13608 800 13638
rect 1577 13635 1643 13638
rect 5758 13636 5764 13700
rect 5828 13698 5834 13700
rect 6085 13698 6151 13701
rect 5828 13696 6151 13698
rect 5828 13640 6090 13696
rect 6146 13640 6151 13696
rect 5828 13638 6151 13640
rect 5828 13636 5834 13638
rect 6085 13635 6151 13638
rect 3545 13632 3861 13633
rect 3545 13568 3551 13632
rect 3615 13568 3631 13632
rect 3695 13568 3711 13632
rect 3775 13568 3791 13632
rect 3855 13568 3861 13632
rect 3545 13567 3861 13568
rect 8743 13632 9059 13633
rect 8743 13568 8749 13632
rect 8813 13568 8829 13632
rect 8893 13568 8909 13632
rect 8973 13568 8989 13632
rect 9053 13568 9059 13632
rect 8743 13567 9059 13568
rect 13941 13632 14257 13633
rect 13941 13568 13947 13632
rect 14011 13568 14027 13632
rect 14091 13568 14107 13632
rect 14171 13568 14187 13632
rect 14251 13568 14257 13632
rect 13941 13567 14257 13568
rect 19139 13632 19455 13633
rect 19139 13568 19145 13632
rect 19209 13568 19225 13632
rect 19289 13568 19305 13632
rect 19369 13568 19385 13632
rect 19449 13568 19455 13632
rect 19139 13567 19455 13568
rect 8661 13426 8727 13429
rect 19517 13426 19583 13429
rect 20805 13426 20871 13429
rect 8661 13424 20871 13426
rect 8661 13368 8666 13424
rect 8722 13368 19522 13424
rect 19578 13368 20810 13424
rect 20866 13368 20871 13424
rect 8661 13366 20871 13368
rect 8661 13363 8727 13366
rect 19517 13363 19583 13366
rect 20805 13363 20871 13366
rect 0 13290 800 13320
rect 1945 13290 2011 13293
rect 0 13288 2011 13290
rect 0 13232 1950 13288
rect 2006 13232 2011 13288
rect 0 13230 2011 13232
rect 0 13200 800 13230
rect 1945 13227 2011 13230
rect 4061 13290 4127 13293
rect 11513 13290 11579 13293
rect 4061 13288 11579 13290
rect 4061 13232 4066 13288
rect 4122 13232 11518 13288
rect 11574 13232 11579 13288
rect 4061 13230 11579 13232
rect 4061 13227 4127 13230
rect 11513 13227 11579 13230
rect 6144 13088 6460 13089
rect 6144 13024 6150 13088
rect 6214 13024 6230 13088
rect 6294 13024 6310 13088
rect 6374 13024 6390 13088
rect 6454 13024 6460 13088
rect 6144 13023 6460 13024
rect 11342 13088 11658 13089
rect 11342 13024 11348 13088
rect 11412 13024 11428 13088
rect 11492 13024 11508 13088
rect 11572 13024 11588 13088
rect 11652 13024 11658 13088
rect 11342 13023 11658 13024
rect 16540 13088 16856 13089
rect 16540 13024 16546 13088
rect 16610 13024 16626 13088
rect 16690 13024 16706 13088
rect 16770 13024 16786 13088
rect 16850 13024 16856 13088
rect 16540 13023 16856 13024
rect 21738 13088 22054 13089
rect 21738 13024 21744 13088
rect 21808 13024 21824 13088
rect 21888 13024 21904 13088
rect 21968 13024 21984 13088
rect 22048 13024 22054 13088
rect 21738 13023 22054 13024
rect 11830 12956 11836 13020
rect 11900 13018 11906 13020
rect 11973 13018 12039 13021
rect 11900 13016 12039 13018
rect 11900 12960 11978 13016
rect 12034 12960 12039 13016
rect 11900 12958 12039 12960
rect 11900 12956 11906 12958
rect 11973 12955 12039 12958
rect 0 12882 800 12912
rect 3417 12882 3483 12885
rect 0 12880 3483 12882
rect 0 12824 3422 12880
rect 3478 12824 3483 12880
rect 0 12822 3483 12824
rect 0 12792 800 12822
rect 3417 12819 3483 12822
rect 5257 12882 5323 12885
rect 17953 12882 18019 12885
rect 5257 12880 18019 12882
rect 5257 12824 5262 12880
rect 5318 12824 17958 12880
rect 18014 12824 18019 12880
rect 5257 12822 18019 12824
rect 5257 12819 5323 12822
rect 17953 12819 18019 12822
rect 5942 12684 5948 12748
rect 6012 12746 6018 12748
rect 6821 12746 6887 12749
rect 6012 12744 6887 12746
rect 6012 12688 6826 12744
rect 6882 12688 6887 12744
rect 6012 12686 6887 12688
rect 6012 12684 6018 12686
rect 6821 12683 6887 12686
rect 7741 12746 7807 12749
rect 14549 12746 14615 12749
rect 16573 12746 16639 12749
rect 7741 12744 16639 12746
rect 7741 12688 7746 12744
rect 7802 12688 14554 12744
rect 14610 12688 16578 12744
rect 16634 12688 16639 12744
rect 7741 12686 16639 12688
rect 7741 12683 7807 12686
rect 14549 12683 14615 12686
rect 16573 12683 16639 12686
rect 12341 12610 12407 12613
rect 12206 12608 12407 12610
rect 12206 12552 12346 12608
rect 12402 12552 12407 12608
rect 12206 12550 12407 12552
rect 3545 12544 3861 12545
rect 0 12474 800 12504
rect 3545 12480 3551 12544
rect 3615 12480 3631 12544
rect 3695 12480 3711 12544
rect 3775 12480 3791 12544
rect 3855 12480 3861 12544
rect 3545 12479 3861 12480
rect 8743 12544 9059 12545
rect 8743 12480 8749 12544
rect 8813 12480 8829 12544
rect 8893 12480 8909 12544
rect 8973 12480 8989 12544
rect 9053 12480 9059 12544
rect 8743 12479 9059 12480
rect 3325 12474 3391 12477
rect 0 12472 3391 12474
rect 0 12416 3330 12472
rect 3386 12416 3391 12472
rect 0 12414 3391 12416
rect 0 12384 800 12414
rect 3325 12411 3391 12414
rect 9489 12474 9555 12477
rect 9622 12474 9628 12476
rect 9489 12472 9628 12474
rect 9489 12416 9494 12472
rect 9550 12416 9628 12472
rect 9489 12414 9628 12416
rect 9489 12411 9555 12414
rect 9622 12412 9628 12414
rect 9692 12412 9698 12476
rect 11789 12474 11855 12477
rect 12206 12474 12266 12550
rect 12341 12547 12407 12550
rect 13941 12544 14257 12545
rect 13941 12480 13947 12544
rect 14011 12480 14027 12544
rect 14091 12480 14107 12544
rect 14171 12480 14187 12544
rect 14251 12480 14257 12544
rect 13941 12479 14257 12480
rect 19139 12544 19455 12545
rect 19139 12480 19145 12544
rect 19209 12480 19225 12544
rect 19289 12480 19305 12544
rect 19369 12480 19385 12544
rect 19449 12480 19455 12544
rect 19139 12479 19455 12480
rect 11789 12472 12266 12474
rect 11789 12416 11794 12472
rect 11850 12416 12266 12472
rect 11789 12414 12266 12416
rect 11789 12411 11855 12414
rect 9949 12338 10015 12341
rect 18965 12338 19031 12341
rect 9949 12336 19031 12338
rect 9949 12280 9954 12336
rect 10010 12280 18970 12336
rect 19026 12280 19031 12336
rect 9949 12278 19031 12280
rect 9949 12275 10015 12278
rect 18965 12275 19031 12278
rect 9489 12202 9555 12205
rect 14733 12202 14799 12205
rect 9489 12200 14799 12202
rect 9489 12144 9494 12200
rect 9550 12144 14738 12200
rect 14794 12144 14799 12200
rect 9489 12142 14799 12144
rect 9489 12139 9555 12142
rect 14733 12139 14799 12142
rect 0 12066 800 12096
rect 1761 12066 1827 12069
rect 0 12064 1827 12066
rect 0 12008 1766 12064
rect 1822 12008 1827 12064
rect 0 12006 1827 12008
rect 0 11976 800 12006
rect 1761 12003 1827 12006
rect 9489 12066 9555 12069
rect 9622 12066 9628 12068
rect 9489 12064 9628 12066
rect 9489 12008 9494 12064
rect 9550 12008 9628 12064
rect 9489 12006 9628 12008
rect 9489 12003 9555 12006
rect 9622 12004 9628 12006
rect 9692 12004 9698 12068
rect 6144 12000 6460 12001
rect 6144 11936 6150 12000
rect 6214 11936 6230 12000
rect 6294 11936 6310 12000
rect 6374 11936 6390 12000
rect 6454 11936 6460 12000
rect 6144 11935 6460 11936
rect 11342 12000 11658 12001
rect 11342 11936 11348 12000
rect 11412 11936 11428 12000
rect 11492 11936 11508 12000
rect 11572 11936 11588 12000
rect 11652 11936 11658 12000
rect 11342 11935 11658 11936
rect 16540 12000 16856 12001
rect 16540 11936 16546 12000
rect 16610 11936 16626 12000
rect 16690 11936 16706 12000
rect 16770 11936 16786 12000
rect 16850 11936 16856 12000
rect 16540 11935 16856 11936
rect 21738 12000 22054 12001
rect 21738 11936 21744 12000
rect 21808 11936 21824 12000
rect 21888 11936 21904 12000
rect 21968 11936 21984 12000
rect 22048 11936 22054 12000
rect 21738 11935 22054 11936
rect 6913 11930 6979 11933
rect 8518 11930 8524 11932
rect 6913 11928 8524 11930
rect 6913 11872 6918 11928
rect 6974 11872 8524 11928
rect 6913 11870 8524 11872
rect 6913 11867 6979 11870
rect 8518 11868 8524 11870
rect 8588 11930 8594 11932
rect 10174 11930 10180 11932
rect 8588 11870 10180 11930
rect 8588 11868 8594 11870
rect 10174 11868 10180 11870
rect 10244 11868 10250 11932
rect 10777 11794 10843 11797
rect 19793 11794 19859 11797
rect 10777 11792 19859 11794
rect 10777 11736 10782 11792
rect 10838 11736 19798 11792
rect 19854 11736 19859 11792
rect 10777 11734 19859 11736
rect 10777 11731 10843 11734
rect 19793 11731 19859 11734
rect 0 11658 800 11688
rect 2865 11658 2931 11661
rect 0 11656 2931 11658
rect 0 11600 2870 11656
rect 2926 11600 2931 11656
rect 0 11598 2931 11600
rect 0 11568 800 11598
rect 2865 11595 2931 11598
rect 3233 11658 3299 11661
rect 5073 11658 5139 11661
rect 12065 11660 12131 11661
rect 12014 11658 12020 11660
rect 3233 11656 5139 11658
rect 3233 11600 3238 11656
rect 3294 11600 5078 11656
rect 5134 11600 5139 11656
rect 3233 11598 5139 11600
rect 11974 11598 12020 11658
rect 12084 11656 12131 11660
rect 12126 11600 12131 11656
rect 3233 11595 3299 11598
rect 5073 11595 5139 11598
rect 12014 11596 12020 11598
rect 12084 11596 12131 11600
rect 12065 11595 12131 11596
rect 3545 11456 3861 11457
rect 3545 11392 3551 11456
rect 3615 11392 3631 11456
rect 3695 11392 3711 11456
rect 3775 11392 3791 11456
rect 3855 11392 3861 11456
rect 3545 11391 3861 11392
rect 8743 11456 9059 11457
rect 8743 11392 8749 11456
rect 8813 11392 8829 11456
rect 8893 11392 8909 11456
rect 8973 11392 8989 11456
rect 9053 11392 9059 11456
rect 8743 11391 9059 11392
rect 13941 11456 14257 11457
rect 13941 11392 13947 11456
rect 14011 11392 14027 11456
rect 14091 11392 14107 11456
rect 14171 11392 14187 11456
rect 14251 11392 14257 11456
rect 13941 11391 14257 11392
rect 19139 11456 19455 11457
rect 19139 11392 19145 11456
rect 19209 11392 19225 11456
rect 19289 11392 19305 11456
rect 19369 11392 19385 11456
rect 19449 11392 19455 11456
rect 19139 11391 19455 11392
rect 11094 11324 11100 11388
rect 11164 11386 11170 11388
rect 11329 11386 11395 11389
rect 11164 11384 11395 11386
rect 11164 11328 11334 11384
rect 11390 11328 11395 11384
rect 11164 11326 11395 11328
rect 11164 11324 11170 11326
rect 11329 11323 11395 11326
rect 0 11250 800 11280
rect 4889 11250 4955 11253
rect 0 11248 4955 11250
rect 0 11192 4894 11248
rect 4950 11192 4955 11248
rect 0 11190 4955 11192
rect 0 11160 800 11190
rect 4889 11187 4955 11190
rect 5073 11250 5139 11253
rect 12249 11250 12315 11253
rect 5073 11248 12315 11250
rect 5073 11192 5078 11248
rect 5134 11192 12254 11248
rect 12310 11192 12315 11248
rect 5073 11190 12315 11192
rect 5073 11187 5139 11190
rect 12249 11187 12315 11190
rect 5625 11116 5691 11117
rect 5574 11052 5580 11116
rect 5644 11114 5691 11116
rect 7741 11114 7807 11117
rect 9806 11114 9812 11116
rect 5644 11112 5736 11114
rect 5686 11056 5736 11112
rect 5644 11054 5736 11056
rect 7741 11112 9812 11114
rect 7741 11056 7746 11112
rect 7802 11056 9812 11112
rect 7741 11054 9812 11056
rect 5644 11052 5691 11054
rect 5625 11051 5691 11052
rect 7741 11051 7807 11054
rect 9806 11052 9812 11054
rect 9876 11052 9882 11116
rect 6144 10912 6460 10913
rect 0 10842 800 10872
rect 6144 10848 6150 10912
rect 6214 10848 6230 10912
rect 6294 10848 6310 10912
rect 6374 10848 6390 10912
rect 6454 10848 6460 10912
rect 6144 10847 6460 10848
rect 11342 10912 11658 10913
rect 11342 10848 11348 10912
rect 11412 10848 11428 10912
rect 11492 10848 11508 10912
rect 11572 10848 11588 10912
rect 11652 10848 11658 10912
rect 11342 10847 11658 10848
rect 16540 10912 16856 10913
rect 16540 10848 16546 10912
rect 16610 10848 16626 10912
rect 16690 10848 16706 10912
rect 16770 10848 16786 10912
rect 16850 10848 16856 10912
rect 16540 10847 16856 10848
rect 21738 10912 22054 10913
rect 21738 10848 21744 10912
rect 21808 10848 21824 10912
rect 21888 10848 21904 10912
rect 21968 10848 21984 10912
rect 22048 10848 22054 10912
rect 21738 10847 22054 10848
rect 4061 10842 4127 10845
rect 0 10840 4127 10842
rect 0 10784 4066 10840
rect 4122 10784 4127 10840
rect 0 10782 4127 10784
rect 0 10752 800 10782
rect 4061 10779 4127 10782
rect 6913 10706 6979 10709
rect 10593 10706 10659 10709
rect 6913 10704 10659 10706
rect 6913 10648 6918 10704
rect 6974 10648 10598 10704
rect 10654 10648 10659 10704
rect 6913 10646 10659 10648
rect 6913 10643 6979 10646
rect 10593 10643 10659 10646
rect 11697 10706 11763 10709
rect 17125 10706 17191 10709
rect 11697 10704 17191 10706
rect 11697 10648 11702 10704
rect 11758 10648 17130 10704
rect 17186 10648 17191 10704
rect 11697 10646 17191 10648
rect 11697 10643 11763 10646
rect 17125 10643 17191 10646
rect 6637 10570 6703 10573
rect 11830 10570 11836 10572
rect 6637 10568 11836 10570
rect 6637 10512 6642 10568
rect 6698 10512 11836 10568
rect 6637 10510 11836 10512
rect 6637 10507 6703 10510
rect 11830 10508 11836 10510
rect 11900 10508 11906 10572
rect 0 10434 800 10464
rect 6085 10434 6151 10437
rect 7230 10434 7236 10436
rect 0 10374 2790 10434
rect 0 10344 800 10374
rect 2730 10162 2790 10374
rect 6085 10432 7236 10434
rect 6085 10376 6090 10432
rect 6146 10376 7236 10432
rect 6085 10374 7236 10376
rect 6085 10371 6151 10374
rect 7230 10372 7236 10374
rect 7300 10372 7306 10436
rect 3545 10368 3861 10369
rect 3545 10304 3551 10368
rect 3615 10304 3631 10368
rect 3695 10304 3711 10368
rect 3775 10304 3791 10368
rect 3855 10304 3861 10368
rect 3545 10303 3861 10304
rect 8743 10368 9059 10369
rect 8743 10304 8749 10368
rect 8813 10304 8829 10368
rect 8893 10304 8909 10368
rect 8973 10304 8989 10368
rect 9053 10304 9059 10368
rect 8743 10303 9059 10304
rect 13941 10368 14257 10369
rect 13941 10304 13947 10368
rect 14011 10304 14027 10368
rect 14091 10304 14107 10368
rect 14171 10304 14187 10368
rect 14251 10304 14257 10368
rect 13941 10303 14257 10304
rect 19139 10368 19455 10369
rect 19139 10304 19145 10368
rect 19209 10304 19225 10368
rect 19289 10304 19305 10368
rect 19369 10304 19385 10368
rect 19449 10304 19455 10368
rect 19139 10303 19455 10304
rect 12341 10298 12407 10301
rect 9262 10296 12407 10298
rect 9262 10240 12346 10296
rect 12402 10240 12407 10296
rect 9262 10238 12407 10240
rect 5165 10162 5231 10165
rect 6269 10162 6335 10165
rect 2730 10102 4170 10162
rect 0 10026 800 10056
rect 3969 10026 4035 10029
rect 0 10024 4035 10026
rect 0 9968 3974 10024
rect 4030 9968 4035 10024
rect 0 9966 4035 9968
rect 0 9936 800 9966
rect 3969 9963 4035 9966
rect 3877 9890 3943 9893
rect 4110 9890 4170 10102
rect 5165 10160 6335 10162
rect 5165 10104 5170 10160
rect 5226 10104 6274 10160
rect 6330 10104 6335 10160
rect 5165 10102 6335 10104
rect 5165 10099 5231 10102
rect 6269 10099 6335 10102
rect 6821 10162 6887 10165
rect 9262 10162 9322 10238
rect 12341 10235 12407 10238
rect 12801 10298 12867 10301
rect 13445 10298 13511 10301
rect 12801 10296 13511 10298
rect 12801 10240 12806 10296
rect 12862 10240 13450 10296
rect 13506 10240 13511 10296
rect 12801 10238 13511 10240
rect 12801 10235 12867 10238
rect 13445 10235 13511 10238
rect 6821 10160 9322 10162
rect 6821 10104 6826 10160
rect 6882 10104 9322 10160
rect 6821 10102 9322 10104
rect 6821 10099 6887 10102
rect 10910 10100 10916 10164
rect 10980 10162 10986 10164
rect 14549 10162 14615 10165
rect 10980 10160 14615 10162
rect 10980 10104 14554 10160
rect 14610 10104 14615 10160
rect 10980 10102 14615 10104
rect 10980 10100 10986 10102
rect 14549 10099 14615 10102
rect 5257 10026 5323 10029
rect 9857 10026 9923 10029
rect 5257 10024 9923 10026
rect 5257 9968 5262 10024
rect 5318 9968 9862 10024
rect 9918 9968 9923 10024
rect 5257 9966 9923 9968
rect 5257 9963 5323 9966
rect 9857 9963 9923 9966
rect 11094 9964 11100 10028
rect 11164 10026 11170 10028
rect 14733 10026 14799 10029
rect 11164 10024 14799 10026
rect 11164 9968 14738 10024
rect 14794 9968 14799 10024
rect 11164 9966 14799 9968
rect 11164 9964 11170 9966
rect 14733 9963 14799 9966
rect 3877 9888 4170 9890
rect 3877 9832 3882 9888
rect 3938 9832 4170 9888
rect 3877 9830 4170 9832
rect 3877 9827 3943 9830
rect 6144 9824 6460 9825
rect 6144 9760 6150 9824
rect 6214 9760 6230 9824
rect 6294 9760 6310 9824
rect 6374 9760 6390 9824
rect 6454 9760 6460 9824
rect 6144 9759 6460 9760
rect 11342 9824 11658 9825
rect 11342 9760 11348 9824
rect 11412 9760 11428 9824
rect 11492 9760 11508 9824
rect 11572 9760 11588 9824
rect 11652 9760 11658 9824
rect 11342 9759 11658 9760
rect 16540 9824 16856 9825
rect 16540 9760 16546 9824
rect 16610 9760 16626 9824
rect 16690 9760 16706 9824
rect 16770 9760 16786 9824
rect 16850 9760 16856 9824
rect 16540 9759 16856 9760
rect 21738 9824 22054 9825
rect 21738 9760 21744 9824
rect 21808 9760 21824 9824
rect 21888 9760 21904 9824
rect 21968 9760 21984 9824
rect 22048 9760 22054 9824
rect 21738 9759 22054 9760
rect 6545 9754 6611 9757
rect 7097 9754 7163 9757
rect 6545 9752 7163 9754
rect 6545 9696 6550 9752
rect 6606 9696 7102 9752
rect 7158 9696 7163 9752
rect 6545 9694 7163 9696
rect 6545 9691 6611 9694
rect 7097 9691 7163 9694
rect 13494 9694 14106 9754
rect 0 9618 800 9648
rect 3785 9618 3851 9621
rect 0 9616 3851 9618
rect 0 9560 3790 9616
rect 3846 9560 3851 9616
rect 0 9558 3851 9560
rect 0 9528 800 9558
rect 3785 9555 3851 9558
rect 5441 9618 5507 9621
rect 6821 9618 6887 9621
rect 10133 9620 10199 9621
rect 10133 9618 10180 9620
rect 5441 9616 6887 9618
rect 5441 9560 5446 9616
rect 5502 9560 6826 9616
rect 6882 9560 6887 9616
rect 5441 9558 6887 9560
rect 10088 9616 10180 9618
rect 10088 9560 10138 9616
rect 10088 9558 10180 9560
rect 5441 9555 5507 9558
rect 6821 9555 6887 9558
rect 10133 9556 10180 9558
rect 10244 9556 10250 9620
rect 10317 9618 10383 9621
rect 13494 9618 13554 9694
rect 13813 9618 13879 9621
rect 10317 9616 13554 9618
rect 10317 9560 10322 9616
rect 10378 9560 13554 9616
rect 10317 9558 13554 9560
rect 13678 9616 13879 9618
rect 13678 9560 13818 9616
rect 13874 9560 13879 9616
rect 13678 9558 13879 9560
rect 14046 9618 14106 9694
rect 16205 9618 16271 9621
rect 14046 9616 16271 9618
rect 14046 9560 16210 9616
rect 16266 9560 16271 9616
rect 14046 9558 16271 9560
rect 10133 9555 10199 9556
rect 10317 9555 10383 9558
rect 4889 9482 4955 9485
rect 5809 9482 5875 9485
rect 4889 9480 5875 9482
rect 4889 9424 4894 9480
rect 4950 9424 5814 9480
rect 5870 9424 5875 9480
rect 4889 9422 5875 9424
rect 4889 9419 4955 9422
rect 5809 9419 5875 9422
rect 7557 9482 7623 9485
rect 13678 9482 13738 9558
rect 13813 9555 13879 9558
rect 16205 9555 16271 9558
rect 7557 9480 13738 9482
rect 7557 9424 7562 9480
rect 7618 9424 13738 9480
rect 7557 9422 13738 9424
rect 13997 9482 14063 9485
rect 17217 9482 17283 9485
rect 13997 9480 17283 9482
rect 13997 9424 14002 9480
rect 14058 9424 17222 9480
rect 17278 9424 17283 9480
rect 13997 9422 17283 9424
rect 7557 9419 7623 9422
rect 13997 9419 14063 9422
rect 17217 9419 17283 9422
rect 5625 9346 5691 9349
rect 6269 9346 6335 9349
rect 13261 9346 13327 9349
rect 5625 9344 6335 9346
rect 5625 9288 5630 9344
rect 5686 9288 6274 9344
rect 6330 9288 6335 9344
rect 5625 9286 6335 9288
rect 5625 9283 5691 9286
rect 6269 9283 6335 9286
rect 12390 9344 13327 9346
rect 12390 9288 13266 9344
rect 13322 9288 13327 9344
rect 12390 9286 13327 9288
rect 3545 9280 3861 9281
rect 0 9210 800 9240
rect 3545 9216 3551 9280
rect 3615 9216 3631 9280
rect 3695 9216 3711 9280
rect 3775 9216 3791 9280
rect 3855 9216 3861 9280
rect 3545 9215 3861 9216
rect 8743 9280 9059 9281
rect 8743 9216 8749 9280
rect 8813 9216 8829 9280
rect 8893 9216 8909 9280
rect 8973 9216 8989 9280
rect 9053 9216 9059 9280
rect 8743 9215 9059 9216
rect 1669 9210 1735 9213
rect 0 9208 1735 9210
rect 0 9152 1674 9208
rect 1730 9152 1735 9208
rect 0 9150 1735 9152
rect 0 9120 800 9150
rect 1669 9147 1735 9150
rect 5073 9210 5139 9213
rect 7465 9210 7531 9213
rect 5073 9208 7531 9210
rect 5073 9152 5078 9208
rect 5134 9152 7470 9208
rect 7526 9152 7531 9208
rect 5073 9150 7531 9152
rect 5073 9147 5139 9150
rect 7465 9147 7531 9150
rect 10593 9210 10659 9213
rect 11513 9210 11579 9213
rect 10593 9208 11579 9210
rect 10593 9152 10598 9208
rect 10654 9152 11518 9208
rect 11574 9152 11579 9208
rect 10593 9150 11579 9152
rect 10593 9147 10659 9150
rect 11513 9147 11579 9150
rect 5257 9074 5323 9077
rect 6085 9074 6151 9077
rect 5257 9072 6151 9074
rect 5257 9016 5262 9072
rect 5318 9016 6090 9072
rect 6146 9016 6151 9072
rect 5257 9014 6151 9016
rect 5257 9011 5323 9014
rect 6085 9011 6151 9014
rect 6821 9074 6887 9077
rect 12390 9074 12450 9286
rect 13261 9283 13327 9286
rect 13941 9280 14257 9281
rect 13941 9216 13947 9280
rect 14011 9216 14027 9280
rect 14091 9216 14107 9280
rect 14171 9216 14187 9280
rect 14251 9216 14257 9280
rect 13941 9215 14257 9216
rect 19139 9280 19455 9281
rect 19139 9216 19145 9280
rect 19209 9216 19225 9280
rect 19289 9216 19305 9280
rect 19369 9216 19385 9280
rect 19449 9216 19455 9280
rect 19139 9215 19455 9216
rect 6821 9072 12450 9074
rect 6821 9016 6826 9072
rect 6882 9016 12450 9072
rect 6821 9014 12450 9016
rect 6821 9011 6887 9014
rect 4337 8938 4403 8941
rect 11329 8938 11395 8941
rect 4337 8936 11395 8938
rect 4337 8880 4342 8936
rect 4398 8880 11334 8936
rect 11390 8880 11395 8936
rect 4337 8878 11395 8880
rect 4337 8875 4403 8878
rect 11329 8875 11395 8878
rect 11513 8938 11579 8941
rect 13537 8938 13603 8941
rect 11513 8936 13603 8938
rect 11513 8880 11518 8936
rect 11574 8880 13542 8936
rect 13598 8880 13603 8936
rect 11513 8878 13603 8880
rect 11513 8875 11579 8878
rect 0 8802 800 8832
rect 1485 8802 1551 8805
rect 0 8800 1551 8802
rect 0 8744 1490 8800
rect 1546 8744 1551 8800
rect 0 8742 1551 8744
rect 0 8712 800 8742
rect 1485 8739 1551 8742
rect 5073 8802 5139 8805
rect 5809 8802 5875 8805
rect 5073 8800 5875 8802
rect 5073 8744 5078 8800
rect 5134 8744 5814 8800
rect 5870 8744 5875 8800
rect 5073 8742 5875 8744
rect 5073 8739 5139 8742
rect 5809 8739 5875 8742
rect 6144 8736 6460 8737
rect 6144 8672 6150 8736
rect 6214 8672 6230 8736
rect 6294 8672 6310 8736
rect 6374 8672 6390 8736
rect 6454 8672 6460 8736
rect 6144 8671 6460 8672
rect 11342 8736 11658 8737
rect 11342 8672 11348 8736
rect 11412 8672 11428 8736
rect 11492 8672 11508 8736
rect 11572 8672 11588 8736
rect 11652 8672 11658 8736
rect 11342 8671 11658 8672
rect 10133 8530 10199 8533
rect 11792 8530 11852 8878
rect 13537 8875 13603 8878
rect 16540 8736 16856 8737
rect 16540 8672 16546 8736
rect 16610 8672 16626 8736
rect 16690 8672 16706 8736
rect 16770 8672 16786 8736
rect 16850 8672 16856 8736
rect 16540 8671 16856 8672
rect 21738 8736 22054 8737
rect 21738 8672 21744 8736
rect 21808 8672 21824 8736
rect 21888 8672 21904 8736
rect 21968 8672 21984 8736
rect 22048 8672 22054 8736
rect 21738 8671 22054 8672
rect 10133 8528 11852 8530
rect 10133 8472 10138 8528
rect 10194 8472 11852 8528
rect 10133 8470 11852 8472
rect 13169 8530 13235 8533
rect 13537 8530 13603 8533
rect 15377 8530 15443 8533
rect 13169 8528 15443 8530
rect 13169 8472 13174 8528
rect 13230 8472 13542 8528
rect 13598 8472 15382 8528
rect 15438 8472 15443 8528
rect 13169 8470 15443 8472
rect 10133 8467 10199 8470
rect 13169 8467 13235 8470
rect 13537 8467 13603 8470
rect 15377 8467 15443 8470
rect 0 8394 800 8424
rect 5533 8394 5599 8397
rect 0 8392 5599 8394
rect 0 8336 5538 8392
rect 5594 8336 5599 8392
rect 0 8334 5599 8336
rect 0 8304 800 8334
rect 5533 8331 5599 8334
rect 9857 8394 9923 8397
rect 12525 8394 12591 8397
rect 9857 8392 12591 8394
rect 9857 8336 9862 8392
rect 9918 8336 12530 8392
rect 12586 8336 12591 8392
rect 9857 8334 12591 8336
rect 9857 8331 9923 8334
rect 12525 8331 12591 8334
rect 13678 8334 14474 8394
rect 11329 8258 11395 8261
rect 13678 8258 13738 8334
rect 11329 8256 13738 8258
rect 11329 8200 11334 8256
rect 11390 8200 13738 8256
rect 11329 8198 13738 8200
rect 14414 8258 14474 8334
rect 18137 8258 18203 8261
rect 18873 8258 18939 8261
rect 14414 8256 18939 8258
rect 14414 8200 18142 8256
rect 18198 8200 18878 8256
rect 18934 8200 18939 8256
rect 14414 8198 18939 8200
rect 11329 8195 11395 8198
rect 18137 8195 18203 8198
rect 18873 8195 18939 8198
rect 3545 8192 3861 8193
rect 3545 8128 3551 8192
rect 3615 8128 3631 8192
rect 3695 8128 3711 8192
rect 3775 8128 3791 8192
rect 3855 8128 3861 8192
rect 3545 8127 3861 8128
rect 8743 8192 9059 8193
rect 8743 8128 8749 8192
rect 8813 8128 8829 8192
rect 8893 8128 8909 8192
rect 8973 8128 8989 8192
rect 9053 8128 9059 8192
rect 8743 8127 9059 8128
rect 13941 8192 14257 8193
rect 13941 8128 13947 8192
rect 14011 8128 14027 8192
rect 14091 8128 14107 8192
rect 14171 8128 14187 8192
rect 14251 8128 14257 8192
rect 13941 8127 14257 8128
rect 19139 8192 19455 8193
rect 19139 8128 19145 8192
rect 19209 8128 19225 8192
rect 19289 8128 19305 8192
rect 19369 8128 19385 8192
rect 19449 8128 19455 8192
rect 19139 8127 19455 8128
rect 9121 8122 9187 8125
rect 13721 8122 13787 8125
rect 9121 8120 13787 8122
rect 9121 8064 9126 8120
rect 9182 8064 13726 8120
rect 13782 8064 13787 8120
rect 9121 8062 13787 8064
rect 9121 8059 9187 8062
rect 13721 8059 13787 8062
rect 0 7986 800 8016
rect 4245 7986 4311 7989
rect 0 7984 4311 7986
rect 0 7928 4250 7984
rect 4306 7928 4311 7984
rect 0 7926 4311 7928
rect 0 7896 800 7926
rect 4245 7923 4311 7926
rect 7189 7986 7255 7989
rect 10501 7986 10567 7989
rect 11329 7986 11395 7989
rect 7189 7984 10567 7986
rect 7189 7928 7194 7984
rect 7250 7928 10506 7984
rect 10562 7928 10567 7984
rect 7189 7926 10567 7928
rect 7189 7923 7255 7926
rect 10501 7923 10567 7926
rect 10734 7984 11395 7986
rect 10734 7928 11334 7984
rect 11390 7928 11395 7984
rect 10734 7926 11395 7928
rect 6361 7850 6427 7853
rect 10593 7850 10659 7853
rect 6361 7848 10659 7850
rect 6361 7792 6366 7848
rect 6422 7792 10598 7848
rect 10654 7792 10659 7848
rect 6361 7790 10659 7792
rect 6361 7787 6427 7790
rect 10593 7787 10659 7790
rect 8334 7652 8340 7716
rect 8404 7714 8410 7716
rect 10734 7714 10794 7926
rect 11329 7923 11395 7926
rect 12525 7986 12591 7989
rect 14273 7986 14339 7989
rect 12525 7984 14339 7986
rect 12525 7928 12530 7984
rect 12586 7928 14278 7984
rect 14334 7928 14339 7984
rect 12525 7926 14339 7928
rect 12525 7923 12591 7926
rect 14273 7923 14339 7926
rect 10869 7850 10935 7853
rect 17769 7850 17835 7853
rect 10869 7848 17835 7850
rect 10869 7792 10874 7848
rect 10930 7792 17774 7848
rect 17830 7792 17835 7848
rect 10869 7790 17835 7792
rect 10869 7787 10935 7790
rect 17769 7787 17835 7790
rect 8404 7654 10794 7714
rect 8404 7652 8410 7654
rect 6144 7648 6460 7649
rect 0 7578 800 7608
rect 6144 7584 6150 7648
rect 6214 7584 6230 7648
rect 6294 7584 6310 7648
rect 6374 7584 6390 7648
rect 6454 7584 6460 7648
rect 6144 7583 6460 7584
rect 11342 7648 11658 7649
rect 11342 7584 11348 7648
rect 11412 7584 11428 7648
rect 11492 7584 11508 7648
rect 11572 7584 11588 7648
rect 11652 7584 11658 7648
rect 11342 7583 11658 7584
rect 16540 7648 16856 7649
rect 16540 7584 16546 7648
rect 16610 7584 16626 7648
rect 16690 7584 16706 7648
rect 16770 7584 16786 7648
rect 16850 7584 16856 7648
rect 16540 7583 16856 7584
rect 21738 7648 22054 7649
rect 21738 7584 21744 7648
rect 21808 7584 21824 7648
rect 21888 7584 21904 7648
rect 21968 7584 21984 7648
rect 22048 7584 22054 7648
rect 21738 7583 22054 7584
rect 3969 7578 4035 7581
rect 0 7576 4035 7578
rect 0 7520 3974 7576
rect 4030 7520 4035 7576
rect 0 7518 4035 7520
rect 0 7488 800 7518
rect 3969 7515 4035 7518
rect 2865 7442 2931 7445
rect 6913 7442 6979 7445
rect 8569 7442 8635 7445
rect 2865 7440 8635 7442
rect 2865 7384 2870 7440
rect 2926 7384 6918 7440
rect 6974 7384 8574 7440
rect 8630 7384 8635 7440
rect 2865 7382 8635 7384
rect 2865 7379 2931 7382
rect 6913 7379 6979 7382
rect 8569 7379 8635 7382
rect 13629 7442 13695 7445
rect 17677 7442 17743 7445
rect 13629 7440 17743 7442
rect 13629 7384 13634 7440
rect 13690 7384 17682 7440
rect 17738 7384 17743 7440
rect 13629 7382 17743 7384
rect 13629 7379 13695 7382
rect 17677 7379 17743 7382
rect 6913 7308 6979 7309
rect 6862 7306 6868 7308
rect 6822 7246 6868 7306
rect 6932 7304 6979 7308
rect 6974 7248 6979 7304
rect 6862 7244 6868 7246
rect 6932 7244 6979 7248
rect 6913 7243 6979 7244
rect 9581 7306 9647 7309
rect 16941 7306 17007 7309
rect 9581 7304 17007 7306
rect 9581 7248 9586 7304
rect 9642 7248 16946 7304
rect 17002 7248 17007 7304
rect 9581 7246 17007 7248
rect 9581 7243 9647 7246
rect 16941 7243 17007 7246
rect 0 7170 800 7200
rect 3417 7170 3483 7173
rect 16389 7170 16455 7173
rect 17953 7170 18019 7173
rect 0 7168 3483 7170
rect 0 7112 3422 7168
rect 3478 7112 3483 7168
rect 0 7110 3483 7112
rect 0 7080 800 7110
rect 3417 7107 3483 7110
rect 15702 7168 18019 7170
rect 15702 7112 16394 7168
rect 16450 7112 17958 7168
rect 18014 7112 18019 7168
rect 15702 7110 18019 7112
rect 3545 7104 3861 7105
rect 3545 7040 3551 7104
rect 3615 7040 3631 7104
rect 3695 7040 3711 7104
rect 3775 7040 3791 7104
rect 3855 7040 3861 7104
rect 3545 7039 3861 7040
rect 8743 7104 9059 7105
rect 8743 7040 8749 7104
rect 8813 7040 8829 7104
rect 8893 7040 8909 7104
rect 8973 7040 8989 7104
rect 9053 7040 9059 7104
rect 8743 7039 9059 7040
rect 13941 7104 14257 7105
rect 13941 7040 13947 7104
rect 14011 7040 14027 7104
rect 14091 7040 14107 7104
rect 14171 7040 14187 7104
rect 14251 7040 14257 7104
rect 13941 7039 14257 7040
rect 12065 7034 12131 7037
rect 10918 7032 12131 7034
rect 10918 6976 12070 7032
rect 12126 6976 12131 7032
rect 10918 6974 12131 6976
rect 6361 6898 6427 6901
rect 6678 6898 6684 6900
rect 6361 6896 6684 6898
rect 6361 6840 6366 6896
rect 6422 6840 6684 6896
rect 6361 6838 6684 6840
rect 6361 6835 6427 6838
rect 6678 6836 6684 6838
rect 6748 6898 6754 6900
rect 7649 6898 7715 6901
rect 6748 6896 7715 6898
rect 6748 6840 7654 6896
rect 7710 6840 7715 6896
rect 6748 6838 7715 6840
rect 6748 6836 6754 6838
rect 7649 6835 7715 6838
rect 8293 6898 8359 6901
rect 10918 6898 10978 6974
rect 12065 6971 12131 6974
rect 8293 6896 10978 6898
rect 8293 6840 8298 6896
rect 8354 6840 10978 6896
rect 8293 6838 10978 6840
rect 11053 6898 11119 6901
rect 15702 6898 15762 7110
rect 16389 7107 16455 7110
rect 17953 7107 18019 7110
rect 19139 7104 19455 7105
rect 19139 7040 19145 7104
rect 19209 7040 19225 7104
rect 19289 7040 19305 7104
rect 19369 7040 19385 7104
rect 19449 7040 19455 7104
rect 19139 7039 19455 7040
rect 11053 6896 15762 6898
rect 11053 6840 11058 6896
rect 11114 6840 15762 6896
rect 11053 6838 15762 6840
rect 8293 6835 8359 6838
rect 11053 6835 11119 6838
rect 0 6762 800 6792
rect 3417 6762 3483 6765
rect 5809 6764 5875 6765
rect 0 6760 3483 6762
rect 0 6704 3422 6760
rect 3478 6704 3483 6760
rect 0 6702 3483 6704
rect 0 6672 800 6702
rect 3417 6699 3483 6702
rect 5758 6700 5764 6764
rect 5828 6762 5875 6764
rect 6821 6762 6887 6765
rect 5828 6760 6887 6762
rect 5870 6704 6826 6760
rect 6882 6704 6887 6760
rect 5828 6702 6887 6704
rect 5828 6700 5875 6702
rect 5809 6699 5875 6700
rect 6821 6699 6887 6702
rect 7189 6762 7255 6765
rect 8109 6762 8175 6765
rect 8569 6764 8635 6765
rect 7189 6760 8175 6762
rect 7189 6704 7194 6760
rect 7250 6704 8114 6760
rect 8170 6704 8175 6760
rect 7189 6702 8175 6704
rect 7189 6699 7255 6702
rect 8109 6699 8175 6702
rect 8518 6700 8524 6764
rect 8588 6762 8635 6764
rect 9581 6762 9647 6765
rect 12014 6762 12020 6764
rect 8588 6760 8680 6762
rect 8630 6704 8680 6760
rect 8588 6702 8680 6704
rect 9581 6760 12020 6762
rect 9581 6704 9586 6760
rect 9642 6704 12020 6760
rect 9581 6702 12020 6704
rect 8588 6700 8635 6702
rect 8569 6699 8635 6700
rect 9581 6699 9647 6702
rect 12014 6700 12020 6702
rect 12084 6700 12090 6764
rect 16941 6762 17007 6765
rect 12390 6760 17007 6762
rect 12390 6704 16946 6760
rect 17002 6704 17007 6760
rect 12390 6702 17007 6704
rect 1669 6626 1735 6629
rect 5717 6626 5783 6629
rect 8385 6626 8451 6629
rect 1669 6624 5783 6626
rect 1669 6568 1674 6624
rect 1730 6568 5722 6624
rect 5778 6568 5783 6624
rect 1669 6566 5783 6568
rect 1669 6563 1735 6566
rect 5717 6563 5783 6566
rect 6686 6624 8451 6626
rect 6686 6568 8390 6624
rect 8446 6568 8451 6624
rect 6686 6566 8451 6568
rect 6144 6560 6460 6561
rect 6144 6496 6150 6560
rect 6214 6496 6230 6560
rect 6294 6496 6310 6560
rect 6374 6496 6390 6560
rect 6454 6496 6460 6560
rect 6144 6495 6460 6496
rect 0 6354 800 6384
rect 3141 6354 3207 6357
rect 0 6352 3207 6354
rect 0 6296 3146 6352
rect 3202 6296 3207 6352
rect 0 6294 3207 6296
rect 0 6264 800 6294
rect 3141 6291 3207 6294
rect 3325 6354 3391 6357
rect 6686 6354 6746 6566
rect 8385 6563 8451 6566
rect 9029 6626 9095 6629
rect 10869 6626 10935 6629
rect 9029 6624 10935 6626
rect 9029 6568 9034 6624
rect 9090 6568 10874 6624
rect 10930 6568 10935 6624
rect 9029 6566 10935 6568
rect 9029 6563 9095 6566
rect 10869 6563 10935 6566
rect 11342 6560 11658 6561
rect 11342 6496 11348 6560
rect 11412 6496 11428 6560
rect 11492 6496 11508 6560
rect 11572 6496 11588 6560
rect 11652 6496 11658 6560
rect 11342 6495 11658 6496
rect 8518 6428 8524 6492
rect 8588 6490 8594 6492
rect 9397 6490 9463 6493
rect 8588 6488 9463 6490
rect 8588 6432 9402 6488
rect 9458 6432 9463 6488
rect 8588 6430 9463 6432
rect 8588 6428 8594 6430
rect 9397 6427 9463 6430
rect 3325 6352 6746 6354
rect 3325 6296 3330 6352
rect 3386 6296 6746 6352
rect 3325 6294 6746 6296
rect 3325 6291 3391 6294
rect 8150 6292 8156 6356
rect 8220 6354 8226 6356
rect 11513 6354 11579 6357
rect 8220 6352 11579 6354
rect 8220 6296 11518 6352
rect 11574 6296 11579 6352
rect 8220 6294 11579 6296
rect 8220 6292 8226 6294
rect 11513 6291 11579 6294
rect 7649 6218 7715 6221
rect 12390 6218 12450 6702
rect 16941 6699 17007 6702
rect 16540 6560 16856 6561
rect 16540 6496 16546 6560
rect 16610 6496 16626 6560
rect 16690 6496 16706 6560
rect 16770 6496 16786 6560
rect 16850 6496 16856 6560
rect 16540 6495 16856 6496
rect 21738 6560 22054 6561
rect 21738 6496 21744 6560
rect 21808 6496 21824 6560
rect 21888 6496 21904 6560
rect 21968 6496 21984 6560
rect 22048 6496 22054 6560
rect 21738 6495 22054 6496
rect 7649 6216 12450 6218
rect 7649 6160 7654 6216
rect 7710 6160 12450 6216
rect 7649 6158 12450 6160
rect 7649 6155 7715 6158
rect 6545 6082 6611 6085
rect 8477 6082 8543 6085
rect 6545 6080 8543 6082
rect 6545 6024 6550 6080
rect 6606 6024 8482 6080
rect 8538 6024 8543 6080
rect 6545 6022 8543 6024
rect 6545 6019 6611 6022
rect 8477 6019 8543 6022
rect 9438 6020 9444 6084
rect 9508 6082 9514 6084
rect 13629 6082 13695 6085
rect 9508 6080 13695 6082
rect 9508 6024 13634 6080
rect 13690 6024 13695 6080
rect 9508 6022 13695 6024
rect 9508 6020 9514 6022
rect 13629 6019 13695 6022
rect 3545 6016 3861 6017
rect 0 5946 800 5976
rect 3545 5952 3551 6016
rect 3615 5952 3631 6016
rect 3695 5952 3711 6016
rect 3775 5952 3791 6016
rect 3855 5952 3861 6016
rect 3545 5951 3861 5952
rect 8743 6016 9059 6017
rect 8743 5952 8749 6016
rect 8813 5952 8829 6016
rect 8893 5952 8909 6016
rect 8973 5952 8989 6016
rect 9053 5952 9059 6016
rect 8743 5951 9059 5952
rect 13941 6016 14257 6017
rect 13941 5952 13947 6016
rect 14011 5952 14027 6016
rect 14091 5952 14107 6016
rect 14171 5952 14187 6016
rect 14251 5952 14257 6016
rect 13941 5951 14257 5952
rect 19139 6016 19455 6017
rect 19139 5952 19145 6016
rect 19209 5952 19225 6016
rect 19289 5952 19305 6016
rect 19369 5952 19385 6016
rect 19449 5952 19455 6016
rect 19139 5951 19455 5952
rect 1393 5946 1459 5949
rect 0 5944 1459 5946
rect 0 5888 1398 5944
rect 1454 5888 1459 5944
rect 0 5886 1459 5888
rect 0 5856 800 5886
rect 1393 5883 1459 5886
rect 6729 5946 6795 5949
rect 7741 5948 7807 5949
rect 9213 5948 9279 5949
rect 7741 5946 7788 5948
rect 6729 5944 7788 5946
rect 6729 5888 6734 5944
rect 6790 5888 7746 5944
rect 6729 5886 7788 5888
rect 6729 5883 6795 5886
rect 7741 5884 7788 5886
rect 7852 5884 7858 5948
rect 9213 5946 9260 5948
rect 9168 5944 9260 5946
rect 9168 5888 9218 5944
rect 9168 5886 9260 5888
rect 9213 5884 9260 5886
rect 9324 5884 9330 5948
rect 10593 5946 10659 5949
rect 11329 5946 11395 5949
rect 10593 5944 11395 5946
rect 10593 5888 10598 5944
rect 10654 5888 11334 5944
rect 11390 5888 11395 5944
rect 10593 5886 11395 5888
rect 7741 5883 7807 5884
rect 9213 5883 9279 5884
rect 10593 5883 10659 5886
rect 11329 5883 11395 5886
rect 11513 5946 11579 5949
rect 12617 5946 12683 5949
rect 11513 5944 12683 5946
rect 11513 5888 11518 5944
rect 11574 5888 12622 5944
rect 12678 5888 12683 5944
rect 11513 5886 12683 5888
rect 11513 5883 11579 5886
rect 12617 5883 12683 5886
rect 5441 5810 5507 5813
rect 11697 5810 11763 5813
rect 5441 5808 11763 5810
rect 5441 5752 5446 5808
rect 5502 5752 11702 5808
rect 11758 5752 11763 5808
rect 5441 5750 11763 5752
rect 5441 5747 5507 5750
rect 11697 5747 11763 5750
rect 12065 5810 12131 5813
rect 15745 5810 15811 5813
rect 12065 5808 15811 5810
rect 12065 5752 12070 5808
rect 12126 5752 15750 5808
rect 15806 5752 15811 5808
rect 12065 5750 15811 5752
rect 12065 5747 12131 5750
rect 15745 5747 15811 5750
rect 21357 5810 21423 5813
rect 22200 5810 23000 5840
rect 21357 5808 23000 5810
rect 21357 5752 21362 5808
rect 21418 5752 23000 5808
rect 21357 5750 23000 5752
rect 21357 5747 21423 5750
rect 22200 5720 23000 5750
rect 9121 5674 9187 5677
rect 7744 5672 9187 5674
rect 7744 5616 9126 5672
rect 9182 5616 9187 5672
rect 7744 5614 9187 5616
rect 0 5538 800 5568
rect 5441 5538 5507 5541
rect 0 5536 5507 5538
rect 0 5480 5446 5536
rect 5502 5480 5507 5536
rect 0 5478 5507 5480
rect 0 5448 800 5478
rect 5441 5475 5507 5478
rect 6821 5538 6887 5541
rect 7744 5538 7804 5614
rect 9121 5611 9187 5614
rect 6821 5536 7804 5538
rect 6821 5480 6826 5536
rect 6882 5480 7804 5536
rect 6821 5478 7804 5480
rect 9397 5538 9463 5541
rect 12433 5538 12499 5541
rect 16389 5538 16455 5541
rect 9397 5536 9644 5538
rect 9397 5480 9402 5536
rect 9458 5480 9644 5536
rect 9397 5478 9644 5480
rect 6821 5475 6887 5478
rect 9397 5475 9463 5478
rect 6144 5472 6460 5473
rect 6144 5408 6150 5472
rect 6214 5408 6230 5472
rect 6294 5408 6310 5472
rect 6374 5408 6390 5472
rect 6454 5408 6460 5472
rect 6144 5407 6460 5408
rect 3969 5402 4035 5405
rect 5625 5402 5691 5405
rect 3969 5400 5691 5402
rect 3969 5344 3974 5400
rect 4030 5344 5630 5400
rect 5686 5344 5691 5400
rect 3969 5342 5691 5344
rect 9584 5402 9644 5478
rect 12433 5536 16455 5538
rect 12433 5480 12438 5536
rect 12494 5480 16394 5536
rect 16450 5480 16455 5536
rect 12433 5478 16455 5480
rect 12433 5475 12499 5478
rect 16389 5475 16455 5478
rect 11342 5472 11658 5473
rect 11342 5408 11348 5472
rect 11412 5408 11428 5472
rect 11492 5408 11508 5472
rect 11572 5408 11588 5472
rect 11652 5408 11658 5472
rect 11342 5407 11658 5408
rect 16540 5472 16856 5473
rect 16540 5408 16546 5472
rect 16610 5408 16626 5472
rect 16690 5408 16706 5472
rect 16770 5408 16786 5472
rect 16850 5408 16856 5472
rect 16540 5407 16856 5408
rect 21738 5472 22054 5473
rect 21738 5408 21744 5472
rect 21808 5408 21824 5472
rect 21888 5408 21904 5472
rect 21968 5408 21984 5472
rect 22048 5408 22054 5472
rect 21738 5407 22054 5408
rect 11053 5402 11119 5405
rect 9584 5400 11119 5402
rect 9584 5344 11058 5400
rect 11114 5344 11119 5400
rect 9584 5342 11119 5344
rect 3969 5339 4035 5342
rect 5625 5339 5691 5342
rect 11053 5339 11119 5342
rect 2037 5266 2103 5269
rect 5073 5266 5139 5269
rect 10777 5266 10843 5269
rect 2037 5264 4906 5266
rect 2037 5208 2042 5264
rect 2098 5208 4906 5264
rect 2037 5206 4906 5208
rect 2037 5203 2103 5206
rect 0 5130 800 5160
rect 3785 5130 3851 5133
rect 0 5128 3851 5130
rect 0 5072 3790 5128
rect 3846 5072 3851 5128
rect 0 5070 3851 5072
rect 4846 5130 4906 5206
rect 5073 5264 10843 5266
rect 5073 5208 5078 5264
rect 5134 5208 10782 5264
rect 10838 5208 10843 5264
rect 5073 5206 10843 5208
rect 5073 5203 5139 5206
rect 10777 5203 10843 5206
rect 11789 5266 11855 5269
rect 13537 5266 13603 5269
rect 11789 5264 13603 5266
rect 11789 5208 11794 5264
rect 11850 5208 13542 5264
rect 13598 5208 13603 5264
rect 11789 5206 13603 5208
rect 11789 5203 11855 5206
rect 13537 5203 13603 5206
rect 5165 5130 5231 5133
rect 9489 5130 9555 5133
rect 10317 5130 10383 5133
rect 4846 5128 8034 5130
rect 4846 5072 5170 5128
rect 5226 5072 8034 5128
rect 4846 5070 8034 5072
rect 0 5040 800 5070
rect 3785 5067 3851 5070
rect 5165 5067 5231 5070
rect 7974 4994 8034 5070
rect 9489 5128 10383 5130
rect 9489 5072 9494 5128
rect 9550 5072 10322 5128
rect 10378 5072 10383 5128
rect 9489 5070 10383 5072
rect 9489 5067 9555 5070
rect 10317 5067 10383 5070
rect 13077 5130 13143 5133
rect 17217 5130 17283 5133
rect 19609 5130 19675 5133
rect 13077 5128 19675 5130
rect 13077 5072 13082 5128
rect 13138 5072 17222 5128
rect 17278 5072 19614 5128
rect 19670 5072 19675 5128
rect 13077 5070 19675 5072
rect 13077 5067 13143 5070
rect 17217 5067 17283 5070
rect 19609 5067 19675 5070
rect 8569 4994 8635 4997
rect 9949 4994 10015 4997
rect 7974 4992 8635 4994
rect 7974 4936 8574 4992
rect 8630 4936 8635 4992
rect 7974 4934 8635 4936
rect 8569 4931 8635 4934
rect 9124 4992 10015 4994
rect 9124 4936 9954 4992
rect 10010 4936 10015 4992
rect 9124 4934 10015 4936
rect 3545 4928 3861 4929
rect 3545 4864 3551 4928
rect 3615 4864 3631 4928
rect 3695 4864 3711 4928
rect 3775 4864 3791 4928
rect 3855 4864 3861 4928
rect 3545 4863 3861 4864
rect 8743 4928 9059 4929
rect 8743 4864 8749 4928
rect 8813 4864 8829 4928
rect 8893 4864 8909 4928
rect 8973 4864 8989 4928
rect 9053 4864 9059 4928
rect 8743 4863 9059 4864
rect 9124 4861 9184 4934
rect 9949 4931 10015 4934
rect 10174 4932 10180 4996
rect 10244 4994 10250 4996
rect 10409 4994 10475 4997
rect 12525 4994 12591 4997
rect 10244 4992 10475 4994
rect 10244 4936 10414 4992
rect 10470 4936 10475 4992
rect 10244 4934 10475 4936
rect 10244 4932 10250 4934
rect 10409 4931 10475 4934
rect 12390 4992 12591 4994
rect 12390 4936 12530 4992
rect 12586 4936 12591 4992
rect 12390 4934 12591 4936
rect 9121 4856 9187 4861
rect 12390 4858 12450 4934
rect 12525 4931 12591 4934
rect 13941 4928 14257 4929
rect 13941 4864 13947 4928
rect 14011 4864 14027 4928
rect 14091 4864 14107 4928
rect 14171 4864 14187 4928
rect 14251 4864 14257 4928
rect 13941 4863 14257 4864
rect 19139 4928 19455 4929
rect 19139 4864 19145 4928
rect 19209 4864 19225 4928
rect 19289 4864 19305 4928
rect 19369 4864 19385 4928
rect 19449 4864 19455 4928
rect 19139 4863 19455 4864
rect 9121 4800 9126 4856
rect 9182 4800 9187 4856
rect 9121 4795 9187 4800
rect 9262 4798 12450 4858
rect 0 4722 800 4752
rect 3969 4722 4035 4725
rect 0 4720 4035 4722
rect 0 4664 3974 4720
rect 4030 4664 4035 4720
rect 0 4662 4035 4664
rect 0 4632 800 4662
rect 3969 4659 4035 4662
rect 4705 4722 4771 4725
rect 8753 4722 8819 4725
rect 9262 4722 9322 4798
rect 4705 4720 8034 4722
rect 4705 4664 4710 4720
rect 4766 4664 8034 4720
rect 4705 4662 8034 4664
rect 4705 4659 4771 4662
rect 7741 4586 7807 4589
rect 5812 4584 7807 4586
rect 5812 4528 7746 4584
rect 7802 4528 7807 4584
rect 5812 4526 7807 4528
rect 7974 4586 8034 4662
rect 8753 4720 9322 4722
rect 8753 4664 8758 4720
rect 8814 4664 9322 4720
rect 8753 4662 9322 4664
rect 8753 4659 8819 4662
rect 9806 4660 9812 4724
rect 9876 4722 9882 4724
rect 14641 4722 14707 4725
rect 9876 4720 14707 4722
rect 9876 4664 14646 4720
rect 14702 4664 14707 4720
rect 9876 4662 14707 4664
rect 9876 4660 9882 4662
rect 14641 4659 14707 4662
rect 8477 4586 8543 4589
rect 7974 4584 8543 4586
rect 7974 4528 8482 4584
rect 8538 4528 8543 4584
rect 7974 4526 8543 4528
rect 0 4314 800 4344
rect 4797 4314 4863 4317
rect 5812 4314 5872 4526
rect 7741 4523 7807 4526
rect 8477 4523 8543 4526
rect 7557 4450 7623 4453
rect 9397 4450 9463 4453
rect 7557 4448 9463 4450
rect 7557 4392 7562 4448
rect 7618 4392 9402 4448
rect 9458 4392 9463 4448
rect 7557 4390 9463 4392
rect 7557 4387 7623 4390
rect 9397 4387 9463 4390
rect 6144 4384 6460 4385
rect 6144 4320 6150 4384
rect 6214 4320 6230 4384
rect 6294 4320 6310 4384
rect 6374 4320 6390 4384
rect 6454 4320 6460 4384
rect 6144 4319 6460 4320
rect 11342 4384 11658 4385
rect 11342 4320 11348 4384
rect 11412 4320 11428 4384
rect 11492 4320 11508 4384
rect 11572 4320 11588 4384
rect 11652 4320 11658 4384
rect 11342 4319 11658 4320
rect 16540 4384 16856 4385
rect 16540 4320 16546 4384
rect 16610 4320 16626 4384
rect 16690 4320 16706 4384
rect 16770 4320 16786 4384
rect 16850 4320 16856 4384
rect 16540 4319 16856 4320
rect 21738 4384 22054 4385
rect 21738 4320 21744 4384
rect 21808 4320 21824 4384
rect 21888 4320 21904 4384
rect 21968 4320 21984 4384
rect 22048 4320 22054 4384
rect 21738 4319 22054 4320
rect 0 4312 5872 4314
rect 0 4256 4802 4312
rect 4858 4256 5872 4312
rect 0 4254 5872 4256
rect 0 4224 800 4254
rect 4797 4251 4863 4254
rect 9673 4178 9739 4181
rect 11053 4178 11119 4181
rect 12709 4178 12775 4181
rect 9673 4176 12775 4178
rect 9673 4120 9678 4176
rect 9734 4120 11058 4176
rect 11114 4120 12714 4176
rect 12770 4120 12775 4176
rect 9673 4118 12775 4120
rect 9673 4115 9739 4118
rect 11053 4115 11119 4118
rect 12709 4115 12775 4118
rect 2497 4042 2563 4045
rect 5717 4042 5783 4045
rect 2497 4040 5783 4042
rect 2497 3984 2502 4040
rect 2558 3984 5722 4040
rect 5778 3984 5783 4040
rect 2497 3982 5783 3984
rect 2497 3979 2563 3982
rect 5717 3979 5783 3982
rect 8109 4042 8175 4045
rect 15193 4042 15259 4045
rect 8109 4040 15259 4042
rect 8109 3984 8114 4040
rect 8170 3984 15198 4040
rect 15254 3984 15259 4040
rect 8109 3982 15259 3984
rect 8109 3979 8175 3982
rect 15193 3979 15259 3982
rect 0 3906 800 3936
rect 3325 3906 3391 3909
rect 0 3904 3391 3906
rect 0 3848 3330 3904
rect 3386 3848 3391 3904
rect 0 3846 3391 3848
rect 0 3816 800 3846
rect 3325 3843 3391 3846
rect 4981 3906 5047 3909
rect 7557 3906 7623 3909
rect 8569 3906 8635 3909
rect 4981 3904 8635 3906
rect 4981 3848 4986 3904
rect 5042 3848 7562 3904
rect 7618 3848 8574 3904
rect 8630 3848 8635 3904
rect 4981 3846 8635 3848
rect 4981 3843 5047 3846
rect 7557 3843 7623 3846
rect 8569 3843 8635 3846
rect 9438 3844 9444 3908
rect 9508 3906 9514 3908
rect 9581 3906 9647 3909
rect 9508 3904 9647 3906
rect 9508 3848 9586 3904
rect 9642 3848 9647 3904
rect 9508 3846 9647 3848
rect 9508 3844 9514 3846
rect 9581 3843 9647 3846
rect 3545 3840 3861 3841
rect 3545 3776 3551 3840
rect 3615 3776 3631 3840
rect 3695 3776 3711 3840
rect 3775 3776 3791 3840
rect 3855 3776 3861 3840
rect 3545 3775 3861 3776
rect 8743 3840 9059 3841
rect 8743 3776 8749 3840
rect 8813 3776 8829 3840
rect 8893 3776 8909 3840
rect 8973 3776 8989 3840
rect 9053 3776 9059 3840
rect 8743 3775 9059 3776
rect 13941 3840 14257 3841
rect 13941 3776 13947 3840
rect 14011 3776 14027 3840
rect 14091 3776 14107 3840
rect 14171 3776 14187 3840
rect 14251 3776 14257 3840
rect 13941 3775 14257 3776
rect 19139 3840 19455 3841
rect 19139 3776 19145 3840
rect 19209 3776 19225 3840
rect 19289 3776 19305 3840
rect 19369 3776 19385 3840
rect 19449 3776 19455 3840
rect 19139 3775 19455 3776
rect 6361 3634 6427 3637
rect 6729 3634 6795 3637
rect 6361 3632 6795 3634
rect 6361 3576 6366 3632
rect 6422 3576 6734 3632
rect 6790 3576 6795 3632
rect 6361 3574 6795 3576
rect 6361 3571 6427 3574
rect 6729 3571 6795 3574
rect 8201 3634 8267 3637
rect 9806 3634 9812 3636
rect 8201 3632 9812 3634
rect 8201 3576 8206 3632
rect 8262 3576 9812 3632
rect 8201 3574 9812 3576
rect 8201 3571 8267 3574
rect 9806 3572 9812 3574
rect 9876 3572 9882 3636
rect 9949 3634 10015 3637
rect 11237 3634 11303 3637
rect 9949 3632 11346 3634
rect 9949 3576 9954 3632
rect 10010 3576 11242 3632
rect 11298 3576 11346 3632
rect 9949 3574 11346 3576
rect 9949 3571 10015 3574
rect 11237 3571 11346 3574
rect 0 3498 800 3528
rect 3233 3498 3299 3501
rect 0 3496 3299 3498
rect 0 3440 3238 3496
rect 3294 3440 3299 3496
rect 0 3438 3299 3440
rect 0 3408 800 3438
rect 3233 3435 3299 3438
rect 5942 3436 5948 3500
rect 6012 3498 6018 3500
rect 11053 3498 11119 3501
rect 6012 3496 11119 3498
rect 6012 3440 11058 3496
rect 11114 3440 11119 3496
rect 6012 3438 11119 3440
rect 11286 3498 11346 3571
rect 15285 3498 15351 3501
rect 11286 3496 15351 3498
rect 11286 3440 15290 3496
rect 15346 3440 15351 3496
rect 11286 3438 15351 3440
rect 6012 3436 6018 3438
rect 11053 3435 11119 3438
rect 15285 3435 15351 3438
rect 8334 3300 8340 3364
rect 8404 3362 8410 3364
rect 9121 3362 9187 3365
rect 8404 3360 9187 3362
rect 8404 3304 9126 3360
rect 9182 3304 9187 3360
rect 8404 3302 9187 3304
rect 8404 3300 8410 3302
rect 9121 3299 9187 3302
rect 6144 3296 6460 3297
rect 6144 3232 6150 3296
rect 6214 3232 6230 3296
rect 6294 3232 6310 3296
rect 6374 3232 6390 3296
rect 6454 3232 6460 3296
rect 6144 3231 6460 3232
rect 11342 3296 11658 3297
rect 11342 3232 11348 3296
rect 11412 3232 11428 3296
rect 11492 3232 11508 3296
rect 11572 3232 11588 3296
rect 11652 3232 11658 3296
rect 11342 3231 11658 3232
rect 16540 3296 16856 3297
rect 16540 3232 16546 3296
rect 16610 3232 16626 3296
rect 16690 3232 16706 3296
rect 16770 3232 16786 3296
rect 16850 3232 16856 3296
rect 16540 3231 16856 3232
rect 21738 3296 22054 3297
rect 21738 3232 21744 3296
rect 21808 3232 21824 3296
rect 21888 3232 21904 3296
rect 21968 3232 21984 3296
rect 22048 3232 22054 3296
rect 21738 3231 22054 3232
rect 5758 3164 5764 3228
rect 5828 3226 5834 3228
rect 5901 3226 5967 3229
rect 5828 3224 5967 3226
rect 5828 3168 5906 3224
rect 5962 3168 5967 3224
rect 5828 3166 5967 3168
rect 5828 3164 5834 3166
rect 5901 3163 5967 3166
rect 6913 3226 6979 3229
rect 11053 3226 11119 3229
rect 6913 3224 11119 3226
rect 6913 3168 6918 3224
rect 6974 3168 11058 3224
rect 11114 3168 11119 3224
rect 6913 3166 11119 3168
rect 6913 3163 6979 3166
rect 11053 3163 11119 3166
rect 0 3090 800 3120
rect 2865 3090 2931 3093
rect 0 3088 2931 3090
rect 0 3032 2870 3088
rect 2926 3032 2931 3088
rect 0 3030 2931 3032
rect 0 3000 800 3030
rect 2865 3027 2931 3030
rect 6545 3090 6611 3093
rect 10593 3090 10659 3093
rect 6545 3088 10659 3090
rect 6545 3032 6550 3088
rect 6606 3032 10598 3088
rect 10654 3032 10659 3088
rect 6545 3030 10659 3032
rect 6545 3027 6611 3030
rect 10593 3027 10659 3030
rect 9673 2954 9739 2957
rect 17677 2954 17743 2957
rect 9673 2952 17743 2954
rect 9673 2896 9678 2952
rect 9734 2896 17682 2952
rect 17738 2896 17743 2952
rect 9673 2894 17743 2896
rect 9673 2891 9739 2894
rect 17677 2891 17743 2894
rect 3545 2752 3861 2753
rect 0 2682 800 2712
rect 3545 2688 3551 2752
rect 3615 2688 3631 2752
rect 3695 2688 3711 2752
rect 3775 2688 3791 2752
rect 3855 2688 3861 2752
rect 3545 2687 3861 2688
rect 8743 2752 9059 2753
rect 8743 2688 8749 2752
rect 8813 2688 8829 2752
rect 8893 2688 8909 2752
rect 8973 2688 8989 2752
rect 9053 2688 9059 2752
rect 8743 2687 9059 2688
rect 13941 2752 14257 2753
rect 13941 2688 13947 2752
rect 14011 2688 14027 2752
rect 14091 2688 14107 2752
rect 14171 2688 14187 2752
rect 14251 2688 14257 2752
rect 13941 2687 14257 2688
rect 19139 2752 19455 2753
rect 19139 2688 19145 2752
rect 19209 2688 19225 2752
rect 19289 2688 19305 2752
rect 19369 2688 19385 2752
rect 19449 2688 19455 2752
rect 19139 2687 19455 2688
rect 3417 2682 3483 2685
rect 0 2680 3483 2682
rect 0 2624 3422 2680
rect 3478 2624 3483 2680
rect 0 2622 3483 2624
rect 0 2592 800 2622
rect 3417 2619 3483 2622
rect 8518 2484 8524 2548
rect 8588 2546 8594 2548
rect 9121 2546 9187 2549
rect 8588 2544 9187 2546
rect 8588 2488 9126 2544
rect 9182 2488 9187 2544
rect 8588 2486 9187 2488
rect 8588 2484 8594 2486
rect 9121 2483 9187 2486
rect 0 2274 800 2304
rect 1669 2274 1735 2277
rect 0 2272 1735 2274
rect 0 2216 1674 2272
rect 1730 2216 1735 2272
rect 0 2214 1735 2216
rect 0 2184 800 2214
rect 1669 2211 1735 2214
rect 6144 2208 6460 2209
rect 6144 2144 6150 2208
rect 6214 2144 6230 2208
rect 6294 2144 6310 2208
rect 6374 2144 6390 2208
rect 6454 2144 6460 2208
rect 6144 2143 6460 2144
rect 11342 2208 11658 2209
rect 11342 2144 11348 2208
rect 11412 2144 11428 2208
rect 11492 2144 11508 2208
rect 11572 2144 11588 2208
rect 11652 2144 11658 2208
rect 11342 2143 11658 2144
rect 16540 2208 16856 2209
rect 16540 2144 16546 2208
rect 16610 2144 16626 2208
rect 16690 2144 16706 2208
rect 16770 2144 16786 2208
rect 16850 2144 16856 2208
rect 16540 2143 16856 2144
rect 21738 2208 22054 2209
rect 21738 2144 21744 2208
rect 21808 2144 21824 2208
rect 21888 2144 21904 2208
rect 21968 2144 21984 2208
rect 22048 2144 22054 2208
rect 21738 2143 22054 2144
rect 0 1866 800 1896
rect 3417 1866 3483 1869
rect 0 1864 3483 1866
rect 0 1808 3422 1864
rect 3478 1808 3483 1864
rect 0 1806 3483 1808
rect 0 1776 800 1806
rect 3417 1803 3483 1806
<< via3 >>
rect 6150 20700 6214 20704
rect 6150 20644 6154 20700
rect 6154 20644 6210 20700
rect 6210 20644 6214 20700
rect 6150 20640 6214 20644
rect 6230 20700 6294 20704
rect 6230 20644 6234 20700
rect 6234 20644 6290 20700
rect 6290 20644 6294 20700
rect 6230 20640 6294 20644
rect 6310 20700 6374 20704
rect 6310 20644 6314 20700
rect 6314 20644 6370 20700
rect 6370 20644 6374 20700
rect 6310 20640 6374 20644
rect 6390 20700 6454 20704
rect 6390 20644 6394 20700
rect 6394 20644 6450 20700
rect 6450 20644 6454 20700
rect 6390 20640 6454 20644
rect 11348 20700 11412 20704
rect 11348 20644 11352 20700
rect 11352 20644 11408 20700
rect 11408 20644 11412 20700
rect 11348 20640 11412 20644
rect 11428 20700 11492 20704
rect 11428 20644 11432 20700
rect 11432 20644 11488 20700
rect 11488 20644 11492 20700
rect 11428 20640 11492 20644
rect 11508 20700 11572 20704
rect 11508 20644 11512 20700
rect 11512 20644 11568 20700
rect 11568 20644 11572 20700
rect 11508 20640 11572 20644
rect 11588 20700 11652 20704
rect 11588 20644 11592 20700
rect 11592 20644 11648 20700
rect 11648 20644 11652 20700
rect 11588 20640 11652 20644
rect 16546 20700 16610 20704
rect 16546 20644 16550 20700
rect 16550 20644 16606 20700
rect 16606 20644 16610 20700
rect 16546 20640 16610 20644
rect 16626 20700 16690 20704
rect 16626 20644 16630 20700
rect 16630 20644 16686 20700
rect 16686 20644 16690 20700
rect 16626 20640 16690 20644
rect 16706 20700 16770 20704
rect 16706 20644 16710 20700
rect 16710 20644 16766 20700
rect 16766 20644 16770 20700
rect 16706 20640 16770 20644
rect 16786 20700 16850 20704
rect 16786 20644 16790 20700
rect 16790 20644 16846 20700
rect 16846 20644 16850 20700
rect 16786 20640 16850 20644
rect 21744 20700 21808 20704
rect 21744 20644 21748 20700
rect 21748 20644 21804 20700
rect 21804 20644 21808 20700
rect 21744 20640 21808 20644
rect 21824 20700 21888 20704
rect 21824 20644 21828 20700
rect 21828 20644 21884 20700
rect 21884 20644 21888 20700
rect 21824 20640 21888 20644
rect 21904 20700 21968 20704
rect 21904 20644 21908 20700
rect 21908 20644 21964 20700
rect 21964 20644 21968 20700
rect 21904 20640 21968 20644
rect 21984 20700 22048 20704
rect 21984 20644 21988 20700
rect 21988 20644 22044 20700
rect 22044 20644 22048 20700
rect 21984 20640 22048 20644
rect 3551 20156 3615 20160
rect 3551 20100 3555 20156
rect 3555 20100 3611 20156
rect 3611 20100 3615 20156
rect 3551 20096 3615 20100
rect 3631 20156 3695 20160
rect 3631 20100 3635 20156
rect 3635 20100 3691 20156
rect 3691 20100 3695 20156
rect 3631 20096 3695 20100
rect 3711 20156 3775 20160
rect 3711 20100 3715 20156
rect 3715 20100 3771 20156
rect 3771 20100 3775 20156
rect 3711 20096 3775 20100
rect 3791 20156 3855 20160
rect 3791 20100 3795 20156
rect 3795 20100 3851 20156
rect 3851 20100 3855 20156
rect 3791 20096 3855 20100
rect 8749 20156 8813 20160
rect 8749 20100 8753 20156
rect 8753 20100 8809 20156
rect 8809 20100 8813 20156
rect 8749 20096 8813 20100
rect 8829 20156 8893 20160
rect 8829 20100 8833 20156
rect 8833 20100 8889 20156
rect 8889 20100 8893 20156
rect 8829 20096 8893 20100
rect 8909 20156 8973 20160
rect 8909 20100 8913 20156
rect 8913 20100 8969 20156
rect 8969 20100 8973 20156
rect 8909 20096 8973 20100
rect 8989 20156 9053 20160
rect 8989 20100 8993 20156
rect 8993 20100 9049 20156
rect 9049 20100 9053 20156
rect 8989 20096 9053 20100
rect 13947 20156 14011 20160
rect 13947 20100 13951 20156
rect 13951 20100 14007 20156
rect 14007 20100 14011 20156
rect 13947 20096 14011 20100
rect 14027 20156 14091 20160
rect 14027 20100 14031 20156
rect 14031 20100 14087 20156
rect 14087 20100 14091 20156
rect 14027 20096 14091 20100
rect 14107 20156 14171 20160
rect 14107 20100 14111 20156
rect 14111 20100 14167 20156
rect 14167 20100 14171 20156
rect 14107 20096 14171 20100
rect 14187 20156 14251 20160
rect 14187 20100 14191 20156
rect 14191 20100 14247 20156
rect 14247 20100 14251 20156
rect 14187 20096 14251 20100
rect 19145 20156 19209 20160
rect 19145 20100 19149 20156
rect 19149 20100 19205 20156
rect 19205 20100 19209 20156
rect 19145 20096 19209 20100
rect 19225 20156 19289 20160
rect 19225 20100 19229 20156
rect 19229 20100 19285 20156
rect 19285 20100 19289 20156
rect 19225 20096 19289 20100
rect 19305 20156 19369 20160
rect 19305 20100 19309 20156
rect 19309 20100 19365 20156
rect 19365 20100 19369 20156
rect 19305 20096 19369 20100
rect 19385 20156 19449 20160
rect 19385 20100 19389 20156
rect 19389 20100 19445 20156
rect 19445 20100 19449 20156
rect 19385 20096 19449 20100
rect 11100 19620 11164 19684
rect 6150 19612 6214 19616
rect 6150 19556 6154 19612
rect 6154 19556 6210 19612
rect 6210 19556 6214 19612
rect 6150 19552 6214 19556
rect 6230 19612 6294 19616
rect 6230 19556 6234 19612
rect 6234 19556 6290 19612
rect 6290 19556 6294 19612
rect 6230 19552 6294 19556
rect 6310 19612 6374 19616
rect 6310 19556 6314 19612
rect 6314 19556 6370 19612
rect 6370 19556 6374 19612
rect 6310 19552 6374 19556
rect 6390 19612 6454 19616
rect 6390 19556 6394 19612
rect 6394 19556 6450 19612
rect 6450 19556 6454 19612
rect 6390 19552 6454 19556
rect 11348 19612 11412 19616
rect 11348 19556 11352 19612
rect 11352 19556 11408 19612
rect 11408 19556 11412 19612
rect 11348 19552 11412 19556
rect 11428 19612 11492 19616
rect 11428 19556 11432 19612
rect 11432 19556 11488 19612
rect 11488 19556 11492 19612
rect 11428 19552 11492 19556
rect 11508 19612 11572 19616
rect 11508 19556 11512 19612
rect 11512 19556 11568 19612
rect 11568 19556 11572 19612
rect 11508 19552 11572 19556
rect 11588 19612 11652 19616
rect 11588 19556 11592 19612
rect 11592 19556 11648 19612
rect 11648 19556 11652 19612
rect 11588 19552 11652 19556
rect 16546 19612 16610 19616
rect 16546 19556 16550 19612
rect 16550 19556 16606 19612
rect 16606 19556 16610 19612
rect 16546 19552 16610 19556
rect 16626 19612 16690 19616
rect 16626 19556 16630 19612
rect 16630 19556 16686 19612
rect 16686 19556 16690 19612
rect 16626 19552 16690 19556
rect 16706 19612 16770 19616
rect 16706 19556 16710 19612
rect 16710 19556 16766 19612
rect 16766 19556 16770 19612
rect 16706 19552 16770 19556
rect 16786 19612 16850 19616
rect 16786 19556 16790 19612
rect 16790 19556 16846 19612
rect 16846 19556 16850 19612
rect 16786 19552 16850 19556
rect 21744 19612 21808 19616
rect 21744 19556 21748 19612
rect 21748 19556 21804 19612
rect 21804 19556 21808 19612
rect 21744 19552 21808 19556
rect 21824 19612 21888 19616
rect 21824 19556 21828 19612
rect 21828 19556 21884 19612
rect 21884 19556 21888 19612
rect 21824 19552 21888 19556
rect 21904 19612 21968 19616
rect 21904 19556 21908 19612
rect 21908 19556 21964 19612
rect 21964 19556 21968 19612
rect 21904 19552 21968 19556
rect 21984 19612 22048 19616
rect 21984 19556 21988 19612
rect 21988 19556 22044 19612
rect 22044 19556 22048 19612
rect 21984 19552 22048 19556
rect 9444 19076 9508 19140
rect 9812 19076 9876 19140
rect 3551 19068 3615 19072
rect 3551 19012 3555 19068
rect 3555 19012 3611 19068
rect 3611 19012 3615 19068
rect 3551 19008 3615 19012
rect 3631 19068 3695 19072
rect 3631 19012 3635 19068
rect 3635 19012 3691 19068
rect 3691 19012 3695 19068
rect 3631 19008 3695 19012
rect 3711 19068 3775 19072
rect 3711 19012 3715 19068
rect 3715 19012 3771 19068
rect 3771 19012 3775 19068
rect 3711 19008 3775 19012
rect 3791 19068 3855 19072
rect 3791 19012 3795 19068
rect 3795 19012 3851 19068
rect 3851 19012 3855 19068
rect 3791 19008 3855 19012
rect 8749 19068 8813 19072
rect 8749 19012 8753 19068
rect 8753 19012 8809 19068
rect 8809 19012 8813 19068
rect 8749 19008 8813 19012
rect 8829 19068 8893 19072
rect 8829 19012 8833 19068
rect 8833 19012 8889 19068
rect 8889 19012 8893 19068
rect 8829 19008 8893 19012
rect 8909 19068 8973 19072
rect 8909 19012 8913 19068
rect 8913 19012 8969 19068
rect 8969 19012 8973 19068
rect 8909 19008 8973 19012
rect 8989 19068 9053 19072
rect 8989 19012 8993 19068
rect 8993 19012 9049 19068
rect 9049 19012 9053 19068
rect 8989 19008 9053 19012
rect 13947 19068 14011 19072
rect 13947 19012 13951 19068
rect 13951 19012 14007 19068
rect 14007 19012 14011 19068
rect 13947 19008 14011 19012
rect 14027 19068 14091 19072
rect 14027 19012 14031 19068
rect 14031 19012 14087 19068
rect 14087 19012 14091 19068
rect 14027 19008 14091 19012
rect 14107 19068 14171 19072
rect 14107 19012 14111 19068
rect 14111 19012 14167 19068
rect 14167 19012 14171 19068
rect 14107 19008 14171 19012
rect 14187 19068 14251 19072
rect 14187 19012 14191 19068
rect 14191 19012 14247 19068
rect 14247 19012 14251 19068
rect 14187 19008 14251 19012
rect 19145 19068 19209 19072
rect 19145 19012 19149 19068
rect 19149 19012 19205 19068
rect 19205 19012 19209 19068
rect 19145 19008 19209 19012
rect 19225 19068 19289 19072
rect 19225 19012 19229 19068
rect 19229 19012 19285 19068
rect 19285 19012 19289 19068
rect 19225 19008 19289 19012
rect 19305 19068 19369 19072
rect 19305 19012 19309 19068
rect 19309 19012 19365 19068
rect 19365 19012 19369 19068
rect 19305 19008 19369 19012
rect 19385 19068 19449 19072
rect 19385 19012 19389 19068
rect 19389 19012 19445 19068
rect 19445 19012 19449 19068
rect 19385 19008 19449 19012
rect 2820 18532 2884 18596
rect 10916 18532 10980 18596
rect 6150 18524 6214 18528
rect 6150 18468 6154 18524
rect 6154 18468 6210 18524
rect 6210 18468 6214 18524
rect 6150 18464 6214 18468
rect 6230 18524 6294 18528
rect 6230 18468 6234 18524
rect 6234 18468 6290 18524
rect 6290 18468 6294 18524
rect 6230 18464 6294 18468
rect 6310 18524 6374 18528
rect 6310 18468 6314 18524
rect 6314 18468 6370 18524
rect 6370 18468 6374 18524
rect 6310 18464 6374 18468
rect 6390 18524 6454 18528
rect 6390 18468 6394 18524
rect 6394 18468 6450 18524
rect 6450 18468 6454 18524
rect 6390 18464 6454 18468
rect 11348 18524 11412 18528
rect 11348 18468 11352 18524
rect 11352 18468 11408 18524
rect 11408 18468 11412 18524
rect 11348 18464 11412 18468
rect 11428 18524 11492 18528
rect 11428 18468 11432 18524
rect 11432 18468 11488 18524
rect 11488 18468 11492 18524
rect 11428 18464 11492 18468
rect 11508 18524 11572 18528
rect 11508 18468 11512 18524
rect 11512 18468 11568 18524
rect 11568 18468 11572 18524
rect 11508 18464 11572 18468
rect 11588 18524 11652 18528
rect 11588 18468 11592 18524
rect 11592 18468 11648 18524
rect 11648 18468 11652 18524
rect 11588 18464 11652 18468
rect 16546 18524 16610 18528
rect 16546 18468 16550 18524
rect 16550 18468 16606 18524
rect 16606 18468 16610 18524
rect 16546 18464 16610 18468
rect 16626 18524 16690 18528
rect 16626 18468 16630 18524
rect 16630 18468 16686 18524
rect 16686 18468 16690 18524
rect 16626 18464 16690 18468
rect 16706 18524 16770 18528
rect 16706 18468 16710 18524
rect 16710 18468 16766 18524
rect 16766 18468 16770 18524
rect 16706 18464 16770 18468
rect 16786 18524 16850 18528
rect 16786 18468 16790 18524
rect 16790 18468 16846 18524
rect 16846 18468 16850 18524
rect 16786 18464 16850 18468
rect 21744 18524 21808 18528
rect 21744 18468 21748 18524
rect 21748 18468 21804 18524
rect 21804 18468 21808 18524
rect 21744 18464 21808 18468
rect 21824 18524 21888 18528
rect 21824 18468 21828 18524
rect 21828 18468 21884 18524
rect 21884 18468 21888 18524
rect 21824 18464 21888 18468
rect 21904 18524 21968 18528
rect 21904 18468 21908 18524
rect 21908 18468 21964 18524
rect 21964 18468 21968 18524
rect 21904 18464 21968 18468
rect 21984 18524 22048 18528
rect 21984 18468 21988 18524
rect 21988 18468 22044 18524
rect 22044 18468 22048 18524
rect 21984 18464 22048 18468
rect 9260 18396 9324 18460
rect 6684 18048 6748 18052
rect 6684 17992 6698 18048
rect 6698 17992 6748 18048
rect 6684 17988 6748 17992
rect 8156 17988 8220 18052
rect 9444 17988 9508 18052
rect 3551 17980 3615 17984
rect 3551 17924 3555 17980
rect 3555 17924 3611 17980
rect 3611 17924 3615 17980
rect 3551 17920 3615 17924
rect 3631 17980 3695 17984
rect 3631 17924 3635 17980
rect 3635 17924 3691 17980
rect 3691 17924 3695 17980
rect 3631 17920 3695 17924
rect 3711 17980 3775 17984
rect 3711 17924 3715 17980
rect 3715 17924 3771 17980
rect 3771 17924 3775 17980
rect 3711 17920 3775 17924
rect 3791 17980 3855 17984
rect 3791 17924 3795 17980
rect 3795 17924 3851 17980
rect 3851 17924 3855 17980
rect 3791 17920 3855 17924
rect 8749 17980 8813 17984
rect 8749 17924 8753 17980
rect 8753 17924 8809 17980
rect 8809 17924 8813 17980
rect 8749 17920 8813 17924
rect 8829 17980 8893 17984
rect 8829 17924 8833 17980
rect 8833 17924 8889 17980
rect 8889 17924 8893 17980
rect 8829 17920 8893 17924
rect 8909 17980 8973 17984
rect 8909 17924 8913 17980
rect 8913 17924 8969 17980
rect 8969 17924 8973 17980
rect 8909 17920 8973 17924
rect 8989 17980 9053 17984
rect 8989 17924 8993 17980
rect 8993 17924 9049 17980
rect 9049 17924 9053 17980
rect 8989 17920 9053 17924
rect 13947 17980 14011 17984
rect 13947 17924 13951 17980
rect 13951 17924 14007 17980
rect 14007 17924 14011 17980
rect 13947 17920 14011 17924
rect 14027 17980 14091 17984
rect 14027 17924 14031 17980
rect 14031 17924 14087 17980
rect 14087 17924 14091 17980
rect 14027 17920 14091 17924
rect 14107 17980 14171 17984
rect 14107 17924 14111 17980
rect 14111 17924 14167 17980
rect 14167 17924 14171 17980
rect 14107 17920 14171 17924
rect 14187 17980 14251 17984
rect 14187 17924 14191 17980
rect 14191 17924 14247 17980
rect 14247 17924 14251 17980
rect 14187 17920 14251 17924
rect 19145 17980 19209 17984
rect 19145 17924 19149 17980
rect 19149 17924 19205 17980
rect 19205 17924 19209 17980
rect 19145 17920 19209 17924
rect 19225 17980 19289 17984
rect 19225 17924 19229 17980
rect 19229 17924 19285 17980
rect 19285 17924 19289 17980
rect 19225 17920 19289 17924
rect 19305 17980 19369 17984
rect 19305 17924 19309 17980
rect 19309 17924 19365 17980
rect 19365 17924 19369 17980
rect 19305 17920 19369 17924
rect 19385 17980 19449 17984
rect 19385 17924 19389 17980
rect 19389 17924 19445 17980
rect 19445 17924 19449 17980
rect 19385 17920 19449 17924
rect 6150 17436 6214 17440
rect 6150 17380 6154 17436
rect 6154 17380 6210 17436
rect 6210 17380 6214 17436
rect 6150 17376 6214 17380
rect 6230 17436 6294 17440
rect 6230 17380 6234 17436
rect 6234 17380 6290 17436
rect 6290 17380 6294 17436
rect 6230 17376 6294 17380
rect 6310 17436 6374 17440
rect 6310 17380 6314 17436
rect 6314 17380 6370 17436
rect 6370 17380 6374 17436
rect 6310 17376 6374 17380
rect 6390 17436 6454 17440
rect 6390 17380 6394 17436
rect 6394 17380 6450 17436
rect 6450 17380 6454 17436
rect 6390 17376 6454 17380
rect 11348 17436 11412 17440
rect 11348 17380 11352 17436
rect 11352 17380 11408 17436
rect 11408 17380 11412 17436
rect 11348 17376 11412 17380
rect 11428 17436 11492 17440
rect 11428 17380 11432 17436
rect 11432 17380 11488 17436
rect 11488 17380 11492 17436
rect 11428 17376 11492 17380
rect 11508 17436 11572 17440
rect 11508 17380 11512 17436
rect 11512 17380 11568 17436
rect 11568 17380 11572 17436
rect 11508 17376 11572 17380
rect 11588 17436 11652 17440
rect 11588 17380 11592 17436
rect 11592 17380 11648 17436
rect 11648 17380 11652 17436
rect 11588 17376 11652 17380
rect 16546 17436 16610 17440
rect 16546 17380 16550 17436
rect 16550 17380 16606 17436
rect 16606 17380 16610 17436
rect 16546 17376 16610 17380
rect 16626 17436 16690 17440
rect 16626 17380 16630 17436
rect 16630 17380 16686 17436
rect 16686 17380 16690 17436
rect 16626 17376 16690 17380
rect 16706 17436 16770 17440
rect 16706 17380 16710 17436
rect 16710 17380 16766 17436
rect 16766 17380 16770 17436
rect 16706 17376 16770 17380
rect 16786 17436 16850 17440
rect 16786 17380 16790 17436
rect 16790 17380 16846 17436
rect 16846 17380 16850 17436
rect 16786 17376 16850 17380
rect 21744 17436 21808 17440
rect 21744 17380 21748 17436
rect 21748 17380 21804 17436
rect 21804 17380 21808 17436
rect 21744 17376 21808 17380
rect 21824 17436 21888 17440
rect 21824 17380 21828 17436
rect 21828 17380 21884 17436
rect 21884 17380 21888 17436
rect 21824 17376 21888 17380
rect 21904 17436 21968 17440
rect 21904 17380 21908 17436
rect 21908 17380 21964 17436
rect 21964 17380 21968 17436
rect 21904 17376 21968 17380
rect 21984 17436 22048 17440
rect 21984 17380 21988 17436
rect 21988 17380 22044 17436
rect 22044 17380 22048 17436
rect 21984 17376 22048 17380
rect 3551 16892 3615 16896
rect 3551 16836 3555 16892
rect 3555 16836 3611 16892
rect 3611 16836 3615 16892
rect 3551 16832 3615 16836
rect 3631 16892 3695 16896
rect 3631 16836 3635 16892
rect 3635 16836 3691 16892
rect 3691 16836 3695 16892
rect 3631 16832 3695 16836
rect 3711 16892 3775 16896
rect 3711 16836 3715 16892
rect 3715 16836 3771 16892
rect 3771 16836 3775 16892
rect 3711 16832 3775 16836
rect 3791 16892 3855 16896
rect 3791 16836 3795 16892
rect 3795 16836 3851 16892
rect 3851 16836 3855 16892
rect 3791 16832 3855 16836
rect 8749 16892 8813 16896
rect 8749 16836 8753 16892
rect 8753 16836 8809 16892
rect 8809 16836 8813 16892
rect 8749 16832 8813 16836
rect 8829 16892 8893 16896
rect 8829 16836 8833 16892
rect 8833 16836 8889 16892
rect 8889 16836 8893 16892
rect 8829 16832 8893 16836
rect 8909 16892 8973 16896
rect 8909 16836 8913 16892
rect 8913 16836 8969 16892
rect 8969 16836 8973 16892
rect 8909 16832 8973 16836
rect 8989 16892 9053 16896
rect 8989 16836 8993 16892
rect 8993 16836 9049 16892
rect 9049 16836 9053 16892
rect 8989 16832 9053 16836
rect 13947 16892 14011 16896
rect 13947 16836 13951 16892
rect 13951 16836 14007 16892
rect 14007 16836 14011 16892
rect 13947 16832 14011 16836
rect 14027 16892 14091 16896
rect 14027 16836 14031 16892
rect 14031 16836 14087 16892
rect 14087 16836 14091 16892
rect 14027 16832 14091 16836
rect 14107 16892 14171 16896
rect 14107 16836 14111 16892
rect 14111 16836 14167 16892
rect 14167 16836 14171 16892
rect 14107 16832 14171 16836
rect 14187 16892 14251 16896
rect 14187 16836 14191 16892
rect 14191 16836 14247 16892
rect 14247 16836 14251 16892
rect 14187 16832 14251 16836
rect 19145 16892 19209 16896
rect 19145 16836 19149 16892
rect 19149 16836 19205 16892
rect 19205 16836 19209 16892
rect 19145 16832 19209 16836
rect 19225 16892 19289 16896
rect 19225 16836 19229 16892
rect 19229 16836 19285 16892
rect 19285 16836 19289 16892
rect 19225 16832 19289 16836
rect 19305 16892 19369 16896
rect 19305 16836 19309 16892
rect 19309 16836 19365 16892
rect 19365 16836 19369 16892
rect 19305 16832 19369 16836
rect 19385 16892 19449 16896
rect 19385 16836 19389 16892
rect 19389 16836 19445 16892
rect 19445 16836 19449 16892
rect 19385 16832 19449 16836
rect 6868 16628 6932 16692
rect 6150 16348 6214 16352
rect 6150 16292 6154 16348
rect 6154 16292 6210 16348
rect 6210 16292 6214 16348
rect 6150 16288 6214 16292
rect 6230 16348 6294 16352
rect 6230 16292 6234 16348
rect 6234 16292 6290 16348
rect 6290 16292 6294 16348
rect 6230 16288 6294 16292
rect 6310 16348 6374 16352
rect 6310 16292 6314 16348
rect 6314 16292 6370 16348
rect 6370 16292 6374 16348
rect 6310 16288 6374 16292
rect 6390 16348 6454 16352
rect 6390 16292 6394 16348
rect 6394 16292 6450 16348
rect 6450 16292 6454 16348
rect 6390 16288 6454 16292
rect 11348 16348 11412 16352
rect 11348 16292 11352 16348
rect 11352 16292 11408 16348
rect 11408 16292 11412 16348
rect 11348 16288 11412 16292
rect 11428 16348 11492 16352
rect 11428 16292 11432 16348
rect 11432 16292 11488 16348
rect 11488 16292 11492 16348
rect 11428 16288 11492 16292
rect 11508 16348 11572 16352
rect 11508 16292 11512 16348
rect 11512 16292 11568 16348
rect 11568 16292 11572 16348
rect 11508 16288 11572 16292
rect 11588 16348 11652 16352
rect 11588 16292 11592 16348
rect 11592 16292 11648 16348
rect 11648 16292 11652 16348
rect 11588 16288 11652 16292
rect 16546 16348 16610 16352
rect 16546 16292 16550 16348
rect 16550 16292 16606 16348
rect 16606 16292 16610 16348
rect 16546 16288 16610 16292
rect 16626 16348 16690 16352
rect 16626 16292 16630 16348
rect 16630 16292 16686 16348
rect 16686 16292 16690 16348
rect 16626 16288 16690 16292
rect 16706 16348 16770 16352
rect 16706 16292 16710 16348
rect 16710 16292 16766 16348
rect 16766 16292 16770 16348
rect 16706 16288 16770 16292
rect 16786 16348 16850 16352
rect 16786 16292 16790 16348
rect 16790 16292 16846 16348
rect 16846 16292 16850 16348
rect 16786 16288 16850 16292
rect 21744 16348 21808 16352
rect 21744 16292 21748 16348
rect 21748 16292 21804 16348
rect 21804 16292 21808 16348
rect 21744 16288 21808 16292
rect 21824 16348 21888 16352
rect 21824 16292 21828 16348
rect 21828 16292 21884 16348
rect 21884 16292 21888 16348
rect 21824 16288 21888 16292
rect 21904 16348 21968 16352
rect 21904 16292 21908 16348
rect 21908 16292 21964 16348
rect 21964 16292 21968 16348
rect 21904 16288 21968 16292
rect 21984 16348 22048 16352
rect 21984 16292 21988 16348
rect 21988 16292 22044 16348
rect 22044 16292 22048 16348
rect 21984 16288 22048 16292
rect 7236 15812 7300 15876
rect 3551 15804 3615 15808
rect 3551 15748 3555 15804
rect 3555 15748 3611 15804
rect 3611 15748 3615 15804
rect 3551 15744 3615 15748
rect 3631 15804 3695 15808
rect 3631 15748 3635 15804
rect 3635 15748 3691 15804
rect 3691 15748 3695 15804
rect 3631 15744 3695 15748
rect 3711 15804 3775 15808
rect 3711 15748 3715 15804
rect 3715 15748 3771 15804
rect 3771 15748 3775 15804
rect 3711 15744 3775 15748
rect 3791 15804 3855 15808
rect 3791 15748 3795 15804
rect 3795 15748 3851 15804
rect 3851 15748 3855 15804
rect 3791 15744 3855 15748
rect 8749 15804 8813 15808
rect 8749 15748 8753 15804
rect 8753 15748 8809 15804
rect 8809 15748 8813 15804
rect 8749 15744 8813 15748
rect 8829 15804 8893 15808
rect 8829 15748 8833 15804
rect 8833 15748 8889 15804
rect 8889 15748 8893 15804
rect 8829 15744 8893 15748
rect 8909 15804 8973 15808
rect 8909 15748 8913 15804
rect 8913 15748 8969 15804
rect 8969 15748 8973 15804
rect 8909 15744 8973 15748
rect 8989 15804 9053 15808
rect 8989 15748 8993 15804
rect 8993 15748 9049 15804
rect 9049 15748 9053 15804
rect 8989 15744 9053 15748
rect 13947 15804 14011 15808
rect 13947 15748 13951 15804
rect 13951 15748 14007 15804
rect 14007 15748 14011 15804
rect 13947 15744 14011 15748
rect 14027 15804 14091 15808
rect 14027 15748 14031 15804
rect 14031 15748 14087 15804
rect 14087 15748 14091 15804
rect 14027 15744 14091 15748
rect 14107 15804 14171 15808
rect 14107 15748 14111 15804
rect 14111 15748 14167 15804
rect 14167 15748 14171 15804
rect 14107 15744 14171 15748
rect 14187 15804 14251 15808
rect 14187 15748 14191 15804
rect 14191 15748 14247 15804
rect 14247 15748 14251 15804
rect 14187 15744 14251 15748
rect 19145 15804 19209 15808
rect 19145 15748 19149 15804
rect 19149 15748 19205 15804
rect 19205 15748 19209 15804
rect 19145 15744 19209 15748
rect 19225 15804 19289 15808
rect 19225 15748 19229 15804
rect 19229 15748 19285 15804
rect 19285 15748 19289 15804
rect 19225 15744 19289 15748
rect 19305 15804 19369 15808
rect 19305 15748 19309 15804
rect 19309 15748 19365 15804
rect 19365 15748 19369 15804
rect 19305 15744 19369 15748
rect 19385 15804 19449 15808
rect 19385 15748 19389 15804
rect 19389 15748 19445 15804
rect 19445 15748 19449 15804
rect 19385 15744 19449 15748
rect 9444 15328 9508 15332
rect 9444 15272 9458 15328
rect 9458 15272 9508 15328
rect 9444 15268 9508 15272
rect 6150 15260 6214 15264
rect 6150 15204 6154 15260
rect 6154 15204 6210 15260
rect 6210 15204 6214 15260
rect 6150 15200 6214 15204
rect 6230 15260 6294 15264
rect 6230 15204 6234 15260
rect 6234 15204 6290 15260
rect 6290 15204 6294 15260
rect 6230 15200 6294 15204
rect 6310 15260 6374 15264
rect 6310 15204 6314 15260
rect 6314 15204 6370 15260
rect 6370 15204 6374 15260
rect 6310 15200 6374 15204
rect 6390 15260 6454 15264
rect 6390 15204 6394 15260
rect 6394 15204 6450 15260
rect 6450 15204 6454 15260
rect 6390 15200 6454 15204
rect 11348 15260 11412 15264
rect 11348 15204 11352 15260
rect 11352 15204 11408 15260
rect 11408 15204 11412 15260
rect 11348 15200 11412 15204
rect 11428 15260 11492 15264
rect 11428 15204 11432 15260
rect 11432 15204 11488 15260
rect 11488 15204 11492 15260
rect 11428 15200 11492 15204
rect 11508 15260 11572 15264
rect 11508 15204 11512 15260
rect 11512 15204 11568 15260
rect 11568 15204 11572 15260
rect 11508 15200 11572 15204
rect 11588 15260 11652 15264
rect 11588 15204 11592 15260
rect 11592 15204 11648 15260
rect 11648 15204 11652 15260
rect 11588 15200 11652 15204
rect 16546 15260 16610 15264
rect 16546 15204 16550 15260
rect 16550 15204 16606 15260
rect 16606 15204 16610 15260
rect 16546 15200 16610 15204
rect 16626 15260 16690 15264
rect 16626 15204 16630 15260
rect 16630 15204 16686 15260
rect 16686 15204 16690 15260
rect 16626 15200 16690 15204
rect 16706 15260 16770 15264
rect 16706 15204 16710 15260
rect 16710 15204 16766 15260
rect 16766 15204 16770 15260
rect 16706 15200 16770 15204
rect 16786 15260 16850 15264
rect 16786 15204 16790 15260
rect 16790 15204 16846 15260
rect 16846 15204 16850 15260
rect 16786 15200 16850 15204
rect 21744 15260 21808 15264
rect 21744 15204 21748 15260
rect 21748 15204 21804 15260
rect 21804 15204 21808 15260
rect 21744 15200 21808 15204
rect 21824 15260 21888 15264
rect 21824 15204 21828 15260
rect 21828 15204 21884 15260
rect 21884 15204 21888 15260
rect 21824 15200 21888 15204
rect 21904 15260 21968 15264
rect 21904 15204 21908 15260
rect 21908 15204 21964 15260
rect 21964 15204 21968 15260
rect 21904 15200 21968 15204
rect 21984 15260 22048 15264
rect 21984 15204 21988 15260
rect 21988 15204 22044 15260
rect 22044 15204 22048 15260
rect 21984 15200 22048 15204
rect 5580 14860 5644 14924
rect 10180 14784 10244 14788
rect 10180 14728 10230 14784
rect 10230 14728 10244 14784
rect 10180 14724 10244 14728
rect 3551 14716 3615 14720
rect 3551 14660 3555 14716
rect 3555 14660 3611 14716
rect 3611 14660 3615 14716
rect 3551 14656 3615 14660
rect 3631 14716 3695 14720
rect 3631 14660 3635 14716
rect 3635 14660 3691 14716
rect 3691 14660 3695 14716
rect 3631 14656 3695 14660
rect 3711 14716 3775 14720
rect 3711 14660 3715 14716
rect 3715 14660 3771 14716
rect 3771 14660 3775 14716
rect 3711 14656 3775 14660
rect 3791 14716 3855 14720
rect 3791 14660 3795 14716
rect 3795 14660 3851 14716
rect 3851 14660 3855 14716
rect 3791 14656 3855 14660
rect 8749 14716 8813 14720
rect 8749 14660 8753 14716
rect 8753 14660 8809 14716
rect 8809 14660 8813 14716
rect 8749 14656 8813 14660
rect 8829 14716 8893 14720
rect 8829 14660 8833 14716
rect 8833 14660 8889 14716
rect 8889 14660 8893 14716
rect 8829 14656 8893 14660
rect 8909 14716 8973 14720
rect 8909 14660 8913 14716
rect 8913 14660 8969 14716
rect 8969 14660 8973 14716
rect 8909 14656 8973 14660
rect 8989 14716 9053 14720
rect 8989 14660 8993 14716
rect 8993 14660 9049 14716
rect 9049 14660 9053 14716
rect 8989 14656 9053 14660
rect 13947 14716 14011 14720
rect 13947 14660 13951 14716
rect 13951 14660 14007 14716
rect 14007 14660 14011 14716
rect 13947 14656 14011 14660
rect 14027 14716 14091 14720
rect 14027 14660 14031 14716
rect 14031 14660 14087 14716
rect 14087 14660 14091 14716
rect 14027 14656 14091 14660
rect 14107 14716 14171 14720
rect 14107 14660 14111 14716
rect 14111 14660 14167 14716
rect 14167 14660 14171 14716
rect 14107 14656 14171 14660
rect 14187 14716 14251 14720
rect 14187 14660 14191 14716
rect 14191 14660 14247 14716
rect 14247 14660 14251 14716
rect 14187 14656 14251 14660
rect 19145 14716 19209 14720
rect 19145 14660 19149 14716
rect 19149 14660 19205 14716
rect 19205 14660 19209 14716
rect 19145 14656 19209 14660
rect 19225 14716 19289 14720
rect 19225 14660 19229 14716
rect 19229 14660 19285 14716
rect 19285 14660 19289 14716
rect 19225 14656 19289 14660
rect 19305 14716 19369 14720
rect 19305 14660 19309 14716
rect 19309 14660 19365 14716
rect 19365 14660 19369 14716
rect 19305 14656 19369 14660
rect 19385 14716 19449 14720
rect 19385 14660 19389 14716
rect 19389 14660 19445 14716
rect 19445 14660 19449 14716
rect 19385 14656 19449 14660
rect 7788 14240 7852 14244
rect 7788 14184 7838 14240
rect 7838 14184 7852 14240
rect 7788 14180 7852 14184
rect 6150 14172 6214 14176
rect 6150 14116 6154 14172
rect 6154 14116 6210 14172
rect 6210 14116 6214 14172
rect 6150 14112 6214 14116
rect 6230 14172 6294 14176
rect 6230 14116 6234 14172
rect 6234 14116 6290 14172
rect 6290 14116 6294 14172
rect 6230 14112 6294 14116
rect 6310 14172 6374 14176
rect 6310 14116 6314 14172
rect 6314 14116 6370 14172
rect 6370 14116 6374 14172
rect 6310 14112 6374 14116
rect 6390 14172 6454 14176
rect 6390 14116 6394 14172
rect 6394 14116 6450 14172
rect 6450 14116 6454 14172
rect 6390 14112 6454 14116
rect 11348 14172 11412 14176
rect 11348 14116 11352 14172
rect 11352 14116 11408 14172
rect 11408 14116 11412 14172
rect 11348 14112 11412 14116
rect 11428 14172 11492 14176
rect 11428 14116 11432 14172
rect 11432 14116 11488 14172
rect 11488 14116 11492 14172
rect 11428 14112 11492 14116
rect 11508 14172 11572 14176
rect 11508 14116 11512 14172
rect 11512 14116 11568 14172
rect 11568 14116 11572 14172
rect 11508 14112 11572 14116
rect 11588 14172 11652 14176
rect 11588 14116 11592 14172
rect 11592 14116 11648 14172
rect 11648 14116 11652 14172
rect 11588 14112 11652 14116
rect 16546 14172 16610 14176
rect 16546 14116 16550 14172
rect 16550 14116 16606 14172
rect 16606 14116 16610 14172
rect 16546 14112 16610 14116
rect 16626 14172 16690 14176
rect 16626 14116 16630 14172
rect 16630 14116 16686 14172
rect 16686 14116 16690 14172
rect 16626 14112 16690 14116
rect 16706 14172 16770 14176
rect 16706 14116 16710 14172
rect 16710 14116 16766 14172
rect 16766 14116 16770 14172
rect 16706 14112 16770 14116
rect 16786 14172 16850 14176
rect 16786 14116 16790 14172
rect 16790 14116 16846 14172
rect 16846 14116 16850 14172
rect 16786 14112 16850 14116
rect 21744 14172 21808 14176
rect 21744 14116 21748 14172
rect 21748 14116 21804 14172
rect 21804 14116 21808 14172
rect 21744 14112 21808 14116
rect 21824 14172 21888 14176
rect 21824 14116 21828 14172
rect 21828 14116 21884 14172
rect 21884 14116 21888 14172
rect 21824 14112 21888 14116
rect 21904 14172 21968 14176
rect 21904 14116 21908 14172
rect 21908 14116 21964 14172
rect 21964 14116 21968 14172
rect 21904 14112 21968 14116
rect 21984 14172 22048 14176
rect 21984 14116 21988 14172
rect 21988 14116 22044 14172
rect 22044 14116 22048 14172
rect 21984 14112 22048 14116
rect 2820 13772 2884 13836
rect 5764 13636 5828 13700
rect 3551 13628 3615 13632
rect 3551 13572 3555 13628
rect 3555 13572 3611 13628
rect 3611 13572 3615 13628
rect 3551 13568 3615 13572
rect 3631 13628 3695 13632
rect 3631 13572 3635 13628
rect 3635 13572 3691 13628
rect 3691 13572 3695 13628
rect 3631 13568 3695 13572
rect 3711 13628 3775 13632
rect 3711 13572 3715 13628
rect 3715 13572 3771 13628
rect 3771 13572 3775 13628
rect 3711 13568 3775 13572
rect 3791 13628 3855 13632
rect 3791 13572 3795 13628
rect 3795 13572 3851 13628
rect 3851 13572 3855 13628
rect 3791 13568 3855 13572
rect 8749 13628 8813 13632
rect 8749 13572 8753 13628
rect 8753 13572 8809 13628
rect 8809 13572 8813 13628
rect 8749 13568 8813 13572
rect 8829 13628 8893 13632
rect 8829 13572 8833 13628
rect 8833 13572 8889 13628
rect 8889 13572 8893 13628
rect 8829 13568 8893 13572
rect 8909 13628 8973 13632
rect 8909 13572 8913 13628
rect 8913 13572 8969 13628
rect 8969 13572 8973 13628
rect 8909 13568 8973 13572
rect 8989 13628 9053 13632
rect 8989 13572 8993 13628
rect 8993 13572 9049 13628
rect 9049 13572 9053 13628
rect 8989 13568 9053 13572
rect 13947 13628 14011 13632
rect 13947 13572 13951 13628
rect 13951 13572 14007 13628
rect 14007 13572 14011 13628
rect 13947 13568 14011 13572
rect 14027 13628 14091 13632
rect 14027 13572 14031 13628
rect 14031 13572 14087 13628
rect 14087 13572 14091 13628
rect 14027 13568 14091 13572
rect 14107 13628 14171 13632
rect 14107 13572 14111 13628
rect 14111 13572 14167 13628
rect 14167 13572 14171 13628
rect 14107 13568 14171 13572
rect 14187 13628 14251 13632
rect 14187 13572 14191 13628
rect 14191 13572 14247 13628
rect 14247 13572 14251 13628
rect 14187 13568 14251 13572
rect 19145 13628 19209 13632
rect 19145 13572 19149 13628
rect 19149 13572 19205 13628
rect 19205 13572 19209 13628
rect 19145 13568 19209 13572
rect 19225 13628 19289 13632
rect 19225 13572 19229 13628
rect 19229 13572 19285 13628
rect 19285 13572 19289 13628
rect 19225 13568 19289 13572
rect 19305 13628 19369 13632
rect 19305 13572 19309 13628
rect 19309 13572 19365 13628
rect 19365 13572 19369 13628
rect 19305 13568 19369 13572
rect 19385 13628 19449 13632
rect 19385 13572 19389 13628
rect 19389 13572 19445 13628
rect 19445 13572 19449 13628
rect 19385 13568 19449 13572
rect 6150 13084 6214 13088
rect 6150 13028 6154 13084
rect 6154 13028 6210 13084
rect 6210 13028 6214 13084
rect 6150 13024 6214 13028
rect 6230 13084 6294 13088
rect 6230 13028 6234 13084
rect 6234 13028 6290 13084
rect 6290 13028 6294 13084
rect 6230 13024 6294 13028
rect 6310 13084 6374 13088
rect 6310 13028 6314 13084
rect 6314 13028 6370 13084
rect 6370 13028 6374 13084
rect 6310 13024 6374 13028
rect 6390 13084 6454 13088
rect 6390 13028 6394 13084
rect 6394 13028 6450 13084
rect 6450 13028 6454 13084
rect 6390 13024 6454 13028
rect 11348 13084 11412 13088
rect 11348 13028 11352 13084
rect 11352 13028 11408 13084
rect 11408 13028 11412 13084
rect 11348 13024 11412 13028
rect 11428 13084 11492 13088
rect 11428 13028 11432 13084
rect 11432 13028 11488 13084
rect 11488 13028 11492 13084
rect 11428 13024 11492 13028
rect 11508 13084 11572 13088
rect 11508 13028 11512 13084
rect 11512 13028 11568 13084
rect 11568 13028 11572 13084
rect 11508 13024 11572 13028
rect 11588 13084 11652 13088
rect 11588 13028 11592 13084
rect 11592 13028 11648 13084
rect 11648 13028 11652 13084
rect 11588 13024 11652 13028
rect 16546 13084 16610 13088
rect 16546 13028 16550 13084
rect 16550 13028 16606 13084
rect 16606 13028 16610 13084
rect 16546 13024 16610 13028
rect 16626 13084 16690 13088
rect 16626 13028 16630 13084
rect 16630 13028 16686 13084
rect 16686 13028 16690 13084
rect 16626 13024 16690 13028
rect 16706 13084 16770 13088
rect 16706 13028 16710 13084
rect 16710 13028 16766 13084
rect 16766 13028 16770 13084
rect 16706 13024 16770 13028
rect 16786 13084 16850 13088
rect 16786 13028 16790 13084
rect 16790 13028 16846 13084
rect 16846 13028 16850 13084
rect 16786 13024 16850 13028
rect 21744 13084 21808 13088
rect 21744 13028 21748 13084
rect 21748 13028 21804 13084
rect 21804 13028 21808 13084
rect 21744 13024 21808 13028
rect 21824 13084 21888 13088
rect 21824 13028 21828 13084
rect 21828 13028 21884 13084
rect 21884 13028 21888 13084
rect 21824 13024 21888 13028
rect 21904 13084 21968 13088
rect 21904 13028 21908 13084
rect 21908 13028 21964 13084
rect 21964 13028 21968 13084
rect 21904 13024 21968 13028
rect 21984 13084 22048 13088
rect 21984 13028 21988 13084
rect 21988 13028 22044 13084
rect 22044 13028 22048 13084
rect 21984 13024 22048 13028
rect 11836 12956 11900 13020
rect 5948 12684 6012 12748
rect 3551 12540 3615 12544
rect 3551 12484 3555 12540
rect 3555 12484 3611 12540
rect 3611 12484 3615 12540
rect 3551 12480 3615 12484
rect 3631 12540 3695 12544
rect 3631 12484 3635 12540
rect 3635 12484 3691 12540
rect 3691 12484 3695 12540
rect 3631 12480 3695 12484
rect 3711 12540 3775 12544
rect 3711 12484 3715 12540
rect 3715 12484 3771 12540
rect 3771 12484 3775 12540
rect 3711 12480 3775 12484
rect 3791 12540 3855 12544
rect 3791 12484 3795 12540
rect 3795 12484 3851 12540
rect 3851 12484 3855 12540
rect 3791 12480 3855 12484
rect 8749 12540 8813 12544
rect 8749 12484 8753 12540
rect 8753 12484 8809 12540
rect 8809 12484 8813 12540
rect 8749 12480 8813 12484
rect 8829 12540 8893 12544
rect 8829 12484 8833 12540
rect 8833 12484 8889 12540
rect 8889 12484 8893 12540
rect 8829 12480 8893 12484
rect 8909 12540 8973 12544
rect 8909 12484 8913 12540
rect 8913 12484 8969 12540
rect 8969 12484 8973 12540
rect 8909 12480 8973 12484
rect 8989 12540 9053 12544
rect 8989 12484 8993 12540
rect 8993 12484 9049 12540
rect 9049 12484 9053 12540
rect 8989 12480 9053 12484
rect 9628 12412 9692 12476
rect 13947 12540 14011 12544
rect 13947 12484 13951 12540
rect 13951 12484 14007 12540
rect 14007 12484 14011 12540
rect 13947 12480 14011 12484
rect 14027 12540 14091 12544
rect 14027 12484 14031 12540
rect 14031 12484 14087 12540
rect 14087 12484 14091 12540
rect 14027 12480 14091 12484
rect 14107 12540 14171 12544
rect 14107 12484 14111 12540
rect 14111 12484 14167 12540
rect 14167 12484 14171 12540
rect 14107 12480 14171 12484
rect 14187 12540 14251 12544
rect 14187 12484 14191 12540
rect 14191 12484 14247 12540
rect 14247 12484 14251 12540
rect 14187 12480 14251 12484
rect 19145 12540 19209 12544
rect 19145 12484 19149 12540
rect 19149 12484 19205 12540
rect 19205 12484 19209 12540
rect 19145 12480 19209 12484
rect 19225 12540 19289 12544
rect 19225 12484 19229 12540
rect 19229 12484 19285 12540
rect 19285 12484 19289 12540
rect 19225 12480 19289 12484
rect 19305 12540 19369 12544
rect 19305 12484 19309 12540
rect 19309 12484 19365 12540
rect 19365 12484 19369 12540
rect 19305 12480 19369 12484
rect 19385 12540 19449 12544
rect 19385 12484 19389 12540
rect 19389 12484 19445 12540
rect 19445 12484 19449 12540
rect 19385 12480 19449 12484
rect 9628 12004 9692 12068
rect 6150 11996 6214 12000
rect 6150 11940 6154 11996
rect 6154 11940 6210 11996
rect 6210 11940 6214 11996
rect 6150 11936 6214 11940
rect 6230 11996 6294 12000
rect 6230 11940 6234 11996
rect 6234 11940 6290 11996
rect 6290 11940 6294 11996
rect 6230 11936 6294 11940
rect 6310 11996 6374 12000
rect 6310 11940 6314 11996
rect 6314 11940 6370 11996
rect 6370 11940 6374 11996
rect 6310 11936 6374 11940
rect 6390 11996 6454 12000
rect 6390 11940 6394 11996
rect 6394 11940 6450 11996
rect 6450 11940 6454 11996
rect 6390 11936 6454 11940
rect 11348 11996 11412 12000
rect 11348 11940 11352 11996
rect 11352 11940 11408 11996
rect 11408 11940 11412 11996
rect 11348 11936 11412 11940
rect 11428 11996 11492 12000
rect 11428 11940 11432 11996
rect 11432 11940 11488 11996
rect 11488 11940 11492 11996
rect 11428 11936 11492 11940
rect 11508 11996 11572 12000
rect 11508 11940 11512 11996
rect 11512 11940 11568 11996
rect 11568 11940 11572 11996
rect 11508 11936 11572 11940
rect 11588 11996 11652 12000
rect 11588 11940 11592 11996
rect 11592 11940 11648 11996
rect 11648 11940 11652 11996
rect 11588 11936 11652 11940
rect 16546 11996 16610 12000
rect 16546 11940 16550 11996
rect 16550 11940 16606 11996
rect 16606 11940 16610 11996
rect 16546 11936 16610 11940
rect 16626 11996 16690 12000
rect 16626 11940 16630 11996
rect 16630 11940 16686 11996
rect 16686 11940 16690 11996
rect 16626 11936 16690 11940
rect 16706 11996 16770 12000
rect 16706 11940 16710 11996
rect 16710 11940 16766 11996
rect 16766 11940 16770 11996
rect 16706 11936 16770 11940
rect 16786 11996 16850 12000
rect 16786 11940 16790 11996
rect 16790 11940 16846 11996
rect 16846 11940 16850 11996
rect 16786 11936 16850 11940
rect 21744 11996 21808 12000
rect 21744 11940 21748 11996
rect 21748 11940 21804 11996
rect 21804 11940 21808 11996
rect 21744 11936 21808 11940
rect 21824 11996 21888 12000
rect 21824 11940 21828 11996
rect 21828 11940 21884 11996
rect 21884 11940 21888 11996
rect 21824 11936 21888 11940
rect 21904 11996 21968 12000
rect 21904 11940 21908 11996
rect 21908 11940 21964 11996
rect 21964 11940 21968 11996
rect 21904 11936 21968 11940
rect 21984 11996 22048 12000
rect 21984 11940 21988 11996
rect 21988 11940 22044 11996
rect 22044 11940 22048 11996
rect 21984 11936 22048 11940
rect 8524 11868 8588 11932
rect 10180 11868 10244 11932
rect 12020 11656 12084 11660
rect 12020 11600 12070 11656
rect 12070 11600 12084 11656
rect 12020 11596 12084 11600
rect 3551 11452 3615 11456
rect 3551 11396 3555 11452
rect 3555 11396 3611 11452
rect 3611 11396 3615 11452
rect 3551 11392 3615 11396
rect 3631 11452 3695 11456
rect 3631 11396 3635 11452
rect 3635 11396 3691 11452
rect 3691 11396 3695 11452
rect 3631 11392 3695 11396
rect 3711 11452 3775 11456
rect 3711 11396 3715 11452
rect 3715 11396 3771 11452
rect 3771 11396 3775 11452
rect 3711 11392 3775 11396
rect 3791 11452 3855 11456
rect 3791 11396 3795 11452
rect 3795 11396 3851 11452
rect 3851 11396 3855 11452
rect 3791 11392 3855 11396
rect 8749 11452 8813 11456
rect 8749 11396 8753 11452
rect 8753 11396 8809 11452
rect 8809 11396 8813 11452
rect 8749 11392 8813 11396
rect 8829 11452 8893 11456
rect 8829 11396 8833 11452
rect 8833 11396 8889 11452
rect 8889 11396 8893 11452
rect 8829 11392 8893 11396
rect 8909 11452 8973 11456
rect 8909 11396 8913 11452
rect 8913 11396 8969 11452
rect 8969 11396 8973 11452
rect 8909 11392 8973 11396
rect 8989 11452 9053 11456
rect 8989 11396 8993 11452
rect 8993 11396 9049 11452
rect 9049 11396 9053 11452
rect 8989 11392 9053 11396
rect 13947 11452 14011 11456
rect 13947 11396 13951 11452
rect 13951 11396 14007 11452
rect 14007 11396 14011 11452
rect 13947 11392 14011 11396
rect 14027 11452 14091 11456
rect 14027 11396 14031 11452
rect 14031 11396 14087 11452
rect 14087 11396 14091 11452
rect 14027 11392 14091 11396
rect 14107 11452 14171 11456
rect 14107 11396 14111 11452
rect 14111 11396 14167 11452
rect 14167 11396 14171 11452
rect 14107 11392 14171 11396
rect 14187 11452 14251 11456
rect 14187 11396 14191 11452
rect 14191 11396 14247 11452
rect 14247 11396 14251 11452
rect 14187 11392 14251 11396
rect 19145 11452 19209 11456
rect 19145 11396 19149 11452
rect 19149 11396 19205 11452
rect 19205 11396 19209 11452
rect 19145 11392 19209 11396
rect 19225 11452 19289 11456
rect 19225 11396 19229 11452
rect 19229 11396 19285 11452
rect 19285 11396 19289 11452
rect 19225 11392 19289 11396
rect 19305 11452 19369 11456
rect 19305 11396 19309 11452
rect 19309 11396 19365 11452
rect 19365 11396 19369 11452
rect 19305 11392 19369 11396
rect 19385 11452 19449 11456
rect 19385 11396 19389 11452
rect 19389 11396 19445 11452
rect 19445 11396 19449 11452
rect 19385 11392 19449 11396
rect 11100 11324 11164 11388
rect 5580 11112 5644 11116
rect 5580 11056 5630 11112
rect 5630 11056 5644 11112
rect 5580 11052 5644 11056
rect 9812 11052 9876 11116
rect 6150 10908 6214 10912
rect 6150 10852 6154 10908
rect 6154 10852 6210 10908
rect 6210 10852 6214 10908
rect 6150 10848 6214 10852
rect 6230 10908 6294 10912
rect 6230 10852 6234 10908
rect 6234 10852 6290 10908
rect 6290 10852 6294 10908
rect 6230 10848 6294 10852
rect 6310 10908 6374 10912
rect 6310 10852 6314 10908
rect 6314 10852 6370 10908
rect 6370 10852 6374 10908
rect 6310 10848 6374 10852
rect 6390 10908 6454 10912
rect 6390 10852 6394 10908
rect 6394 10852 6450 10908
rect 6450 10852 6454 10908
rect 6390 10848 6454 10852
rect 11348 10908 11412 10912
rect 11348 10852 11352 10908
rect 11352 10852 11408 10908
rect 11408 10852 11412 10908
rect 11348 10848 11412 10852
rect 11428 10908 11492 10912
rect 11428 10852 11432 10908
rect 11432 10852 11488 10908
rect 11488 10852 11492 10908
rect 11428 10848 11492 10852
rect 11508 10908 11572 10912
rect 11508 10852 11512 10908
rect 11512 10852 11568 10908
rect 11568 10852 11572 10908
rect 11508 10848 11572 10852
rect 11588 10908 11652 10912
rect 11588 10852 11592 10908
rect 11592 10852 11648 10908
rect 11648 10852 11652 10908
rect 11588 10848 11652 10852
rect 16546 10908 16610 10912
rect 16546 10852 16550 10908
rect 16550 10852 16606 10908
rect 16606 10852 16610 10908
rect 16546 10848 16610 10852
rect 16626 10908 16690 10912
rect 16626 10852 16630 10908
rect 16630 10852 16686 10908
rect 16686 10852 16690 10908
rect 16626 10848 16690 10852
rect 16706 10908 16770 10912
rect 16706 10852 16710 10908
rect 16710 10852 16766 10908
rect 16766 10852 16770 10908
rect 16706 10848 16770 10852
rect 16786 10908 16850 10912
rect 16786 10852 16790 10908
rect 16790 10852 16846 10908
rect 16846 10852 16850 10908
rect 16786 10848 16850 10852
rect 21744 10908 21808 10912
rect 21744 10852 21748 10908
rect 21748 10852 21804 10908
rect 21804 10852 21808 10908
rect 21744 10848 21808 10852
rect 21824 10908 21888 10912
rect 21824 10852 21828 10908
rect 21828 10852 21884 10908
rect 21884 10852 21888 10908
rect 21824 10848 21888 10852
rect 21904 10908 21968 10912
rect 21904 10852 21908 10908
rect 21908 10852 21964 10908
rect 21964 10852 21968 10908
rect 21904 10848 21968 10852
rect 21984 10908 22048 10912
rect 21984 10852 21988 10908
rect 21988 10852 22044 10908
rect 22044 10852 22048 10908
rect 21984 10848 22048 10852
rect 11836 10508 11900 10572
rect 7236 10372 7300 10436
rect 3551 10364 3615 10368
rect 3551 10308 3555 10364
rect 3555 10308 3611 10364
rect 3611 10308 3615 10364
rect 3551 10304 3615 10308
rect 3631 10364 3695 10368
rect 3631 10308 3635 10364
rect 3635 10308 3691 10364
rect 3691 10308 3695 10364
rect 3631 10304 3695 10308
rect 3711 10364 3775 10368
rect 3711 10308 3715 10364
rect 3715 10308 3771 10364
rect 3771 10308 3775 10364
rect 3711 10304 3775 10308
rect 3791 10364 3855 10368
rect 3791 10308 3795 10364
rect 3795 10308 3851 10364
rect 3851 10308 3855 10364
rect 3791 10304 3855 10308
rect 8749 10364 8813 10368
rect 8749 10308 8753 10364
rect 8753 10308 8809 10364
rect 8809 10308 8813 10364
rect 8749 10304 8813 10308
rect 8829 10364 8893 10368
rect 8829 10308 8833 10364
rect 8833 10308 8889 10364
rect 8889 10308 8893 10364
rect 8829 10304 8893 10308
rect 8909 10364 8973 10368
rect 8909 10308 8913 10364
rect 8913 10308 8969 10364
rect 8969 10308 8973 10364
rect 8909 10304 8973 10308
rect 8989 10364 9053 10368
rect 8989 10308 8993 10364
rect 8993 10308 9049 10364
rect 9049 10308 9053 10364
rect 8989 10304 9053 10308
rect 13947 10364 14011 10368
rect 13947 10308 13951 10364
rect 13951 10308 14007 10364
rect 14007 10308 14011 10364
rect 13947 10304 14011 10308
rect 14027 10364 14091 10368
rect 14027 10308 14031 10364
rect 14031 10308 14087 10364
rect 14087 10308 14091 10364
rect 14027 10304 14091 10308
rect 14107 10364 14171 10368
rect 14107 10308 14111 10364
rect 14111 10308 14167 10364
rect 14167 10308 14171 10364
rect 14107 10304 14171 10308
rect 14187 10364 14251 10368
rect 14187 10308 14191 10364
rect 14191 10308 14247 10364
rect 14247 10308 14251 10364
rect 14187 10304 14251 10308
rect 19145 10364 19209 10368
rect 19145 10308 19149 10364
rect 19149 10308 19205 10364
rect 19205 10308 19209 10364
rect 19145 10304 19209 10308
rect 19225 10364 19289 10368
rect 19225 10308 19229 10364
rect 19229 10308 19285 10364
rect 19285 10308 19289 10364
rect 19225 10304 19289 10308
rect 19305 10364 19369 10368
rect 19305 10308 19309 10364
rect 19309 10308 19365 10364
rect 19365 10308 19369 10364
rect 19305 10304 19369 10308
rect 19385 10364 19449 10368
rect 19385 10308 19389 10364
rect 19389 10308 19445 10364
rect 19445 10308 19449 10364
rect 19385 10304 19449 10308
rect 10916 10100 10980 10164
rect 11100 9964 11164 10028
rect 6150 9820 6214 9824
rect 6150 9764 6154 9820
rect 6154 9764 6210 9820
rect 6210 9764 6214 9820
rect 6150 9760 6214 9764
rect 6230 9820 6294 9824
rect 6230 9764 6234 9820
rect 6234 9764 6290 9820
rect 6290 9764 6294 9820
rect 6230 9760 6294 9764
rect 6310 9820 6374 9824
rect 6310 9764 6314 9820
rect 6314 9764 6370 9820
rect 6370 9764 6374 9820
rect 6310 9760 6374 9764
rect 6390 9820 6454 9824
rect 6390 9764 6394 9820
rect 6394 9764 6450 9820
rect 6450 9764 6454 9820
rect 6390 9760 6454 9764
rect 11348 9820 11412 9824
rect 11348 9764 11352 9820
rect 11352 9764 11408 9820
rect 11408 9764 11412 9820
rect 11348 9760 11412 9764
rect 11428 9820 11492 9824
rect 11428 9764 11432 9820
rect 11432 9764 11488 9820
rect 11488 9764 11492 9820
rect 11428 9760 11492 9764
rect 11508 9820 11572 9824
rect 11508 9764 11512 9820
rect 11512 9764 11568 9820
rect 11568 9764 11572 9820
rect 11508 9760 11572 9764
rect 11588 9820 11652 9824
rect 11588 9764 11592 9820
rect 11592 9764 11648 9820
rect 11648 9764 11652 9820
rect 11588 9760 11652 9764
rect 16546 9820 16610 9824
rect 16546 9764 16550 9820
rect 16550 9764 16606 9820
rect 16606 9764 16610 9820
rect 16546 9760 16610 9764
rect 16626 9820 16690 9824
rect 16626 9764 16630 9820
rect 16630 9764 16686 9820
rect 16686 9764 16690 9820
rect 16626 9760 16690 9764
rect 16706 9820 16770 9824
rect 16706 9764 16710 9820
rect 16710 9764 16766 9820
rect 16766 9764 16770 9820
rect 16706 9760 16770 9764
rect 16786 9820 16850 9824
rect 16786 9764 16790 9820
rect 16790 9764 16846 9820
rect 16846 9764 16850 9820
rect 16786 9760 16850 9764
rect 21744 9820 21808 9824
rect 21744 9764 21748 9820
rect 21748 9764 21804 9820
rect 21804 9764 21808 9820
rect 21744 9760 21808 9764
rect 21824 9820 21888 9824
rect 21824 9764 21828 9820
rect 21828 9764 21884 9820
rect 21884 9764 21888 9820
rect 21824 9760 21888 9764
rect 21904 9820 21968 9824
rect 21904 9764 21908 9820
rect 21908 9764 21964 9820
rect 21964 9764 21968 9820
rect 21904 9760 21968 9764
rect 21984 9820 22048 9824
rect 21984 9764 21988 9820
rect 21988 9764 22044 9820
rect 22044 9764 22048 9820
rect 21984 9760 22048 9764
rect 10180 9616 10244 9620
rect 10180 9560 10194 9616
rect 10194 9560 10244 9616
rect 10180 9556 10244 9560
rect 3551 9276 3615 9280
rect 3551 9220 3555 9276
rect 3555 9220 3611 9276
rect 3611 9220 3615 9276
rect 3551 9216 3615 9220
rect 3631 9276 3695 9280
rect 3631 9220 3635 9276
rect 3635 9220 3691 9276
rect 3691 9220 3695 9276
rect 3631 9216 3695 9220
rect 3711 9276 3775 9280
rect 3711 9220 3715 9276
rect 3715 9220 3771 9276
rect 3771 9220 3775 9276
rect 3711 9216 3775 9220
rect 3791 9276 3855 9280
rect 3791 9220 3795 9276
rect 3795 9220 3851 9276
rect 3851 9220 3855 9276
rect 3791 9216 3855 9220
rect 8749 9276 8813 9280
rect 8749 9220 8753 9276
rect 8753 9220 8809 9276
rect 8809 9220 8813 9276
rect 8749 9216 8813 9220
rect 8829 9276 8893 9280
rect 8829 9220 8833 9276
rect 8833 9220 8889 9276
rect 8889 9220 8893 9276
rect 8829 9216 8893 9220
rect 8909 9276 8973 9280
rect 8909 9220 8913 9276
rect 8913 9220 8969 9276
rect 8969 9220 8973 9276
rect 8909 9216 8973 9220
rect 8989 9276 9053 9280
rect 8989 9220 8993 9276
rect 8993 9220 9049 9276
rect 9049 9220 9053 9276
rect 8989 9216 9053 9220
rect 13947 9276 14011 9280
rect 13947 9220 13951 9276
rect 13951 9220 14007 9276
rect 14007 9220 14011 9276
rect 13947 9216 14011 9220
rect 14027 9276 14091 9280
rect 14027 9220 14031 9276
rect 14031 9220 14087 9276
rect 14087 9220 14091 9276
rect 14027 9216 14091 9220
rect 14107 9276 14171 9280
rect 14107 9220 14111 9276
rect 14111 9220 14167 9276
rect 14167 9220 14171 9276
rect 14107 9216 14171 9220
rect 14187 9276 14251 9280
rect 14187 9220 14191 9276
rect 14191 9220 14247 9276
rect 14247 9220 14251 9276
rect 14187 9216 14251 9220
rect 19145 9276 19209 9280
rect 19145 9220 19149 9276
rect 19149 9220 19205 9276
rect 19205 9220 19209 9276
rect 19145 9216 19209 9220
rect 19225 9276 19289 9280
rect 19225 9220 19229 9276
rect 19229 9220 19285 9276
rect 19285 9220 19289 9276
rect 19225 9216 19289 9220
rect 19305 9276 19369 9280
rect 19305 9220 19309 9276
rect 19309 9220 19365 9276
rect 19365 9220 19369 9276
rect 19305 9216 19369 9220
rect 19385 9276 19449 9280
rect 19385 9220 19389 9276
rect 19389 9220 19445 9276
rect 19445 9220 19449 9276
rect 19385 9216 19449 9220
rect 6150 8732 6214 8736
rect 6150 8676 6154 8732
rect 6154 8676 6210 8732
rect 6210 8676 6214 8732
rect 6150 8672 6214 8676
rect 6230 8732 6294 8736
rect 6230 8676 6234 8732
rect 6234 8676 6290 8732
rect 6290 8676 6294 8732
rect 6230 8672 6294 8676
rect 6310 8732 6374 8736
rect 6310 8676 6314 8732
rect 6314 8676 6370 8732
rect 6370 8676 6374 8732
rect 6310 8672 6374 8676
rect 6390 8732 6454 8736
rect 6390 8676 6394 8732
rect 6394 8676 6450 8732
rect 6450 8676 6454 8732
rect 6390 8672 6454 8676
rect 11348 8732 11412 8736
rect 11348 8676 11352 8732
rect 11352 8676 11408 8732
rect 11408 8676 11412 8732
rect 11348 8672 11412 8676
rect 11428 8732 11492 8736
rect 11428 8676 11432 8732
rect 11432 8676 11488 8732
rect 11488 8676 11492 8732
rect 11428 8672 11492 8676
rect 11508 8732 11572 8736
rect 11508 8676 11512 8732
rect 11512 8676 11568 8732
rect 11568 8676 11572 8732
rect 11508 8672 11572 8676
rect 11588 8732 11652 8736
rect 11588 8676 11592 8732
rect 11592 8676 11648 8732
rect 11648 8676 11652 8732
rect 11588 8672 11652 8676
rect 16546 8732 16610 8736
rect 16546 8676 16550 8732
rect 16550 8676 16606 8732
rect 16606 8676 16610 8732
rect 16546 8672 16610 8676
rect 16626 8732 16690 8736
rect 16626 8676 16630 8732
rect 16630 8676 16686 8732
rect 16686 8676 16690 8732
rect 16626 8672 16690 8676
rect 16706 8732 16770 8736
rect 16706 8676 16710 8732
rect 16710 8676 16766 8732
rect 16766 8676 16770 8732
rect 16706 8672 16770 8676
rect 16786 8732 16850 8736
rect 16786 8676 16790 8732
rect 16790 8676 16846 8732
rect 16846 8676 16850 8732
rect 16786 8672 16850 8676
rect 21744 8732 21808 8736
rect 21744 8676 21748 8732
rect 21748 8676 21804 8732
rect 21804 8676 21808 8732
rect 21744 8672 21808 8676
rect 21824 8732 21888 8736
rect 21824 8676 21828 8732
rect 21828 8676 21884 8732
rect 21884 8676 21888 8732
rect 21824 8672 21888 8676
rect 21904 8732 21968 8736
rect 21904 8676 21908 8732
rect 21908 8676 21964 8732
rect 21964 8676 21968 8732
rect 21904 8672 21968 8676
rect 21984 8732 22048 8736
rect 21984 8676 21988 8732
rect 21988 8676 22044 8732
rect 22044 8676 22048 8732
rect 21984 8672 22048 8676
rect 3551 8188 3615 8192
rect 3551 8132 3555 8188
rect 3555 8132 3611 8188
rect 3611 8132 3615 8188
rect 3551 8128 3615 8132
rect 3631 8188 3695 8192
rect 3631 8132 3635 8188
rect 3635 8132 3691 8188
rect 3691 8132 3695 8188
rect 3631 8128 3695 8132
rect 3711 8188 3775 8192
rect 3711 8132 3715 8188
rect 3715 8132 3771 8188
rect 3771 8132 3775 8188
rect 3711 8128 3775 8132
rect 3791 8188 3855 8192
rect 3791 8132 3795 8188
rect 3795 8132 3851 8188
rect 3851 8132 3855 8188
rect 3791 8128 3855 8132
rect 8749 8188 8813 8192
rect 8749 8132 8753 8188
rect 8753 8132 8809 8188
rect 8809 8132 8813 8188
rect 8749 8128 8813 8132
rect 8829 8188 8893 8192
rect 8829 8132 8833 8188
rect 8833 8132 8889 8188
rect 8889 8132 8893 8188
rect 8829 8128 8893 8132
rect 8909 8188 8973 8192
rect 8909 8132 8913 8188
rect 8913 8132 8969 8188
rect 8969 8132 8973 8188
rect 8909 8128 8973 8132
rect 8989 8188 9053 8192
rect 8989 8132 8993 8188
rect 8993 8132 9049 8188
rect 9049 8132 9053 8188
rect 8989 8128 9053 8132
rect 13947 8188 14011 8192
rect 13947 8132 13951 8188
rect 13951 8132 14007 8188
rect 14007 8132 14011 8188
rect 13947 8128 14011 8132
rect 14027 8188 14091 8192
rect 14027 8132 14031 8188
rect 14031 8132 14087 8188
rect 14087 8132 14091 8188
rect 14027 8128 14091 8132
rect 14107 8188 14171 8192
rect 14107 8132 14111 8188
rect 14111 8132 14167 8188
rect 14167 8132 14171 8188
rect 14107 8128 14171 8132
rect 14187 8188 14251 8192
rect 14187 8132 14191 8188
rect 14191 8132 14247 8188
rect 14247 8132 14251 8188
rect 14187 8128 14251 8132
rect 19145 8188 19209 8192
rect 19145 8132 19149 8188
rect 19149 8132 19205 8188
rect 19205 8132 19209 8188
rect 19145 8128 19209 8132
rect 19225 8188 19289 8192
rect 19225 8132 19229 8188
rect 19229 8132 19285 8188
rect 19285 8132 19289 8188
rect 19225 8128 19289 8132
rect 19305 8188 19369 8192
rect 19305 8132 19309 8188
rect 19309 8132 19365 8188
rect 19365 8132 19369 8188
rect 19305 8128 19369 8132
rect 19385 8188 19449 8192
rect 19385 8132 19389 8188
rect 19389 8132 19445 8188
rect 19445 8132 19449 8188
rect 19385 8128 19449 8132
rect 8340 7652 8404 7716
rect 6150 7644 6214 7648
rect 6150 7588 6154 7644
rect 6154 7588 6210 7644
rect 6210 7588 6214 7644
rect 6150 7584 6214 7588
rect 6230 7644 6294 7648
rect 6230 7588 6234 7644
rect 6234 7588 6290 7644
rect 6290 7588 6294 7644
rect 6230 7584 6294 7588
rect 6310 7644 6374 7648
rect 6310 7588 6314 7644
rect 6314 7588 6370 7644
rect 6370 7588 6374 7644
rect 6310 7584 6374 7588
rect 6390 7644 6454 7648
rect 6390 7588 6394 7644
rect 6394 7588 6450 7644
rect 6450 7588 6454 7644
rect 6390 7584 6454 7588
rect 11348 7644 11412 7648
rect 11348 7588 11352 7644
rect 11352 7588 11408 7644
rect 11408 7588 11412 7644
rect 11348 7584 11412 7588
rect 11428 7644 11492 7648
rect 11428 7588 11432 7644
rect 11432 7588 11488 7644
rect 11488 7588 11492 7644
rect 11428 7584 11492 7588
rect 11508 7644 11572 7648
rect 11508 7588 11512 7644
rect 11512 7588 11568 7644
rect 11568 7588 11572 7644
rect 11508 7584 11572 7588
rect 11588 7644 11652 7648
rect 11588 7588 11592 7644
rect 11592 7588 11648 7644
rect 11648 7588 11652 7644
rect 11588 7584 11652 7588
rect 16546 7644 16610 7648
rect 16546 7588 16550 7644
rect 16550 7588 16606 7644
rect 16606 7588 16610 7644
rect 16546 7584 16610 7588
rect 16626 7644 16690 7648
rect 16626 7588 16630 7644
rect 16630 7588 16686 7644
rect 16686 7588 16690 7644
rect 16626 7584 16690 7588
rect 16706 7644 16770 7648
rect 16706 7588 16710 7644
rect 16710 7588 16766 7644
rect 16766 7588 16770 7644
rect 16706 7584 16770 7588
rect 16786 7644 16850 7648
rect 16786 7588 16790 7644
rect 16790 7588 16846 7644
rect 16846 7588 16850 7644
rect 16786 7584 16850 7588
rect 21744 7644 21808 7648
rect 21744 7588 21748 7644
rect 21748 7588 21804 7644
rect 21804 7588 21808 7644
rect 21744 7584 21808 7588
rect 21824 7644 21888 7648
rect 21824 7588 21828 7644
rect 21828 7588 21884 7644
rect 21884 7588 21888 7644
rect 21824 7584 21888 7588
rect 21904 7644 21968 7648
rect 21904 7588 21908 7644
rect 21908 7588 21964 7644
rect 21964 7588 21968 7644
rect 21904 7584 21968 7588
rect 21984 7644 22048 7648
rect 21984 7588 21988 7644
rect 21988 7588 22044 7644
rect 22044 7588 22048 7644
rect 21984 7584 22048 7588
rect 6868 7304 6932 7308
rect 6868 7248 6918 7304
rect 6918 7248 6932 7304
rect 6868 7244 6932 7248
rect 3551 7100 3615 7104
rect 3551 7044 3555 7100
rect 3555 7044 3611 7100
rect 3611 7044 3615 7100
rect 3551 7040 3615 7044
rect 3631 7100 3695 7104
rect 3631 7044 3635 7100
rect 3635 7044 3691 7100
rect 3691 7044 3695 7100
rect 3631 7040 3695 7044
rect 3711 7100 3775 7104
rect 3711 7044 3715 7100
rect 3715 7044 3771 7100
rect 3771 7044 3775 7100
rect 3711 7040 3775 7044
rect 3791 7100 3855 7104
rect 3791 7044 3795 7100
rect 3795 7044 3851 7100
rect 3851 7044 3855 7100
rect 3791 7040 3855 7044
rect 8749 7100 8813 7104
rect 8749 7044 8753 7100
rect 8753 7044 8809 7100
rect 8809 7044 8813 7100
rect 8749 7040 8813 7044
rect 8829 7100 8893 7104
rect 8829 7044 8833 7100
rect 8833 7044 8889 7100
rect 8889 7044 8893 7100
rect 8829 7040 8893 7044
rect 8909 7100 8973 7104
rect 8909 7044 8913 7100
rect 8913 7044 8969 7100
rect 8969 7044 8973 7100
rect 8909 7040 8973 7044
rect 8989 7100 9053 7104
rect 8989 7044 8993 7100
rect 8993 7044 9049 7100
rect 9049 7044 9053 7100
rect 8989 7040 9053 7044
rect 13947 7100 14011 7104
rect 13947 7044 13951 7100
rect 13951 7044 14007 7100
rect 14007 7044 14011 7100
rect 13947 7040 14011 7044
rect 14027 7100 14091 7104
rect 14027 7044 14031 7100
rect 14031 7044 14087 7100
rect 14087 7044 14091 7100
rect 14027 7040 14091 7044
rect 14107 7100 14171 7104
rect 14107 7044 14111 7100
rect 14111 7044 14167 7100
rect 14167 7044 14171 7100
rect 14107 7040 14171 7044
rect 14187 7100 14251 7104
rect 14187 7044 14191 7100
rect 14191 7044 14247 7100
rect 14247 7044 14251 7100
rect 14187 7040 14251 7044
rect 6684 6836 6748 6900
rect 19145 7100 19209 7104
rect 19145 7044 19149 7100
rect 19149 7044 19205 7100
rect 19205 7044 19209 7100
rect 19145 7040 19209 7044
rect 19225 7100 19289 7104
rect 19225 7044 19229 7100
rect 19229 7044 19285 7100
rect 19285 7044 19289 7100
rect 19225 7040 19289 7044
rect 19305 7100 19369 7104
rect 19305 7044 19309 7100
rect 19309 7044 19365 7100
rect 19365 7044 19369 7100
rect 19305 7040 19369 7044
rect 19385 7100 19449 7104
rect 19385 7044 19389 7100
rect 19389 7044 19445 7100
rect 19445 7044 19449 7100
rect 19385 7040 19449 7044
rect 5764 6760 5828 6764
rect 5764 6704 5814 6760
rect 5814 6704 5828 6760
rect 5764 6700 5828 6704
rect 8524 6760 8588 6764
rect 8524 6704 8574 6760
rect 8574 6704 8588 6760
rect 8524 6700 8588 6704
rect 12020 6700 12084 6764
rect 6150 6556 6214 6560
rect 6150 6500 6154 6556
rect 6154 6500 6210 6556
rect 6210 6500 6214 6556
rect 6150 6496 6214 6500
rect 6230 6556 6294 6560
rect 6230 6500 6234 6556
rect 6234 6500 6290 6556
rect 6290 6500 6294 6556
rect 6230 6496 6294 6500
rect 6310 6556 6374 6560
rect 6310 6500 6314 6556
rect 6314 6500 6370 6556
rect 6370 6500 6374 6556
rect 6310 6496 6374 6500
rect 6390 6556 6454 6560
rect 6390 6500 6394 6556
rect 6394 6500 6450 6556
rect 6450 6500 6454 6556
rect 6390 6496 6454 6500
rect 11348 6556 11412 6560
rect 11348 6500 11352 6556
rect 11352 6500 11408 6556
rect 11408 6500 11412 6556
rect 11348 6496 11412 6500
rect 11428 6556 11492 6560
rect 11428 6500 11432 6556
rect 11432 6500 11488 6556
rect 11488 6500 11492 6556
rect 11428 6496 11492 6500
rect 11508 6556 11572 6560
rect 11508 6500 11512 6556
rect 11512 6500 11568 6556
rect 11568 6500 11572 6556
rect 11508 6496 11572 6500
rect 11588 6556 11652 6560
rect 11588 6500 11592 6556
rect 11592 6500 11648 6556
rect 11648 6500 11652 6556
rect 11588 6496 11652 6500
rect 8524 6428 8588 6492
rect 8156 6292 8220 6356
rect 16546 6556 16610 6560
rect 16546 6500 16550 6556
rect 16550 6500 16606 6556
rect 16606 6500 16610 6556
rect 16546 6496 16610 6500
rect 16626 6556 16690 6560
rect 16626 6500 16630 6556
rect 16630 6500 16686 6556
rect 16686 6500 16690 6556
rect 16626 6496 16690 6500
rect 16706 6556 16770 6560
rect 16706 6500 16710 6556
rect 16710 6500 16766 6556
rect 16766 6500 16770 6556
rect 16706 6496 16770 6500
rect 16786 6556 16850 6560
rect 16786 6500 16790 6556
rect 16790 6500 16846 6556
rect 16846 6500 16850 6556
rect 16786 6496 16850 6500
rect 21744 6556 21808 6560
rect 21744 6500 21748 6556
rect 21748 6500 21804 6556
rect 21804 6500 21808 6556
rect 21744 6496 21808 6500
rect 21824 6556 21888 6560
rect 21824 6500 21828 6556
rect 21828 6500 21884 6556
rect 21884 6500 21888 6556
rect 21824 6496 21888 6500
rect 21904 6556 21968 6560
rect 21904 6500 21908 6556
rect 21908 6500 21964 6556
rect 21964 6500 21968 6556
rect 21904 6496 21968 6500
rect 21984 6556 22048 6560
rect 21984 6500 21988 6556
rect 21988 6500 22044 6556
rect 22044 6500 22048 6556
rect 21984 6496 22048 6500
rect 9444 6020 9508 6084
rect 3551 6012 3615 6016
rect 3551 5956 3555 6012
rect 3555 5956 3611 6012
rect 3611 5956 3615 6012
rect 3551 5952 3615 5956
rect 3631 6012 3695 6016
rect 3631 5956 3635 6012
rect 3635 5956 3691 6012
rect 3691 5956 3695 6012
rect 3631 5952 3695 5956
rect 3711 6012 3775 6016
rect 3711 5956 3715 6012
rect 3715 5956 3771 6012
rect 3771 5956 3775 6012
rect 3711 5952 3775 5956
rect 3791 6012 3855 6016
rect 3791 5956 3795 6012
rect 3795 5956 3851 6012
rect 3851 5956 3855 6012
rect 3791 5952 3855 5956
rect 8749 6012 8813 6016
rect 8749 5956 8753 6012
rect 8753 5956 8809 6012
rect 8809 5956 8813 6012
rect 8749 5952 8813 5956
rect 8829 6012 8893 6016
rect 8829 5956 8833 6012
rect 8833 5956 8889 6012
rect 8889 5956 8893 6012
rect 8829 5952 8893 5956
rect 8909 6012 8973 6016
rect 8909 5956 8913 6012
rect 8913 5956 8969 6012
rect 8969 5956 8973 6012
rect 8909 5952 8973 5956
rect 8989 6012 9053 6016
rect 8989 5956 8993 6012
rect 8993 5956 9049 6012
rect 9049 5956 9053 6012
rect 8989 5952 9053 5956
rect 13947 6012 14011 6016
rect 13947 5956 13951 6012
rect 13951 5956 14007 6012
rect 14007 5956 14011 6012
rect 13947 5952 14011 5956
rect 14027 6012 14091 6016
rect 14027 5956 14031 6012
rect 14031 5956 14087 6012
rect 14087 5956 14091 6012
rect 14027 5952 14091 5956
rect 14107 6012 14171 6016
rect 14107 5956 14111 6012
rect 14111 5956 14167 6012
rect 14167 5956 14171 6012
rect 14107 5952 14171 5956
rect 14187 6012 14251 6016
rect 14187 5956 14191 6012
rect 14191 5956 14247 6012
rect 14247 5956 14251 6012
rect 14187 5952 14251 5956
rect 19145 6012 19209 6016
rect 19145 5956 19149 6012
rect 19149 5956 19205 6012
rect 19205 5956 19209 6012
rect 19145 5952 19209 5956
rect 19225 6012 19289 6016
rect 19225 5956 19229 6012
rect 19229 5956 19285 6012
rect 19285 5956 19289 6012
rect 19225 5952 19289 5956
rect 19305 6012 19369 6016
rect 19305 5956 19309 6012
rect 19309 5956 19365 6012
rect 19365 5956 19369 6012
rect 19305 5952 19369 5956
rect 19385 6012 19449 6016
rect 19385 5956 19389 6012
rect 19389 5956 19445 6012
rect 19445 5956 19449 6012
rect 19385 5952 19449 5956
rect 7788 5944 7852 5948
rect 7788 5888 7802 5944
rect 7802 5888 7852 5944
rect 7788 5884 7852 5888
rect 9260 5944 9324 5948
rect 9260 5888 9274 5944
rect 9274 5888 9324 5944
rect 9260 5884 9324 5888
rect 6150 5468 6214 5472
rect 6150 5412 6154 5468
rect 6154 5412 6210 5468
rect 6210 5412 6214 5468
rect 6150 5408 6214 5412
rect 6230 5468 6294 5472
rect 6230 5412 6234 5468
rect 6234 5412 6290 5468
rect 6290 5412 6294 5468
rect 6230 5408 6294 5412
rect 6310 5468 6374 5472
rect 6310 5412 6314 5468
rect 6314 5412 6370 5468
rect 6370 5412 6374 5468
rect 6310 5408 6374 5412
rect 6390 5468 6454 5472
rect 6390 5412 6394 5468
rect 6394 5412 6450 5468
rect 6450 5412 6454 5468
rect 6390 5408 6454 5412
rect 11348 5468 11412 5472
rect 11348 5412 11352 5468
rect 11352 5412 11408 5468
rect 11408 5412 11412 5468
rect 11348 5408 11412 5412
rect 11428 5468 11492 5472
rect 11428 5412 11432 5468
rect 11432 5412 11488 5468
rect 11488 5412 11492 5468
rect 11428 5408 11492 5412
rect 11508 5468 11572 5472
rect 11508 5412 11512 5468
rect 11512 5412 11568 5468
rect 11568 5412 11572 5468
rect 11508 5408 11572 5412
rect 11588 5468 11652 5472
rect 11588 5412 11592 5468
rect 11592 5412 11648 5468
rect 11648 5412 11652 5468
rect 11588 5408 11652 5412
rect 16546 5468 16610 5472
rect 16546 5412 16550 5468
rect 16550 5412 16606 5468
rect 16606 5412 16610 5468
rect 16546 5408 16610 5412
rect 16626 5468 16690 5472
rect 16626 5412 16630 5468
rect 16630 5412 16686 5468
rect 16686 5412 16690 5468
rect 16626 5408 16690 5412
rect 16706 5468 16770 5472
rect 16706 5412 16710 5468
rect 16710 5412 16766 5468
rect 16766 5412 16770 5468
rect 16706 5408 16770 5412
rect 16786 5468 16850 5472
rect 16786 5412 16790 5468
rect 16790 5412 16846 5468
rect 16846 5412 16850 5468
rect 16786 5408 16850 5412
rect 21744 5468 21808 5472
rect 21744 5412 21748 5468
rect 21748 5412 21804 5468
rect 21804 5412 21808 5468
rect 21744 5408 21808 5412
rect 21824 5468 21888 5472
rect 21824 5412 21828 5468
rect 21828 5412 21884 5468
rect 21884 5412 21888 5468
rect 21824 5408 21888 5412
rect 21904 5468 21968 5472
rect 21904 5412 21908 5468
rect 21908 5412 21964 5468
rect 21964 5412 21968 5468
rect 21904 5408 21968 5412
rect 21984 5468 22048 5472
rect 21984 5412 21988 5468
rect 21988 5412 22044 5468
rect 22044 5412 22048 5468
rect 21984 5408 22048 5412
rect 3551 4924 3615 4928
rect 3551 4868 3555 4924
rect 3555 4868 3611 4924
rect 3611 4868 3615 4924
rect 3551 4864 3615 4868
rect 3631 4924 3695 4928
rect 3631 4868 3635 4924
rect 3635 4868 3691 4924
rect 3691 4868 3695 4924
rect 3631 4864 3695 4868
rect 3711 4924 3775 4928
rect 3711 4868 3715 4924
rect 3715 4868 3771 4924
rect 3771 4868 3775 4924
rect 3711 4864 3775 4868
rect 3791 4924 3855 4928
rect 3791 4868 3795 4924
rect 3795 4868 3851 4924
rect 3851 4868 3855 4924
rect 3791 4864 3855 4868
rect 8749 4924 8813 4928
rect 8749 4868 8753 4924
rect 8753 4868 8809 4924
rect 8809 4868 8813 4924
rect 8749 4864 8813 4868
rect 8829 4924 8893 4928
rect 8829 4868 8833 4924
rect 8833 4868 8889 4924
rect 8889 4868 8893 4924
rect 8829 4864 8893 4868
rect 8909 4924 8973 4928
rect 8909 4868 8913 4924
rect 8913 4868 8969 4924
rect 8969 4868 8973 4924
rect 8909 4864 8973 4868
rect 8989 4924 9053 4928
rect 8989 4868 8993 4924
rect 8993 4868 9049 4924
rect 9049 4868 9053 4924
rect 8989 4864 9053 4868
rect 10180 4932 10244 4996
rect 13947 4924 14011 4928
rect 13947 4868 13951 4924
rect 13951 4868 14007 4924
rect 14007 4868 14011 4924
rect 13947 4864 14011 4868
rect 14027 4924 14091 4928
rect 14027 4868 14031 4924
rect 14031 4868 14087 4924
rect 14087 4868 14091 4924
rect 14027 4864 14091 4868
rect 14107 4924 14171 4928
rect 14107 4868 14111 4924
rect 14111 4868 14167 4924
rect 14167 4868 14171 4924
rect 14107 4864 14171 4868
rect 14187 4924 14251 4928
rect 14187 4868 14191 4924
rect 14191 4868 14247 4924
rect 14247 4868 14251 4924
rect 14187 4864 14251 4868
rect 19145 4924 19209 4928
rect 19145 4868 19149 4924
rect 19149 4868 19205 4924
rect 19205 4868 19209 4924
rect 19145 4864 19209 4868
rect 19225 4924 19289 4928
rect 19225 4868 19229 4924
rect 19229 4868 19285 4924
rect 19285 4868 19289 4924
rect 19225 4864 19289 4868
rect 19305 4924 19369 4928
rect 19305 4868 19309 4924
rect 19309 4868 19365 4924
rect 19365 4868 19369 4924
rect 19305 4864 19369 4868
rect 19385 4924 19449 4928
rect 19385 4868 19389 4924
rect 19389 4868 19445 4924
rect 19445 4868 19449 4924
rect 19385 4864 19449 4868
rect 9812 4660 9876 4724
rect 6150 4380 6214 4384
rect 6150 4324 6154 4380
rect 6154 4324 6210 4380
rect 6210 4324 6214 4380
rect 6150 4320 6214 4324
rect 6230 4380 6294 4384
rect 6230 4324 6234 4380
rect 6234 4324 6290 4380
rect 6290 4324 6294 4380
rect 6230 4320 6294 4324
rect 6310 4380 6374 4384
rect 6310 4324 6314 4380
rect 6314 4324 6370 4380
rect 6370 4324 6374 4380
rect 6310 4320 6374 4324
rect 6390 4380 6454 4384
rect 6390 4324 6394 4380
rect 6394 4324 6450 4380
rect 6450 4324 6454 4380
rect 6390 4320 6454 4324
rect 11348 4380 11412 4384
rect 11348 4324 11352 4380
rect 11352 4324 11408 4380
rect 11408 4324 11412 4380
rect 11348 4320 11412 4324
rect 11428 4380 11492 4384
rect 11428 4324 11432 4380
rect 11432 4324 11488 4380
rect 11488 4324 11492 4380
rect 11428 4320 11492 4324
rect 11508 4380 11572 4384
rect 11508 4324 11512 4380
rect 11512 4324 11568 4380
rect 11568 4324 11572 4380
rect 11508 4320 11572 4324
rect 11588 4380 11652 4384
rect 11588 4324 11592 4380
rect 11592 4324 11648 4380
rect 11648 4324 11652 4380
rect 11588 4320 11652 4324
rect 16546 4380 16610 4384
rect 16546 4324 16550 4380
rect 16550 4324 16606 4380
rect 16606 4324 16610 4380
rect 16546 4320 16610 4324
rect 16626 4380 16690 4384
rect 16626 4324 16630 4380
rect 16630 4324 16686 4380
rect 16686 4324 16690 4380
rect 16626 4320 16690 4324
rect 16706 4380 16770 4384
rect 16706 4324 16710 4380
rect 16710 4324 16766 4380
rect 16766 4324 16770 4380
rect 16706 4320 16770 4324
rect 16786 4380 16850 4384
rect 16786 4324 16790 4380
rect 16790 4324 16846 4380
rect 16846 4324 16850 4380
rect 16786 4320 16850 4324
rect 21744 4380 21808 4384
rect 21744 4324 21748 4380
rect 21748 4324 21804 4380
rect 21804 4324 21808 4380
rect 21744 4320 21808 4324
rect 21824 4380 21888 4384
rect 21824 4324 21828 4380
rect 21828 4324 21884 4380
rect 21884 4324 21888 4380
rect 21824 4320 21888 4324
rect 21904 4380 21968 4384
rect 21904 4324 21908 4380
rect 21908 4324 21964 4380
rect 21964 4324 21968 4380
rect 21904 4320 21968 4324
rect 21984 4380 22048 4384
rect 21984 4324 21988 4380
rect 21988 4324 22044 4380
rect 22044 4324 22048 4380
rect 21984 4320 22048 4324
rect 9444 3844 9508 3908
rect 3551 3836 3615 3840
rect 3551 3780 3555 3836
rect 3555 3780 3611 3836
rect 3611 3780 3615 3836
rect 3551 3776 3615 3780
rect 3631 3836 3695 3840
rect 3631 3780 3635 3836
rect 3635 3780 3691 3836
rect 3691 3780 3695 3836
rect 3631 3776 3695 3780
rect 3711 3836 3775 3840
rect 3711 3780 3715 3836
rect 3715 3780 3771 3836
rect 3771 3780 3775 3836
rect 3711 3776 3775 3780
rect 3791 3836 3855 3840
rect 3791 3780 3795 3836
rect 3795 3780 3851 3836
rect 3851 3780 3855 3836
rect 3791 3776 3855 3780
rect 8749 3836 8813 3840
rect 8749 3780 8753 3836
rect 8753 3780 8809 3836
rect 8809 3780 8813 3836
rect 8749 3776 8813 3780
rect 8829 3836 8893 3840
rect 8829 3780 8833 3836
rect 8833 3780 8889 3836
rect 8889 3780 8893 3836
rect 8829 3776 8893 3780
rect 8909 3836 8973 3840
rect 8909 3780 8913 3836
rect 8913 3780 8969 3836
rect 8969 3780 8973 3836
rect 8909 3776 8973 3780
rect 8989 3836 9053 3840
rect 8989 3780 8993 3836
rect 8993 3780 9049 3836
rect 9049 3780 9053 3836
rect 8989 3776 9053 3780
rect 13947 3836 14011 3840
rect 13947 3780 13951 3836
rect 13951 3780 14007 3836
rect 14007 3780 14011 3836
rect 13947 3776 14011 3780
rect 14027 3836 14091 3840
rect 14027 3780 14031 3836
rect 14031 3780 14087 3836
rect 14087 3780 14091 3836
rect 14027 3776 14091 3780
rect 14107 3836 14171 3840
rect 14107 3780 14111 3836
rect 14111 3780 14167 3836
rect 14167 3780 14171 3836
rect 14107 3776 14171 3780
rect 14187 3836 14251 3840
rect 14187 3780 14191 3836
rect 14191 3780 14247 3836
rect 14247 3780 14251 3836
rect 14187 3776 14251 3780
rect 19145 3836 19209 3840
rect 19145 3780 19149 3836
rect 19149 3780 19205 3836
rect 19205 3780 19209 3836
rect 19145 3776 19209 3780
rect 19225 3836 19289 3840
rect 19225 3780 19229 3836
rect 19229 3780 19285 3836
rect 19285 3780 19289 3836
rect 19225 3776 19289 3780
rect 19305 3836 19369 3840
rect 19305 3780 19309 3836
rect 19309 3780 19365 3836
rect 19365 3780 19369 3836
rect 19305 3776 19369 3780
rect 19385 3836 19449 3840
rect 19385 3780 19389 3836
rect 19389 3780 19445 3836
rect 19445 3780 19449 3836
rect 19385 3776 19449 3780
rect 9812 3572 9876 3636
rect 5948 3436 6012 3500
rect 8340 3300 8404 3364
rect 6150 3292 6214 3296
rect 6150 3236 6154 3292
rect 6154 3236 6210 3292
rect 6210 3236 6214 3292
rect 6150 3232 6214 3236
rect 6230 3292 6294 3296
rect 6230 3236 6234 3292
rect 6234 3236 6290 3292
rect 6290 3236 6294 3292
rect 6230 3232 6294 3236
rect 6310 3292 6374 3296
rect 6310 3236 6314 3292
rect 6314 3236 6370 3292
rect 6370 3236 6374 3292
rect 6310 3232 6374 3236
rect 6390 3292 6454 3296
rect 6390 3236 6394 3292
rect 6394 3236 6450 3292
rect 6450 3236 6454 3292
rect 6390 3232 6454 3236
rect 11348 3292 11412 3296
rect 11348 3236 11352 3292
rect 11352 3236 11408 3292
rect 11408 3236 11412 3292
rect 11348 3232 11412 3236
rect 11428 3292 11492 3296
rect 11428 3236 11432 3292
rect 11432 3236 11488 3292
rect 11488 3236 11492 3292
rect 11428 3232 11492 3236
rect 11508 3292 11572 3296
rect 11508 3236 11512 3292
rect 11512 3236 11568 3292
rect 11568 3236 11572 3292
rect 11508 3232 11572 3236
rect 11588 3292 11652 3296
rect 11588 3236 11592 3292
rect 11592 3236 11648 3292
rect 11648 3236 11652 3292
rect 11588 3232 11652 3236
rect 16546 3292 16610 3296
rect 16546 3236 16550 3292
rect 16550 3236 16606 3292
rect 16606 3236 16610 3292
rect 16546 3232 16610 3236
rect 16626 3292 16690 3296
rect 16626 3236 16630 3292
rect 16630 3236 16686 3292
rect 16686 3236 16690 3292
rect 16626 3232 16690 3236
rect 16706 3292 16770 3296
rect 16706 3236 16710 3292
rect 16710 3236 16766 3292
rect 16766 3236 16770 3292
rect 16706 3232 16770 3236
rect 16786 3292 16850 3296
rect 16786 3236 16790 3292
rect 16790 3236 16846 3292
rect 16846 3236 16850 3292
rect 16786 3232 16850 3236
rect 21744 3292 21808 3296
rect 21744 3236 21748 3292
rect 21748 3236 21804 3292
rect 21804 3236 21808 3292
rect 21744 3232 21808 3236
rect 21824 3292 21888 3296
rect 21824 3236 21828 3292
rect 21828 3236 21884 3292
rect 21884 3236 21888 3292
rect 21824 3232 21888 3236
rect 21904 3292 21968 3296
rect 21904 3236 21908 3292
rect 21908 3236 21964 3292
rect 21964 3236 21968 3292
rect 21904 3232 21968 3236
rect 21984 3292 22048 3296
rect 21984 3236 21988 3292
rect 21988 3236 22044 3292
rect 22044 3236 22048 3292
rect 21984 3232 22048 3236
rect 5764 3164 5828 3228
rect 3551 2748 3615 2752
rect 3551 2692 3555 2748
rect 3555 2692 3611 2748
rect 3611 2692 3615 2748
rect 3551 2688 3615 2692
rect 3631 2748 3695 2752
rect 3631 2692 3635 2748
rect 3635 2692 3691 2748
rect 3691 2692 3695 2748
rect 3631 2688 3695 2692
rect 3711 2748 3775 2752
rect 3711 2692 3715 2748
rect 3715 2692 3771 2748
rect 3771 2692 3775 2748
rect 3711 2688 3775 2692
rect 3791 2748 3855 2752
rect 3791 2692 3795 2748
rect 3795 2692 3851 2748
rect 3851 2692 3855 2748
rect 3791 2688 3855 2692
rect 8749 2748 8813 2752
rect 8749 2692 8753 2748
rect 8753 2692 8809 2748
rect 8809 2692 8813 2748
rect 8749 2688 8813 2692
rect 8829 2748 8893 2752
rect 8829 2692 8833 2748
rect 8833 2692 8889 2748
rect 8889 2692 8893 2748
rect 8829 2688 8893 2692
rect 8909 2748 8973 2752
rect 8909 2692 8913 2748
rect 8913 2692 8969 2748
rect 8969 2692 8973 2748
rect 8909 2688 8973 2692
rect 8989 2748 9053 2752
rect 8989 2692 8993 2748
rect 8993 2692 9049 2748
rect 9049 2692 9053 2748
rect 8989 2688 9053 2692
rect 13947 2748 14011 2752
rect 13947 2692 13951 2748
rect 13951 2692 14007 2748
rect 14007 2692 14011 2748
rect 13947 2688 14011 2692
rect 14027 2748 14091 2752
rect 14027 2692 14031 2748
rect 14031 2692 14087 2748
rect 14087 2692 14091 2748
rect 14027 2688 14091 2692
rect 14107 2748 14171 2752
rect 14107 2692 14111 2748
rect 14111 2692 14167 2748
rect 14167 2692 14171 2748
rect 14107 2688 14171 2692
rect 14187 2748 14251 2752
rect 14187 2692 14191 2748
rect 14191 2692 14247 2748
rect 14247 2692 14251 2748
rect 14187 2688 14251 2692
rect 19145 2748 19209 2752
rect 19145 2692 19149 2748
rect 19149 2692 19205 2748
rect 19205 2692 19209 2748
rect 19145 2688 19209 2692
rect 19225 2748 19289 2752
rect 19225 2692 19229 2748
rect 19229 2692 19285 2748
rect 19285 2692 19289 2748
rect 19225 2688 19289 2692
rect 19305 2748 19369 2752
rect 19305 2692 19309 2748
rect 19309 2692 19365 2748
rect 19365 2692 19369 2748
rect 19305 2688 19369 2692
rect 19385 2748 19449 2752
rect 19385 2692 19389 2748
rect 19389 2692 19445 2748
rect 19445 2692 19449 2748
rect 19385 2688 19449 2692
rect 8524 2484 8588 2548
rect 6150 2204 6214 2208
rect 6150 2148 6154 2204
rect 6154 2148 6210 2204
rect 6210 2148 6214 2204
rect 6150 2144 6214 2148
rect 6230 2204 6294 2208
rect 6230 2148 6234 2204
rect 6234 2148 6290 2204
rect 6290 2148 6294 2204
rect 6230 2144 6294 2148
rect 6310 2204 6374 2208
rect 6310 2148 6314 2204
rect 6314 2148 6370 2204
rect 6370 2148 6374 2204
rect 6310 2144 6374 2148
rect 6390 2204 6454 2208
rect 6390 2148 6394 2204
rect 6394 2148 6450 2204
rect 6450 2148 6454 2204
rect 6390 2144 6454 2148
rect 11348 2204 11412 2208
rect 11348 2148 11352 2204
rect 11352 2148 11408 2204
rect 11408 2148 11412 2204
rect 11348 2144 11412 2148
rect 11428 2204 11492 2208
rect 11428 2148 11432 2204
rect 11432 2148 11488 2204
rect 11488 2148 11492 2204
rect 11428 2144 11492 2148
rect 11508 2204 11572 2208
rect 11508 2148 11512 2204
rect 11512 2148 11568 2204
rect 11568 2148 11572 2204
rect 11508 2144 11572 2148
rect 11588 2204 11652 2208
rect 11588 2148 11592 2204
rect 11592 2148 11648 2204
rect 11648 2148 11652 2204
rect 11588 2144 11652 2148
rect 16546 2204 16610 2208
rect 16546 2148 16550 2204
rect 16550 2148 16606 2204
rect 16606 2148 16610 2204
rect 16546 2144 16610 2148
rect 16626 2204 16690 2208
rect 16626 2148 16630 2204
rect 16630 2148 16686 2204
rect 16686 2148 16690 2204
rect 16626 2144 16690 2148
rect 16706 2204 16770 2208
rect 16706 2148 16710 2204
rect 16710 2148 16766 2204
rect 16766 2148 16770 2204
rect 16706 2144 16770 2148
rect 16786 2204 16850 2208
rect 16786 2148 16790 2204
rect 16790 2148 16846 2204
rect 16846 2148 16850 2204
rect 16786 2144 16850 2148
rect 21744 2204 21808 2208
rect 21744 2148 21748 2204
rect 21748 2148 21804 2204
rect 21804 2148 21808 2204
rect 21744 2144 21808 2148
rect 21824 2204 21888 2208
rect 21824 2148 21828 2204
rect 21828 2148 21884 2204
rect 21884 2148 21888 2204
rect 21824 2144 21888 2148
rect 21904 2204 21968 2208
rect 21904 2148 21908 2204
rect 21908 2148 21964 2204
rect 21964 2148 21968 2204
rect 21904 2144 21968 2148
rect 21984 2204 22048 2208
rect 21984 2148 21988 2204
rect 21988 2148 22044 2204
rect 22044 2148 22048 2204
rect 21984 2144 22048 2148
<< metal4 >>
rect 3543 20160 3863 20720
rect 3543 20096 3551 20160
rect 3615 20096 3631 20160
rect 3695 20096 3711 20160
rect 3775 20096 3791 20160
rect 3855 20096 3863 20160
rect 3543 19072 3863 20096
rect 3543 19008 3551 19072
rect 3615 19008 3631 19072
rect 3695 19008 3711 19072
rect 3775 19008 3791 19072
rect 3855 19008 3863 19072
rect 2819 18596 2885 18597
rect 2819 18532 2820 18596
rect 2884 18532 2885 18596
rect 2819 18531 2885 18532
rect 2822 13837 2882 18531
rect 3543 17984 3863 19008
rect 3543 17920 3551 17984
rect 3615 17920 3631 17984
rect 3695 17920 3711 17984
rect 3775 17920 3791 17984
rect 3855 17920 3863 17984
rect 3543 16896 3863 17920
rect 3543 16832 3551 16896
rect 3615 16832 3631 16896
rect 3695 16832 3711 16896
rect 3775 16832 3791 16896
rect 3855 16832 3863 16896
rect 3543 15808 3863 16832
rect 3543 15744 3551 15808
rect 3615 15744 3631 15808
rect 3695 15744 3711 15808
rect 3775 15744 3791 15808
rect 3855 15744 3863 15808
rect 3543 14720 3863 15744
rect 6142 20704 6462 20720
rect 6142 20640 6150 20704
rect 6214 20640 6230 20704
rect 6294 20640 6310 20704
rect 6374 20640 6390 20704
rect 6454 20640 6462 20704
rect 6142 19616 6462 20640
rect 6142 19552 6150 19616
rect 6214 19552 6230 19616
rect 6294 19552 6310 19616
rect 6374 19552 6390 19616
rect 6454 19552 6462 19616
rect 6142 18528 6462 19552
rect 6142 18464 6150 18528
rect 6214 18464 6230 18528
rect 6294 18464 6310 18528
rect 6374 18464 6390 18528
rect 6454 18464 6462 18528
rect 6142 17440 6462 18464
rect 8741 20160 9061 20720
rect 8741 20096 8749 20160
rect 8813 20096 8829 20160
rect 8893 20096 8909 20160
rect 8973 20096 8989 20160
rect 9053 20096 9061 20160
rect 8741 19072 9061 20096
rect 11340 20704 11660 20720
rect 11340 20640 11348 20704
rect 11412 20640 11428 20704
rect 11492 20640 11508 20704
rect 11572 20640 11588 20704
rect 11652 20640 11660 20704
rect 11099 19684 11165 19685
rect 11099 19620 11100 19684
rect 11164 19620 11165 19684
rect 11099 19619 11165 19620
rect 9443 19140 9509 19141
rect 9443 19076 9444 19140
rect 9508 19076 9509 19140
rect 9443 19075 9509 19076
rect 9811 19140 9877 19141
rect 9811 19076 9812 19140
rect 9876 19076 9877 19140
rect 9811 19075 9877 19076
rect 8741 19008 8749 19072
rect 8813 19008 8829 19072
rect 8893 19008 8909 19072
rect 8973 19008 8989 19072
rect 9053 19008 9061 19072
rect 6683 18052 6749 18053
rect 6683 17988 6684 18052
rect 6748 17988 6749 18052
rect 6683 17987 6749 17988
rect 8155 18052 8221 18053
rect 8155 17988 8156 18052
rect 8220 17988 8221 18052
rect 8155 17987 8221 17988
rect 6142 17376 6150 17440
rect 6214 17376 6230 17440
rect 6294 17376 6310 17440
rect 6374 17376 6390 17440
rect 6454 17376 6462 17440
rect 6142 16352 6462 17376
rect 6142 16288 6150 16352
rect 6214 16288 6230 16352
rect 6294 16288 6310 16352
rect 6374 16288 6390 16352
rect 6454 16288 6462 16352
rect 6142 15264 6462 16288
rect 6142 15200 6150 15264
rect 6214 15200 6230 15264
rect 6294 15200 6310 15264
rect 6374 15200 6390 15264
rect 6454 15200 6462 15264
rect 5579 14924 5645 14925
rect 5579 14860 5580 14924
rect 5644 14860 5645 14924
rect 5579 14859 5645 14860
rect 3543 14656 3551 14720
rect 3615 14656 3631 14720
rect 3695 14656 3711 14720
rect 3775 14656 3791 14720
rect 3855 14656 3863 14720
rect 2819 13836 2885 13837
rect 2819 13772 2820 13836
rect 2884 13772 2885 13836
rect 2819 13771 2885 13772
rect 3543 13632 3863 14656
rect 3543 13568 3551 13632
rect 3615 13568 3631 13632
rect 3695 13568 3711 13632
rect 3775 13568 3791 13632
rect 3855 13568 3863 13632
rect 3543 12544 3863 13568
rect 3543 12480 3551 12544
rect 3615 12480 3631 12544
rect 3695 12480 3711 12544
rect 3775 12480 3791 12544
rect 3855 12480 3863 12544
rect 3543 11456 3863 12480
rect 3543 11392 3551 11456
rect 3615 11392 3631 11456
rect 3695 11392 3711 11456
rect 3775 11392 3791 11456
rect 3855 11392 3863 11456
rect 3543 10368 3863 11392
rect 5582 11117 5642 14859
rect 6142 14176 6462 15200
rect 6142 14112 6150 14176
rect 6214 14112 6230 14176
rect 6294 14112 6310 14176
rect 6374 14112 6390 14176
rect 6454 14112 6462 14176
rect 5763 13700 5829 13701
rect 5763 13636 5764 13700
rect 5828 13636 5829 13700
rect 5763 13635 5829 13636
rect 5579 11116 5645 11117
rect 5579 11052 5580 11116
rect 5644 11052 5645 11116
rect 5579 11051 5645 11052
rect 3543 10304 3551 10368
rect 3615 10304 3631 10368
rect 3695 10304 3711 10368
rect 3775 10304 3791 10368
rect 3855 10304 3863 10368
rect 3543 9280 3863 10304
rect 3543 9216 3551 9280
rect 3615 9216 3631 9280
rect 3695 9216 3711 9280
rect 3775 9216 3791 9280
rect 3855 9216 3863 9280
rect 3543 8192 3863 9216
rect 3543 8128 3551 8192
rect 3615 8128 3631 8192
rect 3695 8128 3711 8192
rect 3775 8128 3791 8192
rect 3855 8128 3863 8192
rect 3543 7104 3863 8128
rect 3543 7040 3551 7104
rect 3615 7040 3631 7104
rect 3695 7040 3711 7104
rect 3775 7040 3791 7104
rect 3855 7040 3863 7104
rect 3543 6016 3863 7040
rect 5766 6765 5826 13635
rect 6142 13088 6462 14112
rect 6142 13024 6150 13088
rect 6214 13024 6230 13088
rect 6294 13024 6310 13088
rect 6374 13024 6390 13088
rect 6454 13024 6462 13088
rect 5947 12748 6013 12749
rect 5947 12684 5948 12748
rect 6012 12684 6013 12748
rect 5947 12683 6013 12684
rect 5763 6764 5829 6765
rect 5763 6700 5764 6764
rect 5828 6700 5829 6764
rect 5763 6699 5829 6700
rect 3543 5952 3551 6016
rect 3615 5952 3631 6016
rect 3695 5952 3711 6016
rect 3775 5952 3791 6016
rect 3855 5952 3863 6016
rect 3543 4928 3863 5952
rect 3543 4864 3551 4928
rect 3615 4864 3631 4928
rect 3695 4864 3711 4928
rect 3775 4864 3791 4928
rect 3855 4864 3863 4928
rect 3543 3840 3863 4864
rect 3543 3776 3551 3840
rect 3615 3776 3631 3840
rect 3695 3776 3711 3840
rect 3775 3776 3791 3840
rect 3855 3776 3863 3840
rect 3543 2752 3863 3776
rect 5766 3229 5826 6699
rect 5950 3501 6010 12683
rect 6142 12000 6462 13024
rect 6142 11936 6150 12000
rect 6214 11936 6230 12000
rect 6294 11936 6310 12000
rect 6374 11936 6390 12000
rect 6454 11936 6462 12000
rect 6142 10912 6462 11936
rect 6142 10848 6150 10912
rect 6214 10848 6230 10912
rect 6294 10848 6310 10912
rect 6374 10848 6390 10912
rect 6454 10848 6462 10912
rect 6142 9824 6462 10848
rect 6142 9760 6150 9824
rect 6214 9760 6230 9824
rect 6294 9760 6310 9824
rect 6374 9760 6390 9824
rect 6454 9760 6462 9824
rect 6142 8736 6462 9760
rect 6142 8672 6150 8736
rect 6214 8672 6230 8736
rect 6294 8672 6310 8736
rect 6374 8672 6390 8736
rect 6454 8672 6462 8736
rect 6142 7648 6462 8672
rect 6142 7584 6150 7648
rect 6214 7584 6230 7648
rect 6294 7584 6310 7648
rect 6374 7584 6390 7648
rect 6454 7584 6462 7648
rect 6142 6560 6462 7584
rect 6686 6901 6746 17987
rect 6867 16692 6933 16693
rect 6867 16628 6868 16692
rect 6932 16628 6933 16692
rect 6867 16627 6933 16628
rect 6870 7309 6930 16627
rect 7235 15876 7301 15877
rect 7235 15812 7236 15876
rect 7300 15812 7301 15876
rect 7235 15811 7301 15812
rect 7238 10437 7298 15811
rect 7787 14244 7853 14245
rect 7787 14180 7788 14244
rect 7852 14180 7853 14244
rect 7787 14179 7853 14180
rect 7235 10436 7301 10437
rect 7235 10372 7236 10436
rect 7300 10372 7301 10436
rect 7235 10371 7301 10372
rect 6867 7308 6933 7309
rect 6867 7244 6868 7308
rect 6932 7244 6933 7308
rect 6867 7243 6933 7244
rect 6683 6900 6749 6901
rect 6683 6836 6684 6900
rect 6748 6836 6749 6900
rect 6683 6835 6749 6836
rect 6142 6496 6150 6560
rect 6214 6496 6230 6560
rect 6294 6496 6310 6560
rect 6374 6496 6390 6560
rect 6454 6496 6462 6560
rect 6142 5472 6462 6496
rect 7790 5949 7850 14179
rect 8158 6357 8218 17987
rect 8741 17984 9061 19008
rect 9259 18460 9325 18461
rect 9259 18396 9260 18460
rect 9324 18396 9325 18460
rect 9259 18395 9325 18396
rect 8741 17920 8749 17984
rect 8813 17920 8829 17984
rect 8893 17920 8909 17984
rect 8973 17920 8989 17984
rect 9053 17920 9061 17984
rect 8741 16896 9061 17920
rect 8741 16832 8749 16896
rect 8813 16832 8829 16896
rect 8893 16832 8909 16896
rect 8973 16832 8989 16896
rect 9053 16832 9061 16896
rect 8741 15808 9061 16832
rect 8741 15744 8749 15808
rect 8813 15744 8829 15808
rect 8893 15744 8909 15808
rect 8973 15744 8989 15808
rect 9053 15744 9061 15808
rect 8741 14720 9061 15744
rect 8741 14656 8749 14720
rect 8813 14656 8829 14720
rect 8893 14656 8909 14720
rect 8973 14656 8989 14720
rect 9053 14656 9061 14720
rect 8741 13632 9061 14656
rect 8741 13568 8749 13632
rect 8813 13568 8829 13632
rect 8893 13568 8909 13632
rect 8973 13568 8989 13632
rect 9053 13568 9061 13632
rect 8741 12544 9061 13568
rect 8741 12480 8749 12544
rect 8813 12480 8829 12544
rect 8893 12480 8909 12544
rect 8973 12480 8989 12544
rect 9053 12480 9061 12544
rect 8523 11932 8589 11933
rect 8523 11868 8524 11932
rect 8588 11868 8589 11932
rect 8523 11867 8589 11868
rect 8339 7716 8405 7717
rect 8339 7652 8340 7716
rect 8404 7652 8405 7716
rect 8339 7651 8405 7652
rect 8155 6356 8221 6357
rect 8155 6292 8156 6356
rect 8220 6292 8221 6356
rect 8155 6291 8221 6292
rect 7787 5948 7853 5949
rect 7787 5884 7788 5948
rect 7852 5884 7853 5948
rect 7787 5883 7853 5884
rect 6142 5408 6150 5472
rect 6214 5408 6230 5472
rect 6294 5408 6310 5472
rect 6374 5408 6390 5472
rect 6454 5408 6462 5472
rect 6142 4384 6462 5408
rect 6142 4320 6150 4384
rect 6214 4320 6230 4384
rect 6294 4320 6310 4384
rect 6374 4320 6390 4384
rect 6454 4320 6462 4384
rect 5947 3500 6013 3501
rect 5947 3436 5948 3500
rect 6012 3436 6013 3500
rect 5947 3435 6013 3436
rect 6142 3296 6462 4320
rect 8342 3365 8402 7651
rect 8526 6765 8586 11867
rect 8741 11456 9061 12480
rect 8741 11392 8749 11456
rect 8813 11392 8829 11456
rect 8893 11392 8909 11456
rect 8973 11392 8989 11456
rect 9053 11392 9061 11456
rect 8741 10368 9061 11392
rect 8741 10304 8749 10368
rect 8813 10304 8829 10368
rect 8893 10304 8909 10368
rect 8973 10304 8989 10368
rect 9053 10304 9061 10368
rect 8741 9280 9061 10304
rect 8741 9216 8749 9280
rect 8813 9216 8829 9280
rect 8893 9216 8909 9280
rect 8973 9216 8989 9280
rect 9053 9216 9061 9280
rect 8741 8192 9061 9216
rect 8741 8128 8749 8192
rect 8813 8128 8829 8192
rect 8893 8128 8909 8192
rect 8973 8128 8989 8192
rect 9053 8128 9061 8192
rect 8741 7104 9061 8128
rect 8741 7040 8749 7104
rect 8813 7040 8829 7104
rect 8893 7040 8909 7104
rect 8973 7040 8989 7104
rect 9053 7040 9061 7104
rect 8523 6764 8589 6765
rect 8523 6700 8524 6764
rect 8588 6700 8589 6764
rect 8523 6699 8589 6700
rect 8523 6492 8589 6493
rect 8523 6428 8524 6492
rect 8588 6428 8589 6492
rect 8523 6427 8589 6428
rect 8339 3364 8405 3365
rect 8339 3300 8340 3364
rect 8404 3300 8405 3364
rect 8339 3299 8405 3300
rect 6142 3232 6150 3296
rect 6214 3232 6230 3296
rect 6294 3232 6310 3296
rect 6374 3232 6390 3296
rect 6454 3232 6462 3296
rect 5763 3228 5829 3229
rect 5763 3164 5764 3228
rect 5828 3164 5829 3228
rect 5763 3163 5829 3164
rect 3543 2688 3551 2752
rect 3615 2688 3631 2752
rect 3695 2688 3711 2752
rect 3775 2688 3791 2752
rect 3855 2688 3863 2752
rect 3543 2128 3863 2688
rect 6142 2208 6462 3232
rect 8526 2549 8586 6427
rect 8741 6016 9061 7040
rect 8741 5952 8749 6016
rect 8813 5952 8829 6016
rect 8893 5952 8909 6016
rect 8973 5952 8989 6016
rect 9053 5952 9061 6016
rect 8741 4928 9061 5952
rect 9262 5949 9322 18395
rect 9446 18053 9506 19075
rect 9443 18052 9509 18053
rect 9443 17988 9444 18052
rect 9508 17988 9509 18052
rect 9443 17987 9509 17988
rect 9443 15332 9509 15333
rect 9443 15268 9444 15332
rect 9508 15268 9509 15332
rect 9443 15267 9509 15268
rect 9446 6085 9506 15267
rect 9627 12476 9693 12477
rect 9627 12412 9628 12476
rect 9692 12412 9693 12476
rect 9627 12411 9693 12412
rect 9630 12069 9690 12411
rect 9627 12068 9693 12069
rect 9627 12004 9628 12068
rect 9692 12004 9693 12068
rect 9627 12003 9693 12004
rect 9814 11117 9874 19075
rect 10915 18596 10981 18597
rect 10915 18532 10916 18596
rect 10980 18532 10981 18596
rect 10915 18531 10981 18532
rect 10179 14788 10245 14789
rect 10179 14724 10180 14788
rect 10244 14724 10245 14788
rect 10179 14723 10245 14724
rect 10182 11933 10242 14723
rect 10179 11932 10245 11933
rect 10179 11868 10180 11932
rect 10244 11868 10245 11932
rect 10179 11867 10245 11868
rect 9811 11116 9877 11117
rect 9811 11052 9812 11116
rect 9876 11052 9877 11116
rect 9811 11051 9877 11052
rect 10918 10165 10978 18531
rect 11102 11389 11162 19619
rect 11340 19616 11660 20640
rect 11340 19552 11348 19616
rect 11412 19552 11428 19616
rect 11492 19552 11508 19616
rect 11572 19552 11588 19616
rect 11652 19552 11660 19616
rect 11340 18528 11660 19552
rect 11340 18464 11348 18528
rect 11412 18464 11428 18528
rect 11492 18464 11508 18528
rect 11572 18464 11588 18528
rect 11652 18464 11660 18528
rect 11340 17440 11660 18464
rect 11340 17376 11348 17440
rect 11412 17376 11428 17440
rect 11492 17376 11508 17440
rect 11572 17376 11588 17440
rect 11652 17376 11660 17440
rect 11340 16352 11660 17376
rect 11340 16288 11348 16352
rect 11412 16288 11428 16352
rect 11492 16288 11508 16352
rect 11572 16288 11588 16352
rect 11652 16288 11660 16352
rect 11340 15264 11660 16288
rect 11340 15200 11348 15264
rect 11412 15200 11428 15264
rect 11492 15200 11508 15264
rect 11572 15200 11588 15264
rect 11652 15200 11660 15264
rect 11340 14176 11660 15200
rect 11340 14112 11348 14176
rect 11412 14112 11428 14176
rect 11492 14112 11508 14176
rect 11572 14112 11588 14176
rect 11652 14112 11660 14176
rect 11340 13088 11660 14112
rect 11340 13024 11348 13088
rect 11412 13024 11428 13088
rect 11492 13024 11508 13088
rect 11572 13024 11588 13088
rect 11652 13024 11660 13088
rect 11340 12000 11660 13024
rect 13939 20160 14259 20720
rect 13939 20096 13947 20160
rect 14011 20096 14027 20160
rect 14091 20096 14107 20160
rect 14171 20096 14187 20160
rect 14251 20096 14259 20160
rect 13939 19072 14259 20096
rect 13939 19008 13947 19072
rect 14011 19008 14027 19072
rect 14091 19008 14107 19072
rect 14171 19008 14187 19072
rect 14251 19008 14259 19072
rect 13939 17984 14259 19008
rect 13939 17920 13947 17984
rect 14011 17920 14027 17984
rect 14091 17920 14107 17984
rect 14171 17920 14187 17984
rect 14251 17920 14259 17984
rect 13939 16896 14259 17920
rect 13939 16832 13947 16896
rect 14011 16832 14027 16896
rect 14091 16832 14107 16896
rect 14171 16832 14187 16896
rect 14251 16832 14259 16896
rect 13939 15808 14259 16832
rect 13939 15744 13947 15808
rect 14011 15744 14027 15808
rect 14091 15744 14107 15808
rect 14171 15744 14187 15808
rect 14251 15744 14259 15808
rect 13939 14720 14259 15744
rect 13939 14656 13947 14720
rect 14011 14656 14027 14720
rect 14091 14656 14107 14720
rect 14171 14656 14187 14720
rect 14251 14656 14259 14720
rect 13939 13632 14259 14656
rect 13939 13568 13947 13632
rect 14011 13568 14027 13632
rect 14091 13568 14107 13632
rect 14171 13568 14187 13632
rect 14251 13568 14259 13632
rect 11835 13020 11901 13021
rect 11835 12956 11836 13020
rect 11900 12956 11901 13020
rect 11835 12955 11901 12956
rect 11340 11936 11348 12000
rect 11412 11936 11428 12000
rect 11492 11936 11508 12000
rect 11572 11936 11588 12000
rect 11652 11936 11660 12000
rect 11099 11388 11165 11389
rect 11099 11324 11100 11388
rect 11164 11324 11165 11388
rect 11099 11323 11165 11324
rect 10915 10164 10981 10165
rect 10915 10100 10916 10164
rect 10980 10100 10981 10164
rect 10915 10099 10981 10100
rect 11102 10029 11162 11323
rect 11340 10912 11660 11936
rect 11340 10848 11348 10912
rect 11412 10848 11428 10912
rect 11492 10848 11508 10912
rect 11572 10848 11588 10912
rect 11652 10848 11660 10912
rect 11099 10028 11165 10029
rect 11099 9964 11100 10028
rect 11164 9964 11165 10028
rect 11099 9963 11165 9964
rect 11340 9824 11660 10848
rect 11838 10573 11898 12955
rect 13939 12544 14259 13568
rect 13939 12480 13947 12544
rect 14011 12480 14027 12544
rect 14091 12480 14107 12544
rect 14171 12480 14187 12544
rect 14251 12480 14259 12544
rect 12019 11660 12085 11661
rect 12019 11596 12020 11660
rect 12084 11596 12085 11660
rect 12019 11595 12085 11596
rect 11835 10572 11901 10573
rect 11835 10508 11836 10572
rect 11900 10508 11901 10572
rect 11835 10507 11901 10508
rect 11340 9760 11348 9824
rect 11412 9760 11428 9824
rect 11492 9760 11508 9824
rect 11572 9760 11588 9824
rect 11652 9760 11660 9824
rect 10179 9620 10245 9621
rect 10179 9556 10180 9620
rect 10244 9556 10245 9620
rect 10179 9555 10245 9556
rect 9443 6084 9509 6085
rect 9443 6020 9444 6084
rect 9508 6020 9509 6084
rect 9443 6019 9509 6020
rect 9259 5948 9325 5949
rect 9259 5884 9260 5948
rect 9324 5884 9325 5948
rect 9259 5883 9325 5884
rect 8741 4864 8749 4928
rect 8813 4864 8829 4928
rect 8893 4864 8909 4928
rect 8973 4864 8989 4928
rect 9053 4864 9061 4928
rect 8741 3840 9061 4864
rect 9446 3909 9506 6019
rect 10182 4997 10242 9555
rect 11340 8736 11660 9760
rect 11340 8672 11348 8736
rect 11412 8672 11428 8736
rect 11492 8672 11508 8736
rect 11572 8672 11588 8736
rect 11652 8672 11660 8736
rect 11340 7648 11660 8672
rect 11340 7584 11348 7648
rect 11412 7584 11428 7648
rect 11492 7584 11508 7648
rect 11572 7584 11588 7648
rect 11652 7584 11660 7648
rect 11340 6560 11660 7584
rect 12022 6765 12082 11595
rect 13939 11456 14259 12480
rect 13939 11392 13947 11456
rect 14011 11392 14027 11456
rect 14091 11392 14107 11456
rect 14171 11392 14187 11456
rect 14251 11392 14259 11456
rect 13939 10368 14259 11392
rect 13939 10304 13947 10368
rect 14011 10304 14027 10368
rect 14091 10304 14107 10368
rect 14171 10304 14187 10368
rect 14251 10304 14259 10368
rect 13939 9280 14259 10304
rect 13939 9216 13947 9280
rect 14011 9216 14027 9280
rect 14091 9216 14107 9280
rect 14171 9216 14187 9280
rect 14251 9216 14259 9280
rect 13939 8192 14259 9216
rect 13939 8128 13947 8192
rect 14011 8128 14027 8192
rect 14091 8128 14107 8192
rect 14171 8128 14187 8192
rect 14251 8128 14259 8192
rect 13939 7104 14259 8128
rect 13939 7040 13947 7104
rect 14011 7040 14027 7104
rect 14091 7040 14107 7104
rect 14171 7040 14187 7104
rect 14251 7040 14259 7104
rect 12019 6764 12085 6765
rect 12019 6700 12020 6764
rect 12084 6700 12085 6764
rect 12019 6699 12085 6700
rect 11340 6496 11348 6560
rect 11412 6496 11428 6560
rect 11492 6496 11508 6560
rect 11572 6496 11588 6560
rect 11652 6496 11660 6560
rect 11340 5472 11660 6496
rect 11340 5408 11348 5472
rect 11412 5408 11428 5472
rect 11492 5408 11508 5472
rect 11572 5408 11588 5472
rect 11652 5408 11660 5472
rect 10179 4996 10245 4997
rect 10179 4932 10180 4996
rect 10244 4932 10245 4996
rect 10179 4931 10245 4932
rect 9811 4724 9877 4725
rect 9811 4660 9812 4724
rect 9876 4660 9877 4724
rect 9811 4659 9877 4660
rect 9443 3908 9509 3909
rect 9443 3844 9444 3908
rect 9508 3844 9509 3908
rect 9443 3843 9509 3844
rect 8741 3776 8749 3840
rect 8813 3776 8829 3840
rect 8893 3776 8909 3840
rect 8973 3776 8989 3840
rect 9053 3776 9061 3840
rect 8741 2752 9061 3776
rect 9814 3637 9874 4659
rect 11340 4384 11660 5408
rect 11340 4320 11348 4384
rect 11412 4320 11428 4384
rect 11492 4320 11508 4384
rect 11572 4320 11588 4384
rect 11652 4320 11660 4384
rect 9811 3636 9877 3637
rect 9811 3572 9812 3636
rect 9876 3572 9877 3636
rect 9811 3571 9877 3572
rect 8741 2688 8749 2752
rect 8813 2688 8829 2752
rect 8893 2688 8909 2752
rect 8973 2688 8989 2752
rect 9053 2688 9061 2752
rect 8523 2548 8589 2549
rect 8523 2484 8524 2548
rect 8588 2484 8589 2548
rect 8523 2483 8589 2484
rect 6142 2144 6150 2208
rect 6214 2144 6230 2208
rect 6294 2144 6310 2208
rect 6374 2144 6390 2208
rect 6454 2144 6462 2208
rect 6142 2128 6462 2144
rect 8741 2128 9061 2688
rect 11340 3296 11660 4320
rect 11340 3232 11348 3296
rect 11412 3232 11428 3296
rect 11492 3232 11508 3296
rect 11572 3232 11588 3296
rect 11652 3232 11660 3296
rect 11340 2208 11660 3232
rect 11340 2144 11348 2208
rect 11412 2144 11428 2208
rect 11492 2144 11508 2208
rect 11572 2144 11588 2208
rect 11652 2144 11660 2208
rect 11340 2128 11660 2144
rect 13939 6016 14259 7040
rect 13939 5952 13947 6016
rect 14011 5952 14027 6016
rect 14091 5952 14107 6016
rect 14171 5952 14187 6016
rect 14251 5952 14259 6016
rect 13939 4928 14259 5952
rect 13939 4864 13947 4928
rect 14011 4864 14027 4928
rect 14091 4864 14107 4928
rect 14171 4864 14187 4928
rect 14251 4864 14259 4928
rect 13939 3840 14259 4864
rect 13939 3776 13947 3840
rect 14011 3776 14027 3840
rect 14091 3776 14107 3840
rect 14171 3776 14187 3840
rect 14251 3776 14259 3840
rect 13939 2752 14259 3776
rect 13939 2688 13947 2752
rect 14011 2688 14027 2752
rect 14091 2688 14107 2752
rect 14171 2688 14187 2752
rect 14251 2688 14259 2752
rect 13939 2128 14259 2688
rect 16538 20704 16858 20720
rect 16538 20640 16546 20704
rect 16610 20640 16626 20704
rect 16690 20640 16706 20704
rect 16770 20640 16786 20704
rect 16850 20640 16858 20704
rect 16538 19616 16858 20640
rect 16538 19552 16546 19616
rect 16610 19552 16626 19616
rect 16690 19552 16706 19616
rect 16770 19552 16786 19616
rect 16850 19552 16858 19616
rect 16538 18528 16858 19552
rect 16538 18464 16546 18528
rect 16610 18464 16626 18528
rect 16690 18464 16706 18528
rect 16770 18464 16786 18528
rect 16850 18464 16858 18528
rect 16538 17440 16858 18464
rect 16538 17376 16546 17440
rect 16610 17376 16626 17440
rect 16690 17376 16706 17440
rect 16770 17376 16786 17440
rect 16850 17376 16858 17440
rect 16538 16352 16858 17376
rect 16538 16288 16546 16352
rect 16610 16288 16626 16352
rect 16690 16288 16706 16352
rect 16770 16288 16786 16352
rect 16850 16288 16858 16352
rect 16538 15264 16858 16288
rect 16538 15200 16546 15264
rect 16610 15200 16626 15264
rect 16690 15200 16706 15264
rect 16770 15200 16786 15264
rect 16850 15200 16858 15264
rect 16538 14176 16858 15200
rect 16538 14112 16546 14176
rect 16610 14112 16626 14176
rect 16690 14112 16706 14176
rect 16770 14112 16786 14176
rect 16850 14112 16858 14176
rect 16538 13088 16858 14112
rect 16538 13024 16546 13088
rect 16610 13024 16626 13088
rect 16690 13024 16706 13088
rect 16770 13024 16786 13088
rect 16850 13024 16858 13088
rect 16538 12000 16858 13024
rect 16538 11936 16546 12000
rect 16610 11936 16626 12000
rect 16690 11936 16706 12000
rect 16770 11936 16786 12000
rect 16850 11936 16858 12000
rect 16538 10912 16858 11936
rect 16538 10848 16546 10912
rect 16610 10848 16626 10912
rect 16690 10848 16706 10912
rect 16770 10848 16786 10912
rect 16850 10848 16858 10912
rect 16538 9824 16858 10848
rect 16538 9760 16546 9824
rect 16610 9760 16626 9824
rect 16690 9760 16706 9824
rect 16770 9760 16786 9824
rect 16850 9760 16858 9824
rect 16538 8736 16858 9760
rect 16538 8672 16546 8736
rect 16610 8672 16626 8736
rect 16690 8672 16706 8736
rect 16770 8672 16786 8736
rect 16850 8672 16858 8736
rect 16538 7648 16858 8672
rect 16538 7584 16546 7648
rect 16610 7584 16626 7648
rect 16690 7584 16706 7648
rect 16770 7584 16786 7648
rect 16850 7584 16858 7648
rect 16538 6560 16858 7584
rect 16538 6496 16546 6560
rect 16610 6496 16626 6560
rect 16690 6496 16706 6560
rect 16770 6496 16786 6560
rect 16850 6496 16858 6560
rect 16538 5472 16858 6496
rect 16538 5408 16546 5472
rect 16610 5408 16626 5472
rect 16690 5408 16706 5472
rect 16770 5408 16786 5472
rect 16850 5408 16858 5472
rect 16538 4384 16858 5408
rect 16538 4320 16546 4384
rect 16610 4320 16626 4384
rect 16690 4320 16706 4384
rect 16770 4320 16786 4384
rect 16850 4320 16858 4384
rect 16538 3296 16858 4320
rect 16538 3232 16546 3296
rect 16610 3232 16626 3296
rect 16690 3232 16706 3296
rect 16770 3232 16786 3296
rect 16850 3232 16858 3296
rect 16538 2208 16858 3232
rect 16538 2144 16546 2208
rect 16610 2144 16626 2208
rect 16690 2144 16706 2208
rect 16770 2144 16786 2208
rect 16850 2144 16858 2208
rect 16538 2128 16858 2144
rect 19137 20160 19457 20720
rect 19137 20096 19145 20160
rect 19209 20096 19225 20160
rect 19289 20096 19305 20160
rect 19369 20096 19385 20160
rect 19449 20096 19457 20160
rect 19137 19072 19457 20096
rect 19137 19008 19145 19072
rect 19209 19008 19225 19072
rect 19289 19008 19305 19072
rect 19369 19008 19385 19072
rect 19449 19008 19457 19072
rect 19137 17984 19457 19008
rect 19137 17920 19145 17984
rect 19209 17920 19225 17984
rect 19289 17920 19305 17984
rect 19369 17920 19385 17984
rect 19449 17920 19457 17984
rect 19137 16896 19457 17920
rect 19137 16832 19145 16896
rect 19209 16832 19225 16896
rect 19289 16832 19305 16896
rect 19369 16832 19385 16896
rect 19449 16832 19457 16896
rect 19137 15808 19457 16832
rect 19137 15744 19145 15808
rect 19209 15744 19225 15808
rect 19289 15744 19305 15808
rect 19369 15744 19385 15808
rect 19449 15744 19457 15808
rect 19137 14720 19457 15744
rect 19137 14656 19145 14720
rect 19209 14656 19225 14720
rect 19289 14656 19305 14720
rect 19369 14656 19385 14720
rect 19449 14656 19457 14720
rect 19137 13632 19457 14656
rect 19137 13568 19145 13632
rect 19209 13568 19225 13632
rect 19289 13568 19305 13632
rect 19369 13568 19385 13632
rect 19449 13568 19457 13632
rect 19137 12544 19457 13568
rect 19137 12480 19145 12544
rect 19209 12480 19225 12544
rect 19289 12480 19305 12544
rect 19369 12480 19385 12544
rect 19449 12480 19457 12544
rect 19137 11456 19457 12480
rect 19137 11392 19145 11456
rect 19209 11392 19225 11456
rect 19289 11392 19305 11456
rect 19369 11392 19385 11456
rect 19449 11392 19457 11456
rect 19137 10368 19457 11392
rect 19137 10304 19145 10368
rect 19209 10304 19225 10368
rect 19289 10304 19305 10368
rect 19369 10304 19385 10368
rect 19449 10304 19457 10368
rect 19137 9280 19457 10304
rect 19137 9216 19145 9280
rect 19209 9216 19225 9280
rect 19289 9216 19305 9280
rect 19369 9216 19385 9280
rect 19449 9216 19457 9280
rect 19137 8192 19457 9216
rect 19137 8128 19145 8192
rect 19209 8128 19225 8192
rect 19289 8128 19305 8192
rect 19369 8128 19385 8192
rect 19449 8128 19457 8192
rect 19137 7104 19457 8128
rect 19137 7040 19145 7104
rect 19209 7040 19225 7104
rect 19289 7040 19305 7104
rect 19369 7040 19385 7104
rect 19449 7040 19457 7104
rect 19137 6016 19457 7040
rect 19137 5952 19145 6016
rect 19209 5952 19225 6016
rect 19289 5952 19305 6016
rect 19369 5952 19385 6016
rect 19449 5952 19457 6016
rect 19137 4928 19457 5952
rect 19137 4864 19145 4928
rect 19209 4864 19225 4928
rect 19289 4864 19305 4928
rect 19369 4864 19385 4928
rect 19449 4864 19457 4928
rect 19137 3840 19457 4864
rect 19137 3776 19145 3840
rect 19209 3776 19225 3840
rect 19289 3776 19305 3840
rect 19369 3776 19385 3840
rect 19449 3776 19457 3840
rect 19137 2752 19457 3776
rect 19137 2688 19145 2752
rect 19209 2688 19225 2752
rect 19289 2688 19305 2752
rect 19369 2688 19385 2752
rect 19449 2688 19457 2752
rect 19137 2128 19457 2688
rect 21736 20704 22056 20720
rect 21736 20640 21744 20704
rect 21808 20640 21824 20704
rect 21888 20640 21904 20704
rect 21968 20640 21984 20704
rect 22048 20640 22056 20704
rect 21736 19616 22056 20640
rect 21736 19552 21744 19616
rect 21808 19552 21824 19616
rect 21888 19552 21904 19616
rect 21968 19552 21984 19616
rect 22048 19552 22056 19616
rect 21736 18528 22056 19552
rect 21736 18464 21744 18528
rect 21808 18464 21824 18528
rect 21888 18464 21904 18528
rect 21968 18464 21984 18528
rect 22048 18464 22056 18528
rect 21736 17440 22056 18464
rect 21736 17376 21744 17440
rect 21808 17376 21824 17440
rect 21888 17376 21904 17440
rect 21968 17376 21984 17440
rect 22048 17376 22056 17440
rect 21736 16352 22056 17376
rect 21736 16288 21744 16352
rect 21808 16288 21824 16352
rect 21888 16288 21904 16352
rect 21968 16288 21984 16352
rect 22048 16288 22056 16352
rect 21736 15264 22056 16288
rect 21736 15200 21744 15264
rect 21808 15200 21824 15264
rect 21888 15200 21904 15264
rect 21968 15200 21984 15264
rect 22048 15200 22056 15264
rect 21736 14176 22056 15200
rect 21736 14112 21744 14176
rect 21808 14112 21824 14176
rect 21888 14112 21904 14176
rect 21968 14112 21984 14176
rect 22048 14112 22056 14176
rect 21736 13088 22056 14112
rect 21736 13024 21744 13088
rect 21808 13024 21824 13088
rect 21888 13024 21904 13088
rect 21968 13024 21984 13088
rect 22048 13024 22056 13088
rect 21736 12000 22056 13024
rect 21736 11936 21744 12000
rect 21808 11936 21824 12000
rect 21888 11936 21904 12000
rect 21968 11936 21984 12000
rect 22048 11936 22056 12000
rect 21736 10912 22056 11936
rect 21736 10848 21744 10912
rect 21808 10848 21824 10912
rect 21888 10848 21904 10912
rect 21968 10848 21984 10912
rect 22048 10848 22056 10912
rect 21736 9824 22056 10848
rect 21736 9760 21744 9824
rect 21808 9760 21824 9824
rect 21888 9760 21904 9824
rect 21968 9760 21984 9824
rect 22048 9760 22056 9824
rect 21736 8736 22056 9760
rect 21736 8672 21744 8736
rect 21808 8672 21824 8736
rect 21888 8672 21904 8736
rect 21968 8672 21984 8736
rect 22048 8672 22056 8736
rect 21736 7648 22056 8672
rect 21736 7584 21744 7648
rect 21808 7584 21824 7648
rect 21888 7584 21904 7648
rect 21968 7584 21984 7648
rect 22048 7584 22056 7648
rect 21736 6560 22056 7584
rect 21736 6496 21744 6560
rect 21808 6496 21824 6560
rect 21888 6496 21904 6560
rect 21968 6496 21984 6560
rect 22048 6496 22056 6560
rect 21736 5472 22056 6496
rect 21736 5408 21744 5472
rect 21808 5408 21824 5472
rect 21888 5408 21904 5472
rect 21968 5408 21984 5472
rect 22048 5408 22056 5472
rect 21736 4384 22056 5408
rect 21736 4320 21744 4384
rect 21808 4320 21824 4384
rect 21888 4320 21904 4384
rect 21968 4320 21984 4384
rect 22048 4320 22056 4384
rect 21736 3296 22056 4320
rect 21736 3232 21744 3296
rect 21808 3232 21824 3296
rect 21888 3232 21904 3296
rect 21968 3232 21984 3296
rect 22048 3232 22056 3296
rect 21736 2208 22056 3232
rect 21736 2144 21744 2208
rect 21808 2144 21824 2208
rect 21888 2144 21904 2208
rect 21968 2144 21984 2208
rect 22048 2144 22056 2208
rect 21736 2128 22056 2144
use sky130_fd_sc_hd__diode_2  ANTENNA__079__A dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform 1 0 1656 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__089__A
timestamp 1649977179
transform -1 0 14628 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__091__A
timestamp 1649977179
transform -1 0 11868 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__092__A
timestamp 1649977179
transform -1 0 14996 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__093__A
timestamp 1649977179
transform 1 0 16928 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__095__A
timestamp 1649977179
transform 1 0 16468 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__096__A
timestamp 1649977179
transform -1 0 18400 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__097__A
timestamp 1649977179
transform 1 0 18400 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__099__A
timestamp 1649977179
transform -1 0 19872 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__100__A
timestamp 1649977179
transform -1 0 15732 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__101__A
timestamp 1649977179
transform -1 0 16100 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__103__A
timestamp 1649977179
transform 1 0 18584 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__104__A
timestamp 1649977179
transform -1 0 18032 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__105__A
timestamp 1649977179
transform -1 0 19688 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__109__A
timestamp 1649977179
transform -1 0 8464 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__111__A
timestamp 1649977179
transform -1 0 6992 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__112__A
timestamp 1649977179
transform -1 0 7176 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__113__A
timestamp 1649977179
transform 1 0 9016 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__115__A
timestamp 1649977179
transform 1 0 10212 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__116__A
timestamp 1649977179
transform -1 0 9108 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__117__A
timestamp 1649977179
transform 1 0 10028 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__119__A
timestamp 1649977179
transform -1 0 14812 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__120__A
timestamp 1649977179
transform -1 0 9108 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__121__A
timestamp 1649977179
transform 1 0 8832 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__123__A
timestamp 1649977179
transform 1 0 9476 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__124__A
timestamp 1649977179
transform -1 0 14260 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__125__A
timestamp 1649977179
transform -1 0 16284 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_bottom_track_1.sky130_fd_sc_hd__dfxtp_1_0__CLK
timestamp 1649977179
transform 1 0 21252 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_bottom_track_1.sky130_fd_sc_hd__dfxtp_1_1__CLK
timestamp 1649977179
transform 1 0 14444 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_bottom_track_1.sky130_fd_sc_hd__dfxtp_1_1__D
timestamp 1649977179
transform 1 0 13524 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_bottom_track_1.sky130_fd_sc_hd__dfxtp_1_2__CLK
timestamp 1649977179
transform 1 0 13708 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_bottom_track_1.sky130_fd_sc_hd__dfxtp_1_3__CLK
timestamp 1649977179
transform 1 0 13156 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_bottom_track_3.sky130_fd_sc_hd__dfxtp_1_0__CLK
timestamp 1649977179
transform 1 0 15732 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_bottom_track_3.sky130_fd_sc_hd__dfxtp_1_1__CLK
timestamp 1649977179
transform 1 0 13708 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_bottom_track_3.sky130_fd_sc_hd__dfxtp_1_2__CLK
timestamp 1649977179
transform 1 0 15548 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_bottom_track_3.sky130_fd_sc_hd__dfxtp_1_3__CLK
timestamp 1649977179
transform 1 0 14628 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_bottom_track_5.sky130_fd_sc_hd__dfxtp_1_0__CLK
timestamp 1649977179
transform 1 0 16100 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_bottom_track_5.sky130_fd_sc_hd__dfxtp_1_1__CLK
timestamp 1649977179
transform 1 0 11960 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_bottom_track_5.sky130_fd_sc_hd__dfxtp_1_1__D
timestamp 1649977179
transform -1 0 13892 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_bottom_track_5.sky130_fd_sc_hd__dfxtp_1_2__CLK
timestamp 1649977179
transform 1 0 15916 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_bottom_track_5.sky130_fd_sc_hd__dfxtp_1_3__CLK
timestamp 1649977179
transform 1 0 18952 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_bottom_track_9.sky130_fd_sc_hd__dfxtp_1_0__CLK
timestamp 1649977179
transform 1 0 20792 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_bottom_track_9.sky130_fd_sc_hd__dfxtp_1_1__CLK
timestamp 1649977179
transform 1 0 19412 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_bottom_track_9.sky130_fd_sc_hd__dfxtp_1_2__CLK
timestamp 1649977179
transform 1 0 17848 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_bottom_track_9.sky130_fd_sc_hd__dfxtp_1_2__D
timestamp 1649977179
transform -1 0 18216 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_bottom_track_9.sky130_fd_sc_hd__dfxtp_1_3__CLK
timestamp 1649977179
transform 1 0 17756 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_bottom_track_17.sky130_fd_sc_hd__dfxtp_1_0__CLK
timestamp 1649977179
transform 1 0 21344 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_bottom_track_17.sky130_fd_sc_hd__dfxtp_1_1__CLK
timestamp 1649977179
transform 1 0 13340 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_bottom_track_17.sky130_fd_sc_hd__dfxtp_1_1__D
timestamp 1649977179
transform 1 0 13524 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_bottom_track_17.sky130_fd_sc_hd__dfxtp_1_2__CLK
timestamp 1649977179
transform 1 0 18308 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_bottom_track_25.sky130_fd_sc_hd__dfxtp_1_0__CLK
timestamp 1649977179
transform 1 0 20700 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_bottom_track_25.sky130_fd_sc_hd__dfxtp_1_1__CLK
timestamp 1649977179
transform 1 0 20884 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_bottom_track_25.sky130_fd_sc_hd__dfxtp_1_2__CLK
timestamp 1649977179
transform 1 0 21344 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_bottom_track_33.sky130_fd_sc_hd__dfxtp_1_0__CLK
timestamp 1649977179
transform 1 0 21068 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_bottom_track_33.sky130_fd_sc_hd__dfxtp_1_1__CLK
timestamp 1649977179
transform 1 0 18584 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_bottom_track_33.sky130_fd_sc_hd__dfxtp_1_1__D
timestamp 1649977179
transform 1 0 18768 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_bottom_track_33.sky130_fd_sc_hd__dfxtp_1_2__CLK
timestamp 1649977179
transform 1 0 21068 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_1.sky130_fd_sc_hd__dfxtp_1_0__CLK
timestamp 1649977179
transform 1 0 21436 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_1.sky130_fd_sc_hd__dfxtp_1_1__CLK
timestamp 1649977179
transform 1 0 15916 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_1.sky130_fd_sc_hd__dfxtp_1_1__D
timestamp 1649977179
transform 1 0 16100 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_1.sky130_fd_sc_hd__dfxtp_1_2__CLK
timestamp 1649977179
transform 1 0 18124 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_3.sky130_fd_sc_hd__dfxtp_1_0__CLK
timestamp 1649977179
transform 1 0 18308 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_3.sky130_fd_sc_hd__dfxtp_1_1__CLK
timestamp 1649977179
transform 1 0 13340 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_3.sky130_fd_sc_hd__dfxtp_1_1__D
timestamp 1649977179
transform -1 0 13708 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_3.sky130_fd_sc_hd__dfxtp_1_2__CLK
timestamp 1649977179
transform 1 0 13708 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_5.sky130_fd_sc_hd__dfxtp_1_0__CLK
timestamp 1649977179
transform 1 0 13524 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_5.sky130_fd_sc_hd__dfxtp_1_1__CLK
timestamp 1649977179
transform 1 0 14168 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_5.sky130_fd_sc_hd__dfxtp_1_2__CLK
timestamp 1649977179
transform 1 0 14352 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_7.sky130_fd_sc_hd__dfxtp_1_0__CLK
timestamp 1649977179
transform 1 0 15640 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_7.sky130_fd_sc_hd__dfxtp_1_1__CLK
timestamp 1649977179
transform 1 0 13984 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_7.sky130_fd_sc_hd__dfxtp_1_2__CLK
timestamp 1649977179
transform 1 0 12512 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_9.sky130_fd_sc_hd__dfxtp_1_0__CLK
timestamp 1649977179
transform 1 0 15732 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_9.sky130_fd_sc_hd__dfxtp_1_1__CLK
timestamp 1649977179
transform 1 0 18124 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_9.sky130_fd_sc_hd__dfxtp_1_2__CLK
timestamp 1649977179
transform 1 0 18952 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_11.sky130_fd_sc_hd__dfxtp_1_0__CLK
timestamp 1649977179
transform 1 0 21252 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_11.sky130_fd_sc_hd__dfxtp_1_1__CLK
timestamp 1649977179
transform 1 0 20792 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_11.sky130_fd_sc_hd__dfxtp_1_2__CLK
timestamp 1649977179
transform 1 0 18124 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_13.sky130_fd_sc_hd__dfxtp_1_0__CLK
timestamp 1649977179
transform 1 0 20884 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_13.sky130_fd_sc_hd__dfxtp_1_1__CLK
timestamp 1649977179
transform 1 0 21068 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_13.sky130_fd_sc_hd__dfxtp_1_2__CLK
timestamp 1649977179
transform 1 0 16376 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_15.sky130_fd_sc_hd__dfxtp_1_0__CLK
timestamp 1649977179
transform 1 0 21436 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_15.sky130_fd_sc_hd__dfxtp_1_1__CLK
timestamp 1649977179
transform 1 0 19780 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_15.sky130_fd_sc_hd__dfxtp_1_2__CLK
timestamp 1649977179
transform 1 0 20976 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_17.sky130_fd_sc_hd__dfxtp_1_0__CLK
timestamp 1649977179
transform 1 0 16744 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_17.sky130_fd_sc_hd__dfxtp_1_1__CLK
timestamp 1649977179
transform 1 0 13432 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_19.sky130_fd_sc_hd__dfxtp_1_0__CLK
timestamp 1649977179
transform 1 0 14076 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_19.sky130_fd_sc_hd__dfxtp_1_1__CLK
timestamp 1649977179
transform 1 0 14444 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_21.sky130_fd_sc_hd__dfxtp_1_0__CLK
timestamp 1649977179
transform 1 0 17572 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_21.sky130_fd_sc_hd__dfxtp_1_1__CLK
timestamp 1649977179
transform 1 0 19596 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_23.sky130_fd_sc_hd__dfxtp_1_0__CLK
timestamp 1649977179
transform 1 0 21160 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_23.sky130_fd_sc_hd__dfxtp_1_1__CLK
timestamp 1649977179
transform 1 0 19964 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_25.sky130_fd_sc_hd__dfxtp_1_0__CLK
timestamp 1649977179
transform 1 0 19596 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_25.sky130_fd_sc_hd__dfxtp_1_1__CLK
timestamp 1649977179
transform 1 0 17664 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_29.sky130_fd_sc_hd__dfxtp_1_0__CLK
timestamp 1649977179
transform 1 0 20424 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_29.sky130_fd_sc_hd__dfxtp_1_1__CLK
timestamp 1649977179
transform 1 0 20976 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_31.sky130_fd_sc_hd__dfxtp_1_0__CLK
timestamp 1649977179
transform 1 0 21252 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_31.sky130_fd_sc_hd__dfxtp_1_1__CLK
timestamp 1649977179
transform 1 0 21436 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_33.sky130_fd_sc_hd__dfxtp_1_0__CLK
timestamp 1649977179
transform 1 0 18124 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_33.sky130_fd_sc_hd__dfxtp_1_1__CLK
timestamp 1649977179
transform 1 0 18124 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_35.sky130_fd_sc_hd__dfxtp_1_0__CLK
timestamp 1649977179
transform 1 0 16560 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_35.sky130_fd_sc_hd__dfxtp_1_1__CLK
timestamp 1649977179
transform 1 0 14536 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_37.sky130_fd_sc_hd__dfxtp_1_0__CLK
timestamp 1649977179
transform 1 0 13064 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_37.sky130_fd_sc_hd__dfxtp_1_1__CLK
timestamp 1649977179
transform 1 0 16192 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_39.sky130_fd_sc_hd__dfxtp_1_0__CLK
timestamp 1649977179
transform 1 0 21068 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_39.sky130_fd_sc_hd__dfxtp_1_1__CLK
timestamp 1649977179
transform 1 0 20792 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_track_0.sky130_fd_sc_hd__dfxtp_1_0__CLK
timestamp 1649977179
transform 1 0 21252 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_track_0.sky130_fd_sc_hd__dfxtp_1_0__D
timestamp 1649977179
transform -1 0 21620 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_track_0.sky130_fd_sc_hd__dfxtp_1_1__CLK
timestamp 1649977179
transform 1 0 18124 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_track_0.sky130_fd_sc_hd__dfxtp_1_2__CLK
timestamp 1649977179
transform 1 0 15824 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_track_0.sky130_fd_sc_hd__dfxtp_1_2__D
timestamp 1649977179
transform -1 0 16192 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_track_0.sky130_fd_sc_hd__dfxtp_1_3__CLK
timestamp 1649977179
transform 1 0 14444 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_track_2.sky130_fd_sc_hd__dfxtp_1_0__CLK
timestamp 1649977179
transform 1 0 13248 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_track_2.sky130_fd_sc_hd__dfxtp_1_1__CLK
timestamp 1649977179
transform 1 0 11224 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_track_2.sky130_fd_sc_hd__dfxtp_1_2__CLK
timestamp 1649977179
transform 1 0 13616 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_track_2.sky130_fd_sc_hd__dfxtp_1_3__CLK
timestamp 1649977179
transform 1 0 13524 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_track_4.sky130_fd_sc_hd__dfxtp_1_0__CLK
timestamp 1649977179
transform 1 0 16560 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_track_4.sky130_fd_sc_hd__dfxtp_1_1__CLK
timestamp 1649977179
transform 1 0 13340 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_track_4.sky130_fd_sc_hd__dfxtp_1_1__D
timestamp 1649977179
transform -1 0 13708 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_track_4.sky130_fd_sc_hd__dfxtp_1_2__CLK
timestamp 1649977179
transform 1 0 13708 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_track_4.sky130_fd_sc_hd__dfxtp_1_3__CLK
timestamp 1649977179
transform 1 0 17940 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_track_8.sky130_fd_sc_hd__dfxtp_1_0__CLK
timestamp 1649977179
transform 1 0 19596 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_track_8.sky130_fd_sc_hd__dfxtp_1_1__CLK
timestamp 1649977179
transform 1 0 18216 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_track_8.sky130_fd_sc_hd__dfxtp_1_2__CLK
timestamp 1649977179
transform 1 0 13156 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_track_8.sky130_fd_sc_hd__dfxtp_1_2__D
timestamp 1649977179
transform 1 0 13340 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_track_8.sky130_fd_sc_hd__dfxtp_1_3__CLK
timestamp 1649977179
transform 1 0 20700 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_track_16.sky130_fd_sc_hd__dfxtp_1_0__CLK
timestamp 1649977179
transform 1 0 19320 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_track_16.sky130_fd_sc_hd__dfxtp_1_1__CLK
timestamp 1649977179
transform 1 0 15548 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_track_16.sky130_fd_sc_hd__dfxtp_1_1__D
timestamp 1649977179
transform 1 0 15732 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_track_16.sky130_fd_sc_hd__dfxtp_1_2__CLK
timestamp 1649977179
transform 1 0 13616 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_track_24.sky130_fd_sc_hd__dfxtp_1_0__CLK
timestamp 1649977179
transform 1 0 15916 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_track_24.sky130_fd_sc_hd__dfxtp_1_1__CLK
timestamp 1649977179
transform 1 0 15272 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_track_24.sky130_fd_sc_hd__dfxtp_1_1__D
timestamp 1649977179
transform 1 0 15456 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_track_24.sky130_fd_sc_hd__dfxtp_1_2__CLK
timestamp 1649977179
transform 1 0 18216 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_track_32.sky130_fd_sc_hd__dfxtp_1_0__CLK
timestamp 1649977179
transform 1 0 17572 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_track_32.sky130_fd_sc_hd__dfxtp_1_1__CLK
timestamp 1649977179
transform 1 0 15364 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_track_32.sky130_fd_sc_hd__dfxtp_1_2__CLK
timestamp 1649977179
transform 1 0 18400 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_1.mux_l1_in_0__A0
timestamp 1649977179
transform 1 0 11316 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_1.mux_l1_in_0__A1
timestamp 1649977179
transform 1 0 11132 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_1.mux_l1_in_0__S
timestamp 1649977179
transform 1 0 12328 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_1.mux_l1_in_1__A0
timestamp 1649977179
transform -1 0 10120 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_1.mux_l1_in_1__A1
timestamp 1649977179
transform 1 0 12236 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_1.mux_l1_in_1__S
timestamp 1649977179
transform 1 0 10948 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_1.mux_l1_in_2__A0
timestamp 1649977179
transform 1 0 8464 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_1.mux_l1_in_2__A1
timestamp 1649977179
transform 1 0 8648 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_1.mux_l1_in_2__S
timestamp 1649977179
transform -1 0 10120 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_1.mux_l2_in_1__A0
timestamp 1649977179
transform 1 0 8004 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_1.mux_l2_in_2__A0
timestamp 1649977179
transform 1 0 5244 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_1.mux_l2_in_2__A1
timestamp 1649977179
transform 1 0 5428 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_1.mux_l2_in_3__A1
timestamp 1649977179
transform 1 0 4600 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_3.mux_l1_in_0__A0
timestamp 1649977179
transform 1 0 10580 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_3.mux_l1_in_0__A1
timestamp 1649977179
transform 1 0 9476 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_3.mux_l1_in_1__A0
timestamp 1649977179
transform 1 0 9384 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_3.mux_l1_in_1__A1
timestamp 1649977179
transform -1 0 9752 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_3.mux_l2_in_1__A0
timestamp 1649977179
transform 1 0 4784 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_3.mux_l2_in_1__A1
timestamp 1649977179
transform 1 0 4140 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_3.mux_l2_in_2__A0
timestamp 1649977179
transform -1 0 1564 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_3.mux_l2_in_2__A1
timestamp 1649977179
transform 1 0 1472 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_3.mux_l2_in_3__A1
timestamp 1649977179
transform -1 0 1840 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_5.mux_l1_in_0__A0
timestamp 1649977179
transform 1 0 11684 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_5.mux_l1_in_0__A1
timestamp 1649977179
transform 1 0 11500 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_5.mux_l1_in_0__S
timestamp 1649977179
transform 1 0 13524 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_5.mux_l1_in_1__A0
timestamp 1649977179
transform 1 0 9752 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_5.mux_l1_in_1__A1
timestamp 1649977179
transform 1 0 10580 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_5.mux_l1_in_1__S
timestamp 1649977179
transform -1 0 10948 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_5.mux_l1_in_2__A0
timestamp 1649977179
transform 1 0 6900 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_5.mux_l1_in_2__A1
timestamp 1649977179
transform 1 0 7084 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_5.mux_l1_in_2__S
timestamp 1649977179
transform 1 0 8096 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_5.mux_l1_in_3__A0
timestamp 1649977179
transform 1 0 5888 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_5.mux_l1_in_3__A1
timestamp 1649977179
transform 1 0 6072 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_5.mux_l1_in_3__S
timestamp 1649977179
transform 1 0 7084 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_5.mux_l1_in_4__A0
timestamp 1649977179
transform 1 0 4600 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_5.mux_l1_in_4__A1
timestamp 1649977179
transform 1 0 4784 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_5.mux_l1_in_4__S
timestamp 1649977179
transform -1 0 5980 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_5.mux_l1_in_5__A0
timestamp 1649977179
transform 1 0 4508 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_5.mux_l1_in_5__A1
timestamp 1649977179
transform 1 0 4692 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_5.mux_l1_in_5__S
timestamp 1649977179
transform 1 0 5704 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_5.mux_l1_in_6__A0
timestamp 1649977179
transform -1 0 1564 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_5.mux_l1_in_6__A1
timestamp 1649977179
transform -1 0 1748 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_5.mux_l1_in_6__S
timestamp 1649977179
transform 1 0 3312 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_9.mux_l1_in_0__A0
timestamp 1649977179
transform 1 0 16100 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_9.mux_l1_in_0__A1
timestamp 1649977179
transform -1 0 16468 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_9.mux_l2_in_0__A0
timestamp 1649977179
transform -1 0 16468 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_9.mux_l2_in_0__S
timestamp 1649977179
transform 1 0 17112 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_9.mux_l2_in_1__A0
timestamp 1649977179
transform 1 0 6992 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_9.mux_l2_in_1__A1
timestamp 1649977179
transform 1 0 7176 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_9.mux_l2_in_1__S
timestamp 1649977179
transform 1 0 9016 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_9.mux_l2_in_2__A0
timestamp 1649977179
transform 1 0 3496 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_9.mux_l2_in_2__A1
timestamp 1649977179
transform 1 0 3312 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_9.mux_l2_in_2__S
timestamp 1649977179
transform 1 0 4692 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_9.mux_l2_in_3__A1
timestamp 1649977179
transform -1 0 4048 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_9.mux_l2_in_3__S
timestamp 1649977179
transform 1 0 4876 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_17.mux_l1_in_0__A0
timestamp 1649977179
transform 1 0 12236 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_17.mux_l1_in_0__A1
timestamp 1649977179
transform 1 0 12052 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_17.mux_l1_in_0__S
timestamp 1649977179
transform 1 0 13800 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_17.mux_l1_in_1__A0
timestamp 1649977179
transform 1 0 7360 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_17.mux_l1_in_1__A1
timestamp 1649977179
transform -1 0 7728 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_17.mux_l1_in_1__S
timestamp 1649977179
transform -1 0 8740 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_17.mux_l1_in_2__A0
timestamp 1649977179
transform -1 0 4048 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_17.mux_l1_in_2__A1
timestamp 1649977179
transform 1 0 3680 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_17.mux_l1_in_2__S
timestamp 1649977179
transform 1 0 5244 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_17.mux_l1_in_3__A1
timestamp 1649977179
transform -1 0 3680 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_17.mux_l1_in_3__S
timestamp 1649977179
transform 1 0 4784 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_25.mux_l1_in_0__A0
timestamp 1649977179
transform 1 0 17388 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_25.mux_l1_in_0__A1
timestamp 1649977179
transform 1 0 17204 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_25.mux_l1_in_1__A0
timestamp 1649977179
transform 1 0 8556 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_25.mux_l1_in_1__A1
timestamp 1649977179
transform 1 0 8740 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_25.mux_l1_in_2__A0
timestamp 1649977179
transform 1 0 10856 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_25.mux_l1_in_2__A1
timestamp 1649977179
transform 1 0 10672 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_33.mux_l1_in_0__A0
timestamp 1649977179
transform 1 0 9200 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_33.mux_l1_in_0__A1
timestamp 1649977179
transform 1 0 9016 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_33.mux_l1_in_0__S
timestamp 1649977179
transform 1 0 11040 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_33.mux_l1_in_1__A0
timestamp 1649977179
transform 1 0 3772 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_33.mux_l1_in_1__A1
timestamp 1649977179
transform 1 0 3956 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_33.mux_l1_in_1__S
timestamp 1649977179
transform 1 0 5060 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_33.mux_l1_in_2__A0
timestamp 1649977179
transform -1 0 4600 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_33.mux_l1_in_2__A1
timestamp 1649977179
transform -1 0 4416 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_33.mux_l1_in_2__S
timestamp 1649977179
transform 1 0 5428 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_1.mux_l1_in_0__A0
timestamp 1649977179
transform 1 0 5980 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_1.mux_l1_in_0__A1
timestamp 1649977179
transform 1 0 6164 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_1.mux_l1_in_0__S
timestamp 1649977179
transform 1 0 7176 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_1.mux_l1_in_1__A0
timestamp 1649977179
transform 1 0 4324 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_1.mux_l1_in_1__A1
timestamp 1649977179
transform 1 0 5428 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_1.mux_l1_in_1__S
timestamp 1649977179
transform -1 0 6256 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_1.mux_l1_in_2__A0
timestamp 1649977179
transform 1 0 5888 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_1.mux_l1_in_2__A1
timestamp 1649977179
transform 1 0 6072 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_1.mux_l1_in_2__S
timestamp 1649977179
transform 1 0 7176 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_1.mux_l1_in_3__A1
timestamp 1649977179
transform 1 0 4416 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_1.mux_l1_in_3__S
timestamp 1649977179
transform 1 0 7360 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_3.mux_l1_in_0__A0
timestamp 1649977179
transform -1 0 6256 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_3.mux_l1_in_0__A1
timestamp 1649977179
transform 1 0 5888 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_3.mux_l1_in_0__S
timestamp 1649977179
transform -1 0 7268 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_3.mux_l1_in_1__A0
timestamp 1649977179
transform 1 0 5704 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_3.mux_l1_in_1__A1
timestamp 1649977179
transform 1 0 5888 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_3.mux_l1_in_1__S
timestamp 1649977179
transform 1 0 6900 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_3.mux_l1_in_2__A0
timestamp 1649977179
transform 1 0 6716 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_3.mux_l1_in_2__A1
timestamp 1649977179
transform 1 0 6532 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_3.mux_l1_in_2__S
timestamp 1649977179
transform 1 0 7268 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_3.mux_l1_in_3__A1
timestamp 1649977179
transform 1 0 6072 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_3.mux_l1_in_3__S
timestamp 1649977179
transform 1 0 7268 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_5.mux_l1_in_0__A0
timestamp 1649977179
transform -1 0 6532 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_5.mux_l1_in_0__A1
timestamp 1649977179
transform -1 0 6256 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_5.mux_l1_in_1__A0
timestamp 1649977179
transform 1 0 7544 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_5.mux_l1_in_1__A1
timestamp 1649977179
transform 1 0 7728 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_5.mux_l1_in_2__A0
timestamp 1649977179
transform 1 0 8924 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_5.mux_l1_in_2__A1
timestamp 1649977179
transform 1 0 8556 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_5.mux_l1_in_3__A1
timestamp 1649977179
transform 1 0 7728 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_7.mux_l1_in_0__A0
timestamp 1649977179
transform -1 0 7636 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_7.mux_l1_in_0__A1
timestamp 1649977179
transform -1 0 6440 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_7.mux_l1_in_1__A0
timestamp 1649977179
transform 1 0 8924 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_7.mux_l1_in_1__A1
timestamp 1649977179
transform 1 0 9108 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_7.mux_l1_in_2__A0
timestamp 1649977179
transform 1 0 8648 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_7.mux_l1_in_2__A1
timestamp 1649977179
transform 1 0 8648 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_7.mux_l1_in_3__A1
timestamp 1649977179
transform 1 0 7544 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_9.mux_l1_in_0__A0
timestamp 1649977179
transform 1 0 12052 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_9.mux_l1_in_0__A1
timestamp 1649977179
transform 1 0 11500 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_9.mux_l2_in_0__A0
timestamp 1649977179
transform 1 0 9936 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_9.mux_l2_in_1__A1
timestamp 1649977179
transform 1 0 9476 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_11.mux_l1_in_0__A0
timestamp 1649977179
transform 1 0 14904 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_11.mux_l1_in_0__A1
timestamp 1649977179
transform 1 0 14720 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_11.mux_l2_in_0__A0
timestamp 1649977179
transform -1 0 10120 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_11.mux_l2_in_1__A1
timestamp 1649977179
transform 1 0 10304 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_13.mux_l1_in_0__A0
timestamp 1649977179
transform 1 0 15824 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_13.mux_l1_in_0__A1
timestamp 1649977179
transform 1 0 15640 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_13.mux_l2_in_0__A0
timestamp 1649977179
transform -1 0 11776 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_13.mux_l2_in_1__A1
timestamp 1649977179
transform 1 0 11868 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_15.mux_l1_in_0__A0
timestamp 1649977179
transform 1 0 17664 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_15.mux_l1_in_0__A1
timestamp 1649977179
transform 1 0 17480 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_15.mux_l2_in_0__A0
timestamp 1649977179
transform -1 0 13984 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_15.mux_l2_in_1__A1
timestamp 1649977179
transform 1 0 14352 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_17.mux_l1_in_0__A0
timestamp 1649977179
transform 1 0 9752 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_17.mux_l1_in_0__A1
timestamp 1649977179
transform 1 0 10120 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_17.mux_l1_in_1__A1
timestamp 1649977179
transform 1 0 8556 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_19.mux_l1_in_0__A0
timestamp 1649977179
transform 1 0 9844 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_19.mux_l1_in_0__A1
timestamp 1649977179
transform 1 0 11132 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_19.mux_l1_in_1__A1
timestamp 1649977179
transform 1 0 8096 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_21.mux_l1_in_0__A0
timestamp 1649977179
transform 1 0 11040 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_21.mux_l1_in_0__A1
timestamp 1649977179
transform 1 0 11224 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_21.mux_l1_in_1__A1
timestamp 1649977179
transform 1 0 8372 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_23.mux_l1_in_0__A0
timestamp 1649977179
transform 1 0 10948 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_23.mux_l1_in_0__A1
timestamp 1649977179
transform 1 0 11132 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_23.mux_l1_in_1__A1
timestamp 1649977179
transform 1 0 10304 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_25.mux_l1_in_0__A0
timestamp 1649977179
transform 1 0 11224 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_25.mux_l1_in_0__A1
timestamp 1649977179
transform 1 0 11040 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_25.mux_l1_in_1__A1
timestamp 1649977179
transform 1 0 10304 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_29.mux_l1_in_0__A0
timestamp 1649977179
transform 1 0 10396 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_29.mux_l1_in_0__A1
timestamp 1649977179
transform -1 0 11684 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_31.mux_l1_in_0__A0
timestamp 1649977179
transform 1 0 9384 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_31.mux_l1_in_0__A1
timestamp 1649977179
transform -1 0 11684 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_33.mux_l1_in_0__A0
timestamp 1649977179
transform 1 0 8372 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_33.mux_l1_in_0__A1
timestamp 1649977179
transform -1 0 8740 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_35.mux_l1_in_0__A0
timestamp 1649977179
transform -1 0 7636 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_35.mux_l1_in_0__A1
timestamp 1649977179
transform -1 0 7820 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_37.mux_l1_in_0__A0
timestamp 1649977179
transform 1 0 5704 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_37.mux_l1_in_0__A1
timestamp 1649977179
transform -1 0 6072 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_39.mux_l1_in_0__A0
timestamp 1649977179
transform 1 0 7820 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_39.mux_l1_in_0__A1
timestamp 1649977179
transform -1 0 8188 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_0.mux_l1_in_0__A0
timestamp 1649977179
transform 1 0 4876 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_0.mux_l1_in_0__A1
timestamp 1649977179
transform 1 0 4232 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_0.mux_l1_in_1__A0
timestamp 1649977179
transform 1 0 4048 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_0.mux_l1_in_1__A1
timestamp 1649977179
transform 1 0 4232 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_0.mux_l1_in_2__A0
timestamp 1649977179
transform 1 0 8280 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_0.mux_l1_in_2__A1
timestamp 1649977179
transform 1 0 8740 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_0.mux_l2_in_0__S
timestamp 1649977179
transform -1 0 6532 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_0.mux_l2_in_1__A0
timestamp 1649977179
transform 1 0 11040 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_0.mux_l2_in_1__S
timestamp 1649977179
transform 1 0 10120 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_0.mux_l2_in_2__A0
timestamp 1649977179
transform 1 0 4968 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_0.mux_l2_in_2__A1
timestamp 1649977179
transform 1 0 5152 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_0.mux_l2_in_2__S
timestamp 1649977179
transform -1 0 6532 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_0.mux_l2_in_3__A1
timestamp 1649977179
transform 1 0 4600 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_0.mux_l2_in_3__S
timestamp 1649977179
transform 1 0 5980 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_2.mux_l1_in_0__A0
timestamp 1649977179
transform 1 0 3312 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_2.mux_l1_in_0__A1
timestamp 1649977179
transform 1 0 3496 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_2.mux_l2_in_0__A0
timestamp 1649977179
transform 1 0 4048 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_2.mux_l2_in_1__A0
timestamp 1649977179
transform 1 0 6072 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_2.mux_l2_in_1__A1
timestamp 1649977179
transform -1 0 6072 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_2.mux_l2_in_2__A0
timestamp 1649977179
transform 1 0 7268 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_2.mux_l2_in_2__A1
timestamp 1649977179
transform 1 0 8280 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_2.mux_l2_in_3__A1
timestamp 1649977179
transform 1 0 8740 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_4.mux_l1_in_0__A0
timestamp 1649977179
transform 1 0 4876 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_4.mux_l1_in_0__A1
timestamp 1649977179
transform 1 0 5980 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_4.mux_l1_in_0__S
timestamp 1649977179
transform 1 0 6716 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_4.mux_l1_in_1__A0
timestamp 1649977179
transform 1 0 3772 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_4.mux_l1_in_1__A1
timestamp 1649977179
transform 1 0 3772 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_4.mux_l1_in_1__S
timestamp 1649977179
transform 1 0 4784 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_4.mux_l1_in_2__A0
timestamp 1649977179
transform 1 0 4784 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_4.mux_l1_in_2__A1
timestamp 1649977179
transform 1 0 4968 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_4.mux_l1_in_2__S
timestamp 1649977179
transform 1 0 5980 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_4.mux_l1_in_3__A0
timestamp 1649977179
transform 1 0 3772 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_4.mux_l1_in_3__A1
timestamp 1649977179
transform 1 0 3956 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_4.mux_l1_in_3__S
timestamp 1649977179
transform 1 0 4968 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_4.mux_l1_in_4__A0
timestamp 1649977179
transform 1 0 7360 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_4.mux_l1_in_4__A1
timestamp 1649977179
transform 1 0 8372 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_4.mux_l1_in_4__S
timestamp 1649977179
transform 1 0 8556 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_4.mux_l1_in_5__A0
timestamp 1649977179
transform -1 0 7452 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_4.mux_l1_in_5__A1
timestamp 1649977179
transform 1 0 8464 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_4.mux_l1_in_5__S
timestamp 1649977179
transform 1 0 8556 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_4.mux_l1_in_6__A0
timestamp 1649977179
transform 1 0 3772 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_4.mux_l1_in_6__A1
timestamp 1649977179
transform 1 0 3956 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_4.mux_l1_in_6__S
timestamp 1649977179
transform -1 0 4324 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_8.mux_l1_in_0__A0
timestamp 1649977179
transform 1 0 6532 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_8.mux_l1_in_0__A1
timestamp 1649977179
transform 1 0 6348 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_8.mux_l2_in_0__A0
timestamp 1649977179
transform 1 0 9936 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_8.mux_l2_in_0__S
timestamp 1649977179
transform 1 0 9752 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_8.mux_l2_in_1__A0
timestamp 1649977179
transform -1 0 11684 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_8.mux_l2_in_1__A1
timestamp 1649977179
transform 1 0 9200 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_8.mux_l2_in_1__S
timestamp 1649977179
transform 1 0 10948 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_8.mux_l2_in_2__A0
timestamp 1649977179
transform 1 0 3772 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_8.mux_l2_in_2__A1
timestamp 1649977179
transform 1 0 3588 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_8.mux_l2_in_2__S
timestamp 1649977179
transform -1 0 4324 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_8.mux_l2_in_3__A1
timestamp 1649977179
transform 1 0 4232 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_8.mux_l2_in_3__S
timestamp 1649977179
transform 1 0 5428 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_16.mux_l1_in_0__A0
timestamp 1649977179
transform -1 0 3312 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_16.mux_l1_in_0__A1
timestamp 1649977179
transform 1 0 3312 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_16.mux_l1_in_0__S
timestamp 1649977179
transform 1 0 6072 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_16.mux_l1_in_1__A0
timestamp 1649977179
transform 1 0 10948 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_16.mux_l1_in_1__A1
timestamp 1649977179
transform 1 0 9108 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_16.mux_l1_in_1__S
timestamp 1649977179
transform 1 0 11132 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_16.mux_l1_in_2__A0
timestamp 1649977179
transform 1 0 1656 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_16.mux_l1_in_2__A1
timestamp 1649977179
transform -1 0 1656 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_16.mux_l1_in_2__S
timestamp 1649977179
transform -1 0 3404 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_16.mux_l1_in_3__A1
timestamp 1649977179
transform 1 0 1840 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_16.mux_l1_in_3__S
timestamp 1649977179
transform 1 0 3220 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_24.mux_l1_in_0__A0
timestamp 1649977179
transform 1 0 3496 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_24.mux_l1_in_0__A1
timestamp 1649977179
transform -1 0 2576 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_24.mux_l1_in_0__S
timestamp 1649977179
transform 1 0 3864 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_24.mux_l1_in_1__A0
timestamp 1649977179
transform 1 0 12972 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_24.mux_l1_in_1__A1
timestamp 1649977179
transform 1 0 11316 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_24.mux_l1_in_1__S
timestamp 1649977179
transform 1 0 12328 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_24.mux_l1_in_2__A0
timestamp 1649977179
transform 1 0 1472 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_24.mux_l1_in_2__A1
timestamp 1649977179
transform 1 0 1472 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_24.mux_l1_in_2__S
timestamp 1649977179
transform -1 0 3312 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_24.mux_l1_in_3__A1
timestamp 1649977179
transform 1 0 3220 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_24.mux_l1_in_3__S
timestamp 1649977179
transform 1 0 3956 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_32.mux_l1_in_0__A0
timestamp 1649977179
transform -1 0 4692 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_32.mux_l1_in_0__A1
timestamp 1649977179
transform 1 0 4692 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_32.mux_l1_in_1__A0
timestamp 1649977179
transform 1 0 7176 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_32.mux_l1_in_1__A1
timestamp 1649977179
transform 1 0 8096 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_32.mux_l1_in_2__A0
timestamp 1649977179
transform 1 0 5888 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_32.mux_l1_in_2__A1
timestamp 1649977179
transform 1 0 5704 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_prog_clk_0_FTB00_A
timestamp 1649977179
transform -1 0 20424 0 -1 20672
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3 dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform 1 0 1380 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_15
timestamp 1649977179
transform 1 0 2484 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_27 dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform 1 0 3588 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_29 dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform 1 0 3772 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_37
timestamp 1649977179
transform 1 0 4508 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_53 dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform 1 0 5980 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_0_57 dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform 1 0 6348 0 1 2176
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_67
timestamp 1649977179
transform 1 0 7268 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_79
timestamp 1649977179
transform 1 0 8372 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_98 dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform 1 0 10120 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_102
timestamp 1649977179
transform 1 0 10488 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_107
timestamp 1649977179
transform 1 0 10948 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_111
timestamp 1649977179
transform 1 0 11316 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_113 dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform 1 0 11500 0 1 2176
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_117
timestamp 1649977179
transform 1 0 11868 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_129
timestamp 1649977179
transform 1 0 12972 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_137
timestamp 1649977179
transform 1 0 13708 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_147
timestamp 1649977179
transform 1 0 14628 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_151
timestamp 1649977179
transform 1 0 14996 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_0_159
timestamp 1649977179
transform 1 0 15732 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_163
timestamp 1649977179
transform 1 0 16100 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_167
timestamp 1649977179
transform 1 0 16468 0 1 2176
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_169
timestamp 1649977179
transform 1 0 16652 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_181
timestamp 1649977179
transform 1 0 17756 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_185
timestamp 1649977179
transform 1 0 18124 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_194
timestamp 1649977179
transform 1 0 18952 0 1 2176
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_197
timestamp 1649977179
transform 1 0 19228 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_209
timestamp 1649977179
transform 1 0 20332 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_221
timestamp 1649977179
transform 1 0 21436 0 1 2176
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_1_3
timestamp 1649977179
transform 1 0 1380 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_15
timestamp 1649977179
transform 1 0 2484 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_27
timestamp 1649977179
transform 1 0 3588 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_1_48
timestamp 1649977179
transform 1 0 5520 0 -1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_1_66
timestamp 1649977179
transform 1 0 7176 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_1_78
timestamp 1649977179
transform 1 0 8280 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_1_130
timestamp 1649977179
transform 1 0 13064 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_1_167
timestamp 1649977179
transform 1 0 16468 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_1_177
timestamp 1649977179
transform 1 0 17388 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_1_181
timestamp 1649977179
transform 1 0 17756 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_1_216
timestamp 1649977179
transform 1 0 20976 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_1_222
timestamp 1649977179
transform 1 0 21528 0 -1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_2_3
timestamp 1649977179
transform 1 0 1380 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_15
timestamp 1649977179
transform 1 0 2484 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_2_27
timestamp 1649977179
transform 1 0 3588 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_2_29
timestamp 1649977179
transform 1 0 3772 0 1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_2_67
timestamp 1649977179
transform 1 0 7268 0 1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_2_77
timestamp 1649977179
transform 1 0 8188 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_2_83
timestamp 1649977179
transform 1 0 8740 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_2_94
timestamp 1649977179
transform 1 0 9752 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_2_111
timestamp 1649977179
transform 1 0 11316 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_2_123
timestamp 1649977179
transform 1 0 12420 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_2_138
timestamp 1649977179
transform 1 0 13800 0 1 3264
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_2_141
timestamp 1649977179
transform 1 0 14076 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_153
timestamp 1649977179
transform 1 0 15180 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_2_165
timestamp 1649977179
transform 1 0 16284 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_2_169
timestamp 1649977179
transform 1 0 16652 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_2_179
timestamp 1649977179
transform 1 0 17572 0 1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_2_187
timestamp 1649977179
transform 1 0 18308 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_2_192
timestamp 1649977179
transform 1 0 18768 0 1 3264
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_2_197
timestamp 1649977179
transform 1 0 19228 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_209
timestamp 1649977179
transform 1 0 20332 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_2_221
timestamp 1649977179
transform 1 0 21436 0 1 3264
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_3_3
timestamp 1649977179
transform 1 0 1380 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_15
timestamp 1649977179
transform 1 0 2484 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_27
timestamp 1649977179
transform 1 0 3588 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_3_39
timestamp 1649977179
transform 1 0 4692 0 -1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_3_60
timestamp 1649977179
transform 1 0 6624 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_3_88
timestamp 1649977179
transform 1 0 9200 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_3_111
timestamp 1649977179
transform 1 0 11316 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_3_124
timestamp 1649977179
transform 1 0 12512 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_3_136
timestamp 1649977179
transform 1 0 13616 0 -1 4352
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_3_150
timestamp 1649977179
transform 1 0 14904 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_3_162
timestamp 1649977179
transform 1 0 16008 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_3_167
timestamp 1649977179
transform 1 0 16468 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_3_178
timestamp 1649977179
transform 1 0 17480 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_3_188
timestamp 1649977179
transform 1 0 18400 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_200
timestamp 1649977179
transform 1 0 19504 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_3_212
timestamp 1649977179
transform 1 0 20608 0 -1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_3_220
timestamp 1649977179
transform 1 0 21344 0 -1 4352
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_4_3
timestamp 1649977179
transform 1 0 1380 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_15
timestamp 1649977179
transform 1 0 2484 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_4_27
timestamp 1649977179
transform 1 0 3588 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_4_29
timestamp 1649977179
transform 1 0 3772 0 1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_4_37
timestamp 1649977179
transform 1 0 4508 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_4_42
timestamp 1649977179
transform 1 0 4968 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_4_67
timestamp 1649977179
transform 1 0 7268 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_4_83
timestamp 1649977179
transform 1 0 8740 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_4_85
timestamp 1649977179
transform 1 0 8924 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_4_89
timestamp 1649977179
transform 1 0 9292 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_4_105
timestamp 1649977179
transform 1 0 10764 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_4_113
timestamp 1649977179
transform 1 0 11500 0 1 4352
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_4_123
timestamp 1649977179
transform 1 0 12420 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_4_135
timestamp 1649977179
transform 1 0 13524 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_4_139
timestamp 1649977179
transform 1 0 13892 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_4_141
timestamp 1649977179
transform 1 0 14076 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_4_153
timestamp 1649977179
transform 1 0 15180 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_4_167
timestamp 1649977179
transform 1 0 16468 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_4_185
timestamp 1649977179
transform 1 0 18124 0 1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_4_193
timestamp 1649977179
transform 1 0 18860 0 1 4352
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_4_203
timestamp 1649977179
transform 1 0 19780 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_4_215
timestamp 1649977179
transform 1 0 20884 0 1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_5_3
timestamp 1649977179
transform 1 0 1380 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_5_20
timestamp 1649977179
transform 1 0 2944 0 -1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_5_28
timestamp 1649977179
transform 1 0 3680 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_5_66
timestamp 1649977179
transform 1 0 7176 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_5_110
timestamp 1649977179
transform 1 0 11224 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_5_113
timestamp 1649977179
transform 1 0 11500 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_5_140
timestamp 1649977179
transform 1 0 13984 0 -1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_5_148
timestamp 1649977179
transform 1 0 14720 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_5_166
timestamp 1649977179
transform 1 0 16376 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_5_169
timestamp 1649977179
transform 1 0 16652 0 -1 5440
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_5_176
timestamp 1649977179
transform 1 0 17296 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_188
timestamp 1649977179
transform 1 0 18400 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_200
timestamp 1649977179
transform 1 0 19504 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_5_218
timestamp 1649977179
transform 1 0 21160 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_5_222
timestamp 1649977179
transform 1 0 21528 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_6_5
timestamp 1649977179
transform 1 0 1564 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_6_17
timestamp 1649977179
transform 1 0 2668 0 1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_6_25
timestamp 1649977179
transform 1 0 3404 0 1 5440
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_6_29
timestamp 1649977179
transform 1 0 3772 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_6_67
timestamp 1649977179
transform 1 0 7268 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_6_74
timestamp 1649977179
transform 1 0 7912 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_6_96
timestamp 1649977179
transform 1 0 9936 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_6_100
timestamp 1649977179
transform 1 0 10304 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_6_110
timestamp 1649977179
transform 1 0 11224 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_6_121
timestamp 1649977179
transform 1 0 12236 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_6_139
timestamp 1649977179
transform 1 0 13892 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_6_141
timestamp 1649977179
transform 1 0 14076 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_153
timestamp 1649977179
transform 1 0 15180 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_6_165
timestamp 1649977179
transform 1 0 16284 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_6_186
timestamp 1649977179
transform 1 0 18216 0 1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_6_194
timestamp 1649977179
transform 1 0 18952 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_6_197
timestamp 1649977179
transform 1 0 19228 0 1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_6_214
timestamp 1649977179
transform 1 0 20792 0 1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_6_222
timestamp 1649977179
transform 1 0 21528 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_7_3
timestamp 1649977179
transform 1 0 1380 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_7_15
timestamp 1649977179
transform 1 0 2484 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_7_27
timestamp 1649977179
transform 1 0 3588 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_7_53
timestamp 1649977179
transform 1 0 5980 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_7_59
timestamp 1649977179
transform 1 0 6532 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_7_92
timestamp 1649977179
transform 1 0 9568 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_7_102
timestamp 1649977179
transform 1 0 10488 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_7_118
timestamp 1649977179
transform 1 0 11960 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_7_130
timestamp 1649977179
transform 1 0 13064 0 -1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_7_138
timestamp 1649977179
transform 1 0 13800 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_7_148
timestamp 1649977179
transform 1 0 14720 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_7_160
timestamp 1649977179
transform 1 0 15824 0 -1 6528
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_7_169
timestamp 1649977179
transform 1 0 16652 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_181
timestamp 1649977179
transform 1 0 17756 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_193
timestamp 1649977179
transform 1 0 18860 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_205
timestamp 1649977179
transform 1 0 19964 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_7_217
timestamp 1649977179
transform 1 0 21068 0 -1 6528
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_8_3
timestamp 1649977179
transform 1 0 1380 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_8_15
timestamp 1649977179
transform 1 0 2484 0 1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_8_23
timestamp 1649977179
transform 1 0 3220 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_8_29
timestamp 1649977179
transform 1 0 3772 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_8_41
timestamp 1649977179
transform 1 0 4876 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_49
timestamp 1649977179
transform 1 0 5612 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_8_80
timestamp 1649977179
transform 1 0 8464 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_8_83
timestamp 1649977179
transform 1 0 8740 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_8_107
timestamp 1649977179
transform 1 0 10948 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_113
timestamp 1649977179
transform 1 0 11500 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_8_125
timestamp 1649977179
transform 1 0 12604 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_8_137
timestamp 1649977179
transform 1 0 13708 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_8_152
timestamp 1649977179
transform 1 0 15088 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_164
timestamp 1649977179
transform 1 0 16192 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_176
timestamp 1649977179
transform 1 0 17296 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_8_188
timestamp 1649977179
transform 1 0 18400 0 1 6528
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_8_197
timestamp 1649977179
transform 1 0 19228 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_209
timestamp 1649977179
transform 1 0 20332 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_8_221
timestamp 1649977179
transform 1 0 21436 0 1 6528
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_9_7
timestamp 1649977179
transform 1 0 1748 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_19
timestamp 1649977179
transform 1 0 2852 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_9_31
timestamp 1649977179
transform 1 0 3956 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_9_57
timestamp 1649977179
transform 1 0 6348 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_9_79
timestamp 1649977179
transform 1 0 8372 0 -1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_9_98
timestamp 1649977179
transform 1 0 10120 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_9_111
timestamp 1649977179
transform 1 0 11316 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_9_116
timestamp 1649977179
transform 1 0 11776 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_9_131
timestamp 1649977179
transform 1 0 13156 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_9_161
timestamp 1649977179
transform 1 0 15916 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_9_167
timestamp 1649977179
transform 1 0 16468 0 -1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_9_169
timestamp 1649977179
transform 1 0 16652 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_181
timestamp 1649977179
transform 1 0 17756 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_9_193
timestamp 1649977179
transform 1 0 18860 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_9_197
timestamp 1649977179
transform 1 0 19228 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_9_216
timestamp 1649977179
transform 1 0 20976 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_9_222
timestamp 1649977179
transform 1 0 21528 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_10_3
timestamp 1649977179
transform 1 0 1380 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_10_6
timestamp 1649977179
transform 1 0 1656 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_10_26
timestamp 1649977179
transform 1 0 3496 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_10_29
timestamp 1649977179
transform 1 0 3772 0 1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_10_37
timestamp 1649977179
transform 1 0 4508 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_10_69
timestamp 1649977179
transform 1 0 7452 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_10_72
timestamp 1649977179
transform 1 0 7728 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_10_85
timestamp 1649977179
transform 1 0 8924 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_10_98
timestamp 1649977179
transform 1 0 10120 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_10_102
timestamp 1649977179
transform 1 0 10488 0 1 7616
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_10_126
timestamp 1649977179
transform 1 0 12696 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_10_138
timestamp 1649977179
transform 1 0 13800 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_10_146
timestamp 1649977179
transform 1 0 14536 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_10_150
timestamp 1649977179
transform 1 0 14904 0 1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_10_171
timestamp 1649977179
transform 1 0 16836 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_10_177
timestamp 1649977179
transform 1 0 17388 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_10_191
timestamp 1649977179
transform 1 0 18676 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_10_195
timestamp 1649977179
transform 1 0 19044 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_10_197
timestamp 1649977179
transform 1 0 19228 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_10_201
timestamp 1649977179
transform 1 0 19596 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_10_222
timestamp 1649977179
transform 1 0 21528 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_11_3
timestamp 1649977179
transform 1 0 1380 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_11_25
timestamp 1649977179
transform 1 0 3404 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_11_44
timestamp 1649977179
transform 1 0 5152 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_11_111
timestamp 1649977179
transform 1 0 11316 0 -1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_11_116
timestamp 1649977179
transform 1 0 11776 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_11_128
timestamp 1649977179
transform 1 0 12880 0 -1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_11_136
timestamp 1649977179
transform 1 0 13616 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_11_139
timestamp 1649977179
transform 1 0 13892 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_11_161
timestamp 1649977179
transform 1 0 15916 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_11_167
timestamp 1649977179
transform 1 0 16468 0 -1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_11_169
timestamp 1649977179
transform 1 0 16652 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_11_181
timestamp 1649977179
transform 1 0 17756 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_11_217
timestamp 1649977179
transform 1 0 21068 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_12_3
timestamp 1649977179
transform 1 0 1380 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_12_27
timestamp 1649977179
transform 1 0 3588 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_12_29
timestamp 1649977179
transform 1 0 3772 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_12_36
timestamp 1649977179
transform 1 0 4416 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_12_85
timestamp 1649977179
transform 1 0 8924 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_12_120
timestamp 1649977179
transform 1 0 12144 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_12_139
timestamp 1649977179
transform 1 0 13892 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_12_183
timestamp 1649977179
transform 1 0 17940 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_12_187
timestamp 1649977179
transform 1 0 18308 0 1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_12_195
timestamp 1649977179
transform 1 0 19044 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_12_215
timestamp 1649977179
transform 1 0 20884 0 1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_13_3
timestamp 1649977179
transform 1 0 1380 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_13_12
timestamp 1649977179
transform 1 0 2208 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_13_25
timestamp 1649977179
transform 1 0 3404 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_13_46
timestamp 1649977179
transform 1 0 5336 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_13_49
timestamp 1649977179
transform 1 0 5612 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_13_68
timestamp 1649977179
transform 1 0 7360 0 -1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_13_78
timestamp 1649977179
transform 1 0 8280 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_13_113
timestamp 1649977179
transform 1 0 11500 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_13_117
timestamp 1649977179
transform 1 0 11868 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_13_221
timestamp 1649977179
transform 1 0 21436 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_14_3
timestamp 1649977179
transform 1 0 1380 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_14_7
timestamp 1649977179
transform 1 0 1748 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_14_80
timestamp 1649977179
transform 1 0 8464 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_14_97
timestamp 1649977179
transform 1 0 10028 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_14_102
timestamp 1649977179
transform 1 0 10488 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_14_139
timestamp 1649977179
transform 1 0 13892 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_14_141
timestamp 1649977179
transform 1 0 14076 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_14_197
timestamp 1649977179
transform 1 0 19228 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_14_218
timestamp 1649977179
transform 1 0 21160 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_14_222
timestamp 1649977179
transform 1 0 21528 0 1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_15_3
timestamp 1649977179
transform 1 0 1380 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_15_15
timestamp 1649977179
transform 1 0 2484 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_15_19
timestamp 1649977179
transform 1 0 2852 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_15_23
timestamp 1649977179
transform 1 0 3220 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_15_55
timestamp 1649977179
transform 1 0 6164 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_15_66
timestamp 1649977179
transform 1 0 7176 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_15_96
timestamp 1649977179
transform 1 0 9936 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_15_111
timestamp 1649977179
transform 1 0 11316 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_15_149
timestamp 1649977179
transform 1 0 14812 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_15_189
timestamp 1649977179
transform 1 0 18492 0 -1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_15_197
timestamp 1649977179
transform 1 0 19228 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_15_217
timestamp 1649977179
transform 1 0 21068 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_16_3
timestamp 1649977179
transform 1 0 1380 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_16_7
timestamp 1649977179
transform 1 0 1748 0 1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_16_16
timestamp 1649977179
transform 1 0 2576 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_16_29
timestamp 1649977179
transform 1 0 3772 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_16_33
timestamp 1649977179
transform 1 0 4140 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_16_70
timestamp 1649977179
transform 1 0 7544 0 1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_16_78
timestamp 1649977179
transform 1 0 8280 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_16_94
timestamp 1649977179
transform 1 0 9752 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_16_106
timestamp 1649977179
transform 1 0 10856 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_16_137
timestamp 1649977179
transform 1 0 13708 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_16_141
timestamp 1649977179
transform 1 0 14076 0 1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_16_149
timestamp 1649977179
transform 1 0 14812 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_16_186
timestamp 1649977179
transform 1 0 18216 0 1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_16_194
timestamp 1649977179
transform 1 0 18952 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_16_197
timestamp 1649977179
transform 1 0 19228 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_16_219
timestamp 1649977179
transform 1 0 21252 0 1 10880
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_17_3
timestamp 1649977179
transform 1 0 1380 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_15
timestamp 1649977179
transform 1 0 2484 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_17_27
timestamp 1649977179
transform 1 0 3588 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_17_37
timestamp 1649977179
transform 1 0 4508 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_17_43
timestamp 1649977179
transform 1 0 5060 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_17_49
timestamp 1649977179
transform 1 0 5612 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_17_68
timestamp 1649977179
transform 1 0 7360 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_17_82
timestamp 1649977179
transform 1 0 8648 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_17_88
timestamp 1649977179
transform 1 0 9200 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_17_107
timestamp 1649977179
transform 1 0 10948 0 -1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_17_142
timestamp 1649977179
transform 1 0 14168 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_154
timestamp 1649977179
transform 1 0 15272 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_17_169
timestamp 1649977179
transform 1 0 16652 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_17_172
timestamp 1649977179
transform 1 0 16928 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_17_196
timestamp 1649977179
transform 1 0 19136 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_17_216
timestamp 1649977179
transform 1 0 20976 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_17_222
timestamp 1649977179
transform 1 0 21528 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_18_3
timestamp 1649977179
transform 1 0 1380 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_18_7
timestamp 1649977179
transform 1 0 1748 0 1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_18_12
timestamp 1649977179
transform 1 0 2208 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_18_24
timestamp 1649977179
transform 1 0 3312 0 1 11968
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_18_29
timestamp 1649977179
transform 1 0 3772 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_18_47
timestamp 1649977179
transform 1 0 5428 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_18_58
timestamp 1649977179
transform 1 0 6440 0 1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_18_66
timestamp 1649977179
transform 1 0 7176 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_18_78
timestamp 1649977179
transform 1 0 8280 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_18_83
timestamp 1649977179
transform 1 0 8740 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_18_97
timestamp 1649977179
transform 1 0 10028 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_18_141
timestamp 1649977179
transform 1 0 14076 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_18_146
timestamp 1649977179
transform 1 0 14536 0 1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_18_190
timestamp 1649977179
transform 1 0 18584 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_18_197
timestamp 1649977179
transform 1 0 19228 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_18_221
timestamp 1649977179
transform 1 0 21436 0 1 11968
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_19_3
timestamp 1649977179
transform 1 0 1380 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_19_15
timestamp 1649977179
transform 1 0 2484 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_19_21
timestamp 1649977179
transform 1 0 3036 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_19_28
timestamp 1649977179
transform 1 0 3680 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_19_80
timestamp 1649977179
transform 1 0 8464 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_19_90
timestamp 1649977179
transform 1 0 9384 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_19_105
timestamp 1649977179
transform 1 0 10764 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_19_111
timestamp 1649977179
transform 1 0 11316 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_19_113
timestamp 1649977179
transform 1 0 11500 0 -1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_19_121
timestamp 1649977179
transform 1 0 12236 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_19_160
timestamp 1649977179
transform 1 0 15824 0 -1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_19_219
timestamp 1649977179
transform 1 0 21252 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_19_222
timestamp 1649977179
transform 1 0 21528 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_20_3
timestamp 1649977179
transform 1 0 1380 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_20_7
timestamp 1649977179
transform 1 0 1748 0 1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_20_12
timestamp 1649977179
transform 1 0 2208 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_20_24
timestamp 1649977179
transform 1 0 3312 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_20_29
timestamp 1649977179
transform 1 0 3772 0 1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_20_43
timestamp 1649977179
transform 1 0 5060 0 1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_20_51
timestamp 1649977179
transform 1 0 5796 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_20_85
timestamp 1649977179
transform 1 0 8924 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_20_89
timestamp 1649977179
transform 1 0 9292 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_20_117
timestamp 1649977179
transform 1 0 11868 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_20_123
timestamp 1649977179
transform 1 0 12420 0 1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_20_143
timestamp 1649977179
transform 1 0 14260 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_20_155
timestamp 1649977179
transform 1 0 15364 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_20_181
timestamp 1649977179
transform 1 0 17756 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_20_187
timestamp 1649977179
transform 1 0 18308 0 1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_20_195
timestamp 1649977179
transform 1 0 19044 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_20_197
timestamp 1649977179
transform 1 0 19228 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_20_203
timestamp 1649977179
transform 1 0 19780 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_20_220
timestamp 1649977179
transform 1 0 21344 0 1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_21_3
timestamp 1649977179
transform 1 0 1380 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_15
timestamp 1649977179
transform 1 0 2484 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_21_27
timestamp 1649977179
transform 1 0 3588 0 -1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_21_35
timestamp 1649977179
transform 1 0 4324 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_21_39
timestamp 1649977179
transform 1 0 4692 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_21_51
timestamp 1649977179
transform 1 0 5796 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_21_66
timestamp 1649977179
transform 1 0 7176 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_21_76
timestamp 1649977179
transform 1 0 8096 0 -1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_21_84
timestamp 1649977179
transform 1 0 8832 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_21_111
timestamp 1649977179
transform 1 0 11316 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_21_113
timestamp 1649977179
transform 1 0 11500 0 -1 14144
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_21_139
timestamp 1649977179
transform 1 0 13892 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_21_151
timestamp 1649977179
transform 1 0 14996 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_21_203
timestamp 1649977179
transform 1 0 19780 0 -1 14144
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_22_3
timestamp 1649977179
transform 1 0 1380 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_22_15
timestamp 1649977179
transform 1 0 2484 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_22_21
timestamp 1649977179
transform 1 0 3036 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_22_29
timestamp 1649977179
transform 1 0 3772 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_22_50
timestamp 1649977179
transform 1 0 5704 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_22_61
timestamp 1649977179
transform 1 0 6716 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_22_67
timestamp 1649977179
transform 1 0 7268 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_22_83
timestamp 1649977179
transform 1 0 8740 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_22_85
timestamp 1649977179
transform 1 0 8924 0 1 14144
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_22_105
timestamp 1649977179
transform 1 0 10764 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_22_117
timestamp 1649977179
transform 1 0 11868 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_22_138
timestamp 1649977179
transform 1 0 13800 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_22_141
timestamp 1649977179
transform 1 0 14076 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_22_163
timestamp 1649977179
transform 1 0 16100 0 1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_22_182
timestamp 1649977179
transform 1 0 17848 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_22_194
timestamp 1649977179
transform 1 0 18952 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_22_197
timestamp 1649977179
transform 1 0 19228 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_22_201
timestamp 1649977179
transform 1 0 19596 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_22_220
timestamp 1649977179
transform 1 0 21344 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_23_3
timestamp 1649977179
transform 1 0 1380 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_23_7
timestamp 1649977179
transform 1 0 1748 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_23_12
timestamp 1649977179
transform 1 0 2208 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_23_57
timestamp 1649977179
transform 1 0 6348 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_23_70
timestamp 1649977179
transform 1 0 7544 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_23_100
timestamp 1649977179
transform 1 0 10304 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_23_115
timestamp 1649977179
transform 1 0 11684 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_23_137
timestamp 1649977179
transform 1 0 13708 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_23_157
timestamp 1649977179
transform 1 0 15548 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  FILLER_23_165
timestamp 1649977179
transform 1 0 16284 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_23_187
timestamp 1649977179
transform 1 0 18308 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_24_3
timestamp 1649977179
transform 1 0 1380 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_24_7
timestamp 1649977179
transform 1 0 1748 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_24_20
timestamp 1649977179
transform 1 0 2944 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_24_29
timestamp 1649977179
transform 1 0 3772 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_24_63
timestamp 1649977179
transform 1 0 6900 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_24_80
timestamp 1649977179
transform 1 0 8464 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_24_98
timestamp 1649977179
transform 1 0 10120 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_24_110
timestamp 1649977179
transform 1 0 11224 0 1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_24_136
timestamp 1649977179
transform 1 0 13616 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_24_161
timestamp 1649977179
transform 1 0 15916 0 1 15232
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_24_181
timestamp 1649977179
transform 1 0 17756 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_24_193
timestamp 1649977179
transform 1 0 18860 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_24_197
timestamp 1649977179
transform 1 0 19228 0 1 15232
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_25_3
timestamp 1649977179
transform 1 0 1380 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_25_15
timestamp 1649977179
transform 1 0 2484 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_25_31
timestamp 1649977179
transform 1 0 3956 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_25_36
timestamp 1649977179
transform 1 0 4416 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_25_40
timestamp 1649977179
transform 1 0 4784 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_25_55
timestamp 1649977179
transform 1 0 6164 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_25_68
timestamp 1649977179
transform 1 0 7360 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_25_80
timestamp 1649977179
transform 1 0 8464 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_25_85
timestamp 1649977179
transform 1 0 8924 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_25_115
timestamp 1649977179
transform 1 0 11684 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_25_119
timestamp 1649977179
transform 1 0 12052 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_25_158
timestamp 1649977179
transform 1 0 15640 0 -1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_25_166
timestamp 1649977179
transform 1 0 16376 0 -1 16320
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_25_169
timestamp 1649977179
transform 1 0 16652 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_25_181
timestamp 1649977179
transform 1 0 17756 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_25_200
timestamp 1649977179
transform 1 0 19504 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_25_222
timestamp 1649977179
transform 1 0 21528 0 -1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_26_3
timestamp 1649977179
transform 1 0 1380 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_26_15
timestamp 1649977179
transform 1 0 2484 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_26_42
timestamp 1649977179
transform 1 0 4968 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_26_61
timestamp 1649977179
transform 1 0 6716 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_26_83
timestamp 1649977179
transform 1 0 8740 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_26_85
timestamp 1649977179
transform 1 0 8924 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_26_115
timestamp 1649977179
transform 1 0 11684 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_26_137
timestamp 1649977179
transform 1 0 13708 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_26_141
timestamp 1649977179
transform 1 0 14076 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_26_164
timestamp 1649977179
transform 1 0 16192 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_26_170
timestamp 1649977179
transform 1 0 16744 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_26_189
timestamp 1649977179
transform 1 0 18492 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_26_195
timestamp 1649977179
transform 1 0 19044 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_26_215
timestamp 1649977179
transform 1 0 20884 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_27_3
timestamp 1649977179
transform 1 0 1380 0 -1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_27_55
timestamp 1649977179
transform 1 0 6164 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_27_57
timestamp 1649977179
transform 1 0 6348 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_27_69
timestamp 1649977179
transform 1 0 7452 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_27_109
timestamp 1649977179
transform 1 0 11132 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_27_147
timestamp 1649977179
transform 1 0 14628 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_27_151
timestamp 1649977179
transform 1 0 14996 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_27_187
timestamp 1649977179
transform 1 0 18308 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_27_193
timestamp 1649977179
transform 1 0 18860 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_27_212
timestamp 1649977179
transform 1 0 20608 0 -1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_27_220
timestamp 1649977179
transform 1 0 21344 0 -1 17408
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_28_3
timestamp 1649977179
transform 1 0 1380 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_28_15
timestamp 1649977179
transform 1 0 2484 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_28_21
timestamp 1649977179
transform 1 0 3036 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_28_27
timestamp 1649977179
transform 1 0 3588 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_28_31
timestamp 1649977179
transform 1 0 3956 0 1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_28_39
timestamp 1649977179
transform 1 0 4692 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_28_63
timestamp 1649977179
transform 1 0 6900 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_28_69
timestamp 1649977179
transform 1 0 7452 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_28_82
timestamp 1649977179
transform 1 0 8648 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_28_85
timestamp 1649977179
transform 1 0 8924 0 1 17408
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_28_98
timestamp 1649977179
transform 1 0 10120 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_28_110
timestamp 1649977179
transform 1 0 11224 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_28_114
timestamp 1649977179
transform 1 0 11592 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_28_137
timestamp 1649977179
transform 1 0 13708 0 1 17408
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_28_141
timestamp 1649977179
transform 1 0 14076 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_153
timestamp 1649977179
transform 1 0 15180 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_28_165
timestamp 1649977179
transform 1 0 16284 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_28_187
timestamp 1649977179
transform 1 0 18308 0 1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_28_195
timestamp 1649977179
transform 1 0 19044 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_28_197
timestamp 1649977179
transform 1 0 19228 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_28_221
timestamp 1649977179
transform 1 0 21436 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_29_3
timestamp 1649977179
transform 1 0 1380 0 -1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_29_9
timestamp 1649977179
transform 1 0 1932 0 -1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_29_14
timestamp 1649977179
transform 1 0 2392 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_26
timestamp 1649977179
transform 1 0 3496 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_29_38
timestamp 1649977179
transform 1 0 4600 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_29_55
timestamp 1649977179
transform 1 0 6164 0 -1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_29_57
timestamp 1649977179
transform 1 0 6348 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_29_69
timestamp 1649977179
transform 1 0 7452 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_29_86
timestamp 1649977179
transform 1 0 9016 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_29_100
timestamp 1649977179
transform 1 0 10304 0 -1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_29_108
timestamp 1649977179
transform 1 0 11040 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_29_129
timestamp 1649977179
transform 1 0 12972 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_29_148
timestamp 1649977179
transform 1 0 14720 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_29_219
timestamp 1649977179
transform 1 0 21252 0 -1 18496
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_30_3
timestamp 1649977179
transform 1 0 1380 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_15
timestamp 1649977179
transform 1 0 2484 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_30_27
timestamp 1649977179
transform 1 0 3588 0 1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_30_29
timestamp 1649977179
transform 1 0 3772 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_41
timestamp 1649977179
transform 1 0 4876 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_53
timestamp 1649977179
transform 1 0 5980 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_30_65
timestamp 1649977179
transform 1 0 7084 0 1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_30_73
timestamp 1649977179
transform 1 0 7820 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_30_87
timestamp 1649977179
transform 1 0 9108 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_30_94
timestamp 1649977179
transform 1 0 9752 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_30_139
timestamp 1649977179
transform 1 0 13892 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_30_141
timestamp 1649977179
transform 1 0 14076 0 1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_30_147
timestamp 1649977179
transform 1 0 14628 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_30_166
timestamp 1649977179
transform 1 0 16376 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_30_188
timestamp 1649977179
transform 1 0 18400 0 1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_30_197
timestamp 1649977179
transform 1 0 19228 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_30_218
timestamp 1649977179
transform 1 0 21160 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_30_222
timestamp 1649977179
transform 1 0 21528 0 1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_31_3
timestamp 1649977179
transform 1 0 1380 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_15
timestamp 1649977179
transform 1 0 2484 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_27
timestamp 1649977179
transform 1 0 3588 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_39
timestamp 1649977179
transform 1 0 4692 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_31_51
timestamp 1649977179
transform 1 0 5796 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_31_55
timestamp 1649977179
transform 1 0 6164 0 -1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_31_57
timestamp 1649977179
transform 1 0 6348 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_31_69
timestamp 1649977179
transform 1 0 7452 0 -1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_31_75
timestamp 1649977179
transform 1 0 8004 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_31_92
timestamp 1649977179
transform 1 0 9568 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_31_101
timestamp 1649977179
transform 1 0 10396 0 -1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_31_109
timestamp 1649977179
transform 1 0 11132 0 -1 19584
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_31_147
timestamp 1649977179
transform 1 0 14628 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_31_159
timestamp 1649977179
transform 1 0 15732 0 -1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_31_167
timestamp 1649977179
transform 1 0 16468 0 -1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_31_169
timestamp 1649977179
transform 1 0 16652 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_181
timestamp 1649977179
transform 1 0 17756 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_31_193
timestamp 1649977179
transform 1 0 18860 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_31_197
timestamp 1649977179
transform 1 0 19228 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_31_216
timestamp 1649977179
transform 1 0 20976 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_31_220
timestamp 1649977179
transform 1 0 21344 0 -1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_32_3
timestamp 1649977179
transform 1 0 1380 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_32_15
timestamp 1649977179
transform 1 0 2484 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_32_21
timestamp 1649977179
transform 1 0 3036 0 1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_32_27
timestamp 1649977179
transform 1 0 3588 0 1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_32_29
timestamp 1649977179
transform 1 0 3772 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_41
timestamp 1649977179
transform 1 0 4876 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_32_53
timestamp 1649977179
transform 1 0 5980 0 1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_32_61
timestamp 1649977179
transform 1 0 6716 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_32_107
timestamp 1649977179
transform 1 0 10948 0 1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_32_113
timestamp 1649977179
transform 1 0 11500 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_32_134
timestamp 1649977179
transform 1 0 13432 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_32_139
timestamp 1649977179
transform 1 0 13892 0 1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_32_149
timestamp 1649977179
transform 1 0 14812 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_32_161
timestamp 1649977179
transform 1 0 15916 0 1 19584
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_32_169
timestamp 1649977179
transform 1 0 16652 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_181
timestamp 1649977179
transform 1 0 17756 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_32_193
timestamp 1649977179
transform 1 0 18860 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_32_197
timestamp 1649977179
transform 1 0 19228 0 1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_32_205
timestamp 1649977179
transform 1 0 19964 0 1 19584
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_33_3
timestamp 1649977179
transform 1 0 1380 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_15
timestamp 1649977179
transform 1 0 2484 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_33_27
timestamp 1649977179
transform 1 0 3588 0 -1 20672
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_33_29
timestamp 1649977179
transform 1 0 3772 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_41
timestamp 1649977179
transform 1 0 4876 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_33_53
timestamp 1649977179
transform 1 0 5980 0 -1 20672
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_33_57
timestamp 1649977179
transform 1 0 6348 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_33_69
timestamp 1649977179
transform 1 0 7452 0 -1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_33_77
timestamp 1649977179
transform 1 0 8188 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_33_80
timestamp 1649977179
transform 1 0 8464 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_33_85
timestamp 1649977179
transform 1 0 8924 0 -1 20672
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_33_97
timestamp 1649977179
transform 1 0 10028 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_33_109
timestamp 1649977179
transform 1 0 11132 0 -1 20672
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_33_113
timestamp 1649977179
transform 1 0 11500 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_125
timestamp 1649977179
transform 1 0 12604 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_33_137
timestamp 1649977179
transform 1 0 13708 0 -1 20672
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_33_141
timestamp 1649977179
transform 1 0 14076 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_153
timestamp 1649977179
transform 1 0 15180 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_33_165
timestamp 1649977179
transform 1 0 16284 0 -1 20672
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_33_169
timestamp 1649977179
transform 1 0 16652 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_181
timestamp 1649977179
transform 1 0 17756 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_33_193
timestamp 1649977179
transform 1 0 18860 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_33_197
timestamp 1649977179
transform 1 0 19228 0 -1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_33_205
timestamp 1649977179
transform 1 0 19964 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_33_222
timestamp 1649977179
transform 1 0 21528 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_0
timestamp 1649977179
transform 1 0 1104 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_1
timestamp 1649977179
transform -1 0 21896 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_2
timestamp 1649977179
transform 1 0 1104 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_3
timestamp 1649977179
transform -1 0 21896 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_4
timestamp 1649977179
transform 1 0 1104 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_5
timestamp 1649977179
transform -1 0 21896 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_6
timestamp 1649977179
transform 1 0 1104 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_7
timestamp 1649977179
transform -1 0 21896 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_8
timestamp 1649977179
transform 1 0 1104 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_9
timestamp 1649977179
transform -1 0 21896 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_10
timestamp 1649977179
transform 1 0 1104 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_11
timestamp 1649977179
transform -1 0 21896 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_12
timestamp 1649977179
transform 1 0 1104 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_13
timestamp 1649977179
transform -1 0 21896 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_14
timestamp 1649977179
transform 1 0 1104 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_15
timestamp 1649977179
transform -1 0 21896 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_16
timestamp 1649977179
transform 1 0 1104 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_17
timestamp 1649977179
transform -1 0 21896 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_18
timestamp 1649977179
transform 1 0 1104 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_19
timestamp 1649977179
transform -1 0 21896 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_20
timestamp 1649977179
transform 1 0 1104 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_21
timestamp 1649977179
transform -1 0 21896 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_22
timestamp 1649977179
transform 1 0 1104 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_23
timestamp 1649977179
transform -1 0 21896 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_24
timestamp 1649977179
transform 1 0 1104 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_25
timestamp 1649977179
transform -1 0 21896 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_26
timestamp 1649977179
transform 1 0 1104 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_27
timestamp 1649977179
transform -1 0 21896 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_28
timestamp 1649977179
transform 1 0 1104 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_29
timestamp 1649977179
transform -1 0 21896 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_30
timestamp 1649977179
transform 1 0 1104 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_31
timestamp 1649977179
transform -1 0 21896 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_32
timestamp 1649977179
transform 1 0 1104 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_33
timestamp 1649977179
transform -1 0 21896 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_34
timestamp 1649977179
transform 1 0 1104 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_35
timestamp 1649977179
transform -1 0 21896 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_36
timestamp 1649977179
transform 1 0 1104 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_37
timestamp 1649977179
transform -1 0 21896 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_38
timestamp 1649977179
transform 1 0 1104 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_39
timestamp 1649977179
transform -1 0 21896 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_40
timestamp 1649977179
transform 1 0 1104 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_41
timestamp 1649977179
transform -1 0 21896 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_42
timestamp 1649977179
transform 1 0 1104 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_43
timestamp 1649977179
transform -1 0 21896 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_44
timestamp 1649977179
transform 1 0 1104 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_45
timestamp 1649977179
transform -1 0 21896 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_46
timestamp 1649977179
transform 1 0 1104 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_47
timestamp 1649977179
transform -1 0 21896 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_48
timestamp 1649977179
transform 1 0 1104 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_49
timestamp 1649977179
transform -1 0 21896 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_50
timestamp 1649977179
transform 1 0 1104 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_51
timestamp 1649977179
transform -1 0 21896 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_52
timestamp 1649977179
transform 1 0 1104 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_53
timestamp 1649977179
transform -1 0 21896 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_54
timestamp 1649977179
transform 1 0 1104 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_55
timestamp 1649977179
transform -1 0 21896 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_56
timestamp 1649977179
transform 1 0 1104 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_57
timestamp 1649977179
transform -1 0 21896 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_58
timestamp 1649977179
transform 1 0 1104 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_59
timestamp 1649977179
transform -1 0 21896 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_60
timestamp 1649977179
transform 1 0 1104 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_61
timestamp 1649977179
transform -1 0 21896 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_62
timestamp 1649977179
transform 1 0 1104 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_63
timestamp 1649977179
transform -1 0 21896 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_64
timestamp 1649977179
transform 1 0 1104 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_65
timestamp 1649977179
transform -1 0 21896 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_66
timestamp 1649977179
transform 1 0 1104 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_67
timestamp 1649977179
transform -1 0 21896 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_68 dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform 1 0 3680 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_69
timestamp 1649977179
transform 1 0 6256 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_70
timestamp 1649977179
transform 1 0 8832 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_71
timestamp 1649977179
transform 1 0 11408 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_72
timestamp 1649977179
transform 1 0 13984 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_73
timestamp 1649977179
transform 1 0 16560 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_74
timestamp 1649977179
transform 1 0 19136 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_75
timestamp 1649977179
transform 1 0 6256 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_76
timestamp 1649977179
transform 1 0 11408 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_77
timestamp 1649977179
transform 1 0 16560 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_78
timestamp 1649977179
transform 1 0 3680 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_79
timestamp 1649977179
transform 1 0 8832 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_80
timestamp 1649977179
transform 1 0 13984 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_81
timestamp 1649977179
transform 1 0 19136 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_82
timestamp 1649977179
transform 1 0 6256 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_83
timestamp 1649977179
transform 1 0 11408 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_84
timestamp 1649977179
transform 1 0 16560 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_85
timestamp 1649977179
transform 1 0 3680 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_86
timestamp 1649977179
transform 1 0 8832 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_87
timestamp 1649977179
transform 1 0 13984 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_88
timestamp 1649977179
transform 1 0 19136 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_89
timestamp 1649977179
transform 1 0 6256 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_90
timestamp 1649977179
transform 1 0 11408 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_91
timestamp 1649977179
transform 1 0 16560 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_92
timestamp 1649977179
transform 1 0 3680 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_93
timestamp 1649977179
transform 1 0 8832 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_94
timestamp 1649977179
transform 1 0 13984 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_95
timestamp 1649977179
transform 1 0 19136 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_96
timestamp 1649977179
transform 1 0 6256 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_97
timestamp 1649977179
transform 1 0 11408 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_98
timestamp 1649977179
transform 1 0 16560 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_99
timestamp 1649977179
transform 1 0 3680 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_100
timestamp 1649977179
transform 1 0 8832 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_101
timestamp 1649977179
transform 1 0 13984 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_102
timestamp 1649977179
transform 1 0 19136 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_103
timestamp 1649977179
transform 1 0 6256 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_104
timestamp 1649977179
transform 1 0 11408 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_105
timestamp 1649977179
transform 1 0 16560 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_106
timestamp 1649977179
transform 1 0 3680 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_107
timestamp 1649977179
transform 1 0 8832 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_108
timestamp 1649977179
transform 1 0 13984 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_109
timestamp 1649977179
transform 1 0 19136 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_110
timestamp 1649977179
transform 1 0 6256 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_111
timestamp 1649977179
transform 1 0 11408 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_112
timestamp 1649977179
transform 1 0 16560 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_113
timestamp 1649977179
transform 1 0 3680 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_114
timestamp 1649977179
transform 1 0 8832 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_115
timestamp 1649977179
transform 1 0 13984 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_116
timestamp 1649977179
transform 1 0 19136 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_117
timestamp 1649977179
transform 1 0 6256 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_118
timestamp 1649977179
transform 1 0 11408 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_119
timestamp 1649977179
transform 1 0 16560 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_120
timestamp 1649977179
transform 1 0 3680 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_121
timestamp 1649977179
transform 1 0 8832 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_122
timestamp 1649977179
transform 1 0 13984 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_123
timestamp 1649977179
transform 1 0 19136 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_124
timestamp 1649977179
transform 1 0 6256 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_125
timestamp 1649977179
transform 1 0 11408 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_126
timestamp 1649977179
transform 1 0 16560 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_127
timestamp 1649977179
transform 1 0 3680 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_128
timestamp 1649977179
transform 1 0 8832 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_129
timestamp 1649977179
transform 1 0 13984 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_130
timestamp 1649977179
transform 1 0 19136 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_131
timestamp 1649977179
transform 1 0 6256 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_132
timestamp 1649977179
transform 1 0 11408 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_133
timestamp 1649977179
transform 1 0 16560 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_134
timestamp 1649977179
transform 1 0 3680 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_135
timestamp 1649977179
transform 1 0 8832 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_136
timestamp 1649977179
transform 1 0 13984 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_137
timestamp 1649977179
transform 1 0 19136 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_138
timestamp 1649977179
transform 1 0 6256 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_139
timestamp 1649977179
transform 1 0 11408 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_140
timestamp 1649977179
transform 1 0 16560 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_141
timestamp 1649977179
transform 1 0 3680 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_142
timestamp 1649977179
transform 1 0 8832 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_143
timestamp 1649977179
transform 1 0 13984 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_144
timestamp 1649977179
transform 1 0 19136 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_145
timestamp 1649977179
transform 1 0 6256 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_146
timestamp 1649977179
transform 1 0 11408 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_147
timestamp 1649977179
transform 1 0 16560 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_148
timestamp 1649977179
transform 1 0 3680 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_149
timestamp 1649977179
transform 1 0 8832 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_150
timestamp 1649977179
transform 1 0 13984 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_151
timestamp 1649977179
transform 1 0 19136 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_152
timestamp 1649977179
transform 1 0 6256 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_153
timestamp 1649977179
transform 1 0 11408 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_154
timestamp 1649977179
transform 1 0 16560 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_155
timestamp 1649977179
transform 1 0 3680 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_156
timestamp 1649977179
transform 1 0 8832 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_157
timestamp 1649977179
transform 1 0 13984 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_158
timestamp 1649977179
transform 1 0 19136 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_159
timestamp 1649977179
transform 1 0 6256 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_160
timestamp 1649977179
transform 1 0 11408 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_161
timestamp 1649977179
transform 1 0 16560 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_162
timestamp 1649977179
transform 1 0 3680 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_163
timestamp 1649977179
transform 1 0 8832 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_164
timestamp 1649977179
transform 1 0 13984 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_165
timestamp 1649977179
transform 1 0 19136 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_166
timestamp 1649977179
transform 1 0 6256 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_167
timestamp 1649977179
transform 1 0 11408 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_168
timestamp 1649977179
transform 1 0 16560 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_169
timestamp 1649977179
transform 1 0 3680 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_170
timestamp 1649977179
transform 1 0 8832 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_171
timestamp 1649977179
transform 1 0 13984 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_172
timestamp 1649977179
transform 1 0 19136 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_173
timestamp 1649977179
transform 1 0 6256 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_174
timestamp 1649977179
transform 1 0 11408 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_175
timestamp 1649977179
transform 1 0 16560 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_176
timestamp 1649977179
transform 1 0 3680 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_177
timestamp 1649977179
transform 1 0 8832 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_178
timestamp 1649977179
transform 1 0 13984 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_179
timestamp 1649977179
transform 1 0 19136 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_180
timestamp 1649977179
transform 1 0 6256 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_181
timestamp 1649977179
transform 1 0 11408 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_182
timestamp 1649977179
transform 1 0 16560 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_183
timestamp 1649977179
transform 1 0 3680 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_184
timestamp 1649977179
transform 1 0 8832 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_185
timestamp 1649977179
transform 1 0 13984 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_186
timestamp 1649977179
transform 1 0 19136 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_187
timestamp 1649977179
transform 1 0 3680 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_188
timestamp 1649977179
transform 1 0 6256 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_189
timestamp 1649977179
transform 1 0 8832 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_190
timestamp 1649977179
transform 1 0 11408 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_191
timestamp 1649977179
transform 1 0 13984 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_192
timestamp 1649977179
transform 1 0 16560 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_193
timestamp 1649977179
transform 1 0 19136 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__conb_1  _033_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform 1 0 9752 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _034_
timestamp 1649977179
transform 1 0 8556 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _035_
timestamp 1649977179
transform 1 0 9752 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _036_
timestamp 1649977179
transform -1 0 10304 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _037_
timestamp 1649977179
transform 1 0 11500 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _038_
timestamp 1649977179
transform 1 0 11132 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _039_
timestamp 1649977179
transform 1 0 7268 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _040_
timestamp 1649977179
transform 1 0 11224 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _041_
timestamp 1649977179
transform 1 0 9844 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _042_
timestamp 1649977179
transform -1 0 7084 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _043_
timestamp 1649977179
transform -1 0 5336 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _044_
timestamp 1649977179
transform -1 0 7820 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _045_
timestamp 1649977179
transform 1 0 8740 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _046_
timestamp 1649977179
transform 1 0 9384 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _047_
timestamp 1649977179
transform 1 0 10764 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _048_
timestamp 1649977179
transform -1 0 5612 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _049_
timestamp 1649977179
transform 1 0 2944 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _050_
timestamp 1649977179
transform -1 0 8832 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _051_
timestamp 1649977179
transform -1 0 3680 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _052_
timestamp 1649977179
transform -1 0 7636 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _053_
timestamp 1649977179
transform 1 0 5428 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _054_
timestamp 1649977179
transform 1 0 5152 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _055_
timestamp 1649977179
transform 1 0 5980 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _056_
timestamp 1649977179
transform 1 0 4876 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _057_
timestamp 1649977179
transform -1 0 17296 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _058_
timestamp 1649977179
transform 1 0 2668 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _059_
timestamp 1649977179
transform 1 0 11684 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _060_
timestamp 1649977179
transform 1 0 6348 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _061_
timestamp 1649977179
transform 1 0 5704 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _062_
timestamp 1649977179
transform 1 0 7084 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _063_
timestamp 1649977179
transform 1 0 11500 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _064_
timestamp 1649977179
transform 1 0 12880 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _065_
timestamp 1649977179
transform -1 0 14352 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  _066_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform -1 0 2208 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _067_
timestamp 1649977179
transform -1 0 1840 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _068_
timestamp 1649977179
transform -1 0 2208 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _069_
timestamp 1649977179
transform -1 0 2208 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _070_
timestamp 1649977179
transform -1 0 2392 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _071_
timestamp 1649977179
transform 1 0 2852 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _072_
timestamp 1649977179
transform -1 0 2576 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _073_
timestamp 1649977179
transform -1 0 2208 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _074_
timestamp 1649977179
transform -1 0 2208 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _075_
timestamp 1649977179
transform -1 0 2208 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _076_
timestamp 1649977179
transform -1 0 2944 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _077_
timestamp 1649977179
transform -1 0 2576 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _078_
timestamp 1649977179
transform -1 0 2944 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _079_
timestamp 1649977179
transform -1 0 2208 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _080_
timestamp 1649977179
transform -1 0 3220 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _081_
timestamp 1649977179
transform -1 0 2852 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _082_
timestamp 1649977179
transform -1 0 3036 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _083_
timestamp 1649977179
transform -1 0 2484 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _084_
timestamp 1649977179
transform -1 0 2392 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _085_
timestamp 1649977179
transform -1 0 3036 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _086_
timestamp 1649977179
transform -1 0 13524 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _087_
timestamp 1649977179
transform 1 0 14260 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _088_
timestamp 1649977179
transform 1 0 14076 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _089_
timestamp 1649977179
transform 1 0 14628 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _090_
timestamp 1649977179
transform 1 0 15364 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _091_
timestamp 1649977179
transform 1 0 11868 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _092_
timestamp 1649977179
transform 1 0 14996 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _093_
timestamp 1649977179
transform -1 0 16928 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _094_
timestamp 1649977179
transform 1 0 17020 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _095_
timestamp 1649977179
transform 1 0 16652 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _096_
timestamp 1649977179
transform 1 0 18400 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _097_
timestamp 1649977179
transform 1 0 18584 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _098_
timestamp 1649977179
transform -1 0 20976 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _099_
timestamp 1649977179
transform 1 0 20240 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _100_
timestamp 1649977179
transform 1 0 15732 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _101_
timestamp 1649977179
transform 1 0 16100 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _102_
timestamp 1649977179
transform 1 0 19872 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _103_
timestamp 1649977179
transform 1 0 18768 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _104_
timestamp 1649977179
transform 1 0 18032 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _105_
timestamp 1649977179
transform 1 0 19136 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _106_
timestamp 1649977179
transform -1 0 9844 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _107_
timestamp 1649977179
transform 1 0 10580 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _108_
timestamp 1649977179
transform -1 0 9476 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _109_
timestamp 1649977179
transform 1 0 8464 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _110_
timestamp 1649977179
transform 1 0 10028 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _111_
timestamp 1649977179
transform 1 0 7176 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _112_
timestamp 1649977179
transform 1 0 7544 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _113_
timestamp 1649977179
transform 1 0 9200 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _114_
timestamp 1649977179
transform -1 0 8832 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _115_
timestamp 1649977179
transform 1 0 9660 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _116_
timestamp 1649977179
transform 1 0 9844 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _117_
timestamp 1649977179
transform 1 0 10212 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _118_
timestamp 1649977179
transform -1 0 8832 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _119_
timestamp 1649977179
transform 1 0 14260 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _120_
timestamp 1649977179
transform 1 0 8096 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _121_
timestamp 1649977179
transform 1 0 8096 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _122_
timestamp 1649977179
transform -1 0 10028 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _123_
timestamp 1649977179
transform -1 0 9476 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _124_
timestamp 1649977179
transform 1 0 13524 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _125_
timestamp 1649977179
transform 1 0 16284 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  mem_bottom_track_1.sky130_fd_sc_hd__dfxtp_1_0_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform -1 0 21252 0 1 11968
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_bottom_track_1.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1649977179
transform -1 0 13524 0 1 9792
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_bottom_track_1.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1649977179
transform -1 0 13616 0 -1 9792
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_bottom_track_1.sky130_fd_sc_hd__dfxtp_1_3_
timestamp 1649977179
transform 1 0 11500 0 1 10880
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_bottom_track_3.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1649977179
transform -1 0 15732 0 -1 8704
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_bottom_track_3.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1649977179
transform -1 0 13708 0 1 8704
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_bottom_track_3.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1649977179
transform -1 0 15088 0 -1 9792
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_bottom_track_3.sky130_fd_sc_hd__dfxtp_1_3_
timestamp 1649977179
transform 1 0 12972 0 -1 10880
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_bottom_track_5.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1649977179
transform -1 0 16560 0 -1 9792
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_bottom_track_5.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1649977179
transform -1 0 12052 0 1 9792
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_bottom_track_5.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1649977179
transform 1 0 14076 0 1 8704
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_bottom_track_5.sky130_fd_sc_hd__dfxtp_1_3_
timestamp 1649977179
transform 1 0 17112 0 1 9792
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_bottom_track_9.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1649977179
transform -1 0 20792 0 -1 11968
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_bottom_track_9.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1649977179
transform -1 0 19412 0 -1 8704
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_bottom_track_9.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1649977179
transform -1 0 17848 0 1 10880
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_bottom_track_9.sky130_fd_sc_hd__dfxtp_1_3_
timestamp 1649977179
transform 1 0 16284 0 1 8704
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_bottom_track_17.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1649977179
transform -1 0 21344 0 1 7616
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_bottom_track_17.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1649977179
transform -1 0 12972 0 -1 10880
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_bottom_track_17.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1649977179
transform 1 0 16652 0 -1 10880
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_bottom_track_25.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1649977179
transform -1 0 20700 0 1 8704
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_bottom_track_25.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1649977179
transform 1 0 19412 0 -1 8704
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_bottom_track_25.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1649977179
transform 1 0 19872 0 1 13056
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_bottom_track_33.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1649977179
transform -1 0 21068 0 -1 13056
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_bottom_track_33.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1649977179
transform -1 0 17112 0 1 9792
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_bottom_track_33.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1649977179
transform 1 0 18124 0 -1 9792
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_1.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1649977179
transform -1 0 21620 0 -1 15232
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_1.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1649977179
transform -1 0 15916 0 1 14144
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_1.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1649977179
transform 1 0 16652 0 -1 14144
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_3.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1649977179
transform -1 0 18308 0 1 16320
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_3.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1649977179
transform -1 0 13340 0 1 16320
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_3.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1649977179
transform 1 0 12236 0 -1 14144
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_5.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1649977179
transform -1 0 13524 0 -1 15232
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_5.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1649977179
transform -1 0 14168 0 -1 13056
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_5.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1649977179
transform 1 0 12512 0 1 11968
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_7.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1649977179
transform -1 0 15640 0 -1 13056
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_7.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1649977179
transform -1 0 13984 0 -1 11968
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_7.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1649977179
transform -1 0 12512 0 1 11968
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_9.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1649977179
transform 1 0 14168 0 1 9792
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_9.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1649977179
transform 1 0 15088 0 -1 10880
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_9.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1649977179
transform 1 0 17480 0 -1 11968
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_11.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1649977179
transform 1 0 19596 0 -1 9792
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_11.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1649977179
transform -1 0 20792 0 -1 7616
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_11.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1649977179
transform -1 0 18124 0 -1 9792
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_13.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1649977179
transform -1 0 20884 0 -1 10880
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_13.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1649977179
transform -1 0 21068 0 1 10880
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_13.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1649977179
transform -1 0 16376 0 1 10880
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_15.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1649977179
transform 1 0 20148 0 -1 14144
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_15.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1649977179
transform -1 0 21620 0 1 15232
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_15.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1649977179
transform -1 0 20976 0 1 9792
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_17.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1649977179
transform -1 0 16744 0 1 11968
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_17.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1649977179
transform -1 0 13432 0 1 15232
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_19.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1649977179
transform 1 0 12512 0 1 13056
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_19.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1649977179
transform 1 0 12972 0 -1 17408
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_21.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1649977179
transform 1 0 16100 0 1 15232
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_21.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1649977179
transform 1 0 18124 0 -1 13056
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_23.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1649977179
transform -1 0 21160 0 1 14144
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_23.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1649977179
transform -1 0 20148 0 -1 15232
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_25.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1649977179
transform -1 0 19596 0 -1 14144
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_25.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1649977179
transform -1 0 17664 0 1 14144
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_29.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1649977179
transform 1 0 18952 0 -1 17408
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_29.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1649977179
transform -1 0 20976 0 1 18496
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_31.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1649977179
transform 1 0 19780 0 1 17408
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_31.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1649977179
transform -1 0 21620 0 1 19584
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_33.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1649977179
transform -1 0 18124 0 -1 17408
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_33.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1649977179
transform -1 0 18124 0 -1 18496
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_35.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1649977179
transform -1 0 16560 0 -1 18496
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_35.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1649977179
transform -1 0 14536 0 -1 18496
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_37.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1649977179
transform -1 0 12972 0 -1 19584
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_37.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1649977179
transform 1 0 14720 0 1 18496
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_39.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1649977179
transform 1 0 19596 0 -1 18496
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_39.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1649977179
transform -1 0 20792 0 -1 19584
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_track_0.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1649977179
transform -1 0 21528 0 -1 16320
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_track_0.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1649977179
transform -1 0 18124 0 -1 15232
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_track_0.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1649977179
transform -1 0 15824 0 1 16320
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_track_0.sky130_fd_sc_hd__dfxtp_1_3_
timestamp 1649977179
transform -1 0 14444 0 -1 19584
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_track_2.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1649977179
transform -1 0 13064 0 1 19584
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_track_2.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1649977179
transform -1 0 11868 0 1 18496
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_track_2.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1649977179
transform -1 0 13616 0 -1 16320
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_track_2.sky130_fd_sc_hd__dfxtp_1_3_
timestamp 1649977179
transform 1 0 11684 0 1 17408
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_track_4.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1649977179
transform -1 0 16560 0 -1 17408
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_track_4.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1649977179
transform -1 0 12972 0 -1 18496
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_track_4.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1649977179
transform 1 0 11868 0 1 18496
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_track_4.sky130_fd_sc_hd__dfxtp_1_3_
timestamp 1649977179
transform 1 0 16468 0 1 17408
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_track_8.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1649977179
transform -1 0 19596 0 -1 18496
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_track_8.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1649977179
transform -1 0 18216 0 1 18496
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_track_8.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1649977179
transform -1 0 12972 0 -1 17408
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_track_8.sky130_fd_sc_hd__dfxtp_1_3_
timestamp 1649977179
transform -1 0 20700 0 1 16320
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_track_16.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1649977179
transform -1 0 19320 0 -1 16320
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_track_16.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1649977179
transform -1 0 15548 0 1 15232
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_track_16.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1649977179
transform -1 0 13616 0 1 14144
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_track_24.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1649977179
transform -1 0 16560 0 -1 14144
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_track_24.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1649977179
transform -1 0 15272 0 -1 16320
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_track_24.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1649977179
transform 1 0 16652 0 -1 13056
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_track_32.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1649977179
transform -1 0 17572 0 1 13056
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_track_32.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1649977179
transform -1 0 15364 0 -1 15232
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_track_32.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1649977179
transform 1 0 16744 0 1 11968
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_1.mux_l1_in_0_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform 1 0 11500 0 -1 4352
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_1.mux_l1_in_1_
timestamp 1649977179
transform -1 0 10948 0 1 3264
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_1.mux_l1_in_2_
timestamp 1649977179
transform 1 0 8924 0 1 2176
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_1.mux_l2_in_0_
timestamp 1649977179
transform 1 0 10488 0 -1 4352
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_1.mux_l2_in_1_
timestamp 1649977179
transform -1 0 9016 0 -1 4352
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_1.mux_l2_in_2_
timestamp 1649977179
transform -1 0 6440 0 1 5440
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_1.mux_l2_in_3_
timestamp 1649977179
transform -1 0 5888 0 1 4352
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_1.mux_l3_in_0_
timestamp 1649977179
transform -1 0 11040 0 -1 5440
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_1.mux_l3_in_1_
timestamp 1649977179
transform -1 0 7176 0 -1 5440
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_1.mux_l4_in_0_
timestamp 1649977179
transform -1 0 12420 0 -1 5440
box -38 -48 866 592
use sky130_fd_sc_hd__buf_4  mux_bottom_track_1.sky130_fd_sc_hd__buf_4_0_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform 1 0 13248 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_3.mux_l1_in_0_
timestamp 1649977179
transform 1 0 9660 0 -1 4352
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_3.mux_l1_in_1_
timestamp 1649977179
transform 1 0 9752 0 1 4352
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_3.mux_l2_in_0_
timestamp 1649977179
transform 1 0 9108 0 1 5440
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_3.mux_l2_in_1_
timestamp 1649977179
transform -1 0 5980 0 -1 5440
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_3.mux_l2_in_2_
timestamp 1649977179
transform -1 0 2484 0 -1 6528
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_3.mux_l2_in_3_
timestamp 1649977179
transform -1 0 2668 0 -1 5440
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_3.mux_l3_in_0_
timestamp 1649977179
transform -1 0 8832 0 1 5440
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_3.mux_l3_in_1_
timestamp 1649977179
transform -1 0 5704 0 -1 6528
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_3.mux_l4_in_0_
timestamp 1649977179
transform -1 0 11408 0 -1 6528
box -38 -48 866 592
use sky130_fd_sc_hd__buf_4  mux_bottom_track_3.sky130_fd_sc_hd__buf_4_0_
timestamp 1649977179
transform 1 0 13340 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_5.mux_l1_in_0_
timestamp 1649977179
transform 1 0 12236 0 -1 3264
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_5.mux_l1_in_1_
timestamp 1649977179
transform -1 0 10580 0 -1 3264
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_5.mux_l1_in_2_
timestamp 1649977179
transform 1 0 7268 0 -1 3264
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_5.mux_l1_in_3_
timestamp 1649977179
transform -1 0 7084 0 1 3264
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_5.mux_l1_in_4_
timestamp 1649977179
transform 1 0 4968 0 1 2176
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_5.mux_l1_in_5_
timestamp 1649977179
transform 1 0 4876 0 1 3264
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_5.mux_l1_in_6_
timestamp 1649977179
transform -1 0 2576 0 1 7616
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_5.mux_l2_in_0_
timestamp 1649977179
transform -1 0 11408 0 -1 3264
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_5.mux_l2_in_1_
timestamp 1649977179
transform -1 0 7176 0 -1 3264
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_5.mux_l2_in_2_
timestamp 1649977179
transform -1 0 5520 0 -1 3264
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_5.mux_l2_in_3_
timestamp 1649977179
transform -1 0 6256 0 -1 4352
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_5.mux_l3_in_0_
timestamp 1649977179
transform -1 0 12236 0 1 3264
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_5.mux_l3_in_1_
timestamp 1649977179
transform -1 0 9752 0 1 3264
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_5.mux_l4_in_0_
timestamp 1649977179
transform -1 0 13800 0 1 3264
box -38 -48 866 592
use sky130_fd_sc_hd__buf_4  mux_bottom_track_5.sky130_fd_sc_hd__buf_4_0_
timestamp 1649977179
transform 1 0 13708 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_9.mux_l1_in_0_
timestamp 1649977179
transform 1 0 16652 0 -1 4352
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_9.mux_l2_in_0_
timestamp 1649977179
transform 1 0 15456 0 1 4352
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_9.mux_l2_in_1_
timestamp 1649977179
transform -1 0 8188 0 -1 4352
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_9.mux_l2_in_2_
timestamp 1649977179
transform -1 0 4692 0 1 6528
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_9.mux_l2_in_3_
timestamp 1649977179
transform -1 0 4876 0 -1 6528
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_9.mux_l3_in_0_
timestamp 1649977179
transform 1 0 14996 0 -1 5440
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_9.mux_l3_in_1_
timestamp 1649977179
transform -1 0 10488 0 -1 6528
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_9.mux_l4_in_0_
timestamp 1649977179
transform 1 0 14352 0 1 4352
box -38 -48 866 592
use sky130_fd_sc_hd__buf_4  mux_bottom_track_9.sky130_fd_sc_hd__buf_4_0_
timestamp 1649977179
transform 1 0 14352 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_17.mux_l1_in_0_
timestamp 1649977179
transform -1 0 13248 0 -1 5440
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_17.mux_l1_in_1_
timestamp 1649977179
transform -1 0 8556 0 1 4352
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_17.mux_l1_in_2_
timestamp 1649977179
transform -1 0 5336 0 1 8704
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_17.mux_l1_in_3_
timestamp 1649977179
transform -1 0 4876 0 -1 8704
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_17.mux_l2_in_0_
timestamp 1649977179
transform -1 0 13340 0 1 5440
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_17.mux_l2_in_1_
timestamp 1649977179
transform -1 0 10488 0 -1 8704
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_17.mux_l3_in_0_
timestamp 1649977179
transform -1 0 14720 0 -1 6528
box -38 -48 866 592
use sky130_fd_sc_hd__buf_4  mux_bottom_track_17.sky130_fd_sc_hd__buf_4_0_
timestamp 1649977179
transform 1 0 15824 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_25.mux_l1_in_0_
timestamp 1649977179
transform 1 0 17572 0 -1 4352
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_25.mux_l1_in_1_
timestamp 1649977179
transform -1 0 9752 0 -1 3264
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_25.mux_l1_in_2_
timestamp 1649977179
transform -1 0 11868 0 1 7616
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_25.mux_l2_in_0_
timestamp 1649977179
transform -1 0 18124 0 1 4352
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_25.mux_l2_in_1_
timestamp 1649977179
transform -1 0 18216 0 1 5440
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_25.mux_l3_in_0_
timestamp 1649977179
transform -1 0 20792 0 1 5440
box -38 -48 866 592
use sky130_fd_sc_hd__buf_4  mux_bottom_track_25.sky130_fd_sc_hd__buf_4_0_
timestamp 1649977179
transform 1 0 20608 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_33.mux_l1_in_0_
timestamp 1649977179
transform -1 0 10212 0 -1 5440
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_33.mux_l1_in_1_
timestamp 1649977179
transform -1 0 5152 0 -1 5440
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_33.mux_l1_in_2_
timestamp 1649977179
transform -1 0 5428 0 -1 7616
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_33.mux_l2_in_0_
timestamp 1649977179
transform -1 0 11224 0 1 5440
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_33.mux_l2_in_1_
timestamp 1649977179
transform -1 0 12236 0 1 5440
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_33.mux_l3_in_0_
timestamp 1649977179
transform -1 0 17388 0 1 5440
box -38 -48 866 592
use sky130_fd_sc_hd__buf_4  mux_bottom_track_33.sky130_fd_sc_hd__buf_4_0_
timestamp 1649977179
transform 1 0 19228 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_1.mux_l1_in_0_
timestamp 1649977179
transform 1 0 6348 0 -1 13056
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_1.mux_l1_in_1_
timestamp 1649977179
transform 1 0 5612 0 1 9792
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_1.mux_l1_in_2_
timestamp 1649977179
transform 1 0 6348 0 -1 11968
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_1.mux_l1_in_3_
timestamp 1649977179
transform -1 0 6256 0 1 10880
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_1.mux_l2_in_0_
timestamp 1649977179
transform 1 0 5428 0 -1 13056
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_1.mux_l2_in_1_
timestamp 1649977179
transform 1 0 5612 0 1 11968
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_1.mux_l3_in_0_
timestamp 1649977179
transform 1 0 4600 0 -1 13056
box -38 -48 866 592
use sky130_fd_sc_hd__buf_4  mux_left_track_1.sky130_fd_sc_hd__buf_4_0_
timestamp 1649977179
transform -1 0 3680 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_3.mux_l1_in_0_
timestamp 1649977179
transform 1 0 6256 0 1 4352
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_3.mux_l1_in_1_
timestamp 1649977179
transform 1 0 6440 0 1 6528
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_3.mux_l1_in_2_
timestamp 1649977179
transform 1 0 6440 0 1 7616
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_3.mux_l1_in_3_
timestamp 1649977179
transform 1 0 6440 0 -1 7616
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_3.mux_l2_in_0_
timestamp 1649977179
transform -1 0 6256 0 -1 7616
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_3.mux_l2_in_1_
timestamp 1649977179
transform -1 0 6256 0 -1 8704
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_3.mux_l3_in_0_
timestamp 1649977179
transform 1 0 6164 0 1 8704
box -38 -48 866 592
use sky130_fd_sc_hd__buf_4  mux_left_track_3.sky130_fd_sc_hd__buf_4_0_
timestamp 1649977179
transform -1 0 2852 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_5.mux_l1_in_0_
timestamp 1649977179
transform -1 0 7268 0 1 5440
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_5.mux_l1_in_1_
timestamp 1649977179
transform 1 0 7912 0 -1 6528
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_5.mux_l1_in_2_
timestamp 1649977179
transform 1 0 8740 0 -1 6528
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_5.mux_l1_in_3_
timestamp 1649977179
transform 1 0 7912 0 -1 5440
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_5.mux_l2_in_0_
timestamp 1649977179
transform 1 0 7084 0 -1 6528
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_5.mux_l2_in_1_
timestamp 1649977179
transform 1 0 7544 0 -1 7616
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_5.mux_l3_in_0_
timestamp 1649977179
transform 1 0 6900 0 -1 8704
box -38 -48 866 592
use sky130_fd_sc_hd__buf_4  mux_left_track_5.sky130_fd_sc_hd__buf_4_0_
timestamp 1649977179
transform -1 0 3220 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_7.mux_l1_in_0_
timestamp 1649977179
transform -1 0 8464 0 1 6528
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_7.mux_l1_in_1_
timestamp 1649977179
transform 1 0 9292 0 1 6528
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_7.mux_l1_in_2_
timestamp 1649977179
transform 1 0 8556 0 -1 8704
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_7.mux_l1_in_3_
timestamp 1649977179
transform -1 0 8556 0 -1 8704
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_7.mux_l2_in_0_
timestamp 1649977179
transform 1 0 7820 0 1 7616
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_7.mux_l2_in_1_
timestamp 1649977179
transform 1 0 7820 0 1 8704
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_7.mux_l3_in_0_
timestamp 1649977179
transform 1 0 6992 0 1 8704
box -38 -48 866 592
use sky130_fd_sc_hd__buf_4  mux_left_track_7.sky130_fd_sc_hd__buf_4_0_
timestamp 1649977179
transform -1 0 3588 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_9.mux_l1_in_0_
timestamp 1649977179
transform 1 0 12236 0 -1 6528
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_9.mux_l2_in_0_
timestamp 1649977179
transform -1 0 10948 0 1 6528
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_9.mux_l2_in_1_
timestamp 1649977179
transform -1 0 11316 0 1 8704
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_9.mux_l3_in_0_
timestamp 1649977179
transform 1 0 11316 0 1 8704
box -38 -48 866 592
use sky130_fd_sc_hd__buf_4  mux_left_track_9.sky130_fd_sc_hd__buf_4_0_
timestamp 1649977179
transform -1 0 4416 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_11.mux_l1_in_0_
timestamp 1649977179
transform 1 0 15088 0 -1 7616
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_11.mux_l2_in_0_
timestamp 1649977179
transform -1 0 9936 0 1 7616
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_11.mux_l2_in_1_
timestamp 1649977179
transform 1 0 10488 0 -1 7616
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_11.mux_l3_in_0_
timestamp 1649977179
transform 1 0 9108 0 -1 7616
box -38 -48 866 592
use sky130_fd_sc_hd__buf_4  mux_left_track_11.sky130_fd_sc_hd__buf_4_0_
timestamp 1649977179
transform -1 0 3128 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_13.mux_l1_in_0_
timestamp 1649977179
transform 1 0 16008 0 1 7616
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_13.mux_l2_in_0_
timestamp 1649977179
transform -1 0 12604 0 1 6528
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_13.mux_l2_in_1_
timestamp 1649977179
transform 1 0 12052 0 -1 7616
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_13.mux_l3_in_0_
timestamp 1649977179
transform 1 0 11868 0 1 7616
box -38 -48 866 592
use sky130_fd_sc_hd__buf_4  mux_left_track_13.sky130_fd_sc_hd__buf_4_0_
timestamp 1649977179
transform -1 0 5888 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_15.mux_l1_in_0_
timestamp 1649977179
transform 1 0 17848 0 1 7616
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_15.mux_l2_in_0_
timestamp 1649977179
transform 1 0 14076 0 1 6528
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_15.mux_l2_in_1_
timestamp 1649977179
transform 1 0 14260 0 -1 7616
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_15.mux_l3_in_0_
timestamp 1649977179
transform 1 0 13432 0 -1 7616
box -38 -48 866 592
use sky130_fd_sc_hd__buf_4  mux_left_track_15.sky130_fd_sc_hd__buf_4_0_
timestamp 1649977179
transform -1 0 6440 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_17.mux_l1_in_0_
timestamp 1649977179
transform 1 0 9108 0 -1 10880
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_17.mux_l1_in_1_
timestamp 1649977179
transform -1 0 9752 0 -1 9792
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_17.mux_l2_in_0_
timestamp 1649977179
transform 1 0 8924 0 1 10880
box -38 -48 866 592
use sky130_fd_sc_hd__buf_4  mux_left_track_17.sky130_fd_sc_hd__buf_4_0_
timestamp 1649977179
transform -1 0 4508 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_19.mux_l1_in_0_
timestamp 1649977179
transform 1 0 10028 0 1 10880
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_19.mux_l1_in_1_
timestamp 1649977179
transform -1 0 9108 0 -1 10880
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_19.mux_l2_in_0_
timestamp 1649977179
transform 1 0 8924 0 1 11968
box -38 -48 866 592
use sky130_fd_sc_hd__buf_4  mux_left_track_19.sky130_fd_sc_hd__buf_4_0_
timestamp 1649977179
transform -1 0 4600 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_21.mux_l1_in_0_
timestamp 1649977179
transform 1 0 10212 0 1 11968
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_21.mux_l1_in_1_
timestamp 1649977179
transform 1 0 8556 0 -1 13056
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_21.mux_l2_in_0_
timestamp 1649977179
transform 1 0 8004 0 1 13056
box -38 -48 866 592
use sky130_fd_sc_hd__buf_4  mux_left_track_21.sky130_fd_sc_hd__buf_4_0_
timestamp 1649977179
transform -1 0 5060 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_23.mux_l1_in_0_
timestamp 1649977179
transform 1 0 10120 0 -1 11968
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_23.mux_l1_in_1_
timestamp 1649977179
transform 1 0 10304 0 -1 10880
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_23.mux_l2_in_0_
timestamp 1649977179
transform 1 0 9292 0 -1 11968
box -38 -48 866 592
use sky130_fd_sc_hd__buf_4  mux_left_track_23.sky130_fd_sc_hd__buf_4_0_
timestamp 1649977179
transform -1 0 5428 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_25.mux_l1_in_0_
timestamp 1649977179
transform 1 0 9936 0 -1 9792
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_25.mux_l1_in_1_
timestamp 1649977179
transform 1 0 10488 0 -1 8704
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_25.mux_l2_in_0_
timestamp 1649977179
transform 1 0 9660 0 1 8704
box -38 -48 866 592
use sky130_fd_sc_hd__buf_4  mux_left_track_25.sky130_fd_sc_hd__buf_4_0_
timestamp 1649977179
transform -1 0 5336 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_29.mux_l1_in_0_
timestamp 1649977179
transform 1 0 10580 0 -1 15232
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_29.mux_l2_in_0_
timestamp 1649977179
transform 1 0 10212 0 1 15232
box -38 -48 866 592
use sky130_fd_sc_hd__buf_4  mux_left_track_29.sky130_fd_sc_hd__buf_4_0_
timestamp 1649977179
transform -1 0 3956 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_31.mux_l1_in_0_
timestamp 1649977179
transform -1 0 11132 0 -1 16320
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_31.mux_l2_in_0_
timestamp 1649977179
transform 1 0 10396 0 1 16320
box -38 -48 866 592
use sky130_fd_sc_hd__buf_4  mux_left_track_31.sky130_fd_sc_hd__buf_4_0_
timestamp 1649977179
transform -1 0 3680 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_33.mux_l1_in_0_
timestamp 1649977179
transform 1 0 9568 0 -1 17408
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_33.mux_l2_in_0_
timestamp 1649977179
transform 1 0 8740 0 -1 17408
box -38 -48 866 592
use sky130_fd_sc_hd__buf_4  mux_left_track_33.sky130_fd_sc_hd__buf_4_0_
timestamp 1649977179
transform -1 0 3772 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_35.mux_l1_in_0_
timestamp 1649977179
transform 1 0 7820 0 -1 15232
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_35.mux_l2_in_0_
timestamp 1649977179
transform 1 0 7084 0 1 16320
box -38 -48 866 592
use sky130_fd_sc_hd__buf_4  mux_left_track_35.sky130_fd_sc_hd__buf_4_0_
timestamp 1649977179
transform -1 0 3128 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_37.mux_l1_in_0_
timestamp 1649977179
transform 1 0 6072 0 1 15232
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_37.mux_l2_in_0_
timestamp 1649977179
transform 1 0 5520 0 1 16320
box -38 -48 866 592
use sky130_fd_sc_hd__buf_4  mux_left_track_37.sky130_fd_sc_hd__buf_4_0_
timestamp 1649977179
transform -1 0 3404 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_39.mux_l1_in_0_
timestamp 1649977179
transform 1 0 8188 0 -1 18496
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_39.mux_l2_in_0_
timestamp 1649977179
transform -1 0 8372 0 -1 17408
box -38 -48 866 592
use sky130_fd_sc_hd__buf_4  mux_left_track_39.sky130_fd_sc_hd__buf_4_0_
timestamp 1649977179
transform -1 0 8464 0 1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_0.mux_l1_in_0_
timestamp 1649977179
transform -1 0 6072 0 1 15232
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_0.mux_l1_in_1_
timestamp 1649977179
transform -1 0 5244 0 1 15232
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_0.mux_l1_in_2_
timestamp 1649977179
transform -1 0 8740 0 1 16320
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_0.mux_l2_in_0_
timestamp 1649977179
transform -1 0 6164 0 -1 16320
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_0.mux_l2_in_1_
timestamp 1649977179
transform 1 0 8924 0 1 15232
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_0.mux_l2_in_2_
timestamp 1649977179
transform -1 0 6164 0 1 8704
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_0.mux_l2_in_3_
timestamp 1649977179
transform -1 0 5980 0 -1 10880
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_0.mux_l3_in_0_
timestamp 1649977179
transform -1 0 8280 0 -1 16320
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_0.mux_l3_in_1_
timestamp 1649977179
transform -1 0 7084 0 1 10880
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_0.mux_l4_in_0_
timestamp 1649977179
transform -1 0 8464 0 1 15232
box -38 -48 866 592
use sky130_fd_sc_hd__buf_4  mux_top_track_0.sky130_fd_sc_hd__buf_4_0_
timestamp 1649977179
transform 1 0 9752 0 -1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_2.mux_l1_in_0_
timestamp 1649977179
transform -1 0 4692 0 1 14144
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_2.mux_l2_in_0_
timestamp 1649977179
transform -1 0 5428 0 -1 15232
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_2.mux_l2_in_1_
timestamp 1649977179
transform 1 0 6348 0 -1 14144
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_2.mux_l2_in_2_
timestamp 1649977179
transform -1 0 8280 0 -1 10880
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_2.mux_l2_in_3_
timestamp 1649977179
transform 1 0 8924 0 1 9792
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_2.mux_l3_in_0_
timestamp 1649977179
transform -1 0 6716 0 1 14144
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_2.mux_l3_in_1_
timestamp 1649977179
transform -1 0 8464 0 -1 11968
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_2.mux_l4_in_0_
timestamp 1649977179
transform 1 0 9476 0 -1 15232
box -38 -48 866 592
use sky130_fd_sc_hd__buf_4  mux_top_track_2.sky130_fd_sc_hd__buf_4_0_
timestamp 1649977179
transform -1 0 9752 0 -1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_4.mux_l1_in_0_
timestamp 1649977179
transform 1 0 5888 0 1 17408
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_4.mux_l1_in_1_
timestamp 1649977179
transform -1 0 4784 0 1 16320
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_4.mux_l1_in_2_
timestamp 1649977179
transform 1 0 5152 0 -1 18496
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_4.mux_l1_in_3_
timestamp 1649977179
transform -1 0 4968 0 -1 17408
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_4.mux_l1_in_4_
timestamp 1649977179
transform 1 0 7544 0 1 14144
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_4.mux_l1_in_5_
timestamp 1649977179
transform 1 0 7452 0 1 11968
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_4.mux_l1_in_6_
timestamp 1649977179
transform -1 0 5152 0 -1 10880
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_4.mux_l2_in_0_
timestamp 1649977179
transform -1 0 5980 0 -1 17408
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_4.mux_l2_in_1_
timestamp 1649977179
transform -1 0 5888 0 1 17408
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_4.mux_l2_in_2_
timestamp 1649977179
transform 1 0 7268 0 -1 14144
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_4.mux_l2_in_3_
timestamp 1649977179
transform -1 0 5796 0 -1 14144
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_4.mux_l3_in_0_
timestamp 1649977179
transform -1 0 7452 0 -1 17408
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_4.mux_l3_in_1_
timestamp 1649977179
transform -1 0 7544 0 -1 15232
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_4.mux_l4_in_0_
timestamp 1649977179
transform -1 0 8648 0 1 17408
box -38 -48 866 592
use sky130_fd_sc_hd__buf_4  mux_top_track_4.sky130_fd_sc_hd__buf_4_0_
timestamp 1649977179
transform 1 0 9200 0 1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_8.mux_l1_in_0_
timestamp 1649977179
transform -1 0 7360 0 -1 16320
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_8.mux_l2_in_0_
timestamp 1649977179
transform -1 0 9476 0 -1 15232
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_8.mux_l2_in_1_
timestamp 1649977179
transform -1 0 10396 0 1 16320
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_8.mux_l2_in_2_
timestamp 1649977179
transform -1 0 5336 0 -1 9792
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_8.mux_l2_in_3_
timestamp 1649977179
transform -1 0 5428 0 1 10880
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_8.mux_l3_in_0_
timestamp 1649977179
transform 1 0 9936 0 1 14144
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_8.mux_l3_in_1_
timestamp 1649977179
transform -1 0 7176 0 1 13056
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_8.mux_l4_in_0_
timestamp 1649977179
transform -1 0 9936 0 1 14144
box -38 -48 866 592
use sky130_fd_sc_hd__buf_4  mux_top_track_8.sky130_fd_sc_hd__buf_4_0_
timestamp 1649977179
transform -1 0 10120 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_16.mux_l1_in_0_
timestamp 1649977179
transform -1 0 4600 0 -1 15232
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_16.mux_l1_in_1_
timestamp 1649977179
transform -1 0 10948 0 -1 14144
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_16.mux_l1_in_2_
timestamp 1649977179
transform -1 0 3036 0 1 8704
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_16.mux_l1_in_3_
timestamp 1649977179
transform -1 0 3220 0 1 9792
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_16.mux_l2_in_0_
timestamp 1649977179
transform 1 0 10212 0 1 13056
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_16.mux_l2_in_1_
timestamp 1649977179
transform -1 0 7176 0 -1 10880
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_16.mux_l3_in_0_
timestamp 1649977179
transform 1 0 9936 0 -1 13056
box -38 -48 866 592
use sky130_fd_sc_hd__buf_4  mux_top_track_16.sky130_fd_sc_hd__buf_4_0_
timestamp 1649977179
transform -1 0 9844 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_24.mux_l1_in_0_
timestamp 1649977179
transform -1 0 3772 0 -1 15232
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_24.mux_l1_in_1_
timestamp 1649977179
transform 1 0 11500 0 -1 11968
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_24.mux_l1_in_2_
timestamp 1649977179
transform -1 0 2668 0 -1 8704
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_24.mux_l1_in_3_
timestamp 1649977179
transform -1 0 4600 0 1 9792
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_24.mux_l2_in_0_
timestamp 1649977179
transform 1 0 11040 0 1 13056
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_24.mux_l2_in_1_
timestamp 1649977179
transform -1 0 7268 0 1 9792
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_24.mux_l3_in_0_
timestamp 1649977179
transform 1 0 9384 0 1 13056
box -38 -48 866 592
use sky130_fd_sc_hd__buf_4  mux_top_track_24.sky130_fd_sc_hd__buf_4_0_
timestamp 1649977179
transform -1 0 9568 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_32.mux_l1_in_0_
timestamp 1649977179
transform -1 0 5704 0 1 14144
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_32.mux_l1_in_1_
timestamp 1649977179
transform 1 0 7268 0 1 9792
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_32.mux_l1_in_2_
timestamp 1649977179
transform -1 0 7176 0 -1 9792
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_32.mux_l2_in_0_
timestamp 1649977179
transform -1 0 8004 0 1 13056
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_32.mux_l2_in_1_
timestamp 1649977179
transform -1 0 8464 0 -1 13056
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_32.mux_l3_in_0_
timestamp 1649977179
transform -1 0 10120 0 -1 14144
box -38 -48 866 592
use sky130_fd_sc_hd__buf_4  mux_top_track_32.sky130_fd_sc_hd__buf_4_0_
timestamp 1649977179
transform 1 0 10396 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__buf_8  prog_clk_0_FTB00 dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform 1 0 20424 0 -1 20672
box -38 -48 1142 592
<< labels >>
flabel metal4 s 6142 2128 6462 20720 0 FreeSans 1920 90 0 0 VGND
port 0 nsew ground bidirectional
flabel metal4 s 11340 2128 11660 20720 0 FreeSans 1920 90 0 0 VGND
port 0 nsew ground bidirectional
flabel metal4 s 16538 2128 16858 20720 0 FreeSans 1920 90 0 0 VGND
port 0 nsew ground bidirectional
flabel metal4 s 21736 2128 22056 20720 0 FreeSans 1920 90 0 0 VGND
port 0 nsew ground bidirectional
flabel metal4 s 3543 2128 3863 20720 0 FreeSans 1920 90 0 0 VPWR
port 1 nsew power bidirectional
flabel metal4 s 8741 2128 9061 20720 0 FreeSans 1920 90 0 0 VPWR
port 1 nsew power bidirectional
flabel metal4 s 13939 2128 14259 20720 0 FreeSans 1920 90 0 0 VPWR
port 1 nsew power bidirectional
flabel metal4 s 19137 2128 19457 20720 0 FreeSans 1920 90 0 0 VPWR
port 1 nsew power bidirectional
flabel metal2 s 386 0 442 800 0 FreeSans 224 90 0 0 bottom_left_grid_pin_42_
port 2 nsew signal input
flabel metal2 s 846 0 902 800 0 FreeSans 224 90 0 0 bottom_left_grid_pin_43_
port 3 nsew signal input
flabel metal2 s 1306 0 1362 800 0 FreeSans 224 90 0 0 bottom_left_grid_pin_44_
port 4 nsew signal input
flabel metal2 s 1766 0 1822 800 0 FreeSans 224 90 0 0 bottom_left_grid_pin_45_
port 5 nsew signal input
flabel metal2 s 2226 0 2282 800 0 FreeSans 224 90 0 0 bottom_left_grid_pin_46_
port 6 nsew signal input
flabel metal2 s 2686 0 2742 800 0 FreeSans 224 90 0 0 bottom_left_grid_pin_47_
port 7 nsew signal input
flabel metal2 s 3146 0 3202 800 0 FreeSans 224 90 0 0 bottom_left_grid_pin_48_
port 8 nsew signal input
flabel metal2 s 3606 0 3662 800 0 FreeSans 224 90 0 0 bottom_left_grid_pin_49_
port 9 nsew signal input
flabel metal2 s 22466 0 22522 800 0 FreeSans 224 90 0 0 bottom_right_grid_pin_1_
port 10 nsew signal input
flabel metal3 s 22200 5720 23000 5840 0 FreeSans 480 0 0 0 ccff_head
port 11 nsew signal input
flabel metal3 s 22200 17144 23000 17264 0 FreeSans 480 0 0 0 ccff_tail
port 12 nsew signal tristate
flabel metal3 s 0 5040 800 5160 0 FreeSans 480 0 0 0 chanx_left_in[0]
port 13 nsew signal input
flabel metal3 s 0 9120 800 9240 0 FreeSans 480 0 0 0 chanx_left_in[10]
port 14 nsew signal input
flabel metal3 s 0 9528 800 9648 0 FreeSans 480 0 0 0 chanx_left_in[11]
port 15 nsew signal input
flabel metal3 s 0 9936 800 10056 0 FreeSans 480 0 0 0 chanx_left_in[12]
port 16 nsew signal input
flabel metal3 s 0 10344 800 10464 0 FreeSans 480 0 0 0 chanx_left_in[13]
port 17 nsew signal input
flabel metal3 s 0 10752 800 10872 0 FreeSans 480 0 0 0 chanx_left_in[14]
port 18 nsew signal input
flabel metal3 s 0 11160 800 11280 0 FreeSans 480 0 0 0 chanx_left_in[15]
port 19 nsew signal input
flabel metal3 s 0 11568 800 11688 0 FreeSans 480 0 0 0 chanx_left_in[16]
port 20 nsew signal input
flabel metal3 s 0 11976 800 12096 0 FreeSans 480 0 0 0 chanx_left_in[17]
port 21 nsew signal input
flabel metal3 s 0 12384 800 12504 0 FreeSans 480 0 0 0 chanx_left_in[18]
port 22 nsew signal input
flabel metal3 s 0 12792 800 12912 0 FreeSans 480 0 0 0 chanx_left_in[19]
port 23 nsew signal input
flabel metal3 s 0 5448 800 5568 0 FreeSans 480 0 0 0 chanx_left_in[1]
port 24 nsew signal input
flabel metal3 s 0 5856 800 5976 0 FreeSans 480 0 0 0 chanx_left_in[2]
port 25 nsew signal input
flabel metal3 s 0 6264 800 6384 0 FreeSans 480 0 0 0 chanx_left_in[3]
port 26 nsew signal input
flabel metal3 s 0 6672 800 6792 0 FreeSans 480 0 0 0 chanx_left_in[4]
port 27 nsew signal input
flabel metal3 s 0 7080 800 7200 0 FreeSans 480 0 0 0 chanx_left_in[5]
port 28 nsew signal input
flabel metal3 s 0 7488 800 7608 0 FreeSans 480 0 0 0 chanx_left_in[6]
port 29 nsew signal input
flabel metal3 s 0 7896 800 8016 0 FreeSans 480 0 0 0 chanx_left_in[7]
port 30 nsew signal input
flabel metal3 s 0 8304 800 8424 0 FreeSans 480 0 0 0 chanx_left_in[8]
port 31 nsew signal input
flabel metal3 s 0 8712 800 8832 0 FreeSans 480 0 0 0 chanx_left_in[9]
port 32 nsew signal input
flabel metal3 s 0 13200 800 13320 0 FreeSans 480 0 0 0 chanx_left_out[0]
port 33 nsew signal tristate
flabel metal3 s 0 17280 800 17400 0 FreeSans 480 0 0 0 chanx_left_out[10]
port 34 nsew signal tristate
flabel metal3 s 0 17688 800 17808 0 FreeSans 480 0 0 0 chanx_left_out[11]
port 35 nsew signal tristate
flabel metal3 s 0 18096 800 18216 0 FreeSans 480 0 0 0 chanx_left_out[12]
port 36 nsew signal tristate
flabel metal3 s 0 18504 800 18624 0 FreeSans 480 0 0 0 chanx_left_out[13]
port 37 nsew signal tristate
flabel metal3 s 0 18912 800 19032 0 FreeSans 480 0 0 0 chanx_left_out[14]
port 38 nsew signal tristate
flabel metal3 s 0 19320 800 19440 0 FreeSans 480 0 0 0 chanx_left_out[15]
port 39 nsew signal tristate
flabel metal3 s 0 19728 800 19848 0 FreeSans 480 0 0 0 chanx_left_out[16]
port 40 nsew signal tristate
flabel metal3 s 0 20136 800 20256 0 FreeSans 480 0 0 0 chanx_left_out[17]
port 41 nsew signal tristate
flabel metal3 s 0 20544 800 20664 0 FreeSans 480 0 0 0 chanx_left_out[18]
port 42 nsew signal tristate
flabel metal3 s 0 20952 800 21072 0 FreeSans 480 0 0 0 chanx_left_out[19]
port 43 nsew signal tristate
flabel metal3 s 0 13608 800 13728 0 FreeSans 480 0 0 0 chanx_left_out[1]
port 44 nsew signal tristate
flabel metal3 s 0 14016 800 14136 0 FreeSans 480 0 0 0 chanx_left_out[2]
port 45 nsew signal tristate
flabel metal3 s 0 14424 800 14544 0 FreeSans 480 0 0 0 chanx_left_out[3]
port 46 nsew signal tristate
flabel metal3 s 0 14832 800 14952 0 FreeSans 480 0 0 0 chanx_left_out[4]
port 47 nsew signal tristate
flabel metal3 s 0 15240 800 15360 0 FreeSans 480 0 0 0 chanx_left_out[5]
port 48 nsew signal tristate
flabel metal3 s 0 15648 800 15768 0 FreeSans 480 0 0 0 chanx_left_out[6]
port 49 nsew signal tristate
flabel metal3 s 0 16056 800 16176 0 FreeSans 480 0 0 0 chanx_left_out[7]
port 50 nsew signal tristate
flabel metal3 s 0 16464 800 16584 0 FreeSans 480 0 0 0 chanx_left_out[8]
port 51 nsew signal tristate
flabel metal3 s 0 16872 800 16992 0 FreeSans 480 0 0 0 chanx_left_out[9]
port 52 nsew signal tristate
flabel metal2 s 4066 0 4122 800 0 FreeSans 224 90 0 0 chany_bottom_in[0]
port 53 nsew signal input
flabel metal2 s 8666 0 8722 800 0 FreeSans 224 90 0 0 chany_bottom_in[10]
port 54 nsew signal input
flabel metal2 s 9126 0 9182 800 0 FreeSans 224 90 0 0 chany_bottom_in[11]
port 55 nsew signal input
flabel metal2 s 9586 0 9642 800 0 FreeSans 224 90 0 0 chany_bottom_in[12]
port 56 nsew signal input
flabel metal2 s 10046 0 10102 800 0 FreeSans 224 90 0 0 chany_bottom_in[13]
port 57 nsew signal input
flabel metal2 s 10506 0 10562 800 0 FreeSans 224 90 0 0 chany_bottom_in[14]
port 58 nsew signal input
flabel metal2 s 10966 0 11022 800 0 FreeSans 224 90 0 0 chany_bottom_in[15]
port 59 nsew signal input
flabel metal2 s 11426 0 11482 800 0 FreeSans 224 90 0 0 chany_bottom_in[16]
port 60 nsew signal input
flabel metal2 s 11886 0 11942 800 0 FreeSans 224 90 0 0 chany_bottom_in[17]
port 61 nsew signal input
flabel metal2 s 12346 0 12402 800 0 FreeSans 224 90 0 0 chany_bottom_in[18]
port 62 nsew signal input
flabel metal2 s 12806 0 12862 800 0 FreeSans 224 90 0 0 chany_bottom_in[19]
port 63 nsew signal input
flabel metal2 s 4526 0 4582 800 0 FreeSans 224 90 0 0 chany_bottom_in[1]
port 64 nsew signal input
flabel metal2 s 4986 0 5042 800 0 FreeSans 224 90 0 0 chany_bottom_in[2]
port 65 nsew signal input
flabel metal2 s 5446 0 5502 800 0 FreeSans 224 90 0 0 chany_bottom_in[3]
port 66 nsew signal input
flabel metal2 s 5906 0 5962 800 0 FreeSans 224 90 0 0 chany_bottom_in[4]
port 67 nsew signal input
flabel metal2 s 6366 0 6422 800 0 FreeSans 224 90 0 0 chany_bottom_in[5]
port 68 nsew signal input
flabel metal2 s 6826 0 6882 800 0 FreeSans 224 90 0 0 chany_bottom_in[6]
port 69 nsew signal input
flabel metal2 s 7286 0 7342 800 0 FreeSans 224 90 0 0 chany_bottom_in[7]
port 70 nsew signal input
flabel metal2 s 7746 0 7802 800 0 FreeSans 224 90 0 0 chany_bottom_in[8]
port 71 nsew signal input
flabel metal2 s 8206 0 8262 800 0 FreeSans 224 90 0 0 chany_bottom_in[9]
port 72 nsew signal input
flabel metal2 s 13266 0 13322 800 0 FreeSans 224 90 0 0 chany_bottom_out[0]
port 73 nsew signal tristate
flabel metal2 s 17866 0 17922 800 0 FreeSans 224 90 0 0 chany_bottom_out[10]
port 74 nsew signal tristate
flabel metal2 s 18326 0 18382 800 0 FreeSans 224 90 0 0 chany_bottom_out[11]
port 75 nsew signal tristate
flabel metal2 s 18786 0 18842 800 0 FreeSans 224 90 0 0 chany_bottom_out[12]
port 76 nsew signal tristate
flabel metal2 s 19246 0 19302 800 0 FreeSans 224 90 0 0 chany_bottom_out[13]
port 77 nsew signal tristate
flabel metal2 s 19706 0 19762 800 0 FreeSans 224 90 0 0 chany_bottom_out[14]
port 78 nsew signal tristate
flabel metal2 s 20166 0 20222 800 0 FreeSans 224 90 0 0 chany_bottom_out[15]
port 79 nsew signal tristate
flabel metal2 s 20626 0 20682 800 0 FreeSans 224 90 0 0 chany_bottom_out[16]
port 80 nsew signal tristate
flabel metal2 s 21086 0 21142 800 0 FreeSans 224 90 0 0 chany_bottom_out[17]
port 81 nsew signal tristate
flabel metal2 s 21546 0 21602 800 0 FreeSans 224 90 0 0 chany_bottom_out[18]
port 82 nsew signal tristate
flabel metal2 s 22006 0 22062 800 0 FreeSans 224 90 0 0 chany_bottom_out[19]
port 83 nsew signal tristate
flabel metal2 s 13726 0 13782 800 0 FreeSans 224 90 0 0 chany_bottom_out[1]
port 84 nsew signal tristate
flabel metal2 s 14186 0 14242 800 0 FreeSans 224 90 0 0 chany_bottom_out[2]
port 85 nsew signal tristate
flabel metal2 s 14646 0 14702 800 0 FreeSans 224 90 0 0 chany_bottom_out[3]
port 86 nsew signal tristate
flabel metal2 s 15106 0 15162 800 0 FreeSans 224 90 0 0 chany_bottom_out[4]
port 87 nsew signal tristate
flabel metal2 s 15566 0 15622 800 0 FreeSans 224 90 0 0 chany_bottom_out[5]
port 88 nsew signal tristate
flabel metal2 s 16026 0 16082 800 0 FreeSans 224 90 0 0 chany_bottom_out[6]
port 89 nsew signal tristate
flabel metal2 s 16486 0 16542 800 0 FreeSans 224 90 0 0 chany_bottom_out[7]
port 90 nsew signal tristate
flabel metal2 s 16946 0 17002 800 0 FreeSans 224 90 0 0 chany_bottom_out[8]
port 91 nsew signal tristate
flabel metal2 s 17406 0 17462 800 0 FreeSans 224 90 0 0 chany_bottom_out[9]
port 92 nsew signal tristate
flabel metal2 s 3882 22200 3938 23000 0 FreeSans 224 90 0 0 chany_top_in[0]
port 93 nsew signal input
flabel metal2 s 8482 22200 8538 23000 0 FreeSans 224 90 0 0 chany_top_in[10]
port 94 nsew signal input
flabel metal2 s 8942 22200 8998 23000 0 FreeSans 224 90 0 0 chany_top_in[11]
port 95 nsew signal input
flabel metal2 s 9402 22200 9458 23000 0 FreeSans 224 90 0 0 chany_top_in[12]
port 96 nsew signal input
flabel metal2 s 9862 22200 9918 23000 0 FreeSans 224 90 0 0 chany_top_in[13]
port 97 nsew signal input
flabel metal2 s 10322 22200 10378 23000 0 FreeSans 224 90 0 0 chany_top_in[14]
port 98 nsew signal input
flabel metal2 s 10782 22200 10838 23000 0 FreeSans 224 90 0 0 chany_top_in[15]
port 99 nsew signal input
flabel metal2 s 11242 22200 11298 23000 0 FreeSans 224 90 0 0 chany_top_in[16]
port 100 nsew signal input
flabel metal2 s 11702 22200 11758 23000 0 FreeSans 224 90 0 0 chany_top_in[17]
port 101 nsew signal input
flabel metal2 s 12162 22200 12218 23000 0 FreeSans 224 90 0 0 chany_top_in[18]
port 102 nsew signal input
flabel metal2 s 12622 22200 12678 23000 0 FreeSans 224 90 0 0 chany_top_in[19]
port 103 nsew signal input
flabel metal2 s 4342 22200 4398 23000 0 FreeSans 224 90 0 0 chany_top_in[1]
port 104 nsew signal input
flabel metal2 s 4802 22200 4858 23000 0 FreeSans 224 90 0 0 chany_top_in[2]
port 105 nsew signal input
flabel metal2 s 5262 22200 5318 23000 0 FreeSans 224 90 0 0 chany_top_in[3]
port 106 nsew signal input
flabel metal2 s 5722 22200 5778 23000 0 FreeSans 224 90 0 0 chany_top_in[4]
port 107 nsew signal input
flabel metal2 s 6182 22200 6238 23000 0 FreeSans 224 90 0 0 chany_top_in[5]
port 108 nsew signal input
flabel metal2 s 6642 22200 6698 23000 0 FreeSans 224 90 0 0 chany_top_in[6]
port 109 nsew signal input
flabel metal2 s 7102 22200 7158 23000 0 FreeSans 224 90 0 0 chany_top_in[7]
port 110 nsew signal input
flabel metal2 s 7562 22200 7618 23000 0 FreeSans 224 90 0 0 chany_top_in[8]
port 111 nsew signal input
flabel metal2 s 8022 22200 8078 23000 0 FreeSans 224 90 0 0 chany_top_in[9]
port 112 nsew signal input
flabel metal2 s 13082 22200 13138 23000 0 FreeSans 224 90 0 0 chany_top_out[0]
port 113 nsew signal tristate
flabel metal2 s 17682 22200 17738 23000 0 FreeSans 224 90 0 0 chany_top_out[10]
port 114 nsew signal tristate
flabel metal2 s 18142 22200 18198 23000 0 FreeSans 224 90 0 0 chany_top_out[11]
port 115 nsew signal tristate
flabel metal2 s 18602 22200 18658 23000 0 FreeSans 224 90 0 0 chany_top_out[12]
port 116 nsew signal tristate
flabel metal2 s 19062 22200 19118 23000 0 FreeSans 224 90 0 0 chany_top_out[13]
port 117 nsew signal tristate
flabel metal2 s 19522 22200 19578 23000 0 FreeSans 224 90 0 0 chany_top_out[14]
port 118 nsew signal tristate
flabel metal2 s 19982 22200 20038 23000 0 FreeSans 224 90 0 0 chany_top_out[15]
port 119 nsew signal tristate
flabel metal2 s 20442 22200 20498 23000 0 FreeSans 224 90 0 0 chany_top_out[16]
port 120 nsew signal tristate
flabel metal2 s 20902 22200 20958 23000 0 FreeSans 224 90 0 0 chany_top_out[17]
port 121 nsew signal tristate
flabel metal2 s 21362 22200 21418 23000 0 FreeSans 224 90 0 0 chany_top_out[18]
port 122 nsew signal tristate
flabel metal2 s 21822 22200 21878 23000 0 FreeSans 224 90 0 0 chany_top_out[19]
port 123 nsew signal tristate
flabel metal2 s 13542 22200 13598 23000 0 FreeSans 224 90 0 0 chany_top_out[1]
port 124 nsew signal tristate
flabel metal2 s 14002 22200 14058 23000 0 FreeSans 224 90 0 0 chany_top_out[2]
port 125 nsew signal tristate
flabel metal2 s 14462 22200 14518 23000 0 FreeSans 224 90 0 0 chany_top_out[3]
port 126 nsew signal tristate
flabel metal2 s 14922 22200 14978 23000 0 FreeSans 224 90 0 0 chany_top_out[4]
port 127 nsew signal tristate
flabel metal2 s 15382 22200 15438 23000 0 FreeSans 224 90 0 0 chany_top_out[5]
port 128 nsew signal tristate
flabel metal2 s 15842 22200 15898 23000 0 FreeSans 224 90 0 0 chany_top_out[6]
port 129 nsew signal tristate
flabel metal2 s 16302 22200 16358 23000 0 FreeSans 224 90 0 0 chany_top_out[7]
port 130 nsew signal tristate
flabel metal2 s 16762 22200 16818 23000 0 FreeSans 224 90 0 0 chany_top_out[8]
port 131 nsew signal tristate
flabel metal2 s 17222 22200 17278 23000 0 FreeSans 224 90 0 0 chany_top_out[9]
port 132 nsew signal tristate
flabel metal3 s 0 1776 800 1896 0 FreeSans 480 0 0 0 left_bottom_grid_pin_34_
port 133 nsew signal input
flabel metal3 s 0 2184 800 2304 0 FreeSans 480 0 0 0 left_bottom_grid_pin_35_
port 134 nsew signal input
flabel metal3 s 0 2592 800 2712 0 FreeSans 480 0 0 0 left_bottom_grid_pin_36_
port 135 nsew signal input
flabel metal3 s 0 3000 800 3120 0 FreeSans 480 0 0 0 left_bottom_grid_pin_37_
port 136 nsew signal input
flabel metal3 s 0 3408 800 3528 0 FreeSans 480 0 0 0 left_bottom_grid_pin_38_
port 137 nsew signal input
flabel metal3 s 0 3816 800 3936 0 FreeSans 480 0 0 0 left_bottom_grid_pin_39_
port 138 nsew signal input
flabel metal3 s 0 4224 800 4344 0 FreeSans 480 0 0 0 left_bottom_grid_pin_40_
port 139 nsew signal input
flabel metal3 s 0 4632 800 4752 0 FreeSans 480 0 0 0 left_bottom_grid_pin_41_
port 140 nsew signal input
flabel metal2 s 22282 22200 22338 23000 0 FreeSans 224 90 0 0 prog_clk_0_N_in
port 141 nsew signal input
flabel metal2 s 202 22200 258 23000 0 FreeSans 224 90 0 0 top_left_grid_pin_42_
port 142 nsew signal input
flabel metal2 s 662 22200 718 23000 0 FreeSans 224 90 0 0 top_left_grid_pin_43_
port 143 nsew signal input
flabel metal2 s 1122 22200 1178 23000 0 FreeSans 224 90 0 0 top_left_grid_pin_44_
port 144 nsew signal input
flabel metal2 s 1582 22200 1638 23000 0 FreeSans 224 90 0 0 top_left_grid_pin_45_
port 145 nsew signal input
flabel metal2 s 2042 22200 2098 23000 0 FreeSans 224 90 0 0 top_left_grid_pin_46_
port 146 nsew signal input
flabel metal2 s 2502 22200 2558 23000 0 FreeSans 224 90 0 0 top_left_grid_pin_47_
port 147 nsew signal input
flabel metal2 s 2962 22200 3018 23000 0 FreeSans 224 90 0 0 top_left_grid_pin_48_
port 148 nsew signal input
flabel metal2 s 3422 22200 3478 23000 0 FreeSans 224 90 0 0 top_left_grid_pin_49_
port 149 nsew signal input
flabel metal2 s 22742 22200 22798 23000 0 FreeSans 224 90 0 0 top_right_grid_pin_1_
port 150 nsew signal input
<< properties >>
string FIXED_BBOX 0 0 23000 23000
<< end >>
