* NGSPICE file created from sb_2__0_.ext - technology: sky130A

* Black-box entry subcircuit for sky130_fd_sc_hd__fill_2 abstract view
.subckt sky130_fd_sc_hd__fill_2 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_12 abstract view
.subckt sky130_fd_sc_hd__decap_12 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dfxtp_1 abstract view
.subckt sky130_fd_sc_hd__dfxtp_1 CLK D VGND VNB VPB VPWR Q
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_8 abstract view
.subckt sky130_fd_sc_hd__decap_8 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_3 abstract view
.subckt sky130_fd_sc_hd__decap_3 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__diode_2 abstract view
.subckt sky130_fd_sc_hd__diode_2 DIODE VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__conb_1 abstract view
.subckt sky130_fd_sc_hd__conb_1 VGND VNB VPB VPWR HI LO
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_4 abstract view
.subckt sky130_fd_sc_hd__decap_4 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_2 abstract view
.subckt sky130_fd_sc_hd__clkbuf_2 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__tapvpwrvgnd_1 abstract view
.subckt sky130_fd_sc_hd__tapvpwrvgnd_1 VGND VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_6 abstract view
.subckt sky130_fd_sc_hd__decap_6 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__fill_1 abstract view
.subckt sky130_fd_sc_hd__fill_1 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_1 abstract view
.subckt sky130_fd_sc_hd__clkbuf_1 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__mux2_1 abstract view
.subckt sky130_fd_sc_hd__mux2_1 A0 A1 S VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_16 abstract view
.subckt sky130_fd_sc_hd__clkbuf_16 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__buf_8 abstract view
.subckt sky130_fd_sc_hd__buf_8 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__buf_1 abstract view
.subckt sky130_fd_sc_hd__buf_1 A VGND VNB VPB VPWR X
.ends

.subckt sb_2__0_ ccff_head ccff_tail chanx_left_in[0] chanx_left_in[10] chanx_left_in[11]
+ chanx_left_in[12] chanx_left_in[13] chanx_left_in[14] chanx_left_in[15] chanx_left_in[16]
+ chanx_left_in[17] chanx_left_in[18] chanx_left_in[19] chanx_left_in[1] chanx_left_in[2]
+ chanx_left_in[3] chanx_left_in[4] chanx_left_in[5] chanx_left_in[6] chanx_left_in[7]
+ chanx_left_in[8] chanx_left_in[9] chanx_left_out[0] chanx_left_out[10] chanx_left_out[11]
+ chanx_left_out[12] chanx_left_out[13] chanx_left_out[14] chanx_left_out[15] chanx_left_out[16]
+ chanx_left_out[17] chanx_left_out[18] chanx_left_out[19] chanx_left_out[1] chanx_left_out[2]
+ chanx_left_out[3] chanx_left_out[4] chanx_left_out[5] chanx_left_out[6] chanx_left_out[7]
+ chanx_left_out[8] chanx_left_out[9] chany_top_in[0] chany_top_in[10] chany_top_in[11]
+ chany_top_in[12] chany_top_in[13] chany_top_in[14] chany_top_in[15] chany_top_in[16]
+ chany_top_in[17] chany_top_in[18] chany_top_in[19] chany_top_in[1] chany_top_in[2]
+ chany_top_in[3] chany_top_in[4] chany_top_in[5] chany_top_in[6] chany_top_in[7]
+ chany_top_in[8] chany_top_in[9] chany_top_out[0] chany_top_out[10] chany_top_out[11]
+ chany_top_out[12] chany_top_out[13] chany_top_out[14] chany_top_out[15] chany_top_out[16]
+ chany_top_out[17] chany_top_out[18] chany_top_out[19] chany_top_out[1] chany_top_out[2]
+ chany_top_out[3] chany_top_out[4] chany_top_out[5] chany_top_out[6] chany_top_out[7]
+ chany_top_out[8] chany_top_out[9] left_bottom_grid_pin_11_ left_bottom_grid_pin_13_
+ left_bottom_grid_pin_15_ left_bottom_grid_pin_17_ left_bottom_grid_pin_1_ left_bottom_grid_pin_3_
+ left_bottom_grid_pin_5_ left_bottom_grid_pin_7_ left_bottom_grid_pin_9_ prog_clk_0_N_in
+ top_left_grid_pin_42_ top_left_grid_pin_43_ top_left_grid_pin_44_ top_left_grid_pin_45_
+ top_left_grid_pin_46_ top_left_grid_pin_47_ top_left_grid_pin_48_ top_left_grid_pin_49_
+ top_right_grid_pin_1_ VPWR VGND
XFILLER_22_144 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_26_30 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_9_115 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xmem_left_track_17.sky130_fd_sc_hd__dfxtp_1_0_ clkbuf_3_3_0_mem_left_track_1.prog_clk/X
+ mux_left_track_15.mux_l2_in_0_/S VGND VGND VPWR VPWR mux_left_track_17.mux_l1_in_0_/S
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_8_192 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_12_10 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_12_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_12_87 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_5_151 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_5_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_mux_top_track_0.mux_l1_in_0__A0 input53/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_062_ VGND VGND VPWR VPWR _062_/HI _062_/LO sky130_fd_sc_hd__conb_1
XANTENNA_input55_A top_left_grid_pin_46_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_9_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_21_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_18_20 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_7_213 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_11_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_045_ VGND VGND VPWR VPWR _045_/HI _045_/LO sky130_fd_sc_hd__conb_1
XFILLER_20_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_20_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_20_87 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_20_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_input18_A chanx_left_in[6] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_6_78 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_19_172 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_1_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_17_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_25_131 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_15_76 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xoutput75 _072_/X VGND VGND VPWR VPWR chanx_left_out[4] sky130_fd_sc_hd__clkbuf_2
Xoutput64 _080_/X VGND VGND VPWR VPWR chanx_left_out[12] sky130_fd_sc_hd__clkbuf_2
Xoutput86 _102_/X VGND VGND VPWR VPWR chany_top_out[14] sky130_fd_sc_hd__clkbuf_2
Xoutput97 _094_/X VGND VGND VPWR VPWR chany_top_out[6] sky130_fd_sc_hd__clkbuf_2
XPHY_170 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_192 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_181 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_22_101 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_22_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_9_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_13_101 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_26_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_9_127 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_3_13 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_5_196 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_5_163 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA_mux_top_track_0.mux_l1_in_0__A1 input51/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_23_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_23_43 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_2_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_23_76 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_061_ VGND VGND VPWR VPWR _061_/HI _061_/LO sky130_fd_sc_hd__conb_1
XFILLER_2_144 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_input48_A left_bottom_grid_pin_5_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_25 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_9_89 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_9_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_20_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmux_left_track_9.sky130_fd_sc_hd__buf_4_0_ mux_left_track_9.mux_l2_in_0_/X VGND VGND
+ VPWR VPWR _072_/A sky130_fd_sc_hd__clkbuf_1
XFILLER_18_10 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_044_ VGND VGND VPWR VPWR _044_/HI _044_/LO sky130_fd_sc_hd__conb_1
XFILLER_20_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_20_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmux_left_track_31.sky130_fd_sc_hd__buf_4_0_ mux_left_track_31.mux_l2_in_0_/X VGND
+ VGND VPWR VPWR _083_/A sky130_fd_sc_hd__clkbuf_1
Xmux_top_track_10.mux_l2_in_0_ _043_/HI mux_top_track_10.mux_l1_in_0_/X mux_top_track_10.mux_l2_in_0_/S
+ VGND VGND VPWR VPWR mux_top_track_10.mux_l2_in_0_/X sky130_fd_sc_hd__mux2_1
Xmem_left_track_35.sky130_fd_sc_hd__dfxtp_1_1_ clkbuf_3_2_0_mem_left_track_1.prog_clk/X
+ mux_left_track_35.mux_l1_in_0_/S VGND VGND VPWR VPWR mux_left_track_35.mux_l2_in_0_/S
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_25_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xoutput76 _073_/X VGND VGND VPWR VPWR chanx_left_out[5] sky130_fd_sc_hd__clkbuf_2
Xoutput65 _081_/X VGND VGND VPWR VPWR chanx_left_out[13] sky130_fd_sc_hd__clkbuf_2
Xoutput98 _095_/X VGND VGND VPWR VPWR chany_top_out[7] sky130_fd_sc_hd__clkbuf_2
Xoutput87 _103_/X VGND VGND VPWR VPWR chany_top_out[15] sky130_fd_sc_hd__clkbuf_2
XANTENNA_input30_A chany_top_in[17] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_193 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_160 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_171 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_31_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_31_146 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_31_157 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_182 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_31_168 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xmux_left_track_25.sky130_fd_sc_hd__buf_4_0_ mux_left_track_25.mux_l2_in_0_/X VGND
+ VGND VPWR VPWR _080_/A sky130_fd_sc_hd__clkbuf_1
XFILLER_22_179 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_9_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_13_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_26_87 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_26_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_3_58 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_5_6 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmux_left_track_19.sky130_fd_sc_hd__buf_4_0_ mux_left_track_19.mux_l2_in_0_/X VGND
+ VGND VPWR VPWR _077_/A sky130_fd_sc_hd__clkbuf_1
Xmux_left_track_7.mux_l3_in_0_ mux_left_track_7.mux_l2_in_1_/X mux_left_track_7.mux_l2_in_0_/X
+ mux_left_track_7.mux_l3_in_0_/S VGND VGND VPWR VPWR mux_left_track_7.mux_l3_in_0_/X
+ sky130_fd_sc_hd__mux2_1
Xclkbuf_0_mem_left_track_1.prog_clk prog_clk_0_FTB00/X VGND VGND VPWR VPWR clkbuf_0_mem_left_track_1.prog_clk/X
+ sky130_fd_sc_hd__clkbuf_16
Xmem_top_track_10.sky130_fd_sc_hd__dfxtp_1_1_ clkbuf_3_4_0_mem_left_track_1.prog_clk/X
+ mux_top_track_10.mux_l1_in_0_/S VGND VGND VPWR VPWR mux_top_track_10.mux_l2_in_0_/S
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_23_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_3_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_2_156 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_2_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_060_ VGND VGND VPWR VPWR _060_/HI _060_/LO sky130_fd_sc_hd__conb_1
XFILLER_0_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_59 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xclkbuf_2_0_0_mem_left_track_1.prog_clk clkbuf_2_1_0_mem_left_track_1.prog_clk/A VGND
+ VGND VPWR VPWR clkbuf_3_1_0_mem_left_track_1.prog_clk/A sky130_fd_sc_hd__clkbuf_1
XFILLER_7_204 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmux_left_track_7.mux_l2_in_1_ _040_/HI input44/X mux_left_track_7.mux_l2_in_1_/S
+ VGND VGND VPWR VPWR mux_left_track_7.mux_l2_in_1_/X sky130_fd_sc_hd__mux2_1
X_043_ VGND VGND VPWR VPWR _043_/HI _043_/LO sky130_fd_sc_hd__conb_1
XFILLER_22_9 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_29_108 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_20_23 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_28_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_28_174 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_29_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_29_76 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_29_87 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_29_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmem_left_track_35.sky130_fd_sc_hd__dfxtp_1_0_ clkbuf_3_2_0_mem_left_track_1.prog_clk/X
+ mux_left_track_33.mux_l2_in_0_/S VGND VGND VPWR VPWR mux_left_track_35.mux_l1_in_0_/S
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_15_34 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_15_45 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_31_33 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_31_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xoutput77 _074_/X VGND VGND VPWR VPWR chanx_left_out[6] sky130_fd_sc_hd__clkbuf_2
Xoutput66 _082_/X VGND VGND VPWR VPWR chanx_left_out[14] sky130_fd_sc_hd__clkbuf_2
Xoutput99 _096_/X VGND VGND VPWR VPWR chany_top_out[8] sky130_fd_sc_hd__clkbuf_2
Xoutput88 _104_/X VGND VGND VPWR VPWR chany_top_out[16] sky130_fd_sc_hd__clkbuf_2
XANTENNA_input23_A chany_top_in[10] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_16_144 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_150 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_161 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_172 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_31_136 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_183 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_output91_A _107_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xmux_top_track_10.mux_l1_in_0_ input8/X input52/X mux_top_track_10.mux_l1_in_0_/S
+ VGND VGND VPWR VPWR mux_top_track_10.mux_l1_in_0_/X sky130_fd_sc_hd__mux2_1
XANTENNA_mux_top_track_2.mux_l1_in_1__A0 input58/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xmux_top_track_22.mux_l2_in_0_ _050_/HI mux_top_track_22.mux_l1_in_0_/X mux_top_track_22.mux_l2_in_0_/S
+ VGND VGND VPWR VPWR mux_top_track_22.mux_l2_in_0_/X sky130_fd_sc_hd__mux2_1
XFILLER_12_180 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xclkbuf_2_3_0_mem_left_track_1.prog_clk clkbuf_2_3_0_mem_left_track_1.prog_clk/A VGND
+ VGND VPWR VPWR clkbuf_3_7_0_mem_left_track_1.prog_clk/A sky130_fd_sc_hd__clkbuf_1
XFILLER_12_24 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xmux_left_track_15.mux_l2_in_0_ _059_/HI mux_left_track_15.mux_l1_in_0_/X mux_left_track_15.mux_l2_in_0_/S
+ VGND VGND VPWR VPWR mux_left_track_15.mux_l2_in_0_/X sky130_fd_sc_hd__mux2_1
Xmem_top_track_10.sky130_fd_sc_hd__dfxtp_1_0_ clkbuf_3_1_0_mem_left_track_1.prog_clk/X
+ mux_top_track_8.mux_l2_in_0_/S VGND VGND VPWR VPWR mux_top_track_10.mux_l1_in_0_/S
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_2_168 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_2_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xprog_clk_0_FTB00 prog_clk_0_N_in VGND VGND VPWR VPWR prog_clk_0_FTB00/X sky130_fd_sc_hd__buf_8
XFILLER_9_58 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_9_47 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_9_36 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_9_25 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_29_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_20_201 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_18_89 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xmux_left_track_7.mux_l2_in_0_ mux_left_track_7.mux_l1_in_1_/X mux_left_track_7.mux_l1_in_0_/X
+ mux_left_track_7.mux_l2_in_1_/S VGND VGND VPWR VPWR mux_left_track_7.mux_l2_in_0_/X
+ sky130_fd_sc_hd__mux2_1
X_042_ VGND VGND VPWR VPWR _042_/HI _042_/LO sky130_fd_sc_hd__conb_1
XANTENNA_input53_A top_left_grid_pin_44_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_1_70 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xmux_top_track_0.mux_l3_in_0_ mux_top_track_0.mux_l2_in_1_/X mux_top_track_0.mux_l2_in_0_/X
+ mux_top_track_0.mux_l3_in_0_/S VGND VGND VPWR VPWR mux_top_track_0.mux_l3_in_0_/X
+ sky130_fd_sc_hd__mux2_1
XFILLER_20_13 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_28_131 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_28_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_13_6 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmem_top_track_16.sky130_fd_sc_hd__dfxtp_1_1_ clkbuf_3_7_0_mem_left_track_1.prog_clk/X
+ mux_top_track_16.mux_l1_in_0_/S VGND VGND VPWR VPWR mux_top_track_16.mux_l2_in_0_/S
+ sky130_fd_sc_hd__dfxtp_1
Xmux_left_track_7.mux_l1_in_1_ input42/X input49/X mux_left_track_7.mux_l1_in_1_/S
+ VGND VGND VPWR VPWR mux_left_track_7.mux_l1_in_1_/X sky130_fd_sc_hd__mux2_1
XFILLER_25_112 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_31_67 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xoutput78 _075_/X VGND VGND VPWR VPWR chanx_left_out[7] sky130_fd_sc_hd__clkbuf_2
Xoutput67 _083_/X VGND VGND VPWR VPWR chanx_left_out[15] sky130_fd_sc_hd__clkbuf_2
Xoutput89 _105_/X VGND VGND VPWR VPWR chany_top_out[17] sky130_fd_sc_hd__clkbuf_2
XANTENNA_input16_A chanx_left_in[4] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_140 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_151 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_162 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_173 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_184 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xmux_top_track_0.mux_l2_in_1_ _042_/HI mux_top_track_0.mux_l1_in_2_/X mux_top_track_0.mux_l2_in_1_/S
+ VGND VGND VPWR VPWR mux_top_track_0.mux_l2_in_1_/X sky130_fd_sc_hd__mux2_1
XANTENNA_mux_left_track_1.mux_l1_in_1__A0 input50/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_input8_A chanx_left_in[15] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mux_top_track_2.mux_l1_in_1__A1 input56/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_13_115 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_26_67 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_26_78 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_21_170 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xmux_top_track_22.sky130_fd_sc_hd__buf_4_0_ mux_top_track_22.mux_l2_in_0_/X VGND VGND
+ VPWR VPWR _099_/A sky130_fd_sc_hd__clkbuf_1
XFILLER_12_192 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xmux_top_track_0.mux_l1_in_2_ input2/X input59/X mux_top_track_0.mux_l1_in_2_/S VGND
+ VGND VPWR VPWR mux_top_track_0.mux_l1_in_2_/X sky130_fd_sc_hd__mux2_1
XFILLER_32_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmux_top_track_22.mux_l1_in_0_ input21/X input58/X mux_top_track_22.mux_l1_in_0_/S
+ VGND VGND VPWR VPWR mux_top_track_22.mux_l1_in_0_/X sky130_fd_sc_hd__mux2_1
Xmux_top_track_16.sky130_fd_sc_hd__buf_4_0_ mux_top_track_16.mux_l2_in_0_/X VGND VGND
+ VPWR VPWR _096_/A sky130_fd_sc_hd__clkbuf_1
XFILLER_9_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_14_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_13_90 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_20_213 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xmux_left_track_15.mux_l1_in_0_ input49/X input26/X mux_left_track_15.mux_l1_in_0_/S
+ VGND VGND VPWR VPWR mux_left_track_15.mux_l1_in_0_/X sky130_fd_sc_hd__mux2_1
XFILLER_18_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_18_79 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_041_ VGND VGND VPWR VPWR _041_/HI _041_/LO sky130_fd_sc_hd__conb_1
XANTENNA_input46_A left_bottom_grid_pin_1_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xmux_left_track_27.mux_l2_in_0_ _065_/HI mux_left_track_27.mux_l1_in_0_/X mux_left_track_27.mux_l2_in_0_/S
+ VGND VGND VPWR VPWR mux_left_track_27.mux_l2_in_0_/X sky130_fd_sc_hd__mux2_1
XFILLER_1_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_20_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_3_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xmem_top_track_16.sky130_fd_sc_hd__dfxtp_1_0_ clkbuf_3_5_0_mem_left_track_1.prog_clk/X
+ mux_top_track_14.mux_l2_in_0_/S VGND VGND VPWR VPWR mux_top_track_16.mux_l1_in_0_/S
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_20_8 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmux_left_track_7.mux_l1_in_0_ input47/X input30/X mux_left_track_7.mux_l1_in_1_/S
+ VGND VGND VPWR VPWR mux_left_track_7.mux_l1_in_0_/X sky130_fd_sc_hd__mux2_1
XFILLER_25_102 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_25_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_33_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_15_58 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_25_168 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xmux_top_track_0.sky130_fd_sc_hd__buf_4_0_ mux_top_track_0.mux_l3_in_0_/X VGND VGND
+ VPWR VPWR _088_/A sky130_fd_sc_hd__clkbuf_1
Xoutput79 _076_/X VGND VGND VPWR VPWR chanx_left_out[8] sky130_fd_sc_hd__clkbuf_2
Xoutput68 _084_/X VGND VGND VPWR VPWR chanx_left_out[16] sky130_fd_sc_hd__clkbuf_2
XPHY_130 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_141 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_152 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_31_127 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_163 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_174 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_185 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xmux_top_track_0.mux_l2_in_0_ mux_top_track_0.mux_l1_in_1_/X mux_top_track_0.mux_l1_in_0_/X
+ mux_top_track_0.mux_l2_in_1_/S VGND VGND VPWR VPWR mux_top_track_0.mux_l2_in_0_/X
+ sky130_fd_sc_hd__mux2_1
XFILLER_15_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_22_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_7_70 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_30_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_mux_left_track_1.mux_l1_in_1__A1 input48/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_13_127 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_26_35 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_3_17 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_mux_top_track_22.mux_l1_in_0__A0 input21/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_12_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmux_top_track_0.mux_l1_in_1_ input57/X input55/X mux_top_track_0.mux_l1_in_2_/S VGND
+ VGND VPWR VPWR mux_top_track_0.mux_l1_in_1_/X sky130_fd_sc_hd__mux2_1
Xmem_left_track_21.sky130_fd_sc_hd__dfxtp_1_1_ clkbuf_3_3_0_mem_left_track_1.prog_clk/X
+ mux_left_track_21.mux_l1_in_0_/S VGND VGND VPWR VPWR mux_left_track_21.mux_l2_in_0_/S
+ sky130_fd_sc_hd__dfxtp_1
XANTENNA_mux_top_track_14.mux_l1_in_0__A1 input54/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_23_14 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_23_211 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_23_58 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_23_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_mux_top_track_6.mux_l1_in_0__A0 input54/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_18_25 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_1_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_040_ VGND VGND VPWR VPWR _040_/HI _040_/LO sky130_fd_sc_hd__conb_1
XANTENNA_input39_A chany_top_in[7] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_1_94 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_29_35 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_28_188 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_6_28 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_19_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_19_144 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_19_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_19_188 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_19_199 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_25_158 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xmux_left_track_27.mux_l1_in_0_ input47/X input39/X mux_left_track_27.mux_l1_in_0_/S
+ VGND VGND VPWR VPWR mux_left_track_27.mux_l1_in_0_/X sky130_fd_sc_hd__mux2_1
XFILLER_31_58 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xoutput69 _085_/X VGND VGND VPWR VPWR chanx_left_out[17] sky130_fd_sc_hd__clkbuf_2
XPHY_120 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_16_136 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_131 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_142 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_153 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_164 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_175 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_31_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmux_left_track_39.mux_l2_in_0_ _038_/HI mux_left_track_39.mux_l1_in_0_/X output60/A
+ VGND VGND VPWR VPWR mux_left_track_39.mux_l2_in_0_/X sky130_fd_sc_hd__mux2_1
XPHY_186 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_0 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_11_5 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_30_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_30_183 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_7_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_26_14 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_13_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_26_25 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_26_58 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_21_172 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_3_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_input21_A chanx_left_in[9] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mux_top_track_22.mux_l1_in_0__A1 input58/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_27_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_mux_left_track_15.mux_l1_in_0__A0 input49/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xmux_top_track_0.mux_l1_in_0_ input53/X input51/X mux_top_track_0.mux_l1_in_2_/S VGND
+ VGND VPWR VPWR mux_top_track_0.mux_l1_in_0_/X sky130_fd_sc_hd__mux2_1
Xmem_left_track_21.sky130_fd_sc_hd__dfxtp_1_0_ clkbuf_3_2_0_mem_left_track_1.prog_clk/X
+ mux_left_track_19.mux_l2_in_0_/S VGND VGND VPWR VPWR mux_left_track_21.mux_l1_in_0_/S
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_14_201 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_mux_top_track_6.mux_l1_in_0__A1 input52/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_18_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_18_48 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_27_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_099_ _099_/A VGND VGND VPWR VPWR _099_/X sky130_fd_sc_hd__clkbuf_1
Xmem_left_track_27.sky130_fd_sc_hd__dfxtp_1_1_ clkbuf_3_0_0_mem_left_track_1.prog_clk/X
+ mux_left_track_27.mux_l1_in_0_/S VGND VGND VPWR VPWR mux_left_track_27.mux_l2_in_0_/S
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_20_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_28_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_input51_A top_left_grid_pin_42_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_19_101 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_19_112 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_19_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_15_16 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_15_49 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_25_115 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_25_126 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_31_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_31_37 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_16_115 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_187 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_110 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_121 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_132 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_143 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_154 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_165 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_176 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_21_92 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_1 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_7_94 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_26_48 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_input14_A chanx_left_in[2] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_8_144 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_8_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_12_140 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_16_92 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xclkbuf_1_0_0_mem_left_track_1.prog_clk clkbuf_0_mem_left_track_1.prog_clk/X VGND
+ VGND VPWR VPWR clkbuf_2_1_0_mem_left_track_1.prog_clk/A sky130_fd_sc_hd__clkbuf_1
XFILLER_12_28 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_input6_A chanx_left_in[13] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xmux_left_track_39.mux_l1_in_0_ input44/X input33/X mux_left_track_39.mux_l1_in_0_/S
+ VGND VGND VPWR VPWR mux_left_track_39.mux_l1_in_0_/X sky130_fd_sc_hd__mux2_1
XFILLER_17_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_27_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_4_180 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_14_213 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_1_172 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_7_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_24_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_098_ _098_/A VGND VGND VPWR VPWR _098_/X sky130_fd_sc_hd__clkbuf_1
Xmem_left_track_27.sky130_fd_sc_hd__dfxtp_1_0_ clkbuf_3_0_0_mem_left_track_1.prog_clk/X
+ mux_left_track_25.mux_l2_in_0_/S VGND VGND VPWR VPWR mux_left_track_27.mux_l1_in_0_/S
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_29_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_28_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_28_146 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_input44_A left_bottom_grid_pin_15_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mux_left_track_31.mux_l1_in_0__A0 input49/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_19_70 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_33_160 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_204 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_100 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_188 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_111 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_122 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_133 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_144 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_155 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_166 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_177 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_22_119 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_30_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmux_left_track_5.sky130_fd_sc_hd__buf_4_0_ mux_left_track_5.mux_l3_in_0_/X VGND VGND
+ VPWR VPWR _070_/A sky130_fd_sc_hd__clkbuf_1
XFILLER_16_60 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_16_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_8_156 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_8_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_32_92 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_5_115 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xmem_left_track_1.sky130_fd_sc_hd__dfxtp_1_2_ clkbuf_3_0_0_mem_left_track_1.prog_clk/X
+ mux_left_track_1.mux_l2_in_1_/S VGND VGND VPWR VPWR mux_left_track_1.mux_l3_in_0_/S
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_32_203 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_4_192 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_4_30 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_3_9 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_9_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_1_151 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_1_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xmux_left_track_21.sky130_fd_sc_hd__buf_4_0_ mux_left_track_21.mux_l2_in_0_/X VGND
+ VGND VPWR VPWR _078_/A sky130_fd_sc_hd__clkbuf_1
X_097_ _097_/A VGND VGND VPWR VPWR _097_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_20_18 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_29_49 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmem_top_track_4.sky130_fd_sc_hd__dfxtp_1_2_ clkbuf_3_6_0_mem_left_track_1.prog_clk/X
+ mux_top_track_4.mux_l2_in_1_/S VGND VGND VPWR VPWR mux_top_track_4.mux_l3_in_0_/S
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_28_103 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_28_136 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_28_158 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_28_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmux_left_track_15.sky130_fd_sc_hd__buf_4_0_ mux_left_track_15.mux_l2_in_0_/X VGND
+ VGND VPWR VPWR _075_/A sky130_fd_sc_hd__clkbuf_1
XANTENNA_mux_top_track_24.mux_l1_in_1__A1 input20/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_10_84 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_input37_A chany_top_in[5] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_19_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_32_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_33_172 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_216 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_101 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_112 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_123 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_134 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_31_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_189 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_145 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_156 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_24_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_167 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_178 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xmux_left_track_3.mux_l3_in_0_ mux_left_track_3.mux_l2_in_1_/X mux_left_track_3.mux_l2_in_0_/X
+ mux_left_track_3.mux_l3_in_0_/S VGND VGND VPWR VPWR mux_left_track_3.mux_l3_in_0_/X
+ sky130_fd_sc_hd__mux2_1
XPHY_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_15_172 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_30_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_13_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_21_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_12_120 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_16_50 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_8_168 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_8_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA_mux_left_track_7.mux_l1_in_1__A0 input42/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_5_127 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xmem_left_track_1.sky130_fd_sc_hd__dfxtp_1_1_ clkbuf_3_0_0_mem_left_track_1.prog_clk/X
+ mux_left_track_1.mux_l1_in_2_/S VGND VGND VPWR VPWR mux_left_track_1.mux_l2_in_1_/S
+ sky130_fd_sc_hd__dfxtp_1
Xmux_left_track_3.mux_l2_in_1_ _067_/HI input44/X mux_left_track_3.mux_l2_in_1_/S
+ VGND VGND VPWR VPWR mux_left_track_3.mux_l2_in_1_/X sky130_fd_sc_hd__mux2_1
XFILLER_27_60 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_32_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_4_42 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_13_73 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_1_163 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_1_196 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_29_9 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_6_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_096_ _096_/A VGND VGND VPWR VPWR _096_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_1_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmem_left_track_7.sky130_fd_sc_hd__dfxtp_1_2_ clkbuf_3_0_0_mem_left_track_1.prog_clk/X
+ mux_left_track_7.mux_l2_in_1_/S VGND VGND VPWR VPWR mux_left_track_7.mux_l3_in_0_/S
+ sky130_fd_sc_hd__dfxtp_1
Xmux_top_track_16.mux_l2_in_0_ _046_/HI mux_top_track_16.mux_l1_in_0_/X mux_top_track_16.mux_l2_in_0_/S
+ VGND VGND VPWR VPWR mux_top_track_16.mux_l2_in_0_/X sky130_fd_sc_hd__mux2_1
XFILLER_29_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xmem_top_track_4.sky130_fd_sc_hd__dfxtp_1_1_ clkbuf_3_6_0_mem_left_track_1.prog_clk/X
+ mux_top_track_4.mux_l1_in_2_/S VGND VGND VPWR VPWR mux_top_track_4.mux_l2_in_1_/S
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_10_30 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_19_104 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_19_115 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_27_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_079_ _079_/A VGND VGND VPWR VPWR _079_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_25_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_18_192 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_33_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_33_140 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_102 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_113 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_124 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_135 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_146 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_157 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xmux_left_track_11.mux_l2_in_0_ _057_/HI mux_left_track_11.mux_l1_in_0_/X mux_left_track_11.mux_l2_in_0_/S
+ VGND VGND VPWR VPWR mux_left_track_11.mux_l2_in_0_/X sky130_fd_sc_hd__mux2_1
XFILLER_21_73 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_168 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_179 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xmem_top_track_20.sky130_fd_sc_hd__dfxtp_1_1_ clkbuf_3_7_0_mem_left_track_1.prog_clk/X
+ mux_top_track_20.mux_l1_in_0_/S VGND VGND VPWR VPWR mux_top_track_20.mux_l2_in_0_/S
+ sky130_fd_sc_hd__dfxtp_1
Xmux_left_track_37.sky130_fd_sc_hd__buf_4_0_ mux_left_track_37.mux_l2_in_0_/X VGND
+ VGND VPWR VPWR _086_/A sky130_fd_sc_hd__clkbuf_1
XPHY_4 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_15_151 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_30_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_30_132 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_21_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_21_176 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_12_132 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA_mux_left_track_7.mux_l1_in_1__A1 input49/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xmem_left_track_13.sky130_fd_sc_hd__dfxtp_1_1_ clkbuf_3_3_0_mem_left_track_1.prog_clk/X
+ mux_left_track_13.mux_l1_in_0_/S VGND VGND VPWR VPWR mux_left_track_13.mux_l2_in_0_/S
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_5_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_5_106 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xmem_left_track_1.sky130_fd_sc_hd__dfxtp_1_0_ clkbuf_3_5_0_mem_left_track_1.prog_clk/X
+ mux_top_track_26.mux_l2_in_0_/S VGND VGND VPWR VPWR mux_left_track_1.mux_l1_in_2_/S
+ sky130_fd_sc_hd__dfxtp_1
Xmux_left_track_3.mux_l2_in_0_ mux_left_track_3.mux_l1_in_1_/X mux_left_track_3.mux_l1_in_0_/X
+ mux_left_track_3.mux_l2_in_1_/S VGND VGND VPWR VPWR mux_left_track_3.mux_l2_in_0_/X
+ sky130_fd_sc_hd__mux2_1
Xclkbuf_3_2_0_mem_left_track_1.prog_clk clkbuf_3_3_0_mem_left_track_1.prog_clk/A VGND
+ VGND VPWR VPWR clkbuf_3_2_0_mem_left_track_1.prog_clk/X sky130_fd_sc_hd__clkbuf_1
XANTENNA_input12_A chanx_left_in[19] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_4_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_4_87 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_input4_A chanx_left_in[11] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_13_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xmux_left_track_3.mux_l1_in_1_ input42/X input49/X mux_left_track_3.mux_l1_in_1_/S
+ VGND VGND VPWR VPWR mux_left_track_3.mux_l1_in_1_/X sky130_fd_sc_hd__mux2_1
XFILLER_11_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_6_201 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_095_ _095_/A VGND VGND VPWR VPWR _095_/X sky130_fd_sc_hd__clkbuf_1
Xmem_left_track_7.sky130_fd_sc_hd__dfxtp_1_1_ clkbuf_3_1_0_mem_left_track_1.prog_clk/X
+ mux_left_track_7.mux_l1_in_1_/S VGND VGND VPWR VPWR mux_left_track_7.mux_l2_in_1_/S
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_1_33 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xmem_top_track_4.sky130_fd_sc_hd__dfxtp_1_0_ clkbuf_3_7_0_mem_left_track_1.prog_clk/X
+ mux_top_track_2.mux_l3_in_0_/S VGND VGND VPWR VPWR mux_top_track_4.mux_l1_in_2_/S
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_19_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__106__A _106_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_078_ _078_/A VGND VGND VPWR VPWR _078_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_33_152 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xmux_top_track_12.sky130_fd_sc_hd__buf_4_0_ mux_top_track_12.mux_l2_in_0_/X VGND VGND
+ VPWR VPWR _094_/A sky130_fd_sc_hd__clkbuf_1
XFILLER_33_196 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_16_119 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_103 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_114 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_125 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_136 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_147 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_24_130 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_24_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_24_152 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_158 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_169 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_21_30 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_input42_A left_bottom_grid_pin_11_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xclkbuf_3_5_0_mem_left_track_1.prog_clk clkbuf_3_5_0_mem_left_track_1.prog_clk/A VGND
+ VGND VPWR VPWR clkbuf_3_5_0_mem_left_track_1.prog_clk/X sky130_fd_sc_hd__clkbuf_1
Xmux_top_track_16.mux_l1_in_0_ input5/X input55/X mux_top_track_16.mux_l1_in_0_/S
+ VGND VGND VPWR VPWR mux_top_track_16.mux_l1_in_0_/X sky130_fd_sc_hd__mux2_1
Xmem_top_track_20.sky130_fd_sc_hd__dfxtp_1_0_ clkbuf_3_7_0_mem_left_track_1.prog_clk/X
+ mux_top_track_18.mux_l2_in_0_/S VGND VGND VPWR VPWR mux_top_track_20.mux_l1_in_0_/S
+ sky130_fd_sc_hd__dfxtp_1
XPHY_5 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_7_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_7_10 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_30_188 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_26_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_21_155 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_21_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_16_30 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_16_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_12_144 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_32_73 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_32_84 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmem_left_track_13.sky130_fd_sc_hd__dfxtp_1_0_ clkbuf_3_4_0_mem_left_track_1.prog_clk/X
+ mux_left_track_11.mux_l2_in_0_/S VGND VGND VPWR VPWR mux_left_track_13.mux_l1_in_0_/S
+ sky130_fd_sc_hd__dfxtp_1
Xmux_left_track_11.mux_l1_in_0_ input47/X input28/X mux_left_track_11.mux_l1_in_0_/S
+ VGND VGND VPWR VPWR mux_left_track_11.mux_l1_in_0_/X sky130_fd_sc_hd__mux2_1
XFILLER_26_203 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmux_left_track_23.mux_l2_in_0_ _063_/HI mux_left_track_23.mux_l1_in_0_/X mux_left_track_23.mux_l2_in_0_/S
+ VGND VGND VPWR VPWR mux_left_track_23.mux_l2_in_0_/X sky130_fd_sc_hd__mux2_1
XFILLER_4_99 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_4_66 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_4_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmem_top_track_26.sky130_fd_sc_hd__dfxtp_1_1_ clkbuf_3_5_0_mem_left_track_1.prog_clk/X
+ mux_top_track_26.mux_l1_in_0_/S VGND VGND VPWR VPWR mux_top_track_26.mux_l2_in_0_/S
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_13_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_9_210 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xmux_left_track_3.mux_l1_in_0_ input47/X input32/X mux_left_track_3.mux_l1_in_1_/S
+ VGND VGND VPWR VPWR mux_left_track_3.mux_l1_in_0_/X sky130_fd_sc_hd__mux2_1
XFILLER_1_9 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmem_left_track_19.sky130_fd_sc_hd__dfxtp_1_1_ clkbuf_3_3_0_mem_left_track_1.prog_clk/X
+ mux_left_track_19.mux_l1_in_0_/S VGND VGND VPWR VPWR mux_left_track_19.mux_l2_in_0_/S
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_24_30 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_24_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xmux_top_track_6.mux_l3_in_0_ mux_top_track_6.mux_l2_in_1_/X mux_top_track_6.mux_l2_in_0_/X
+ mux_top_track_6.mux_l3_in_0_/S VGND VGND VPWR VPWR mux_top_track_6.mux_l3_in_0_/X
+ sky130_fd_sc_hd__mux2_1
X_094_ _094_/A VGND VGND VPWR VPWR _094_/X sky130_fd_sc_hd__clkbuf_1
Xmem_left_track_7.sky130_fd_sc_hd__dfxtp_1_0_ clkbuf_3_1_0_mem_left_track_1.prog_clk/X
+ mux_left_track_5.mux_l3_in_0_/S VGND VGND VPWR VPWR mux_left_track_7.mux_l1_in_1_/S
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_1_45 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_10_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_10_87 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_27_172 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_077_ _077_/A VGND VGND VPWR VPWR _077_/X sky130_fd_sc_hd__clkbuf_1
XPHY_104 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_115 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_126 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_137 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xmux_top_track_6.mux_l2_in_1_ _054_/HI input10/X mux_top_track_6.mux_l2_in_1_/S VGND
+ VGND VPWR VPWR mux_top_track_6.mux_l2_in_1_/X sky130_fd_sc_hd__mux2_1
XPHY_148 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_24_175 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_159 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_input35_A chany_top_in[3] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_6 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_15_164 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_7_22 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_30_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_30_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_16_64 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_12_156 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_mux_left_track_29.mux_l1_in_0__A0 input48/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_32_30 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_32_96 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_4_78 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xmem_top_track_26.sky130_fd_sc_hd__dfxtp_1_0_ clkbuf_3_5_0_mem_left_track_1.prog_clk/X
+ mux_top_track_24.mux_l2_in_0_/S VGND VGND VPWR VPWR mux_top_track_26.mux_l1_in_0_/S
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_9_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xmux_left_track_23.mux_l1_in_0_ input44/X input41/X mux_left_track_23.mux_l1_in_0_/S
+ VGND VGND VPWR VPWR mux_left_track_23.mux_l1_in_0_/X sky130_fd_sc_hd__mux2_1
Xmem_left_track_19.sky130_fd_sc_hd__dfxtp_1_0_ clkbuf_3_3_0_mem_left_track_1.prog_clk/X
+ mux_left_track_17.mux_l2_in_0_/S VGND VGND VPWR VPWR mux_left_track_19.mux_l1_in_0_/S
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_10_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_24_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_6_214 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_093_ _093_/A VGND VGND VPWR VPWR _093_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_27_9 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmux_left_track_35.mux_l2_in_0_ _036_/HI mux_left_track_35.mux_l1_in_0_/X mux_left_track_35.mux_l2_in_0_/S
+ VGND VGND VPWR VPWR mux_left_track_35.mux_l2_in_0_/X sky130_fd_sc_hd__mux2_1
Xinput1 ccff_head VGND VGND VPWR VPWR input1/X sky130_fd_sc_hd__clkbuf_1
XFILLER_10_66 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_19_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_27_140 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_076_ _076_/A VGND VGND VPWR VPWR _076_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_18_5 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_18_162 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_18_173 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xmem_left_track_31.sky130_fd_sc_hd__dfxtp_1_1_ clkbuf_3_2_0_mem_left_track_1.prog_clk/X
+ mux_left_track_31.mux_l1_in_0_/S VGND VGND VPWR VPWR mux_left_track_31.mux_l2_in_0_/S
+ sky130_fd_sc_hd__dfxtp_1
XPHY_105 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_116 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_mux_left_track_37.mux_l1_in_0__A0 input43/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xmux_top_track_6.mux_l2_in_0_ mux_top_track_6.mux_l1_in_1_/X mux_top_track_6.mux_l1_in_0_/X
+ mux_top_track_6.mux_l2_in_1_/S VGND VGND VPWR VPWR mux_top_track_6.mux_l2_in_0_/X
+ sky130_fd_sc_hd__mux2_1
XPHY_127 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_138 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_149 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_24_198 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_input28_A chany_top_in[15] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_30_146 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_7_34 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_30_157 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_23_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_059_ VGND VGND VPWR VPWR _059_/HI _059_/LO sky130_fd_sc_hd__conb_1
XFILLER_21_179 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_16_87 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_16_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_12_168 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_32_64 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmux_top_track_6.sky130_fd_sc_hd__buf_4_0_ mux_top_track_6.mux_l3_in_0_/X VGND VGND
+ VPWR VPWR _091_/A sky130_fd_sc_hd__clkbuf_1
XFILLER_7_172 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xmux_top_track_6.mux_l1_in_1_ input58/X input56/X mux_top_track_6.mux_l1_in_1_/S VGND
+ VGND VPWR VPWR mux_top_track_6.mux_l1_in_1_/X sky130_fd_sc_hd__mux2_1
XFILLER_17_216 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_27_86 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_13_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_13_33 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_input10_A chanx_left_in[17] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_input2_A chanx_left_in[0] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_24_76 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_24_87 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_24_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_input58_A top_left_grid_pin_49_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_092_ _092_/A VGND VGND VPWR VPWR _092_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_1_25 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_1_58 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xinput2 chanx_left_in[0] VGND VGND VPWR VPWR input2/X sky130_fd_sc_hd__buf_1
XFILLER_28_108 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_19_10 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_19_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_19_108 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_075_ _075_/A VGND VGND VPWR VPWR _075_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_33_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_33_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_33_144 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_33_122 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmem_left_track_31.sky130_fd_sc_hd__dfxtp_1_0_ clkbuf_3_2_0_mem_left_track_1.prog_clk/X
+ mux_left_track_29.mux_l2_in_0_/S VGND VGND VPWR VPWR mux_left_track_31.mux_l1_in_0_/S
+ sky130_fd_sc_hd__dfxtp_1
XPHY_106 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_117 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_mux_top_track_10.mux_l1_in_0__A1 input52/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_128 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_139 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_24_122 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmux_left_track_35.mux_l1_in_0_ input42/X input35/X mux_left_track_35.mux_l1_in_0_/S
+ VGND VGND VPWR VPWR mux_left_track_35.mux_l1_in_0_/X sky130_fd_sc_hd__mux2_1
XFILLER_21_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_8 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_15_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_30_114 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_30_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_30_136 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_7_46 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_058_ VGND VGND VPWR VPWR _058_/HI _058_/LO sky130_fd_sc_hd__conb_1
XANTENNA_mux_top_track_2.mux_l1_in_0__A0 input54/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_16_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_32_87 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_input40_A chany_top_in[8] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_7_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_7_151 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xmux_top_track_6.mux_l1_in_0_ input54/X input52/X mux_top_track_6.mux_l1_in_1_/S VGND
+ VGND VPWR VPWR mux_top_track_6.mux_l1_in_0_/X sky130_fd_sc_hd__mux2_1
Xmem_left_track_37.sky130_fd_sc_hd__dfxtp_1_1_ clkbuf_3_2_0_mem_left_track_1.prog_clk/X
+ mux_left_track_37.mux_l1_in_0_/S VGND VGND VPWR VPWR mux_left_track_37.mux_l2_in_0_/S
+ sky130_fd_sc_hd__dfxtp_1
XANTENNA_mux_top_track_0.mux_l1_in_2__A0 input2/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_32_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_13_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xmux_left_track_1.sky130_fd_sc_hd__buf_4_0_ mux_left_track_1.mux_l3_in_0_/X VGND VGND
+ VPWR VPWR _068_/A sky130_fd_sc_hd__clkbuf_1
XFILLER_10_201 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_091_ _091_/A VGND VGND VPWR VPWR _091_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_1_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xinput3 chanx_left_in[10] VGND VGND VPWR VPWR input3/X sky130_fd_sc_hd__buf_1
XFILLER_10_13 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_3_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_19_88 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_074_ _074_/A VGND VGND VPWR VPWR _074_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_32_9 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_33_134 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_18_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xmem_top_track_12.sky130_fd_sc_hd__dfxtp_1_1_ clkbuf_3_4_0_mem_left_track_1.prog_clk/X
+ mux_top_track_12.mux_l1_in_0_/S VGND VGND VPWR VPWR mux_top_track_12.mux_l2_in_0_/S
+ sky130_fd_sc_hd__dfxtp_1
XPHY_107 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_118 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_129 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_24_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xclkbuf_2_2_0_mem_left_track_1.prog_clk clkbuf_2_3_0_mem_left_track_1.prog_clk/A VGND
+ VGND VPWR VPWR clkbuf_3_5_0_mem_left_track_1.prog_clk/A sky130_fd_sc_hd__clkbuf_1
XPHY_9 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_15_112 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_7_58 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_057_ VGND VGND VPWR VPWR _057_/HI _057_/LO sky130_fd_sc_hd__conb_1
XFILLER_21_115 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xinput50 left_bottom_grid_pin_9_ VGND VGND VPWR VPWR input50/X sky130_fd_sc_hd__clkbuf_2
XFILLER_21_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_mux_top_track_2.mux_l1_in_0__A1 input52/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_16_23 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_prog_clk_0_FTB00_A prog_clk_0_N_in VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_20_170 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_input33_A chany_top_in[1] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_7_163 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_7_196 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_26_207 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xmux_left_track_11.sky130_fd_sc_hd__buf_4_0_ mux_left_track_11.mux_l2_in_0_/X VGND
+ VGND VPWR VPWR _073_/A sky130_fd_sc_hd__clkbuf_1
Xmem_left_track_37.sky130_fd_sc_hd__dfxtp_1_0_ clkbuf_3_2_0_mem_left_track_1.prog_clk/X
+ mux_left_track_35.mux_l2_in_0_/S VGND VGND VPWR VPWR mux_left_track_37.mux_l1_in_0_/S
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_27_33 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_27_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_27_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_4_144 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_4_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_4_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_31_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_22_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_8_6 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_10_213 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_090_ _090_/A VGND VGND VPWR VPWR _090_/X sky130_fd_sc_hd__clkbuf_1
Xinput4 chanx_left_in[11] VGND VGND VPWR VPWR input4/X sky130_fd_sc_hd__buf_1
XFILLER_27_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_27_198 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_073_ _073_/A VGND VGND VPWR VPWR _073_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_25_9 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_33_146 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmem_top_track_12.sky130_fd_sc_hd__dfxtp_1_0_ clkbuf_3_4_0_mem_left_track_1.prog_clk/X
+ mux_top_track_10.mux_l2_in_0_/S VGND VGND VPWR VPWR mux_top_track_12.mux_l1_in_0_/S
+ sky130_fd_sc_hd__dfxtp_1
XPHY_108 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_119 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_24_146 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_24_157 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_24_179 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_21_35 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_30_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_056_ VGND VGND VPWR VPWR _056_/HI _056_/LO sky130_fd_sc_hd__conb_1
Xinput40 chany_top_in[8] VGND VGND VPWR VPWR input40/X sky130_fd_sc_hd__clkbuf_1
Xinput51 top_left_grid_pin_42_ VGND VGND VPWR VPWR input51/X sky130_fd_sc_hd__clkbuf_2
XFILLER_29_205 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_16_46 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_input26_A chany_top_in[13] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_039_ VGND VGND VPWR VPWR _039_/HI _039_/LO sky130_fd_sc_hd__conb_1
XFILLER_21_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_26_219 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xmem_top_track_18.sky130_fd_sc_hd__dfxtp_1_1_ clkbuf_3_7_0_mem_left_track_1.prog_clk/X
+ mux_top_track_18.mux_l1_in_0_/S VGND VGND VPWR VPWR mux_top_track_18.mux_l2_in_0_/S
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_17_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_4_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_4_156 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_4_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmux_top_track_12.mux_l2_in_0_ _044_/HI mux_top_track_12.mux_l1_in_0_/X mux_top_track_12.mux_l2_in_0_/S
+ VGND VGND VPWR VPWR mux_top_track_12.mux_l2_in_0_/X sky130_fd_sc_hd__mux2_1
XFILLER_13_58 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_13_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_1_115 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xmux_left_track_33.sky130_fd_sc_hd__buf_4_0_ mux_left_track_33.mux_l2_in_0_/X VGND
+ VGND VPWR VPWR _084_/A sky130_fd_sc_hd__clkbuf_1
XFILLER_0_170 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_5_70 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_24_24 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_24_35 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_6_218 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xinput5 chanx_left_in[12] VGND VGND VPWR VPWR input5/X sky130_fd_sc_hd__buf_1
Xmux_left_track_27.sky130_fd_sc_hd__buf_4_0_ mux_left_track_27.mux_l2_in_0_/X VGND
+ VGND VPWR VPWR _081_/A sky130_fd_sc_hd__clkbuf_1
XFILLER_10_48 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_27_144 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_27_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_2_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_072_ _072_/A VGND VGND VPWR VPWR _072_/X sky130_fd_sc_hd__clkbuf_1
XANTENNA_input56_A top_left_grid_pin_47_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_33_114 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_18_144 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_24_103 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_109 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_21_14 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_21_25 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_21_58 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_21_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_15_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_055_ VGND VGND VPWR VPWR _055_/HI _055_/LO sky130_fd_sc_hd__conb_1
XFILLER_23_180 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_16_6 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xinput41 chany_top_in[9] VGND VGND VPWR VPWR input41/X sky130_fd_sc_hd__clkbuf_1
Xinput30 chany_top_in[17] VGND VGND VPWR VPWR input30/X sky130_fd_sc_hd__buf_1
Xinput52 top_left_grid_pin_43_ VGND VGND VPWR VPWR input52/X sky130_fd_sc_hd__clkbuf_2
XFILLER_29_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_32_35 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_32_46 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_input19_A chanx_left_in[7] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_107_ _107_/A VGND VGND VPWR VPWR _107_/X sky130_fd_sc_hd__buf_1
XFILLER_11_172 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_038_ VGND VGND VPWR VPWR _038_/HI _038_/LO sky130_fd_sc_hd__conb_1
XFILLER_8_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xmem_top_track_18.sky130_fd_sc_hd__dfxtp_1_0_ clkbuf_3_7_0_mem_left_track_1.prog_clk/X
+ mux_top_track_16.mux_l2_in_0_/S VGND VGND VPWR VPWR mux_top_track_18.mux_l1_in_0_/S
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_4_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_4_168 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_31_201 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_22_201 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_13_37 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_1_127 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_5_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_24_14 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_24_58 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_1_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmux_top_track_12.mux_l1_in_0_ input7/X input53/X mux_top_track_12.mux_l1_in_0_/S
+ VGND VGND VPWR VPWR mux_top_track_12.mux_l1_in_0_/X sky130_fd_sc_hd__mux2_1
Xinput6 chanx_left_in[13] VGND VGND VPWR VPWR input6/X sky130_fd_sc_hd__buf_1
Xmux_top_track_24.mux_l2_in_0_ mux_top_track_24.mux_l1_in_1_/X mux_top_track_24.mux_l1_in_0_/X
+ mux_top_track_24.mux_l2_in_0_/S VGND VGND VPWR VPWR mux_top_track_24.mux_l2_in_0_/X
+ sky130_fd_sc_hd__mux2_1
XFILLER_10_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_mux_left_track_3.mux_l1_in_1__A0 input42/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_19_36 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_19_58 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xmem_left_track_23.sky130_fd_sc_hd__dfxtp_1_1_ clkbuf_3_2_0_mem_left_track_1.prog_clk/X
+ mux_left_track_23.mux_l1_in_0_/S VGND VGND VPWR VPWR mux_left_track_23.mux_l2_in_0_/S
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_27_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_071_ _071_/A VGND VGND VPWR VPWR _071_/X sky130_fd_sc_hd__clkbuf_1
XANTENNA_input49_A left_bottom_grid_pin_7_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_18_112 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_18_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_18_134 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_33_104 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_90 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_24_126 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmux_left_track_17.mux_l2_in_0_ _060_/HI mux_left_track_17.mux_l1_in_0_/X mux_left_track_17.mux_l2_in_0_/S
+ VGND VGND VPWR VPWR mux_left_track_17.mux_l2_in_0_/X sky130_fd_sc_hd__mux2_1
XFILLER_15_115 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_054_ VGND VGND VPWR VPWR _054_/HI _054_/LO sky130_fd_sc_hd__conb_1
Xmux_top_track_24.mux_l1_in_1_ _051_/HI input20/X mux_top_track_24.mux_l1_in_1_/S
+ VGND VGND VPWR VPWR mux_top_track_24.mux_l1_in_1_/X sky130_fd_sc_hd__mux2_1
XFILLER_30_9 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_mux_top_track_16.mux_l1_in_0__A0 input5/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xinput20 chanx_left_in[8] VGND VGND VPWR VPWR input20/X sky130_fd_sc_hd__buf_1
Xinput31 chany_top_in[18] VGND VGND VPWR VPWR input31/X sky130_fd_sc_hd__buf_1
Xinput42 left_bottom_grid_pin_11_ VGND VGND VPWR VPWR input42/X sky130_fd_sc_hd__clkbuf_2
Xinput53 top_left_grid_pin_44_ VGND VGND VPWR VPWR input53/X sky130_fd_sc_hd__clkbuf_2
XFILLER_20_140 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_20_162 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_32_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_11_151 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_106_ _106_/A VGND VGND VPWR VPWR _106_/X sky130_fd_sc_hd__buf_1
XFILLER_11_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_037_ VGND VGND VPWR VPWR _037_/HI _037_/LO sky130_fd_sc_hd__conb_1
Xmux_left_track_9.mux_l2_in_0_ mux_left_track_9.mux_l1_in_1_/X mux_left_track_9.mux_l1_in_0_/X
+ mux_left_track_9.mux_l2_in_0_/S VGND VGND VPWR VPWR mux_left_track_9.mux_l2_in_0_/X
+ sky130_fd_sc_hd__mux2_1
Xmux_top_track_2.mux_l3_in_0_ mux_top_track_2.mux_l2_in_1_/X mux_top_track_2.mux_l2_in_0_/X
+ mux_top_track_2.mux_l3_in_0_/S VGND VGND VPWR VPWR mux_top_track_2.mux_l3_in_0_/X
+ sky130_fd_sc_hd__mux2_1
XANTENNA_input31_A chany_top_in[18] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_16_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_17_91 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_22_213 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_1_106 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_1_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xmux_left_track_9.mux_l1_in_1_ _041_/HI input45/X mux_left_track_9.mux_l1_in_1_/S
+ VGND VGND VPWR VPWR mux_left_track_9.mux_l1_in_1_/X sky130_fd_sc_hd__mux2_1
XFILLER_5_94 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_5_50 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_6_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_6_6 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmux_top_track_2.mux_l2_in_1_ _048_/HI input12/X mux_top_track_2.mux_l2_in_1_/S VGND
+ VGND VPWR VPWR mux_top_track_2.mux_l2_in_1_/X sky130_fd_sc_hd__mux2_1
XFILLER_14_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xinput7 chanx_left_in[14] VGND VGND VPWR VPWR input7/X sky130_fd_sc_hd__buf_1
XFILLER_10_17 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_mux_left_track_3.mux_l1_in_1__A1 input49/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_19_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xmem_left_track_23.sky130_fd_sc_hd__dfxtp_1_0_ clkbuf_3_2_0_mem_left_track_1.prog_clk/X
+ mux_left_track_21.mux_l2_in_0_/S VGND VGND VPWR VPWR mux_left_track_23.mux_l1_in_0_/S
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_27_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_070_ _070_/A VGND VGND VPWR VPWR _070_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_2_201 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xmux_top_track_24.sky130_fd_sc_hd__buf_4_0_ mux_top_track_24.mux_l2_in_0_/X VGND VGND
+ VPWR VPWR _100_/A sky130_fd_sc_hd__clkbuf_1
XPHY_91 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_80 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_25_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_32_171 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_32_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_053_ VGND VGND VPWR VPWR _053_/HI _053_/LO sky130_fd_sc_hd__conb_1
Xmux_top_track_24.mux_l1_in_0_ input59/X input51/X mux_top_track_24.mux_l1_in_1_/S
+ VGND VGND VPWR VPWR mux_top_track_24.mux_l1_in_0_/X sky130_fd_sc_hd__mux2_1
XFILLER_23_9 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xinput54 top_left_grid_pin_45_ VGND VGND VPWR VPWR input54/X sky130_fd_sc_hd__clkbuf_2
Xinput43 left_bottom_grid_pin_13_ VGND VGND VPWR VPWR input43/X sky130_fd_sc_hd__clkbuf_2
Xinput21 chanx_left_in[9] VGND VGND VPWR VPWR input21/X sky130_fd_sc_hd__buf_1
Xinput10 chanx_left_in[17] VGND VGND VPWR VPWR input10/X sky130_fd_sc_hd__clkbuf_1
Xinput32 chany_top_in[19] VGND VGND VPWR VPWR input32/X sky130_fd_sc_hd__buf_1
XFILLER_12_108 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_16_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_20_130 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xmux_top_track_18.sky130_fd_sc_hd__buf_4_0_ mux_top_track_18.mux_l2_in_0_/X VGND VGND
+ VPWR VPWR _097_/A sky130_fd_sc_hd__clkbuf_1
XFILLER_20_174 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_105_ _105_/A VGND VGND VPWR VPWR _105_/X sky130_fd_sc_hd__buf_1
XFILLER_11_163 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_11_196 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xmem_left_track_29.sky130_fd_sc_hd__dfxtp_1_1_ clkbuf_3_2_0_mem_left_track_1.prog_clk/X
+ mux_left_track_29.mux_l1_in_0_/S VGND VGND VPWR VPWR mux_left_track_29.mux_l2_in_0_/S
+ sky130_fd_sc_hd__dfxtp_1
Xmux_left_track_17.mux_l1_in_0_ input50/X input25/X mux_left_track_17.mux_l1_in_0_/S
+ VGND VGND VPWR VPWR mux_left_track_17.mux_l1_in_0_/X sky130_fd_sc_hd__mux2_1
X_036_ VGND VGND VPWR VPWR _036_/HI _036_/LO sky130_fd_sc_hd__conb_1
Xmux_left_track_29.mux_l2_in_0_ _066_/HI mux_left_track_29.mux_l1_in_0_/X mux_left_track_29.mux_l2_in_0_/S
+ VGND VGND VPWR VPWR mux_left_track_29.mux_l2_in_0_/X sky130_fd_sc_hd__mux2_1
XFILLER_25_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_27_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_input24_A chany_top_in[11] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xmux_left_track_31.mux_l2_in_0_ _034_/HI mux_left_track_31.mux_l1_in_0_/X mux_left_track_31.mux_l2_in_0_/S
+ VGND VGND VPWR VPWR mux_left_track_31.mux_l2_in_0_/X sky130_fd_sc_hd__mux2_1
Xmux_left_track_9.mux_l1_in_0_ input46/X input29/X mux_left_track_9.mux_l1_in_1_/S
+ VGND VGND VPWR VPWR mux_left_track_9.mux_l1_in_0_/X sky130_fd_sc_hd__mux2_1
Xmux_top_track_2.mux_l2_in_0_ mux_top_track_2.mux_l1_in_1_/X mux_top_track_2.mux_l1_in_0_/X
+ mux_top_track_2.mux_l2_in_1_/S VGND VGND VPWR VPWR mux_top_track_2.mux_l2_in_0_/X
+ sky130_fd_sc_hd__mux2_1
Xmux_top_track_2.sky130_fd_sc_hd__buf_4_0_ mux_top_track_2.mux_l3_in_0_/X VGND VGND
+ VPWR VPWR _089_/A sky130_fd_sc_hd__clkbuf_1
XFILLER_5_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xinput8 chanx_left_in[15] VGND VGND VPWR VPWR input8/X sky130_fd_sc_hd__clkbuf_1
XFILLER_27_136 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_27_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_2_213 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xmem_top_track_0.sky130_fd_sc_hd__dfxtp_1_2_ clkbuf_3_6_0_mem_left_track_1.prog_clk/X
+ mux_top_track_0.mux_l2_in_1_/S VGND VGND VPWR VPWR mux_top_track_0.mux_l3_in_0_/S
+ sky130_fd_sc_hd__dfxtp_1
XANTENNA_mux_top_track_24.mux_l1_in_0__A1 input51/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_33_128 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_33_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_18_103 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_92 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_81 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_70 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_30 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xmux_top_track_2.mux_l1_in_1_ input58/X input56/X mux_top_track_2.mux_l1_in_1_/S VGND
+ VGND VPWR VPWR mux_top_track_2.mux_l1_in_1_/X sky130_fd_sc_hd__mux2_1
XFILLER_32_150 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_32_183 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_mux_left_track_17.mux_l1_in_0__A0 input50/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_052_ VGND VGND VPWR VPWR _052_/HI _052_/LO sky130_fd_sc_hd__conb_1
XANTENNA_input54_A top_left_grid_pin_45_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xinput22 chany_top_in[0] VGND VGND VPWR VPWR input22/X sky130_fd_sc_hd__clkbuf_1
Xinput44 left_bottom_grid_pin_15_ VGND VGND VPWR VPWR input44/X sky130_fd_sc_hd__clkbuf_2
Xinput11 chanx_left_in[18] VGND VGND VPWR VPWR input11/X sky130_fd_sc_hd__buf_1
Xinput55 top_left_grid_pin_46_ VGND VGND VPWR VPWR input55/X sky130_fd_sc_hd__buf_1
Xinput33 chany_top_in[1] VGND VGND VPWR VPWR input33/X sky130_fd_sc_hd__clkbuf_1
XFILLER_32_16 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_32_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmem_left_track_29.sky130_fd_sc_hd__dfxtp_1_0_ clkbuf_3_0_0_mem_left_track_1.prog_clk/X
+ mux_left_track_27.mux_l2_in_0_/S VGND VGND VPWR VPWR mux_left_track_29.mux_l1_in_0_/S
+ sky130_fd_sc_hd__dfxtp_1
X_104_ _104_/A VGND VGND VPWR VPWR _104_/X sky130_fd_sc_hd__buf_1
X_035_ VGND VGND VPWR VPWR _035_/HI _035_/LO sky130_fd_sc_hd__conb_1
XANTENNA_mux_top_track_8.mux_l1_in_0__A1 input51/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_14_6 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_input17_A chanx_left_in[5] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_16_201 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_13_18 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_13_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_input9_A chanx_left_in[16] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xmux_left_track_29.mux_l1_in_0_ input48/X input38/X mux_left_track_29.mux_l1_in_0_/S
+ VGND VGND VPWR VPWR mux_left_track_29.mux_l1_in_0_/X sky130_fd_sc_hd__mux2_1
XFILLER_24_28 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xmux_left_track_31.mux_l1_in_0_ input49/X input37/X mux_left_track_31.mux_l1_in_0_/S
+ VGND VGND VPWR VPWR mux_left_track_31.mux_l1_in_0_/X sky130_fd_sc_hd__mux2_1
XFILLER_14_61 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xinput9 chanx_left_in[16] VGND VGND VPWR VPWR input9/X sky130_fd_sc_hd__clkbuf_1
Xmem_left_track_3.sky130_fd_sc_hd__dfxtp_1_2_ clkbuf_3_0_0_mem_left_track_1.prog_clk/X
+ mux_left_track_3.mux_l2_in_1_/S VGND VGND VPWR VPWR mux_left_track_3.mux_l3_in_0_/S
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_27_104 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_27_148 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xmem_top_track_0.sky130_fd_sc_hd__dfxtp_1_1_ clkbuf_3_4_0_mem_left_track_1.prog_clk/X
+ mux_top_track_0.mux_l1_in_2_/S VGND VGND VPWR VPWR mux_top_track_0.mux_l2_in_1_/S
+ sky130_fd_sc_hd__dfxtp_1
XPHY_82 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_71 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_60 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_93 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_42 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xmux_top_track_2.mux_l1_in_0_ input54/X input52/X mux_top_track_2.mux_l1_in_1_/S VGND
+ VGND VPWR VPWR mux_top_track_2.mux_l1_in_0_/X sky130_fd_sc_hd__mux2_1
XFILLER_17_170 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_15_107 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_051_ VGND VGND VPWR VPWR _051_/HI _051_/LO sky130_fd_sc_hd__conb_1
XANTENNA_input47_A left_bottom_grid_pin_3_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xinput45 left_bottom_grid_pin_17_ VGND VGND VPWR VPWR input45/X sky130_fd_sc_hd__clkbuf_2
Xinput12 chanx_left_in[19] VGND VGND VPWR VPWR input12/X sky130_fd_sc_hd__buf_1
Xinput34 chany_top_in[2] VGND VGND VPWR VPWR input34/X sky130_fd_sc_hd__clkbuf_1
Xinput56 top_left_grid_pin_47_ VGND VGND VPWR VPWR input56/X sky130_fd_sc_hd__clkbuf_2
Xinput23 chany_top_in[10] VGND VGND VPWR VPWR input23/X sky130_fd_sc_hd__clkbuf_1
XFILLER_20_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_28_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_103_ _103_/A VGND VGND VPWR VPWR _103_/X sky130_fd_sc_hd__buf_1
XFILLER_22_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_034_ VGND VGND VPWR VPWR _034_/HI _034_/LO sky130_fd_sc_hd__conb_1
Xmem_top_track_6.sky130_fd_sc_hd__dfxtp_1_2_ clkbuf_3_6_0_mem_left_track_1.prog_clk/X
+ mux_top_track_6.mux_l2_in_1_/S VGND VGND VPWR VPWR mux_top_track_6.mux_l3_in_0_/S
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_8_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_8_30 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_6_180 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_25_202 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_16_213 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_17_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_33_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_33_71 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_31_205 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_3_172 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_mux_left_track_5.mux_l1_in_2__A1 input43/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_175 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_mux_left_track_33.mux_l1_in_0__A0 input50/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_28_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_30_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xmem_left_track_3.sky130_fd_sc_hd__dfxtp_1_1_ clkbuf_3_0_0_mem_left_track_1.prog_clk/X
+ mux_left_track_3.mux_l1_in_1_/S VGND VGND VPWR VPWR mux_left_track_3.mux_l2_in_1_/S
+ sky130_fd_sc_hd__dfxtp_1
Xmem_top_track_0.sky130_fd_sc_hd__dfxtp_1_0_ clkbuf_3_5_0_mem_left_track_1.prog_clk/X
+ input1/X VGND VGND VPWR VPWR mux_top_track_0.mux_l1_in_2_/S sky130_fd_sc_hd__dfxtp_1
XFILLER_4_6 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_33_108 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_94 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_83 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_72 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_50 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_26_160 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_61 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_output60_A output60/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_2_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_2_87 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_21_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xoutput100 _097_/X VGND VGND VPWR VPWR chany_top_out[9] sky130_fd_sc_hd__clkbuf_2
XFILLER_23_174 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_050_ VGND VGND VPWR VPWR _050_/HI _050_/LO sky130_fd_sc_hd__conb_1
XFILLER_2_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xinput13 chanx_left_in[1] VGND VGND VPWR VPWR _107_/A sky130_fd_sc_hd__buf_1
XFILLER_14_152 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xclkbuf_3_1_0_mem_left_track_1.prog_clk clkbuf_3_1_0_mem_left_track_1.prog_clk/A VGND
+ VGND VPWR VPWR clkbuf_3_1_0_mem_left_track_1.prog_clk/X sky130_fd_sc_hd__clkbuf_1
Xinput24 chany_top_in[11] VGND VGND VPWR VPWR input24/X sky130_fd_sc_hd__clkbuf_1
Xinput46 left_bottom_grid_pin_1_ VGND VGND VPWR VPWR input46/X sky130_fd_sc_hd__clkbuf_2
Xinput57 top_left_grid_pin_48_ VGND VGND VPWR VPWR input57/X sky130_fd_sc_hd__buf_1
Xinput35 chany_top_in[3] VGND VGND VPWR VPWR input35/X sky130_fd_sc_hd__clkbuf_1
XFILLER_20_144 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_20_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_20_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_20_188 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_11_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_102_ _102_/A VGND VGND VPWR VPWR _102_/X sky130_fd_sc_hd__buf_1
XFILLER_7_115 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_22_73 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_19_211 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_21_9 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmem_top_track_6.sky130_fd_sc_hd__dfxtp_1_1_ clkbuf_3_3_0_mem_left_track_1.prog_clk/X
+ mux_top_track_6.mux_l1_in_1_/S VGND VGND VPWR VPWR mux_top_track_6.mux_l2_in_1_/S
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_8_64 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_6_192 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_17_73 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__104__A _104_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_3_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_3_151 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_12_5 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmem_top_track_22.sky130_fd_sc_hd__dfxtp_1_1_ clkbuf_3_7_0_mem_left_track_1.prog_clk/X
+ mux_top_track_22.mux_l1_in_0_/S VGND VGND VPWR VPWR mux_top_track_22.mux_l2_in_0_/S
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_187 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_28_61 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_input22_A chany_top_in[0] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_8_210 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_5_10 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_output90_A _106_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_24_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_14_30 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_14_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_14_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xmem_left_track_15.sky130_fd_sc_hd__dfxtp_1_1_ clkbuf_3_3_0_mem_left_track_1.prog_clk/X
+ mux_left_track_15.mux_l1_in_0_/S VGND VGND VPWR VPWR mux_left_track_15.mux_l2_in_0_/S
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_30_40 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmem_left_track_3.sky130_fd_sc_hd__dfxtp_1_0_ clkbuf_3_0_0_mem_left_track_1.prog_clk/X
+ mux_left_track_1.mux_l3_in_0_/S VGND VGND VPWR VPWR mux_left_track_3.mux_l1_in_1_/S
+ sky130_fd_sc_hd__dfxtp_1
Xclkbuf_3_4_0_mem_left_track_1.prog_clk clkbuf_3_5_0_mem_left_track_1.prog_clk/A VGND
+ VGND VPWR VPWR clkbuf_3_4_0_mem_left_track_1.prog_clk/X sky130_fd_sc_hd__clkbuf_1
XFILLER_19_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_27_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xmux_left_track_7.sky130_fd_sc_hd__buf_4_0_ mux_left_track_7.mux_l3_in_0_/X VGND VGND
+ VPWR VPWR _071_/A sky130_fd_sc_hd__clkbuf_1
XFILLER_18_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_95 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_84 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_73 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_40 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_26_150 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_2_66 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_2_99 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_17_150 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_17_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_32_120 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_32_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xinput25 chany_top_in[12] VGND VGND VPWR VPWR input25/X sky130_fd_sc_hd__clkbuf_1
XANTENNA__107__A _107_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xinput14 chanx_left_in[2] VGND VGND VPWR VPWR _106_/A sky130_fd_sc_hd__buf_1
XFILLER_14_142 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_14_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xinput36 chany_top_in[4] VGND VGND VPWR VPWR input36/X sky130_fd_sc_hd__clkbuf_1
Xinput58 top_left_grid_pin_49_ VGND VGND VPWR VPWR input58/X sky130_fd_sc_hd__clkbuf_2
Xinput47 left_bottom_grid_pin_3_ VGND VGND VPWR VPWR input47/X sky130_fd_sc_hd__clkbuf_2
XFILLER_28_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmem_left_track_9.sky130_fd_sc_hd__dfxtp_1_1_ clkbuf_3_1_0_mem_left_track_1.prog_clk/X
+ mux_left_track_9.mux_l1_in_1_/S VGND VGND VPWR VPWR mux_left_track_9.mux_l2_in_0_/S
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_28_201 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_7_127 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_22_30 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_101_ _101_/A VGND VGND VPWR VPWR _101_/X sky130_fd_sc_hd__clkbuf_1
XANTENNA_input52_A top_left_grid_pin_43_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xmem_top_track_6.sky130_fd_sc_hd__dfxtp_1_0_ clkbuf_3_6_0_mem_left_track_1.prog_clk/X
+ mux_top_track_4.mux_l3_in_0_/S VGND VGND VPWR VPWR mux_top_track_6.mux_l1_in_1_/S
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_8_87 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_8_76 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_8_10 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xmux_left_track_23.sky130_fd_sc_hd__buf_4_0_ mux_left_track_23.mux_l2_in_0_/X VGND
+ VGND VPWR VPWR _079_/A sky130_fd_sc_hd__clkbuf_1
XFILLER_3_196 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_3_163 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xmem_top_track_22.sky130_fd_sc_hd__dfxtp_1_0_ clkbuf_3_7_0_mem_left_track_1.prog_clk/X
+ mux_top_track_20.mux_l2_in_0_/S VGND VGND VPWR VPWR mux_top_track_22.mux_l1_in_0_/S
+ sky130_fd_sc_hd__dfxtp_1
Xclkbuf_3_7_0_mem_left_track_1.prog_clk clkbuf_3_7_0_mem_left_track_1.prog_clk/A VGND
+ VGND VPWR VPWR clkbuf_3_7_0_mem_left_track_1.prog_clk/X sky130_fd_sc_hd__clkbuf_1
XFILLER_0_100 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xmux_left_track_17.sky130_fd_sc_hd__buf_4_0_ mux_left_track_17.mux_l2_in_0_/X VGND
+ VGND VPWR VPWR _076_/A sky130_fd_sc_hd__clkbuf_1
XANTENNA_input15_A chanx_left_in[3] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_199 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_8_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xmux_left_track_5.mux_l3_in_0_ mux_left_track_5.mux_l2_in_1_/X mux_left_track_5.mux_l2_in_0_/X
+ mux_left_track_5.mux_l3_in_0_/S VGND VGND VPWR VPWR mux_left_track_5.mux_l3_in_0_/X
+ sky130_fd_sc_hd__mux2_1
XANTENNA_input7_A chanx_left_in[14] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xmem_left_track_15.sky130_fd_sc_hd__dfxtp_1_0_ clkbuf_3_3_0_mem_left_track_1.prog_clk/X
+ mux_left_track_13.mux_l2_in_0_/S VGND VGND VPWR VPWR mux_left_track_15.mux_l1_in_0_/S
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_30_30 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_30_63 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_30 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_96 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_85 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_74 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_25_63 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_52 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_63 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_2_23 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_2_78 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_32_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_32_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmux_left_track_5.mux_l2_in_1_ _039_/HI mux_left_track_5.mux_l1_in_2_/X mux_left_track_5.mux_l2_in_1_/S
+ VGND VGND VPWR VPWR mux_left_track_5.mux_l2_in_1_/X sky130_fd_sc_hd__mux2_1
XFILLER_11_10 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_11_76 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_11_87 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xinput59 top_right_grid_pin_1_ VGND VGND VPWR VPWR input59/X sky130_fd_sc_hd__clkbuf_2
Xinput15 chanx_left_in[3] VGND VGND VPWR VPWR _105_/A sky130_fd_sc_hd__buf_1
Xinput48 left_bottom_grid_pin_5_ VGND VGND VPWR VPWR input48/X sky130_fd_sc_hd__clkbuf_2
Xinput37 chany_top_in[5] VGND VGND VPWR VPWR input37/X sky130_fd_sc_hd__clkbuf_1
Xinput26 chany_top_in[13] VGND VGND VPWR VPWR input26/X sky130_fd_sc_hd__clkbuf_1
XFILLER_20_102 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xmem_left_track_9.sky130_fd_sc_hd__dfxtp_1_0_ clkbuf_3_1_0_mem_left_track_1.prog_clk/X
+ mux_left_track_7.mux_l3_in_0_/S VGND VGND VPWR VPWR mux_left_track_9.mux_l1_in_1_/S
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_28_213 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_7_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_7_106 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_100_ _100_/A VGND VGND VPWR VPWR _100_/X sky130_fd_sc_hd__clkbuf_1
XANTENNA_input45_A left_bottom_grid_pin_17_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xmux_left_track_5.mux_l1_in_2_ input45/X input43/X mux_left_track_5.mux_l1_in_2_/S
+ VGND VGND VPWR VPWR mux_left_track_5.mux_l1_in_2_/X sky130_fd_sc_hd__mux2_1
XFILLER_8_33 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_8_22 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_8_99 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_8_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_17_20 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_33_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_33_30 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmux_top_track_18.mux_l2_in_0_ _047_/HI mux_top_track_18.mux_l1_in_0_/X mux_top_track_18.mux_l2_in_0_/S
+ VGND VGND VPWR VPWR mux_top_track_18.mux_l2_in_0_/X sky130_fd_sc_hd__mux2_1
Xmux_top_track_20.mux_l2_in_0_ _049_/HI mux_top_track_20.mux_l1_in_0_/X mux_top_track_20.mux_l2_in_0_/S
+ VGND VGND VPWR VPWR mux_top_track_20.mux_l2_in_0_/X sky130_fd_sc_hd__mux2_1
XFILLER_13_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_0_112 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_28_30 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_8_201 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_5_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xmux_left_track_13.mux_l2_in_0_ _058_/HI mux_left_track_13.mux_l1_in_0_/X mux_left_track_13.mux_l2_in_0_/S
+ VGND VGND VPWR VPWR mux_left_track_13.mux_l2_in_0_/X sky130_fd_sc_hd__mux2_1
XFILLER_14_87 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_30_20 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmux_left_track_39.sky130_fd_sc_hd__buf_4_0_ mux_left_track_39.mux_l2_in_0_/X VGND
+ VGND VPWR VPWR _087_/A sky130_fd_sc_hd__clkbuf_1
XFILLER_29_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_20 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_31 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_18_108 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_42 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_26_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_64 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_97 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_86 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_75 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_174 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_17_196 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_32_144 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_32_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_32_188 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmux_left_track_5.mux_l2_in_0_ mux_left_track_5.mux_l1_in_1_/X mux_left_track_5.mux_l1_in_0_/X
+ mux_left_track_5.mux_l2_in_1_/S VGND VGND VPWR VPWR mux_left_track_5.mux_l2_in_0_/X
+ sky130_fd_sc_hd__mux2_1
XFILLER_23_199 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_11_99 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_14_122 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_14_144 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_14_155 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_14_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xinput16 chanx_left_in[4] VGND VGND VPWR VPWR _104_/A sky130_fd_sc_hd__buf_1
Xinput49 left_bottom_grid_pin_7_ VGND VGND VPWR VPWR input49/X sky130_fd_sc_hd__clkbuf_2
Xinput38 chany_top_in[6] VGND VGND VPWR VPWR input38/X sky130_fd_sc_hd__clkbuf_1
Xinput27 chany_top_in[14] VGND VGND VPWR VPWR input27/X sky130_fd_sc_hd__clkbuf_1
XFILLER_20_158 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_input38_A chany_top_in[6] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xmux_left_track_5.mux_l1_in_1_ input50/X input48/X mux_left_track_5.mux_l1_in_2_/S
+ VGND VGND VPWR VPWR mux_left_track_5.mux_l1_in_1_/X sky130_fd_sc_hd__mux2_1
XFILLER_8_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_10_180 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_33_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_25_206 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_17_10 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmux_top_track_20.sky130_fd_sc_hd__buf_4_0_ mux_top_track_20.mux_l2_in_0_/X VGND VGND
+ VPWR VPWR _098_/A sky130_fd_sc_hd__clkbuf_1
XFILLER_33_86 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xmem_left_track_33.sky130_fd_sc_hd__dfxtp_1_1_ clkbuf_3_2_0_mem_left_track_1.prog_clk/X
+ mux_left_track_33.mux_l1_in_0_/S VGND VGND VPWR VPWR mux_left_track_33.mux_l2_in_0_/S
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_146 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xmux_top_track_14.sky130_fd_sc_hd__buf_4_0_ mux_top_track_14.mux_l2_in_0_/X VGND VGND
+ VPWR VPWR _095_/A sky130_fd_sc_hd__clkbuf_1
Xmux_top_track_18.mux_l1_in_0_ input4/X input56/X mux_top_track_18.mux_l1_in_0_/S
+ VGND VGND VPWR VPWR mux_top_track_18.mux_l1_in_0_/X sky130_fd_sc_hd__mux2_1
XFILLER_14_66 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_30_87 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_input20_A chanx_left_in[8] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_29_172 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmux_top_track_20.mux_l1_in_0_ input3/X input57/X mux_top_track_20.mux_l1_in_0_/S
+ VGND VGND VPWR VPWR mux_top_track_20.mux_l1_in_0_/X sky130_fd_sc_hd__mux2_1
XFILLER_27_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_98 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_10 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_87 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_76 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_43 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_25_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_26_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_25_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xmux_left_track_13.mux_l1_in_0_ input48/X input27/X mux_left_track_13.mux_l1_in_0_/S
+ VGND VGND VPWR VPWR mux_left_track_13.mux_l1_in_0_/X sky130_fd_sc_hd__mux2_1
XFILLER_32_134 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmux_left_track_25.mux_l2_in_0_ mux_left_track_25.mux_l1_in_1_/X mux_left_track_25.mux_l1_in_0_/X
+ mux_left_track_25.mux_l2_in_0_/S VGND VGND VPWR VPWR mux_left_track_25.mux_l2_in_0_/X
+ sky130_fd_sc_hd__mux2_1
XFILLER_23_112 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_11_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_14_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_14_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xinput17 chanx_left_in[5] VGND VGND VPWR VPWR _103_/A sky130_fd_sc_hd__buf_1
Xinput39 chany_top_in[7] VGND VGND VPWR VPWR input39/X sky130_fd_sc_hd__clkbuf_1
Xinput28 chany_top_in[15] VGND VGND VPWR VPWR input28/X sky130_fd_sc_hd__clkbuf_1
XFILLER_9_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_20_115 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_20_126 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_11_115 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_22_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmux_left_track_5.mux_l1_in_0_ input46/X input31/X mux_left_track_5.mux_l1_in_2_/S
+ VGND VGND VPWR VPWR mux_left_track_5.mux_l1_in_0_/X sky130_fd_sc_hd__mux2_1
XFILLER_10_192 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xmux_left_track_25.mux_l1_in_1_ _064_/HI input45/X mux_left_track_25.mux_l1_in_1_/S
+ VGND VGND VPWR VPWR mux_left_track_25.mux_l1_in_1_/X sky130_fd_sc_hd__mux2_1
X_089_ _089_/A VGND VGND VPWR VPWR _089_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_26_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_25_218 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_17_33 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_17_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_17_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_33_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_33_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmem_left_track_33.sky130_fd_sc_hd__dfxtp_1_0_ clkbuf_3_2_0_mem_left_track_1.prog_clk/X
+ mux_left_track_31.mux_l2_in_0_/S VGND VGND VPWR VPWR mux_left_track_33.mux_l1_in_0_/S
+ sky130_fd_sc_hd__dfxtp_1
XANTENNA_input50_A left_bottom_grid_pin_9_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_30_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_21_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_158 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_28_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_12_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_28_87 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_28_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_5_58 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_5_14 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_10_6 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_5_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_input13_A chanx_left_in[1] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xclkbuf_2_1_0_mem_left_track_1.prog_clk clkbuf_2_1_0_mem_left_track_1.prog_clk/A VGND
+ VGND VPWR VPWR clkbuf_3_3_0_mem_left_track_1.prog_clk/A sky130_fd_sc_hd__clkbuf_1
XFILLER_29_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmem_left_track_39.sky130_fd_sc_hd__dfxtp_1_1_ clkbuf_3_2_0_mem_left_track_1.prog_clk/X
+ mux_left_track_39.mux_l1_in_0_/S VGND VGND VPWR VPWR output60/A sky130_fd_sc_hd__dfxtp_1
XANTENNA_input5_A chanx_left_in[12] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_26_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_99 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_88 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_77 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_22 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_33 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_66 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_1_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_2_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_32_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_23_146 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_23_157 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xinput18 chanx_left_in[6] VGND VGND VPWR VPWR _102_/A sky130_fd_sc_hd__buf_1
Xinput29 chany_top_in[16] VGND VGND VPWR VPWR input29/X sky130_fd_sc_hd__buf_1
XFILLER_9_172 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_20_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_11_127 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_22_78 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_22_89 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xmux_left_track_25.mux_l1_in_0_ input46/X input40/X mux_left_track_25.mux_l1_in_1_/S
+ VGND VGND VPWR VPWR mux_left_track_25.mux_l1_in_0_/X sky130_fd_sc_hd__mux2_1
X_088_ _088_/A VGND VGND VPWR VPWR _088_/X sky130_fd_sc_hd__clkbuf_1
Xmux_left_track_37.mux_l2_in_0_ _037_/HI mux_left_track_37.mux_l1_in_0_/X mux_left_track_37.mux_l2_in_0_/S
+ VGND VGND VPWR VPWR mux_left_track_37.mux_l2_in_0_/X sky130_fd_sc_hd__mux2_1
Xmem_top_track_14.sky130_fd_sc_hd__dfxtp_1_1_ clkbuf_3_4_0_mem_left_track_1.prog_clk/X
+ mux_top_track_14.mux_l1_in_0_/S VGND VGND VPWR VPWR mux_top_track_14.mux_l2_in_0_/S
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_33_99 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_33_88 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_33_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_input43_A left_bottom_grid_pin_13_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mux_top_track_20.mux_l1_in_0__A0 input3/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_5_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xmux_top_track_8.mux_l2_in_0_ mux_top_track_8.mux_l1_in_1_/X mux_top_track_8.mux_l1_in_0_/X
+ mux_top_track_8.mux_l2_in_0_/S VGND VGND VPWR VPWR mux_top_track_8.mux_l2_in_0_/X
+ sky130_fd_sc_hd__mux2_1
XANTENNA_mux_top_track_12.mux_l1_in_0__A1 input53/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_14_24 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_30_67 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_30_78 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmem_left_track_39.sky130_fd_sc_hd__dfxtp_1_0_ clkbuf_3_2_0_mem_left_track_1.prog_clk/X
+ mux_left_track_37.mux_l2_in_0_/S VGND VGND VPWR VPWR mux_left_track_39.mux_l1_in_0_/S
+ sky130_fd_sc_hd__dfxtp_1
XANTENNA_mux_top_track_4.mux_l1_in_0__A0 input53/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_12 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_67 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_89 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_78 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_23 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_34 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_45 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_25_34 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xmux_top_track_8.mux_l1_in_1_ _055_/HI input9/X mux_top_track_8.mux_l1_in_1_/S VGND
+ VGND VPWR VPWR mux_top_track_8.mux_l1_in_1_/X sky130_fd_sc_hd__mux2_1
XFILLER_17_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xmux_top_track_8.sky130_fd_sc_hd__buf_4_0_ mux_top_track_8.mux_l2_in_0_/X VGND VGND
+ VPWR VPWR _092_/A sky130_fd_sc_hd__clkbuf_1
XFILLER_32_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_23_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_11_58 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_2_9 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xinput19 chanx_left_in[7] VGND VGND VPWR VPWR input19/X sky130_fd_sc_hd__buf_1
XFILLER_9_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_9_151 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_3_70 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_11_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_087_ _087_/A VGND VGND VPWR VPWR _087_/X sky130_fd_sc_hd__clkbuf_1
Xmem_top_track_14.sky130_fd_sc_hd__dfxtp_1_0_ clkbuf_3_4_0_mem_left_track_1.prog_clk/X
+ mux_top_track_12.mux_l2_in_0_/S VGND VGND VPWR VPWR mux_top_track_14.mux_l1_in_0_/S
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_33_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_33_45 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_input36_A chany_top_in[4] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_30_201 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_31_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_71 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_0_127 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_28_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_12_201 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_mux_left_track_13.mux_l1_in_0__A0 input48/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_5_38 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xmux_left_track_37.mux_l1_in_0_ input43/X input34/X mux_left_track_37.mux_l1_in_0_/S
+ VGND VGND VPWR VPWR mux_left_track_37.mux_l1_in_0_/X sky130_fd_sc_hd__mux2_1
XFILLER_5_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_30_35 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_mux_top_track_4.mux_l1_in_0__A1 input51/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_13 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_24 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_35 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_46 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_25_24 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_68 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_79 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_25_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xmux_top_track_8.mux_l1_in_0_ input59/X input51/X mux_top_track_8.mux_l1_in_1_/S VGND
+ VGND VPWR VPWR mux_top_track_8.mux_l1_in_0_/X sky130_fd_sc_hd__mux2_1
XFILLER_32_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_15_90 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_31_192 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_11_48 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_14_126 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_28_9 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_9_163 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_3_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_6_144 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_6_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_086_ _086_/A VGND VGND VPWR VPWR _086_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_19_5 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_33_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_33_210 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xmux_left_track_3.sky130_fd_sc_hd__buf_4_0_ mux_left_track_3.mux_l3_in_0_/X VGND VGND
+ VPWR VPWR _069_/A sky130_fd_sc_hd__clkbuf_1
XANTENNA_mux_left_track_21.mux_l1_in_0__A0 input43/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_17_58 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_17_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_24_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_input29_A chany_top_in[16] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_30_213 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_069_ _069_/A VGND VGND VPWR VPWR _069_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_2_180 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_24_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_28_35 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_8_206 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_12_213 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_30_25 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_30_58 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_14 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_69 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_25 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_36 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_47 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_25_14 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_25_58 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_26_146 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_26_179 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_58 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_17_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_input11_A chanx_left_in[18] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_15_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xoutput90 _106_/X VGND VGND VPWR VPWR chany_top_out[18] sky130_fd_sc_hd__clkbuf_2
XFILLER_31_182 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_input3_A chanx_left_in[10] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mux_left_track_1.mux_l1_in_2__A1 input43/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xmux_left_track_13.sky130_fd_sc_hd__buf_4_0_ mux_left_track_13.mux_l2_in_0_/X VGND
+ VGND VPWR VPWR _074_/A sky130_fd_sc_hd__clkbuf_1
XFILLER_14_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_14_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_22_171 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_input59_A top_right_grid_pin_1_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_3_94 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_22_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_22_48 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_8_28 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_6_156 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_6_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_12_92 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmem_left_track_25.sky130_fd_sc_hd__dfxtp_1_1_ clkbuf_3_0_0_mem_left_track_1.prog_clk/X
+ mux_left_track_25.mux_l1_in_1_/S VGND VGND VPWR VPWR mux_left_track_25.mux_l2_in_0_/S
+ sky130_fd_sc_hd__dfxtp_1
X_085_ _085_/A VGND VGND VPWR VPWR _085_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_33_200 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_17_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_17_48 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xmux_left_track_1.mux_l3_in_0_ mux_left_track_1.mux_l2_in_1_/X mux_left_track_1.mux_l2_in_0_/X
+ mux_left_track_1.mux_l3_in_0_/S VGND VGND VPWR VPWR mux_left_track_1.mux_l3_in_0_/X
+ sky130_fd_sc_hd__mux2_1
XFILLER_3_115 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_15_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_2_192 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_068_ _068_/A VGND VGND VPWR VPWR _068_/X sky130_fd_sc_hd__clkbuf_1
XANTENNA_mux_top_track_6.mux_l1_in_1__A0 input58/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_9_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_input41_A chany_top_in[9] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xmux_left_track_1.mux_l2_in_1_ _056_/HI mux_left_track_1.mux_l1_in_2_/X mux_left_track_1.mux_l2_in_1_/S
+ VGND VGND VPWR VPWR mux_left_track_1.mux_l2_in_1_/X sky130_fd_sc_hd__mux2_1
XFILLER_30_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_29_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_4_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_26_103 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_37 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_48 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_59 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_2_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_32_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xmux_left_track_1.mux_l1_in_2_ input45/X input43/X mux_left_track_1.mux_l1_in_2_/S
+ VGND VGND VPWR VPWR mux_left_track_1.mux_l1_in_2_/X sky130_fd_sc_hd__mux2_1
XFILLER_31_91 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xoutput91 _107_/X VGND VGND VPWR VPWR chany_top_out[19] sky130_fd_sc_hd__clkbuf_2
Xoutput80 _077_/X VGND VGND VPWR VPWR chanx_left_out[9] sky130_fd_sc_hd__clkbuf_2
XFILLER_16_180 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_23_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_23_128 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_31_172 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmux_top_track_14.mux_l2_in_0_ _045_/HI mux_top_track_14.mux_l1_in_0_/X mux_top_track_14.mux_l2_in_0_/S
+ VGND VGND VPWR VPWR mux_top_track_14.mux_l2_in_0_/X sky130_fd_sc_hd__mux2_1
XFILLER_9_198 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_13_172 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_22_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_9 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_10_142 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_6_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xmux_left_track_35.sky130_fd_sc_hd__buf_4_0_ mux_left_track_35.mux_l2_in_0_/X VGND
+ VGND VPWR VPWR _085_/A sky130_fd_sc_hd__clkbuf_1
XFILLER_6_168 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xmem_left_track_25.sky130_fd_sc_hd__dfxtp_1_0_ clkbuf_3_0_0_mem_left_track_1.prog_clk/X
+ mux_left_track_23.mux_l2_in_0_/S VGND VGND VPWR VPWR mux_left_track_25.mux_l1_in_1_/S
+ sky130_fd_sc_hd__dfxtp_1
X_084_ _084_/A VGND VGND VPWR VPWR _084_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_33_9 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_mux_left_track_39.mux_l2_in_0__S output60/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_24_201 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_33_59 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_33_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_3_127 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xclkbuf_1_1_0_mem_left_track_1.prog_clk clkbuf_0_mem_left_track_1.prog_clk/X VGND
+ VGND VPWR VPWR clkbuf_2_3_0_mem_left_track_1.prog_clk/A sky130_fd_sc_hd__clkbuf_1
X_067_ VGND VGND VPWR VPWR _067_/HI _067_/LO sky130_fd_sc_hd__conb_1
XANTENNA_mux_left_track_5.mux_l1_in_1__A0 input50/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mux_top_track_6.mux_l1_in_1__A1 input56/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xmux_left_track_29.sky130_fd_sc_hd__buf_4_0_ mux_left_track_29.mux_l2_in_0_/X VGND
+ VGND VPWR VPWR _082_/A sky130_fd_sc_hd__clkbuf_1
XFILLER_28_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_input34_A chany_top_in[2] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xmux_left_track_1.mux_l2_in_0_ mux_left_track_1.mux_l1_in_1_/X mux_left_track_1.mux_l1_in_0_/X
+ mux_left_track_1.mux_l2_in_1_/S VGND VGND VPWR VPWR mux_left_track_1.mux_l2_in_0_/X
+ sky130_fd_sc_hd__mux2_1
XFILLER_14_28 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_29_112 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_29_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_20_60 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_mux_top_track_18.mux_l1_in_0__A0 input4/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_26_126 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_26_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_16 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_38 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_49 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_9_6 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_32_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmux_left_track_1.mux_l1_in_1_ input50/X input48/X mux_left_track_1.mux_l1_in_2_/S
+ VGND VGND VPWR VPWR mux_left_track_1.mux_l1_in_1_/X sky130_fd_sc_hd__mux2_1
Xoutput70 _086_/X VGND VGND VPWR VPWR chanx_left_out[18] sky130_fd_sc_hd__clkbuf_2
Xoutput92 _089_/X VGND VGND VPWR VPWR chany_top_out[1] sky130_fd_sc_hd__clkbuf_2
Xoutput81 _088_/X VGND VGND VPWR VPWR chany_top_out[0] sky130_fd_sc_hd__clkbuf_2
XFILLER_16_192 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_31_151 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_11_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_14_118 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_13_151 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_13_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_3_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xmux_top_track_10.sky130_fd_sc_hd__buf_4_0_ mux_top_track_10.mux_l2_in_0_/X VGND VGND
+ VPWR VPWR _093_/A sky130_fd_sc_hd__clkbuf_1
XFILLER_27_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_10_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_12_50 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_083_ _083_/A VGND VGND VPWR VPWR _083_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_18_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_26_9 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmem_top_track_2.sky130_fd_sc_hd__dfxtp_1_2_ clkbuf_3_7_0_mem_left_track_1.prog_clk/X
+ mux_top_track_2.mux_l2_in_1_/S VGND VGND VPWR VPWR mux_top_track_2.mux_l3_in_0_/S
+ sky130_fd_sc_hd__dfxtp_1
Xmux_top_track_14.mux_l1_in_0_ input6/X input54/X mux_top_track_14.mux_l1_in_0_/S
+ VGND VGND VPWR VPWR mux_top_track_14.mux_l1_in_0_/X sky130_fd_sc_hd__mux2_1
XFILLER_24_213 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_33_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_3_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_3_106 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_15_202 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xmux_top_track_26.mux_l2_in_0_ _052_/HI mux_top_track_26.mux_l1_in_0_/X mux_top_track_26.mux_l2_in_0_/S
+ VGND VGND VPWR VPWR mux_top_track_26.mux_l2_in_0_/X sky130_fd_sc_hd__mux2_1
X_066_ VGND VGND VPWR VPWR _066_/HI _066_/LO sky130_fd_sc_hd__conb_1
XFILLER_17_5 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_mux_left_track_5.mux_l1_in_1__A1 input48/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_28_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmux_left_track_19.mux_l2_in_0_ _061_/HI mux_left_track_19.mux_l1_in_0_/X mux_left_track_19.mux_l2_in_0_/S
+ VGND VGND VPWR VPWR mux_left_track_19.mux_l2_in_0_/X sky130_fd_sc_hd__mux2_1
XFILLER_18_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_input27_A chany_top_in[14] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_049_ VGND VGND VPWR VPWR _049_/HI _049_/LO sky130_fd_sc_hd__conb_1
XFILLER_22_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmux_left_track_21.mux_l2_in_0_ _062_/HI mux_left_track_21.mux_l1_in_0_/X mux_left_track_21.mux_l2_in_0_/S
+ VGND VGND VPWR VPWR mux_left_track_21.mux_l2_in_0_/X sky130_fd_sc_hd__mux2_1
XFILLER_29_157 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_29_168 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_4_201 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_mux_top_track_18.mux_l1_in_0__A1 input56/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_29_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_6_30 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_17 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_28 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xmux_left_track_1.mux_l1_in_0_ input46/X input22/X mux_left_track_1.mux_l1_in_2_/S
+ VGND VGND VPWR VPWR mux_left_track_1.mux_l1_in_0_/X sky130_fd_sc_hd__mux2_1
Xoutput82 _098_/X VGND VGND VPWR VPWR chany_top_out[10] sky130_fd_sc_hd__clkbuf_2
Xoutput93 _090_/X VGND VGND VPWR VPWR chany_top_out[2] sky130_fd_sc_hd__clkbuf_2
Xoutput71 _087_/X VGND VGND VPWR VPWR chanx_left_out[19] sky130_fd_sc_hd__clkbuf_2
Xoutput60 output60/A VGND VGND VPWR VPWR ccff_tail sky130_fd_sc_hd__clkbuf_2
XFILLER_31_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_31_163 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmux_top_track_4.mux_l3_in_0_ mux_top_track_4.mux_l2_in_1_/X mux_top_track_4.mux_l2_in_0_/X
+ mux_top_track_4.mux_l3_in_0_/S VGND VGND VPWR VPWR mux_top_track_4.mux_l3_in_0_/X
+ sky130_fd_sc_hd__mux2_1
XFILLER_22_130 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_22_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_13_163 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_13_196 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_3_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_input1_A ccff_head VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xmem_left_track_5.sky130_fd_sc_hd__dfxtp_1_2_ clkbuf_3_1_0_mem_left_track_1.prog_clk/X
+ mux_left_track_5.mux_l2_in_1_/S VGND VGND VPWR VPWR mux_left_track_5.mux_l3_in_0_/S
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_10_144 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_10_122 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_12_40 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_12_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_082_ _082_/A VGND VGND VPWR VPWR _082_/X sky130_fd_sc_hd__clkbuf_1
XANTENNA_input57_A top_left_grid_pin_48_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xmux_top_track_4.mux_l2_in_1_ _053_/HI mux_top_track_4.mux_l1_in_2_/X mux_top_track_4.mux_l2_in_1_/S
+ VGND VGND VPWR VPWR mux_top_track_4.mux_l2_in_1_/X sky130_fd_sc_hd__mux2_1
Xmem_top_track_2.sky130_fd_sc_hd__dfxtp_1_1_ clkbuf_3_6_0_mem_left_track_1.prog_clk/X
+ mux_top_track_2.mux_l1_in_1_/S VGND VGND VPWR VPWR mux_top_track_2.mux_l2_in_1_/S
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_15_214 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_065_ VGND VGND VPWR VPWR _065_/HI _065_/LO sky130_fd_sc_hd__conb_1
XFILLER_23_94 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_9_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_9_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_9_63 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_9_52 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_28_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_mux_top_track_26.mux_l1_in_0__A1 input52/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xmux_top_track_4.mux_l1_in_2_ input11/X input59/X mux_top_track_4.mux_l1_in_2_/S VGND
+ VGND VPWR VPWR mux_top_track_4.mux_l1_in_2_/X sky130_fd_sc_hd__mux2_1
XFILLER_7_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmux_top_track_26.sky130_fd_sc_hd__buf_4_0_ mux_top_track_26.mux_l2_in_0_/X VGND VGND
+ VPWR VPWR _101_/A sky130_fd_sc_hd__clkbuf_1
X_048_ VGND VGND VPWR VPWR _048_/HI _048_/LO sky130_fd_sc_hd__conb_1
XANTENNA_mux_left_track_19.mux_l1_in_0__A0 input42/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xmux_top_track_26.mux_l1_in_0_ input19/X input52/X mux_top_track_26.mux_l1_in_0_/S
+ VGND VGND VPWR VPWR mux_top_track_26.mux_l1_in_0_/X sky130_fd_sc_hd__mux2_1
XFILLER_29_103 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_4_213 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_20_73 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_20_84 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmem_left_track_11.sky130_fd_sc_hd__dfxtp_1_1_ clkbuf_3_3_0_mem_left_track_1.prog_clk/X
+ mux_left_track_11.mux_l1_in_0_/S VGND VGND VPWR VPWR mux_left_track_11.mux_l2_in_0_/S
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_29_60 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_29_71 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_6_42 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_18 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xclkbuf_3_0_0_mem_left_track_1.prog_clk clkbuf_3_1_0_mem_left_track_1.prog_clk/A VGND
+ VGND VPWR VPWR clkbuf_3_0_0_mem_left_track_1.prog_clk/X sky130_fd_sc_hd__clkbuf_1
XFILLER_25_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmux_left_track_19.mux_l1_in_0_ input42/X input24/X mux_left_track_19.mux_l1_in_0_/S
+ VGND VGND VPWR VPWR mux_left_track_19.mux_l1_in_0_/X sky130_fd_sc_hd__mux2_1
XFILLER_17_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_17_128 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_17_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_25_172 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_25_183 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_15_95 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xoutput83 _099_/X VGND VGND VPWR VPWR chany_top_out[11] sky130_fd_sc_hd__clkbuf_2
Xoutput94 _091_/X VGND VGND VPWR VPWR chany_top_out[3] sky130_fd_sc_hd__clkbuf_2
Xoutput61 _068_/X VGND VGND VPWR VPWR chanx_left_out[0] sky130_fd_sc_hd__clkbuf_2
Xoutput72 _069_/X VGND VGND VPWR VPWR chanx_left_out[1] sky130_fd_sc_hd__clkbuf_2
Xmux_left_track_21.mux_l1_in_0_ input43/X input23/X mux_left_track_21.mux_l1_in_0_/S
+ VGND VGND VPWR VPWR mux_left_track_21.mux_l1_in_0_/X sky130_fd_sc_hd__mux2_1
XFILLER_31_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmux_left_track_33.mux_l2_in_0_ _035_/HI mux_left_track_33.mux_l1_in_0_/X mux_left_track_33.mux_l2_in_0_/S
+ VGND VGND VPWR VPWR mux_left_track_33.mux_l2_in_0_/X sky130_fd_sc_hd__mux2_1
XFILLER_22_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_22_175 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_22_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_9_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_26_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xmem_left_track_5.sky130_fd_sc_hd__dfxtp_1_1_ clkbuf_3_0_0_mem_left_track_1.prog_clk/X
+ mux_left_track_5.mux_l1_in_2_/S VGND VGND VPWR VPWR mux_left_track_5.mux_l2_in_1_/S
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_10_134 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_10_156 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_12_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_12_96 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_081_ _081_/A VGND VGND VPWR VPWR _081_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_18_201 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_33_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_33_204 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmem_top_track_2.sky130_fd_sc_hd__dfxtp_1_0_ clkbuf_3_6_0_mem_left_track_1.prog_clk/X
+ mux_top_track_0.mux_l3_in_0_/S VGND VGND VPWR VPWR mux_top_track_2.mux_l1_in_1_/S
+ sky130_fd_sc_hd__dfxtp_1
Xmux_top_track_4.mux_l2_in_0_ mux_top_track_4.mux_l1_in_1_/X mux_top_track_4.mux_l1_in_0_/X
+ mux_top_track_4.mux_l2_in_1_/S VGND VGND VPWR VPWR mux_top_track_4.mux_l2_in_0_/X
+ sky130_fd_sc_hd__mux2_1
Xmux_top_track_4.sky130_fd_sc_hd__buf_4_0_ mux_top_track_4.mux_l3_in_0_/X VGND VGND
+ VPWR VPWR _090_/A sky130_fd_sc_hd__clkbuf_1
X_064_ VGND VGND VPWR VPWR _064_/HI _064_/LO sky130_fd_sc_hd__conb_1
XFILLER_31_9 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_0_88 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xclkbuf_3_3_0_mem_left_track_1.prog_clk clkbuf_3_3_0_mem_left_track_1.prog_clk/A VGND
+ VGND VPWR VPWR clkbuf_3_3_0_mem_left_track_1.prog_clk/X sky130_fd_sc_hd__clkbuf_1
Xmux_top_track_4.mux_l1_in_1_ input57/X input55/X mux_top_track_4.mux_l1_in_2_/S VGND
+ VGND VPWR VPWR mux_top_track_4.mux_l1_in_1_/X sky130_fd_sc_hd__mux2_1
XFILLER_18_84 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__105__A _105_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_047_ VGND VGND VPWR VPWR _047_/HI _047_/LO sky130_fd_sc_hd__conb_1
Xmem_top_track_8.sky130_fd_sc_hd__dfxtp_1_1_ clkbuf_3_1_0_mem_left_track_1.prog_clk/X
+ mux_top_track_8.mux_l1_in_1_/S VGND VGND VPWR VPWR mux_top_track_8.mux_l2_in_0_/S
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_29_115 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_29_126 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_29_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xmem_left_track_11.sky130_fd_sc_hd__dfxtp_1_0_ clkbuf_3_1_0_mem_left_track_1.prog_clk/X
+ mux_left_track_9.mux_l2_in_0_/S VGND VGND VPWR VPWR mux_left_track_11.mux_l1_in_0_/S
+ sky130_fd_sc_hd__dfxtp_1
XANTENNA_input32_A chany_top_in[19] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_6_87 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_6_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_6_10 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_25_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmem_top_track_24.sky130_fd_sc_hd__dfxtp_1_1_ clkbuf_3_5_0_mem_left_track_1.prog_clk/X
+ mux_top_track_24.mux_l1_in_1_/S VGND VGND VPWR VPWR mux_top_track_24.mux_l2_in_0_/S
+ sky130_fd_sc_hd__dfxtp_1
Xoutput84 _100_/X VGND VGND VPWR VPWR chany_top_out[12] sky130_fd_sc_hd__clkbuf_2
Xoutput95 _092_/X VGND VGND VPWR VPWR chany_top_out[4] sky130_fd_sc_hd__clkbuf_2
Xoutput73 _070_/X VGND VGND VPWR VPWR chanx_left_out[2] sky130_fd_sc_hd__clkbuf_2
Xoutput62 _078_/X VGND VGND VPWR VPWR chanx_left_out[10] sky130_fd_sc_hd__clkbuf_2
XFILLER_16_162 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_190 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_31_132 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_31_187 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_7_6 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_26_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmem_left_track_17.sky130_fd_sc_hd__dfxtp_1_1_ clkbuf_3_3_0_mem_left_track_1.prog_clk/X
+ mux_left_track_17.mux_l1_in_0_/S VGND VGND VPWR VPWR mux_left_track_17.mux_l2_in_0_/S
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_8_180 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xmem_left_track_5.sky130_fd_sc_hd__dfxtp_1_0_ clkbuf_3_0_0_mem_left_track_1.prog_clk/X
+ mux_left_track_3.mux_l3_in_0_/S VGND VGND VPWR VPWR mux_left_track_5.mux_l1_in_2_/S
+ sky130_fd_sc_hd__dfxtp_1
XANTENNA_mux_left_track_35.mux_l1_in_0__A0 input42/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_10_168 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_12_20 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_080_ _080_/A VGND VGND VPWR VPWR _080_/X sky130_fd_sc_hd__clkbuf_1
Xclkbuf_3_6_0_mem_left_track_1.prog_clk clkbuf_3_7_0_mem_left_track_1.prog_clk/A VGND
+ VGND VPWR VPWR clkbuf_3_6_0_mem_left_track_1.prog_clk/X sky130_fd_sc_hd__clkbuf_1
Xmux_left_track_33.mux_l1_in_0_ input50/X input36/X mux_left_track_33.mux_l1_in_0_/S
+ VGND VGND VPWR VPWR mux_left_track_33.mux_l1_in_0_/X sky130_fd_sc_hd__mux2_1
XFILLER_5_172 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_063_ VGND VGND VPWR VPWR _063_/HI _063_/LO sky130_fd_sc_hd__conb_1
XFILLER_0_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_24_9 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_18_30 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmux_top_track_4.mux_l1_in_0_ input53/X input51/X mux_top_track_4.mux_l1_in_2_/S VGND
+ VGND VPWR VPWR mux_top_track_4.mux_l1_in_0_/X sky130_fd_sc_hd__mux2_1
X_046_ VGND VGND VPWR VPWR _046_/HI _046_/LO sky130_fd_sc_hd__conb_1
XFILLER_15_5 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmem_top_track_8.sky130_fd_sc_hd__dfxtp_1_0_ clkbuf_3_4_0_mem_left_track_1.prog_clk/X
+ mux_top_track_6.mux_l3_in_0_/S VGND VGND VPWR VPWR mux_top_track_8.mux_l1_in_1_/S
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_28_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_input25_A chany_top_in[12] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_6_99 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_6_66 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_6_22 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_20_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_15_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xmem_top_track_24.sky130_fd_sc_hd__dfxtp_1_0_ clkbuf_3_5_0_mem_left_track_1.prog_clk/X
+ mux_top_track_22.mux_l2_in_0_/S VGND VGND VPWR VPWR mux_top_track_24.mux_l1_in_1_/S
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_31_63 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_31_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xoutput85 _101_/X VGND VGND VPWR VPWR chany_top_out[13] sky130_fd_sc_hd__clkbuf_2
Xoutput74 _071_/X VGND VGND VPWR VPWR chanx_left_out[3] sky130_fd_sc_hd__clkbuf_2
Xoutput63 _079_/X VGND VGND VPWR VPWR chanx_left_out[11] sky130_fd_sc_hd__clkbuf_2
Xoutput96 _093_/X VGND VGND VPWR VPWR chany_top_out[5] sky130_fd_sc_hd__clkbuf_2
XFILLER_16_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_31_122 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_191 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_180 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_31_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
.ends

